VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_256x64m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_256x64m4w8   ;
    SIZE 690.120 BY 291.640 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 286.710 0.000 286.850 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 292.810 0.000 292.950 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 298.910 0.000 299.050 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 305.010 0.000 305.150 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 311.110 0.000 311.250 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 317.210 0.000 317.350 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 323.310 0.000 323.450 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 329.410 0.000 329.550 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 335.510 0.000 335.650 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 341.610 0.000 341.750 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 347.710 0.000 347.850 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 353.810 0.000 353.950 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 359.910 0.000 360.050 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 366.010 0.000 366.150 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 372.110 0.000 372.250 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 378.210 0.000 378.350 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 384.310 0.000 384.450 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 390.410 0.000 390.550 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 396.510 0.000 396.650 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 402.610 0.000 402.750 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 408.710 0.000 408.850 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 414.810 0.000 414.950 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 420.910 0.000 421.050 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 427.010 0.000 427.150 0.140 ; 
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 433.110 0.000 433.250 0.140 ; 
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 439.210 0.000 439.350 0.140 ; 
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 445.310 0.000 445.450 0.140 ; 
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 451.410 0.000 451.550 0.140 ; 
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 457.510 0.000 457.650 0.140 ; 
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 463.610 0.000 463.750 0.140 ; 
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 469.710 0.000 469.850 0.140 ; 
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 475.810 0.000 475.950 0.140 ; 
        END 
    END dout[31] 
    PIN dout[32] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 481.910 0.000 482.050 0.140 ; 
        END 
    END dout[32] 
    PIN dout[33] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 488.010 0.000 488.150 0.140 ; 
        END 
    END dout[33] 
    PIN dout[34] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 494.110 0.000 494.250 0.140 ; 
        END 
    END dout[34] 
    PIN dout[35] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 500.210 0.000 500.350 0.140 ; 
        END 
    END dout[35] 
    PIN dout[36] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 506.310 0.000 506.450 0.140 ; 
        END 
    END dout[36] 
    PIN dout[37] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 512.410 0.000 512.550 0.140 ; 
        END 
    END dout[37] 
    PIN dout[38] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 518.510 0.000 518.650 0.140 ; 
        END 
    END dout[38] 
    PIN dout[39] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 524.610 0.000 524.750 0.140 ; 
        END 
    END dout[39] 
    PIN dout[40] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 530.710 0.000 530.850 0.140 ; 
        END 
    END dout[40] 
    PIN dout[41] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 536.810 0.000 536.950 0.140 ; 
        END 
    END dout[41] 
    PIN dout[42] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 542.910 0.000 543.050 0.140 ; 
        END 
    END dout[42] 
    PIN dout[43] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 549.010 0.000 549.150 0.140 ; 
        END 
    END dout[43] 
    PIN dout[44] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 555.110 0.000 555.250 0.140 ; 
        END 
    END dout[44] 
    PIN dout[45] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 561.210 0.000 561.350 0.140 ; 
        END 
    END dout[45] 
    PIN dout[46] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 567.310 0.000 567.450 0.140 ; 
        END 
    END dout[46] 
    PIN dout[47] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 573.410 0.000 573.550 0.140 ; 
        END 
    END dout[47] 
    PIN dout[48] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 579.510 0.000 579.650 0.140 ; 
        END 
    END dout[48] 
    PIN dout[49] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 585.610 0.000 585.750 0.140 ; 
        END 
    END dout[49] 
    PIN dout[50] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 591.710 0.000 591.850 0.140 ; 
        END 
    END dout[50] 
    PIN dout[51] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 597.810 0.000 597.950 0.140 ; 
        END 
    END dout[51] 
    PIN dout[52] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 603.910 0.000 604.050 0.140 ; 
        END 
    END dout[52] 
    PIN dout[53] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 610.010 0.000 610.150 0.140 ; 
        END 
    END dout[53] 
    PIN dout[54] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 616.110 0.000 616.250 0.140 ; 
        END 
    END dout[54] 
    PIN dout[55] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 622.210 0.000 622.350 0.140 ; 
        END 
    END dout[55] 
    PIN dout[56] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 628.310 0.000 628.450 0.140 ; 
        END 
    END dout[56] 
    PIN dout[57] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 634.410 0.000 634.550 0.140 ; 
        END 
    END dout[57] 
    PIN dout[58] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 640.510 0.000 640.650 0.140 ; 
        END 
    END dout[58] 
    PIN dout[59] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 646.610 0.000 646.750 0.140 ; 
        END 
    END dout[59] 
    PIN dout[60] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 652.710 0.000 652.850 0.140 ; 
        END 
    END dout[60] 
    PIN dout[61] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 658.810 0.000 658.950 0.140 ; 
        END 
    END dout[61] 
    PIN dout[62] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 664.910 0.000 665.050 0.140 ; 
        END 
    END dout[62] 
    PIN dout[63] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 671.010 0.000 671.150 0.140 ; 
        END 
    END dout[63] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 286.290 0.000 286.430 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 292.390 0.000 292.530 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 298.490 0.000 298.630 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 304.590 0.000 304.730 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 310.690 0.000 310.830 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 316.790 0.000 316.930 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 322.890 0.000 323.030 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 328.990 0.000 329.130 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 335.090 0.000 335.230 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 341.190 0.000 341.330 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 347.290 0.000 347.430 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 353.390 0.000 353.530 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 359.490 0.000 359.630 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 365.590 0.000 365.730 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 371.690 0.000 371.830 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 377.790 0.000 377.930 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 383.890 0.000 384.030 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 389.990 0.000 390.130 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 396.090 0.000 396.230 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 402.190 0.000 402.330 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 408.290 0.000 408.430 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 414.390 0.000 414.530 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 420.490 0.000 420.630 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 426.590 0.000 426.730 0.140 ; 
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 432.690 0.000 432.830 0.140 ; 
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 438.790 0.000 438.930 0.140 ; 
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 444.890 0.000 445.030 0.140 ; 
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 450.990 0.000 451.130 0.140 ; 
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 457.090 0.000 457.230 0.140 ; 
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 463.190 0.000 463.330 0.140 ; 
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 469.290 0.000 469.430 0.140 ; 
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 475.390 0.000 475.530 0.140 ; 
        END 
    END din[31] 
    PIN din[32] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 481.490 0.000 481.630 0.140 ; 
        END 
    END din[32] 
    PIN din[33] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 487.590 0.000 487.730 0.140 ; 
        END 
    END din[33] 
    PIN din[34] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 493.690 0.000 493.830 0.140 ; 
        END 
    END din[34] 
    PIN din[35] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 499.790 0.000 499.930 0.140 ; 
        END 
    END din[35] 
    PIN din[36] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 505.890 0.000 506.030 0.140 ; 
        END 
    END din[36] 
    PIN din[37] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 511.990 0.000 512.130 0.140 ; 
        END 
    END din[37] 
    PIN din[38] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 518.090 0.000 518.230 0.140 ; 
        END 
    END din[38] 
    PIN din[39] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 524.190 0.000 524.330 0.140 ; 
        END 
    END din[39] 
    PIN din[40] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 530.290 0.000 530.430 0.140 ; 
        END 
    END din[40] 
    PIN din[41] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 536.390 0.000 536.530 0.140 ; 
        END 
    END din[41] 
    PIN din[42] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 542.490 0.000 542.630 0.140 ; 
        END 
    END din[42] 
    PIN din[43] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 548.590 0.000 548.730 0.140 ; 
        END 
    END din[43] 
    PIN din[44] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 554.690 0.000 554.830 0.140 ; 
        END 
    END din[44] 
    PIN din[45] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 560.790 0.000 560.930 0.140 ; 
        END 
    END din[45] 
    PIN din[46] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 566.890 0.000 567.030 0.140 ; 
        END 
    END din[46] 
    PIN din[47] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 572.990 0.000 573.130 0.140 ; 
        END 
    END din[47] 
    PIN din[48] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 579.090 0.000 579.230 0.140 ; 
        END 
    END din[48] 
    PIN din[49] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 585.190 0.000 585.330 0.140 ; 
        END 
    END din[49] 
    PIN din[50] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 591.290 0.000 591.430 0.140 ; 
        END 
    END din[50] 
    PIN din[51] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 597.390 0.000 597.530 0.140 ; 
        END 
    END din[51] 
    PIN din[52] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 603.490 0.000 603.630 0.140 ; 
        END 
    END din[52] 
    PIN din[53] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 609.590 0.000 609.730 0.140 ; 
        END 
    END din[53] 
    PIN din[54] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 615.690 0.000 615.830 0.140 ; 
        END 
    END din[54] 
    PIN din[55] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 621.790 0.000 621.930 0.140 ; 
        END 
    END din[55] 
    PIN din[56] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 627.890 0.000 628.030 0.140 ; 
        END 
    END din[56] 
    PIN din[57] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 633.990 0.000 634.130 0.140 ; 
        END 
    END din[57] 
    PIN din[58] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 640.090 0.000 640.230 0.140 ; 
        END 
    END din[58] 
    PIN din[59] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 646.190 0.000 646.330 0.140 ; 
        END 
    END din[59] 
    PIN din[60] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 652.290 0.000 652.430 0.140 ; 
        END 
    END din[60] 
    PIN din[61] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 658.390 0.000 658.530 0.140 ; 
        END 
    END din[61] 
    PIN din[62] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 664.490 0.000 664.630 0.140 ; 
        END 
    END din[62] 
    PIN din[63] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 670.590 0.000 670.730 0.140 ; 
        END 
    END din[63] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 285.940 0.000 286.080 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 334.740 0.000 334.880 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 383.540 0.000 383.680 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 432.340 0.000 432.480 0.140 ; 
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 481.140 0.000 481.280 0.140 ; 
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 529.940 0.000 530.080 0.140 ; 
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 578.740 0.000 578.880 0.140 ; 
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 627.540 0.000 627.680 0.140 ; 
        END 
    END wmask[7] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 244.600 0.000 244.920 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 238.480 0.000 238.800 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 232.360 0.000 232.680 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 226.240 0.000 226.560 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 220.120 0.000 220.440 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 214.000 0.000 214.320 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 207.880 0.000 208.200 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 201.760 0.000 202.080 0.320 ; 
        END 
    END addr[7] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 256.840 0.000 257.160 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.842300 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 250.720 0.000 251.040 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 41.292000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 259.560 0.000 259.880 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 45.198000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 260.240 0.000 260.560 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 285.720 6.240 ; 
                RECT 671.640 5.920 689.960 6.240 ; 
                RECT 0.160 7.280 689.960 7.600 ; 
                RECT 0.160 8.640 689.960 8.960 ; 
                RECT 0.160 10.000 259.200 10.320 ; 
                RECT 628.120 10.000 689.960 10.320 ; 
                RECT 0.160 11.360 275.520 11.680 ; 
                RECT 680.480 11.360 689.960 11.680 ; 
                RECT 0.160 12.720 275.520 13.040 ; 
                RECT 680.480 12.720 689.960 13.040 ; 
                RECT 0.160 14.080 198.000 14.400 ; 
                RECT 260.920 14.080 275.520 14.400 ; 
                RECT 680.480 14.080 689.960 14.400 ; 
                RECT 0.160 15.440 275.520 15.760 ; 
                RECT 680.480 15.440 689.960 15.760 ; 
                RECT 0.160 16.800 275.520 17.120 ; 
                RECT 680.480 16.800 689.960 17.120 ; 
                RECT 0.160 18.160 198.000 18.480 ; 
                RECT 260.240 18.160 275.520 18.480 ; 
                RECT 680.480 18.160 689.960 18.480 ; 
                RECT 0.160 19.520 275.520 19.840 ; 
                RECT 680.480 19.520 689.960 19.840 ; 
                RECT 0.160 20.880 275.520 21.200 ; 
                RECT 680.480 20.880 689.960 21.200 ; 
                RECT 0.160 22.240 275.520 22.560 ; 
                RECT 680.480 22.240 689.960 22.560 ; 
                RECT 0.160 23.600 275.520 23.920 ; 
                RECT 680.480 23.600 689.960 23.920 ; 
                RECT 0.160 24.960 275.520 25.280 ; 
                RECT 680.480 24.960 689.960 25.280 ; 
                RECT 0.160 26.320 275.520 26.640 ; 
                RECT 680.480 26.320 689.960 26.640 ; 
                RECT 0.160 27.680 274.840 28.000 ; 
                RECT 680.480 27.680 689.960 28.000 ; 
                RECT 0.160 29.040 275.520 29.360 ; 
                RECT 680.480 29.040 689.960 29.360 ; 
                RECT 0.160 30.400 275.520 30.720 ; 
                RECT 680.480 30.400 689.960 30.720 ; 
                RECT 0.160 31.760 275.520 32.080 ; 
                RECT 680.480 31.760 689.960 32.080 ; 
                RECT 0.160 33.120 275.520 33.440 ; 
                RECT 680.480 33.120 689.960 33.440 ; 
                RECT 0.160 34.480 168.080 34.800 ; 
                RECT 237.800 34.480 275.520 34.800 ; 
                RECT 680.480 34.480 689.960 34.800 ; 
                RECT 0.160 35.840 166.720 36.160 ; 
                RECT 243.920 35.840 275.520 36.160 ; 
                RECT 680.480 35.840 689.960 36.160 ; 
                RECT 0.160 37.200 147.000 37.520 ; 
                RECT 260.920 37.200 275.520 37.520 ; 
                RECT 680.480 37.200 689.960 37.520 ; 
                RECT 0.160 38.560 146.320 38.880 ; 
                RECT 256.840 38.560 275.520 38.880 ; 
                RECT 680.480 38.560 689.960 38.880 ; 
                RECT 0.160 39.920 275.520 40.240 ; 
                RECT 680.480 39.920 689.960 40.240 ; 
                RECT 0.160 41.280 275.520 41.600 ; 
                RECT 680.480 41.280 689.960 41.600 ; 
                RECT 0.160 42.640 275.520 42.960 ; 
                RECT 680.480 42.640 689.960 42.960 ; 
                RECT 0.160 44.000 275.520 44.320 ; 
                RECT 680.480 44.000 689.960 44.320 ; 
                RECT 0.160 45.360 142.240 45.680 ; 
                RECT 153.480 45.360 275.520 45.680 ; 
                RECT 680.480 45.360 689.960 45.680 ; 
                RECT 0.160 46.720 143.600 47.040 ; 
                RECT 149.400 46.720 157.200 47.040 ; 
                RECT 159.600 46.720 275.520 47.040 ; 
                RECT 680.480 46.720 689.960 47.040 ; 
                RECT 0.160 48.080 144.960 48.400 ; 
                RECT 148.720 48.080 275.520 48.400 ; 
                RECT 680.480 48.080 689.960 48.400 ; 
                RECT 0.160 49.440 151.760 49.760 ; 
                RECT 158.920 49.440 275.520 49.760 ; 
                RECT 680.480 49.440 689.960 49.760 ; 
                RECT 0.160 50.800 154.480 51.120 ; 
                RECT 160.280 50.800 275.520 51.120 ; 
                RECT 680.480 50.800 689.960 51.120 ; 
                RECT 0.160 52.160 144.280 52.480 ; 
                RECT 153.480 52.160 275.520 52.480 ; 
                RECT 680.480 52.160 689.960 52.480 ; 
                RECT 0.160 53.520 147.680 53.840 ; 
                RECT 152.800 53.520 253.080 53.840 ; 
                RECT 258.880 53.520 275.520 53.840 ; 
                RECT 680.480 53.520 689.960 53.840 ; 
                RECT 0.160 54.880 253.080 55.200 ; 
                RECT 680.480 54.880 689.960 55.200 ; 
                RECT 0.160 56.240 143.600 56.560 ; 
                RECT 153.480 56.240 253.080 56.560 ; 
                RECT 680.480 56.240 689.960 56.560 ; 
                RECT 0.160 57.600 150.400 57.920 ; 
                RECT 158.920 57.600 253.080 57.920 ; 
                RECT 258.880 57.600 275.520 57.920 ; 
                RECT 680.480 57.600 689.960 57.920 ; 
                RECT 0.160 58.960 253.080 59.280 ; 
                RECT 258.880 58.960 275.520 59.280 ; 
                RECT 680.480 58.960 689.960 59.280 ; 
                RECT 0.160 60.320 151.760 60.640 ; 
                RECT 157.560 60.320 275.520 60.640 ; 
                RECT 680.480 60.320 689.960 60.640 ; 
                RECT 0.160 61.680 154.480 62.000 ; 
                RECT 159.600 61.680 275.520 62.000 ; 
                RECT 680.480 61.680 689.960 62.000 ; 
                RECT 0.160 63.040 148.360 63.360 ; 
                RECT 153.480 63.040 275.520 63.360 ; 
                RECT 680.480 63.040 689.960 63.360 ; 
                RECT 0.160 64.400 177.600 64.720 ; 
                RECT 258.200 64.400 275.520 64.720 ; 
                RECT 680.480 64.400 689.960 64.720 ; 
                RECT 0.160 65.760 141.560 66.080 ; 
                RECT 165.040 65.760 167.400 66.080 ; 
                RECT 171.840 65.760 177.600 66.080 ; 
                RECT 258.200 65.760 275.520 66.080 ; 
                RECT 680.480 65.760 689.960 66.080 ; 
                RECT 0.160 67.120 151.760 67.440 ; 
                RECT 159.600 67.120 168.760 67.440 ; 
                RECT 171.160 67.120 177.600 67.440 ; 
                RECT 267.720 67.120 275.520 67.440 ; 
                RECT 680.480 67.120 689.960 67.440 ; 
                RECT 0.160 68.480 150.400 68.800 ; 
                RECT 153.480 68.480 159.920 68.800 ; 
                RECT 167.080 68.480 177.600 68.800 ; 
                RECT 267.720 68.480 275.520 68.800 ; 
                RECT 680.480 68.480 689.960 68.800 ; 
                RECT 0.160 69.840 142.240 70.160 ; 
                RECT 156.200 69.840 177.600 70.160 ; 
                RECT 267.720 69.840 275.520 70.160 ; 
                RECT 680.480 69.840 689.960 70.160 ; 
                RECT 0.160 71.200 151.080 71.520 ; 
                RECT 159.600 71.200 177.600 71.520 ; 
                RECT 266.360 71.200 275.520 71.520 ; 
                RECT 680.480 71.200 689.960 71.520 ; 
                RECT 0.160 72.560 149.040 72.880 ; 
                RECT 152.800 72.560 177.600 72.880 ; 
                RECT 267.720 72.560 275.520 72.880 ; 
                RECT 680.480 72.560 689.960 72.880 ; 
                RECT 0.160 73.920 144.280 74.240 ; 
                RECT 148.720 73.920 151.760 74.240 ; 
                RECT 160.280 73.920 177.600 74.240 ; 
                RECT 258.200 73.920 275.520 74.240 ; 
                RECT 680.480 73.920 689.960 74.240 ; 
                RECT 0.160 75.280 147.000 75.600 ; 
                RECT 150.760 75.280 177.600 75.600 ; 
                RECT 270.440 75.280 275.520 75.600 ; 
                RECT 680.480 75.280 689.960 75.600 ; 
                RECT 0.160 76.640 143.600 76.960 ; 
                RECT 147.360 76.640 177.600 76.960 ; 
                RECT 270.440 76.640 275.520 76.960 ; 
                RECT 680.480 76.640 689.960 76.960 ; 
                RECT 0.160 78.000 147.680 78.320 ; 
                RECT 153.480 78.000 177.600 78.320 ; 
                RECT 269.080 78.000 275.520 78.320 ; 
                RECT 680.480 78.000 689.960 78.320 ; 
                RECT 0.160 79.360 143.600 79.680 ; 
                RECT 158.920 79.360 177.600 79.680 ; 
                RECT 270.440 79.360 275.520 79.680 ; 
                RECT 680.480 79.360 689.960 79.680 ; 
                RECT 0.160 80.720 150.400 81.040 ; 
                RECT 152.800 80.720 177.600 81.040 ; 
                RECT 270.440 80.720 275.520 81.040 ; 
                RECT 680.480 80.720 689.960 81.040 ; 
                RECT 0.160 82.080 177.600 82.400 ; 
                RECT 258.200 82.080 275.520 82.400 ; 
                RECT 680.480 82.080 689.960 82.400 ; 
                RECT 0.160 83.440 151.760 83.760 ; 
                RECT 153.480 83.440 177.600 83.760 ; 
                RECT 273.160 83.440 275.520 83.760 ; 
                RECT 680.480 83.440 689.960 83.760 ; 
                RECT 0.160 84.800 142.240 85.120 ; 
                RECT 152.800 84.800 177.600 85.120 ; 
                RECT 271.800 84.800 275.520 85.120 ; 
                RECT 680.480 84.800 689.960 85.120 ; 
                RECT 0.160 86.160 147.680 86.480 ; 
                RECT 159.600 86.160 177.600 86.480 ; 
                RECT 273.160 86.160 275.520 86.480 ; 
                RECT 680.480 86.160 689.960 86.480 ; 
                RECT 0.160 87.520 145.640 87.840 ; 
                RECT 153.480 87.520 177.600 87.840 ; 
                RECT 273.160 87.520 275.520 87.840 ; 
                RECT 680.480 87.520 689.960 87.840 ; 
                RECT 0.160 88.880 151.080 89.200 ; 
                RECT 153.480 88.880 177.600 89.200 ; 
                RECT 273.160 88.880 275.520 89.200 ; 
                RECT 680.480 88.880 689.960 89.200 ; 
                RECT 0.160 90.240 177.600 90.560 ; 
                RECT 271.800 90.240 275.520 90.560 ; 
                RECT 680.480 90.240 689.960 90.560 ; 
                RECT 0.160 91.600 177.600 91.920 ; 
                RECT 258.200 91.600 275.520 91.920 ; 
                RECT 680.480 91.600 689.960 91.920 ; 
                RECT 0.160 92.960 138.840 93.280 ; 
                RECT 156.200 92.960 177.600 93.280 ; 
                RECT 680.480 92.960 689.960 93.280 ; 
                RECT 0.160 94.320 177.600 94.640 ; 
                RECT 680.480 94.320 689.960 94.640 ; 
                RECT 0.160 95.680 177.600 96.000 ; 
                RECT 680.480 95.680 689.960 96.000 ; 
                RECT 0.160 97.040 147.680 97.360 ; 
                RECT 159.600 97.040 177.600 97.360 ; 
                RECT 680.480 97.040 689.960 97.360 ; 
                RECT 0.160 98.400 154.480 98.720 ; 
                RECT 161.640 98.400 177.600 98.720 ; 
                RECT 680.480 98.400 689.960 98.720 ; 
                RECT 0.160 99.760 177.600 100.080 ; 
                RECT 258.200 99.760 275.520 100.080 ; 
                RECT 680.480 99.760 689.960 100.080 ; 
                RECT 0.160 101.120 275.520 101.440 ; 
                RECT 680.480 101.120 689.960 101.440 ; 
                RECT 0.160 102.480 141.560 102.800 ; 
                RECT 147.360 102.480 275.520 102.800 ; 
                RECT 680.480 102.480 689.960 102.800 ; 
                RECT 0.160 103.840 261.920 104.160 ; 
                RECT 680.480 103.840 689.960 104.160 ; 
                RECT 0.160 105.200 272.800 105.520 ; 
                RECT 680.480 105.200 689.960 105.520 ; 
                RECT 0.160 106.560 157.200 106.880 ; 
                RECT 160.280 106.560 166.040 106.880 ; 
                RECT 202.440 106.560 205.480 106.880 ; 
                RECT 258.200 106.560 270.080 106.880 ; 
                RECT 680.480 106.560 689.960 106.880 ; 
                RECT 0.160 107.920 120.480 108.240 ; 
                RECT 139.200 107.920 205.480 108.240 ; 
                RECT 258.200 107.920 267.360 108.240 ; 
                RECT 680.480 107.920 689.960 108.240 ; 
                RECT 0.160 109.280 120.480 109.600 ; 
                RECT 139.200 109.280 205.480 109.600 ; 
                RECT 258.200 109.280 264.640 109.600 ; 
                RECT 680.480 109.280 689.960 109.600 ; 
                RECT 0.160 110.640 120.480 110.960 ; 
                RECT 139.200 110.640 205.480 110.960 ; 
                RECT 258.200 110.640 264.640 110.960 ; 
                RECT 680.480 110.640 689.960 110.960 ; 
                RECT 0.160 112.000 120.480 112.320 ; 
                RECT 139.200 112.000 144.280 112.320 ; 
                RECT 149.400 112.000 205.480 112.320 ; 
                RECT 258.200 112.000 275.520 112.320 ; 
                RECT 680.480 112.000 689.960 112.320 ; 
                RECT 0.160 113.360 120.480 113.680 ; 
                RECT 139.200 113.360 275.520 113.680 ; 
                RECT 680.480 113.360 689.960 113.680 ; 
                RECT 0.160 114.720 120.480 115.040 ; 
                RECT 139.200 114.720 147.680 115.040 ; 
                RECT 158.920 114.720 275.520 115.040 ; 
                RECT 680.480 114.720 689.960 115.040 ; 
                RECT 0.160 116.080 120.480 116.400 ; 
                RECT 139.200 116.080 275.520 116.400 ; 
                RECT 680.480 116.080 689.960 116.400 ; 
                RECT 0.160 117.440 120.480 117.760 ; 
                RECT 139.200 117.440 275.520 117.760 ; 
                RECT 680.480 117.440 689.960 117.760 ; 
                RECT 0.160 118.800 120.480 119.120 ; 
                RECT 139.880 118.800 143.600 119.120 ; 
                RECT 146.680 118.800 202.760 119.120 ; 
                RECT 258.200 118.800 275.520 119.120 ; 
                RECT 680.480 118.800 689.960 119.120 ; 
                RECT 0.160 120.160 120.480 120.480 ; 
                RECT 139.200 120.160 144.280 120.480 ; 
                RECT 149.400 120.160 202.760 120.480 ; 
                RECT 258.200 120.160 275.520 120.480 ; 
                RECT 680.480 120.160 689.960 120.480 ; 
                RECT 0.160 121.520 120.480 121.840 ; 
                RECT 139.200 121.520 202.760 121.840 ; 
                RECT 258.200 121.520 275.520 121.840 ; 
                RECT 680.480 121.520 689.960 121.840 ; 
                RECT 0.160 122.880 120.480 123.200 ; 
                RECT 139.200 122.880 202.760 123.200 ; 
                RECT 258.200 122.880 275.520 123.200 ; 
                RECT 680.480 122.880 689.960 123.200 ; 
                RECT 0.160 124.240 120.480 124.560 ; 
                RECT 139.200 124.240 202.760 124.560 ; 
                RECT 258.200 124.240 266.000 124.560 ; 
                RECT 680.480 124.240 689.960 124.560 ; 
                RECT 0.160 125.600 120.480 125.920 ; 
                RECT 139.200 125.600 202.760 125.920 ; 
                RECT 258.200 125.600 266.000 125.920 ; 
                RECT 680.480 125.600 689.960 125.920 ; 
                RECT 0.160 126.960 120.480 127.280 ; 
                RECT 139.200 126.960 202.760 127.280 ; 
                RECT 258.200 126.960 268.720 127.280 ; 
                RECT 680.480 126.960 689.960 127.280 ; 
                RECT 0.160 128.320 120.480 128.640 ; 
                RECT 139.200 128.320 202.760 128.640 ; 
                RECT 258.200 128.320 271.440 128.640 ; 
                RECT 680.480 128.320 689.960 128.640 ; 
                RECT 0.160 129.680 120.480 130.000 ; 
                RECT 139.200 129.680 202.760 130.000 ; 
                RECT 680.480 129.680 689.960 130.000 ; 
                RECT 0.160 131.040 120.480 131.360 ; 
                RECT 139.200 131.040 145.640 131.360 ; 
                RECT 149.400 131.040 202.760 131.360 ; 
                RECT 680.480 131.040 689.960 131.360 ; 
                RECT 0.160 132.400 202.760 132.720 ; 
                RECT 258.200 132.400 275.520 132.720 ; 
                RECT 680.480 132.400 689.960 132.720 ; 
                RECT 0.160 133.760 202.760 134.080 ; 
                RECT 258.200 133.760 275.520 134.080 ; 
                RECT 680.480 133.760 689.960 134.080 ; 
                RECT 0.160 135.120 147.680 135.440 ; 
                RECT 153.480 135.120 202.760 135.440 ; 
                RECT 258.200 135.120 275.520 135.440 ; 
                RECT 680.480 135.120 689.960 135.440 ; 
                RECT 0.160 136.480 102.120 136.800 ; 
                RECT 120.840 136.480 126.600 136.800 ; 
                RECT 133.760 136.480 202.760 136.800 ; 
                RECT 258.200 136.480 275.520 136.800 ; 
                RECT 680.480 136.480 689.960 136.800 ; 
                RECT 0.160 137.840 102.120 138.160 ; 
                RECT 138.520 137.840 202.760 138.160 ; 
                RECT 258.200 137.840 275.520 138.160 ; 
                RECT 680.480 137.840 689.960 138.160 ; 
                RECT 0.160 139.200 102.120 139.520 ; 
                RECT 138.520 139.200 202.760 139.520 ; 
                RECT 680.480 139.200 689.960 139.520 ; 
                RECT 0.160 140.560 102.120 140.880 ; 
                RECT 120.840 140.560 126.600 140.880 ; 
                RECT 133.760 140.560 146.320 140.880 ; 
                RECT 152.120 140.560 202.760 140.880 ; 
                RECT 680.480 140.560 689.960 140.880 ; 
                RECT 0.160 141.920 100.760 142.240 ; 
                RECT 133.080 141.920 202.760 142.240 ; 
                RECT 258.200 141.920 689.960 142.240 ; 
                RECT 0.160 143.280 132.720 143.600 ; 
                RECT 199.720 143.280 689.960 143.600 ; 
                RECT 0.160 144.640 272.800 144.960 ; 
                RECT 682.520 144.640 689.960 144.960 ; 
                RECT 0.160 146.000 272.800 146.320 ; 
                RECT 682.520 146.000 689.960 146.320 ; 
                RECT 0.160 147.360 272.800 147.680 ; 
                RECT 682.520 147.360 689.960 147.680 ; 
                RECT 0.160 148.720 26.640 149.040 ; 
                RECT 33.120 148.720 34.800 149.040 ; 
                RECT 47.400 148.720 80.360 149.040 ; 
                RECT 682.520 148.720 689.960 149.040 ; 
                RECT 0.160 150.080 24.600 150.400 ; 
                RECT 46.720 150.080 64.040 150.400 ; 
                RECT 69.840 150.080 80.360 150.400 ; 
                RECT 682.520 150.080 689.960 150.400 ; 
                RECT 0.160 151.440 24.600 151.760 ; 
                RECT 45.360 151.440 59.960 151.760 ; 
                RECT 69.840 151.440 80.360 151.760 ; 
                RECT 682.520 151.440 689.960 151.760 ; 
                RECT 0.160 152.800 24.600 153.120 ; 
                RECT 35.160 152.800 59.960 153.120 ; 
                RECT 69.840 152.800 80.360 153.120 ; 
                RECT 682.520 152.800 689.960 153.120 ; 
                RECT 0.160 154.160 59.960 154.480 ; 
                RECT 69.840 154.160 80.360 154.480 ; 
                RECT 682.520 154.160 689.960 154.480 ; 
                RECT 0.160 155.520 24.600 155.840 ; 
                RECT 35.160 155.520 59.960 155.840 ; 
                RECT 69.840 155.520 80.360 155.840 ; 
                RECT 682.520 155.520 689.960 155.840 ; 
                RECT 0.160 156.880 24.600 157.200 ; 
                RECT 35.160 156.880 80.360 157.200 ; 
                RECT 682.520 156.880 689.960 157.200 ; 
                RECT 0.160 158.240 59.960 158.560 ; 
                RECT 69.840 158.240 80.360 158.560 ; 
                RECT 682.520 158.240 689.960 158.560 ; 
                RECT 0.160 159.600 59.960 159.920 ; 
                RECT 69.840 159.600 80.360 159.920 ; 
                RECT 682.520 159.600 689.960 159.920 ; 
                RECT 0.160 160.960 59.960 161.280 ; 
                RECT 69.840 160.960 80.360 161.280 ; 
                RECT 682.520 160.960 689.960 161.280 ; 
                RECT 0.160 162.320 17.800 162.640 ; 
                RECT 20.200 162.320 33.440 162.640 ; 
                RECT 35.840 162.320 59.960 162.640 ; 
                RECT 69.840 162.320 80.360 162.640 ; 
                RECT 682.520 162.320 689.960 162.640 ; 
                RECT 0.160 163.680 17.120 164.000 ; 
                RECT 20.200 163.680 33.440 164.000 ; 
                RECT 36.520 163.680 59.960 164.000 ; 
                RECT 69.840 163.680 80.360 164.000 ; 
                RECT 682.520 163.680 689.960 164.000 ; 
                RECT 0.160 165.040 16.440 165.360 ; 
                RECT 20.200 165.040 80.360 165.360 ; 
                RECT 682.520 165.040 689.960 165.360 ; 
                RECT 0.160 166.400 15.760 166.720 ; 
                RECT 20.200 166.400 60.640 166.720 ; 
                RECT 69.840 166.400 80.360 166.720 ; 
                RECT 682.520 166.400 689.960 166.720 ; 
                RECT 0.160 167.760 59.960 168.080 ; 
                RECT 69.840 167.760 80.360 168.080 ; 
                RECT 682.520 167.760 689.960 168.080 ; 
                RECT 0.160 169.120 15.080 169.440 ; 
                RECT 20.200 169.120 59.960 169.440 ; 
                RECT 69.840 169.120 80.360 169.440 ; 
                RECT 682.520 169.120 689.960 169.440 ; 
                RECT 0.160 170.480 14.400 170.800 ; 
                RECT 20.200 170.480 59.960 170.800 ; 
                RECT 69.840 170.480 80.360 170.800 ; 
                RECT 682.520 170.480 689.960 170.800 ; 
                RECT 0.160 171.840 59.960 172.160 ; 
                RECT 69.840 171.840 80.360 172.160 ; 
                RECT 682.520 171.840 689.960 172.160 ; 
                RECT 0.160 173.200 13.720 173.520 ; 
                RECT 20.200 173.200 80.360 173.520 ; 
                RECT 682.520 173.200 689.960 173.520 ; 
                RECT 0.160 174.560 13.040 174.880 ; 
                RECT 20.200 174.560 33.440 174.880 ; 
                RECT 38.560 174.560 59.960 174.880 ; 
                RECT 69.840 174.560 80.360 174.880 ; 
                RECT 682.520 174.560 689.960 174.880 ; 
                RECT 0.160 175.920 59.960 176.240 ; 
                RECT 69.840 175.920 80.360 176.240 ; 
                RECT 682.520 175.920 689.960 176.240 ; 
                RECT 0.160 177.280 12.360 177.600 ; 
                RECT 20.200 177.280 33.440 177.600 ; 
                RECT 37.880 177.280 59.960 177.600 ; 
                RECT 69.840 177.280 80.360 177.600 ; 
                RECT 682.520 177.280 689.960 177.600 ; 
                RECT 0.160 178.640 11.680 178.960 ; 
                RECT 20.200 178.640 33.440 178.960 ; 
                RECT 37.200 178.640 59.960 178.960 ; 
                RECT 69.840 178.640 80.360 178.960 ; 
                RECT 682.520 178.640 689.960 178.960 ; 
                RECT 0.160 180.000 11.000 180.320 ; 
                RECT 20.200 180.000 33.440 180.320 ; 
                RECT 36.520 180.000 59.960 180.320 ; 
                RECT 69.160 180.000 80.360 180.320 ; 
                RECT 682.520 180.000 689.960 180.320 ; 
                RECT 0.160 181.360 10.320 181.680 ; 
                RECT 20.200 181.360 64.040 181.680 ; 
                RECT 69.840 181.360 80.360 181.680 ; 
                RECT 682.520 181.360 689.960 181.680 ; 
                RECT 0.160 182.720 61.320 183.040 ; 
                RECT 69.840 182.720 80.360 183.040 ; 
                RECT 682.520 182.720 689.960 183.040 ; 
                RECT 0.160 184.080 61.320 184.400 ; 
                RECT 69.840 184.080 80.360 184.400 ; 
                RECT 682.520 184.080 689.960 184.400 ; 
                RECT 0.160 185.440 61.320 185.760 ; 
                RECT 69.840 185.440 80.360 185.760 ; 
                RECT 682.520 185.440 689.960 185.760 ; 
                RECT 0.160 186.800 61.320 187.120 ; 
                RECT 69.840 186.800 80.360 187.120 ; 
                RECT 682.520 186.800 689.960 187.120 ; 
                RECT 0.160 188.160 38.200 188.480 ; 
                RECT 47.400 188.160 80.360 188.480 ; 
                RECT 682.520 188.160 689.960 188.480 ; 
                RECT 0.160 189.520 36.840 189.840 ; 
                RECT 46.720 189.520 66.080 189.840 ; 
                RECT 69.840 189.520 80.360 189.840 ; 
                RECT 682.520 189.520 689.960 189.840 ; 
                RECT 0.160 190.880 35.480 191.200 ; 
                RECT 45.360 190.880 59.960 191.200 ; 
                RECT 69.840 190.880 80.360 191.200 ; 
                RECT 682.520 190.880 689.960 191.200 ; 
                RECT 0.160 192.240 59.960 192.560 ; 
                RECT 69.840 192.240 80.360 192.560 ; 
                RECT 682.520 192.240 689.960 192.560 ; 
                RECT 0.160 193.600 59.960 193.920 ; 
                RECT 69.840 193.600 80.360 193.920 ; 
                RECT 682.520 193.600 689.960 193.920 ; 
                RECT 0.160 194.960 59.960 195.280 ; 
                RECT 69.840 194.960 80.360 195.280 ; 
                RECT 682.520 194.960 689.960 195.280 ; 
                RECT 0.160 196.320 59.960 196.640 ; 
                RECT 62.360 196.320 80.360 196.640 ; 
                RECT 682.520 196.320 689.960 196.640 ; 
                RECT 0.160 197.680 61.320 198.000 ; 
                RECT 69.840 197.680 80.360 198.000 ; 
                RECT 682.520 197.680 689.960 198.000 ; 
                RECT 0.160 199.040 59.960 199.360 ; 
                RECT 69.840 199.040 80.360 199.360 ; 
                RECT 682.520 199.040 689.960 199.360 ; 
                RECT 0.160 200.400 59.960 200.720 ; 
                RECT 69.840 200.400 80.360 200.720 ; 
                RECT 682.520 200.400 689.960 200.720 ; 
                RECT 0.160 201.760 59.960 202.080 ; 
                RECT 69.840 201.760 80.360 202.080 ; 
                RECT 682.520 201.760 689.960 202.080 ; 
                RECT 0.160 203.120 59.960 203.440 ; 
                RECT 69.840 203.120 80.360 203.440 ; 
                RECT 682.520 203.120 689.960 203.440 ; 
                RECT 0.160 204.480 80.360 204.800 ; 
                RECT 682.520 204.480 689.960 204.800 ; 
                RECT 0.160 205.840 61.320 206.160 ; 
                RECT 69.840 205.840 80.360 206.160 ; 
                RECT 682.520 205.840 689.960 206.160 ; 
                RECT 0.160 207.200 59.960 207.520 ; 
                RECT 69.840 207.200 80.360 207.520 ; 
                RECT 682.520 207.200 689.960 207.520 ; 
                RECT 0.160 208.560 59.960 208.880 ; 
                RECT 69.840 208.560 80.360 208.880 ; 
                RECT 682.520 208.560 689.960 208.880 ; 
                RECT 0.160 209.920 59.960 210.240 ; 
                RECT 69.840 209.920 80.360 210.240 ; 
                RECT 682.520 209.920 689.960 210.240 ; 
                RECT 0.160 211.280 59.960 211.600 ; 
                RECT 69.840 211.280 80.360 211.600 ; 
                RECT 682.520 211.280 689.960 211.600 ; 
                RECT 0.160 212.640 80.360 212.960 ; 
                RECT 682.520 212.640 689.960 212.960 ; 
                RECT 0.160 214.000 59.960 214.320 ; 
                RECT 69.840 214.000 80.360 214.320 ; 
                RECT 682.520 214.000 689.960 214.320 ; 
                RECT 0.160 215.360 59.960 215.680 ; 
                RECT 69.840 215.360 80.360 215.680 ; 
                RECT 682.520 215.360 689.960 215.680 ; 
                RECT 0.160 216.720 59.960 217.040 ; 
                RECT 69.840 216.720 80.360 217.040 ; 
                RECT 682.520 216.720 689.960 217.040 ; 
                RECT 0.160 218.080 59.960 218.400 ; 
                RECT 69.840 218.080 80.360 218.400 ; 
                RECT 682.520 218.080 689.960 218.400 ; 
                RECT 0.160 219.440 59.960 219.760 ; 
                RECT 69.840 219.440 80.360 219.760 ; 
                RECT 682.520 219.440 689.960 219.760 ; 
                RECT 0.160 220.800 80.360 221.120 ; 
                RECT 682.520 220.800 689.960 221.120 ; 
                RECT 0.160 222.160 62.000 222.480 ; 
                RECT 69.840 222.160 80.360 222.480 ; 
                RECT 682.520 222.160 689.960 222.480 ; 
                RECT 0.160 223.520 62.000 223.840 ; 
                RECT 69.840 223.520 80.360 223.840 ; 
                RECT 682.520 223.520 689.960 223.840 ; 
                RECT 0.160 224.880 62.000 225.200 ; 
                RECT 69.840 224.880 80.360 225.200 ; 
                RECT 682.520 224.880 689.960 225.200 ; 
                RECT 0.160 226.240 62.000 226.560 ; 
                RECT 69.840 226.240 80.360 226.560 ; 
                RECT 682.520 226.240 689.960 226.560 ; 
                RECT 0.160 227.600 80.360 227.920 ; 
                RECT 682.520 227.600 689.960 227.920 ; 
                RECT 0.160 228.960 64.040 229.280 ; 
                RECT 69.840 228.960 80.360 229.280 ; 
                RECT 682.520 228.960 689.960 229.280 ; 
                RECT 0.160 230.320 62.680 230.640 ; 
                RECT 69.840 230.320 80.360 230.640 ; 
                RECT 682.520 230.320 689.960 230.640 ; 
                RECT 0.160 231.680 62.680 232.000 ; 
                RECT 69.840 231.680 80.360 232.000 ; 
                RECT 682.520 231.680 689.960 232.000 ; 
                RECT 0.160 233.040 62.680 233.360 ; 
                RECT 69.840 233.040 80.360 233.360 ; 
                RECT 682.520 233.040 689.960 233.360 ; 
                RECT 0.160 234.400 62.680 234.720 ; 
                RECT 69.840 234.400 80.360 234.720 ; 
                RECT 682.520 234.400 689.960 234.720 ; 
                RECT 0.160 235.760 80.360 236.080 ; 
                RECT 682.520 235.760 689.960 236.080 ; 
                RECT 0.160 237.120 66.080 237.440 ; 
                RECT 69.840 237.120 80.360 237.440 ; 
                RECT 682.520 237.120 689.960 237.440 ; 
                RECT 0.160 238.480 66.080 238.800 ; 
                RECT 69.840 238.480 80.360 238.800 ; 
                RECT 682.520 238.480 689.960 238.800 ; 
                RECT 0.160 239.840 62.680 240.160 ; 
                RECT 69.840 239.840 80.360 240.160 ; 
                RECT 682.520 239.840 689.960 240.160 ; 
                RECT 0.160 241.200 62.680 241.520 ; 
                RECT 69.840 241.200 80.360 241.520 ; 
                RECT 682.520 241.200 689.960 241.520 ; 
                RECT 0.160 242.560 62.680 242.880 ; 
                RECT 69.840 242.560 80.360 242.880 ; 
                RECT 682.520 242.560 689.960 242.880 ; 
                RECT 0.160 243.920 80.360 244.240 ; 
                RECT 682.520 243.920 689.960 244.240 ; 
                RECT 0.160 245.280 62.680 245.600 ; 
                RECT 69.840 245.280 80.360 245.600 ; 
                RECT 682.520 245.280 689.960 245.600 ; 
                RECT 0.160 246.640 62.680 246.960 ; 
                RECT 69.840 246.640 80.360 246.960 ; 
                RECT 682.520 246.640 689.960 246.960 ; 
                RECT 0.160 248.000 64.720 248.320 ; 
                RECT 69.840 248.000 80.360 248.320 ; 
                RECT 682.520 248.000 689.960 248.320 ; 
                RECT 0.160 249.360 62.680 249.680 ; 
                RECT 69.840 249.360 80.360 249.680 ; 
                RECT 682.520 249.360 689.960 249.680 ; 
                RECT 0.160 250.720 62.680 251.040 ; 
                RECT 69.840 250.720 80.360 251.040 ; 
                RECT 682.520 250.720 689.960 251.040 ; 
                RECT 0.160 252.080 80.360 252.400 ; 
                RECT 682.520 252.080 689.960 252.400 ; 
                RECT 0.160 253.440 62.680 253.760 ; 
                RECT 69.840 253.440 80.360 253.760 ; 
                RECT 682.520 253.440 689.960 253.760 ; 
                RECT 0.160 254.800 62.680 255.120 ; 
                RECT 69.840 254.800 80.360 255.120 ; 
                RECT 682.520 254.800 689.960 255.120 ; 
                RECT 0.160 256.160 62.680 256.480 ; 
                RECT 69.840 256.160 80.360 256.480 ; 
                RECT 682.520 256.160 689.960 256.480 ; 
                RECT 0.160 257.520 67.440 257.840 ; 
                RECT 69.840 257.520 80.360 257.840 ; 
                RECT 682.520 257.520 689.960 257.840 ; 
                RECT 0.160 258.880 62.680 259.200 ; 
                RECT 69.840 258.880 80.360 259.200 ; 
                RECT 682.520 258.880 689.960 259.200 ; 
                RECT 0.160 260.240 80.360 260.560 ; 
                RECT 682.520 260.240 689.960 260.560 ; 
                RECT 0.160 261.600 63.360 261.920 ; 
                RECT 69.840 261.600 80.360 261.920 ; 
                RECT 682.520 261.600 689.960 261.920 ; 
                RECT 0.160 262.960 63.360 263.280 ; 
                RECT 69.840 262.960 80.360 263.280 ; 
                RECT 682.520 262.960 689.960 263.280 ; 
                RECT 0.160 264.320 63.360 264.640 ; 
                RECT 69.840 264.320 80.360 264.640 ; 
                RECT 682.520 264.320 689.960 264.640 ; 
                RECT 0.160 265.680 63.360 266.000 ; 
                RECT 69.840 265.680 80.360 266.000 ; 
                RECT 682.520 265.680 689.960 266.000 ; 
                RECT 0.160 267.040 80.360 267.360 ; 
                RECT 682.520 267.040 689.960 267.360 ; 
                RECT 0.160 268.400 66.080 268.720 ; 
                RECT 69.840 268.400 80.360 268.720 ; 
                RECT 682.520 268.400 689.960 268.720 ; 
                RECT 0.160 269.760 63.360 270.080 ; 
                RECT 69.840 269.760 80.360 270.080 ; 
                RECT 682.520 269.760 689.960 270.080 ; 
                RECT 0.160 271.120 63.360 271.440 ; 
                RECT 69.840 271.120 80.360 271.440 ; 
                RECT 682.520 271.120 689.960 271.440 ; 
                RECT 0.160 272.480 63.360 272.800 ; 
                RECT 69.840 272.480 80.360 272.800 ; 
                RECT 682.520 272.480 689.960 272.800 ; 
                RECT 0.160 273.840 63.360 274.160 ; 
                RECT 69.840 273.840 80.360 274.160 ; 
                RECT 682.520 273.840 689.960 274.160 ; 
                RECT 0.160 275.200 80.360 275.520 ; 
                RECT 682.520 275.200 689.960 275.520 ; 
                RECT 0.160 276.560 80.360 276.880 ; 
                RECT 682.520 276.560 689.960 276.880 ; 
                RECT 0.160 277.920 272.800 278.240 ; 
                RECT 682.520 277.920 689.960 278.240 ; 
                RECT 0.160 279.280 272.800 279.600 ; 
                RECT 682.520 279.280 689.960 279.600 ; 
                RECT 0.160 280.640 689.960 280.960 ; 
                RECT 0.160 282.000 689.960 282.320 ; 
                RECT 0.160 283.360 689.960 283.680 ; 
                RECT 0.160 284.720 689.960 285.040 ; 
                RECT 0.160 286.080 689.960 286.400 ; 
                RECT 0.160 0.160 689.960 1.520 ; 
                RECT 0.160 290.120 689.960 291.480 ; 
                RECT 276.940 32.275 282.740 33.645 ; 
                RECT 672.840 32.275 678.640 33.645 ; 
                RECT 276.940 37.795 282.740 39.535 ; 
                RECT 672.840 37.795 678.640 39.535 ; 
                RECT 276.940 43.640 282.740 45.210 ; 
                RECT 672.840 43.640 678.640 45.210 ; 
                RECT 276.940 49.230 282.740 50.800 ; 
                RECT 672.840 49.230 678.640 50.800 ; 
                RECT 276.940 84.710 678.640 86.800 ; 
                RECT 276.940 69.130 678.640 69.930 ; 
                RECT 276.940 90.135 678.640 90.425 ; 
                RECT 276.940 113.775 678.640 115.575 ; 
                RECT 276.940 57.660 678.640 59.460 ; 
                RECT 276.940 134.765 678.640 137.365 ; 
                RECT 276.940 72.140 678.640 72.940 ; 
                RECT 276.940 77.030 678.640 77.830 ; 
                RECT 276.940 16.520 678.640 18.320 ; 
                RECT 84.730 148.435 86.650 276.415 ; 
                RECT 88.570 148.435 90.490 276.415 ; 
                RECT 100.765 148.435 102.685 276.415 ; 
                RECT 104.605 148.435 106.525 276.415 ; 
                RECT 108.445 148.435 110.365 276.415 ; 
                RECT 112.285 148.435 114.205 276.415 ; 
                RECT 133.600 148.435 135.520 276.415 ; 
                RECT 137.440 148.435 139.360 276.415 ; 
                RECT 141.280 148.435 143.200 276.415 ; 
                RECT 145.120 148.435 147.040 276.415 ; 
                RECT 148.960 148.435 150.880 276.415 ; 
                RECT 152.800 148.435 154.720 276.415 ; 
                RECT 156.640 148.435 158.560 276.415 ; 
                RECT 160.480 148.435 162.400 276.415 ; 
                RECT 199.005 148.435 200.925 276.415 ; 
                RECT 202.845 148.435 204.765 276.415 ; 
                RECT 206.685 148.435 208.605 276.415 ; 
                RECT 210.525 148.435 212.445 276.415 ; 
                RECT 214.365 148.435 216.285 276.415 ; 
                RECT 218.205 148.435 220.125 276.415 ; 
                RECT 222.045 148.435 223.965 276.415 ; 
                RECT 225.885 148.435 227.805 276.415 ; 
                RECT 229.725 148.435 231.645 276.415 ; 
                RECT 233.565 148.435 235.485 276.415 ; 
                RECT 237.405 148.435 239.325 276.415 ; 
                RECT 241.245 148.435 243.165 276.415 ; 
                RECT 245.085 148.435 247.005 276.415 ; 
                RECT 248.925 148.435 250.845 276.415 ; 
                RECT 252.765 148.435 254.685 276.415 ; 
                RECT 256.605 148.435 258.525 276.415 ; 
                RECT 260.445 148.435 262.365 276.415 ; 
                RECT 264.285 148.435 266.205 276.415 ; 
                RECT 268.125 148.435 270.045 276.415 ; 
                RECT 181.055 64.700 182.975 100.100 ; 
                RECT 187.575 64.700 189.115 100.100 ; 
                RECT 195.435 64.700 197.355 100.100 ; 
                RECT 206.955 64.700 208.875 100.100 ; 
                RECT 210.795 64.700 212.715 100.100 ; 
                RECT 214.635 64.700 216.555 100.100 ; 
                RECT 232.480 64.700 234.400 100.100 ; 
                RECT 236.320 64.700 238.240 100.100 ; 
                RECT 240.160 64.700 242.080 100.100 ; 
                RECT 244.000 64.700 245.920 100.100 ; 
                RECT 247.840 64.700 249.760 100.100 ; 
                RECT 251.680 64.700 253.600 100.100 ; 
                RECT 255.520 64.700 257.440 100.100 ; 
                RECT 206.620 118.840 208.540 141.800 ; 
                RECT 213.595 118.840 215.515 141.800 ; 
                RECT 220.225 118.840 221.975 141.800 ; 
                RECT 229.480 118.840 231.400 141.800 ; 
                RECT 243.810 118.840 245.730 141.800 ; 
                RECT 247.650 118.840 249.570 141.800 ; 
                RECT 251.490 118.840 253.410 141.800 ; 
                RECT 255.330 118.840 257.250 141.800 ; 
                RECT 208.615 106.100 210.365 112.840 ; 
                RECT 218.085 106.100 220.005 112.840 ; 
                RECT 236.100 106.100 238.020 112.840 ; 
                RECT 239.940 106.100 241.860 112.840 ; 
                RECT 243.780 106.100 245.700 112.840 ; 
                RECT 247.620 106.100 249.540 112.840 ; 
                RECT 251.460 106.100 253.380 112.840 ; 
                RECT 255.300 106.100 257.220 112.840 ; 
                RECT 256.535 53.540 258.285 58.700 ; 
                RECT 25.030 150.705 34.190 151.455 ; 
                RECT 25.030 155.460 34.190 157.380 ; 
                RECT 121.800 138.490 137.840 139.290 ; 
                RECT 102.600 139.200 119.840 140.890 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 285.720 5.560 ; 
                RECT 671.640 5.240 687.240 5.560 ; 
                RECT 2.880 6.600 687.240 6.920 ; 
                RECT 2.880 7.960 687.240 8.280 ; 
                RECT 2.880 9.320 259.880 9.640 ; 
                RECT 281.320 9.320 687.240 9.640 ; 
                RECT 2.880 10.680 275.520 11.000 ; 
                RECT 680.480 10.680 687.240 11.000 ; 
                RECT 2.880 12.040 275.520 12.360 ; 
                RECT 680.480 12.040 687.240 12.360 ; 
                RECT 2.880 13.400 198.000 13.720 ; 
                RECT 260.920 13.400 275.520 13.720 ; 
                RECT 680.480 13.400 687.240 13.720 ; 
                RECT 2.880 14.760 275.520 15.080 ; 
                RECT 680.480 14.760 687.240 15.080 ; 
                RECT 2.880 16.120 275.520 16.440 ; 
                RECT 680.480 16.120 687.240 16.440 ; 
                RECT 2.880 17.480 198.000 17.800 ; 
                RECT 260.240 17.480 275.520 17.800 ; 
                RECT 680.480 17.480 687.240 17.800 ; 
                RECT 2.880 18.840 275.520 19.160 ; 
                RECT 680.480 18.840 687.240 19.160 ; 
                RECT 2.880 20.200 275.520 20.520 ; 
                RECT 680.480 20.200 687.240 20.520 ; 
                RECT 2.880 21.560 275.520 21.880 ; 
                RECT 680.480 21.560 687.240 21.880 ; 
                RECT 2.880 22.920 275.520 23.240 ; 
                RECT 680.480 22.920 687.240 23.240 ; 
                RECT 2.880 24.280 275.520 24.600 ; 
                RECT 680.480 24.280 687.240 24.600 ; 
                RECT 2.880 25.640 275.520 25.960 ; 
                RECT 680.480 25.640 687.240 25.960 ; 
                RECT 2.880 27.000 275.520 27.320 ; 
                RECT 680.480 27.000 687.240 27.320 ; 
                RECT 2.880 28.360 274.840 28.680 ; 
                RECT 680.480 28.360 687.240 28.680 ; 
                RECT 2.880 29.720 275.520 30.040 ; 
                RECT 680.480 29.720 687.240 30.040 ; 
                RECT 2.880 31.080 275.520 31.400 ; 
                RECT 680.480 31.080 687.240 31.400 ; 
                RECT 2.880 32.440 275.520 32.760 ; 
                RECT 680.480 32.440 687.240 32.760 ; 
                RECT 2.880 33.800 168.760 34.120 ; 
                RECT 239.160 33.800 275.520 34.120 ; 
                RECT 680.480 33.800 687.240 34.120 ; 
                RECT 2.880 35.160 167.400 35.480 ; 
                RECT 245.280 35.160 275.520 35.480 ; 
                RECT 680.480 35.160 687.240 35.480 ; 
                RECT 2.880 36.520 144.280 36.840 ; 
                RECT 260.240 36.520 275.520 36.840 ; 
                RECT 680.480 36.520 687.240 36.840 ; 
                RECT 2.880 37.880 144.960 38.200 ; 
                RECT 250.720 37.880 275.520 38.200 ; 
                RECT 680.480 37.880 687.240 38.200 ; 
                RECT 2.880 39.240 275.520 39.560 ; 
                RECT 680.480 39.240 687.240 39.560 ; 
                RECT 2.880 40.600 275.520 40.920 ; 
                RECT 680.480 40.600 687.240 40.920 ; 
                RECT 2.880 41.960 275.520 42.280 ; 
                RECT 680.480 41.960 687.240 42.280 ; 
                RECT 2.880 43.320 275.520 43.640 ; 
                RECT 680.480 43.320 687.240 43.640 ; 
                RECT 2.880 44.680 142.240 45.000 ; 
                RECT 153.480 44.680 275.520 45.000 ; 
                RECT 680.480 44.680 687.240 45.000 ; 
                RECT 2.880 46.040 143.600 46.360 ; 
                RECT 146.000 46.040 275.520 46.360 ; 
                RECT 680.480 46.040 687.240 46.360 ; 
                RECT 2.880 47.400 144.960 47.720 ; 
                RECT 149.400 47.400 157.200 47.720 ; 
                RECT 159.600 47.400 275.520 47.720 ; 
                RECT 680.480 47.400 687.240 47.720 ; 
                RECT 2.880 48.760 144.960 49.080 ; 
                RECT 148.720 48.760 275.520 49.080 ; 
                RECT 680.480 48.760 687.240 49.080 ; 
                RECT 2.880 50.120 151.760 50.440 ; 
                RECT 160.280 50.120 275.520 50.440 ; 
                RECT 680.480 50.120 687.240 50.440 ; 
                RECT 2.880 51.480 147.000 51.800 ; 
                RECT 153.480 51.480 275.520 51.800 ; 
                RECT 680.480 51.480 687.240 51.800 ; 
                RECT 2.880 52.840 144.280 53.160 ; 
                RECT 153.480 52.840 275.520 53.160 ; 
                RECT 680.480 52.840 687.240 53.160 ; 
                RECT 2.880 54.200 253.080 54.520 ; 
                RECT 258.880 54.200 275.520 54.520 ; 
                RECT 680.480 54.200 687.240 54.520 ; 
                RECT 2.880 55.560 143.600 55.880 ; 
                RECT 153.480 55.560 253.080 55.880 ; 
                RECT 680.480 55.560 687.240 55.880 ; 
                RECT 2.880 56.920 151.760 57.240 ; 
                RECT 158.920 56.920 253.080 57.240 ; 
                RECT 680.480 56.920 687.240 57.240 ; 
                RECT 2.880 58.280 150.400 58.600 ; 
                RECT 153.480 58.280 165.360 58.600 ; 
                RECT 258.880 58.280 275.520 58.600 ; 
                RECT 680.480 58.280 687.240 58.600 ; 
                RECT 2.880 59.640 275.520 59.960 ; 
                RECT 680.480 59.640 687.240 59.960 ; 
                RECT 2.880 61.000 151.760 61.320 ; 
                RECT 159.600 61.000 275.520 61.320 ; 
                RECT 680.480 61.000 687.240 61.320 ; 
                RECT 2.880 62.360 148.360 62.680 ; 
                RECT 153.480 62.360 275.520 62.680 ; 
                RECT 680.480 62.360 687.240 62.680 ; 
                RECT 2.880 63.720 150.400 64.040 ; 
                RECT 153.480 63.720 275.520 64.040 ; 
                RECT 680.480 63.720 687.240 64.040 ; 
                RECT 2.880 65.080 154.480 65.400 ; 
                RECT 172.520 65.080 177.600 65.400 ; 
                RECT 258.200 65.080 275.520 65.400 ; 
                RECT 680.480 65.080 687.240 65.400 ; 
                RECT 2.880 66.440 141.560 66.760 ; 
                RECT 159.600 66.440 168.080 66.760 ; 
                RECT 171.160 66.440 177.600 66.760 ; 
                RECT 267.720 66.440 275.520 66.760 ; 
                RECT 680.480 66.440 687.240 66.760 ; 
                RECT 2.880 67.800 159.920 68.120 ; 
                RECT 166.400 67.800 177.600 68.120 ; 
                RECT 267.720 67.800 275.520 68.120 ; 
                RECT 680.480 67.800 687.240 68.120 ; 
                RECT 2.880 69.160 150.400 69.480 ; 
                RECT 153.480 69.160 163.320 69.480 ; 
                RECT 167.080 69.160 177.600 69.480 ; 
                RECT 266.360 69.160 275.520 69.480 ; 
                RECT 680.480 69.160 687.240 69.480 ; 
                RECT 2.880 70.520 142.240 70.840 ; 
                RECT 156.200 70.520 177.600 70.840 ; 
                RECT 267.720 70.520 275.520 70.840 ; 
                RECT 680.480 70.520 687.240 70.840 ; 
                RECT 2.880 71.880 151.080 72.200 ; 
                RECT 159.600 71.880 177.600 72.200 ; 
                RECT 267.720 71.880 275.520 72.200 ; 
                RECT 680.480 71.880 687.240 72.200 ; 
                RECT 2.880 73.240 149.040 73.560 ; 
                RECT 160.280 73.240 177.600 73.560 ; 
                RECT 266.360 73.240 275.520 73.560 ; 
                RECT 680.480 73.240 687.240 73.560 ; 
                RECT 2.880 74.600 144.280 74.920 ; 
                RECT 150.760 74.600 177.600 74.920 ; 
                RECT 270.440 74.600 275.520 74.920 ; 
                RECT 680.480 74.600 687.240 74.920 ; 
                RECT 2.880 75.960 177.600 76.280 ; 
                RECT 269.080 75.960 275.520 76.280 ; 
                RECT 680.480 75.960 687.240 76.280 ; 
                RECT 2.880 77.320 143.600 77.640 ; 
                RECT 147.360 77.320 177.600 77.640 ; 
                RECT 270.440 77.320 275.520 77.640 ; 
                RECT 680.480 77.320 687.240 77.640 ; 
                RECT 2.880 78.680 143.600 79.000 ; 
                RECT 153.480 78.680 177.600 79.000 ; 
                RECT 270.440 78.680 275.520 79.000 ; 
                RECT 680.480 78.680 687.240 79.000 ; 
                RECT 2.880 80.040 147.680 80.360 ; 
                RECT 158.920 80.040 177.600 80.360 ; 
                RECT 269.080 80.040 275.520 80.360 ; 
                RECT 680.480 80.040 687.240 80.360 ; 
                RECT 2.880 81.400 150.400 81.720 ; 
                RECT 152.800 81.400 177.600 81.720 ; 
                RECT 270.440 81.400 275.520 81.720 ; 
                RECT 680.480 81.400 687.240 81.720 ; 
                RECT 2.880 82.760 151.760 83.080 ; 
                RECT 153.480 82.760 177.600 83.080 ; 
                RECT 258.200 82.760 275.520 83.080 ; 
                RECT 680.480 82.760 687.240 83.080 ; 
                RECT 2.880 84.120 177.600 84.440 ; 
                RECT 273.160 84.120 275.520 84.440 ; 
                RECT 680.480 84.120 687.240 84.440 ; 
                RECT 2.880 85.480 142.240 85.800 ; 
                RECT 159.600 85.480 177.600 85.800 ; 
                RECT 273.160 85.480 275.520 85.800 ; 
                RECT 680.480 85.480 687.240 85.800 ; 
                RECT 2.880 86.840 145.640 87.160 ; 
                RECT 153.480 86.840 157.200 87.160 ; 
                RECT 159.600 86.840 177.600 87.160 ; 
                RECT 258.200 86.840 275.520 87.160 ; 
                RECT 680.480 86.840 687.240 87.160 ; 
                RECT 2.880 88.200 151.080 88.520 ; 
                RECT 153.480 88.200 177.600 88.520 ; 
                RECT 271.800 88.200 275.520 88.520 ; 
                RECT 680.480 88.200 687.240 88.520 ; 
                RECT 2.880 89.560 177.600 89.880 ; 
                RECT 273.160 89.560 275.520 89.880 ; 
                RECT 680.480 89.560 687.240 89.880 ; 
                RECT 2.880 90.920 177.600 91.240 ; 
                RECT 258.200 90.920 275.520 91.240 ; 
                RECT 680.480 90.920 687.240 91.240 ; 
                RECT 2.880 92.280 138.840 92.600 ; 
                RECT 152.120 92.280 177.600 92.600 ; 
                RECT 680.480 92.280 687.240 92.600 ; 
                RECT 2.880 93.640 149.040 93.960 ; 
                RECT 156.200 93.640 177.600 93.960 ; 
                RECT 680.480 93.640 687.240 93.960 ; 
                RECT 2.880 95.000 177.600 95.320 ; 
                RECT 680.480 95.000 687.240 95.320 ; 
                RECT 2.880 96.360 177.600 96.680 ; 
                RECT 680.480 96.360 687.240 96.680 ; 
                RECT 2.880 97.720 147.680 98.040 ; 
                RECT 161.640 97.720 177.600 98.040 ; 
                RECT 680.480 97.720 687.240 98.040 ; 
                RECT 2.880 99.080 177.600 99.400 ; 
                RECT 680.480 99.080 687.240 99.400 ; 
                RECT 2.880 100.440 177.600 100.760 ; 
                RECT 258.200 100.440 275.520 100.760 ; 
                RECT 680.480 100.440 687.240 100.760 ; 
                RECT 2.880 101.800 144.280 102.120 ; 
                RECT 147.360 101.800 275.520 102.120 ; 
                RECT 680.480 101.800 687.240 102.120 ; 
                RECT 2.880 103.160 141.560 103.480 ; 
                RECT 146.000 103.160 275.520 103.480 ; 
                RECT 680.480 103.160 687.240 103.480 ; 
                RECT 2.880 104.520 261.920 104.840 ; 
                RECT 680.480 104.520 687.240 104.840 ; 
                RECT 2.880 105.880 157.200 106.200 ; 
                RECT 160.280 105.880 205.480 106.200 ; 
                RECT 258.200 105.880 272.800 106.200 ; 
                RECT 680.480 105.880 687.240 106.200 ; 
                RECT 2.880 107.240 205.480 107.560 ; 
                RECT 258.200 107.240 270.080 107.560 ; 
                RECT 680.480 107.240 687.240 107.560 ; 
                RECT 2.880 108.600 120.480 108.920 ; 
                RECT 139.200 108.600 205.480 108.920 ; 
                RECT 258.200 108.600 267.360 108.920 ; 
                RECT 680.480 108.600 687.240 108.920 ; 
                RECT 2.880 109.960 120.480 110.280 ; 
                RECT 139.200 109.960 205.480 110.280 ; 
                RECT 258.200 109.960 264.640 110.280 ; 
                RECT 680.480 109.960 687.240 110.280 ; 
                RECT 2.880 111.320 120.480 111.640 ; 
                RECT 139.200 111.320 144.280 111.640 ; 
                RECT 149.400 111.320 205.480 111.640 ; 
                RECT 258.200 111.320 275.520 111.640 ; 
                RECT 680.480 111.320 687.240 111.640 ; 
                RECT 2.880 112.680 120.480 113.000 ; 
                RECT 139.200 112.680 205.480 113.000 ; 
                RECT 258.200 112.680 275.520 113.000 ; 
                RECT 680.480 112.680 687.240 113.000 ; 
                RECT 2.880 114.040 120.480 114.360 ; 
                RECT 139.200 114.040 147.680 114.360 ; 
                RECT 158.920 114.040 275.520 114.360 ; 
                RECT 680.480 114.040 687.240 114.360 ; 
                RECT 2.880 115.400 120.480 115.720 ; 
                RECT 139.200 115.400 275.520 115.720 ; 
                RECT 680.480 115.400 687.240 115.720 ; 
                RECT 2.880 116.760 120.480 117.080 ; 
                RECT 139.200 116.760 275.520 117.080 ; 
                RECT 680.480 116.760 687.240 117.080 ; 
                RECT 2.880 118.120 120.480 118.440 ; 
                RECT 139.200 118.120 143.600 118.440 ; 
                RECT 146.680 118.120 275.520 118.440 ; 
                RECT 680.480 118.120 687.240 118.440 ; 
                RECT 2.880 119.480 120.480 119.800 ; 
                RECT 139.880 119.480 144.280 119.800 ; 
                RECT 149.400 119.480 202.760 119.800 ; 
                RECT 258.200 119.480 275.520 119.800 ; 
                RECT 680.480 119.480 687.240 119.800 ; 
                RECT 2.880 120.840 120.480 121.160 ; 
                RECT 139.200 120.840 202.760 121.160 ; 
                RECT 258.200 120.840 275.520 121.160 ; 
                RECT 680.480 120.840 687.240 121.160 ; 
                RECT 2.880 122.200 120.480 122.520 ; 
                RECT 139.200 122.200 202.760 122.520 ; 
                RECT 258.200 122.200 275.520 122.520 ; 
                RECT 680.480 122.200 687.240 122.520 ; 
                RECT 2.880 123.560 120.480 123.880 ; 
                RECT 139.200 123.560 202.760 123.880 ; 
                RECT 258.200 123.560 275.520 123.880 ; 
                RECT 680.480 123.560 687.240 123.880 ; 
                RECT 2.880 124.920 120.480 125.240 ; 
                RECT 139.200 124.920 202.760 125.240 ; 
                RECT 258.200 124.920 266.000 125.240 ; 
                RECT 680.480 124.920 687.240 125.240 ; 
                RECT 2.880 126.280 120.480 126.600 ; 
                RECT 139.200 126.280 202.760 126.600 ; 
                RECT 258.200 126.280 268.720 126.600 ; 
                RECT 680.480 126.280 687.240 126.600 ; 
                RECT 2.880 127.640 120.480 127.960 ; 
                RECT 139.200 127.640 202.760 127.960 ; 
                RECT 258.200 127.640 271.440 127.960 ; 
                RECT 680.480 127.640 687.240 127.960 ; 
                RECT 2.880 129.000 120.480 129.320 ; 
                RECT 139.200 129.000 202.760 129.320 ; 
                RECT 258.200 129.000 274.160 129.320 ; 
                RECT 680.480 129.000 687.240 129.320 ; 
                RECT 2.880 130.360 120.480 130.680 ; 
                RECT 139.200 130.360 145.640 130.680 ; 
                RECT 149.400 130.360 202.760 130.680 ; 
                RECT 680.480 130.360 687.240 130.680 ; 
                RECT 2.880 131.720 120.480 132.040 ; 
                RECT 139.200 131.720 202.760 132.040 ; 
                RECT 258.200 131.720 275.520 132.040 ; 
                RECT 680.480 131.720 687.240 132.040 ; 
                RECT 2.880 133.080 202.760 133.400 ; 
                RECT 258.200 133.080 275.520 133.400 ; 
                RECT 680.480 133.080 687.240 133.400 ; 
                RECT 2.880 134.440 202.760 134.760 ; 
                RECT 258.200 134.440 275.520 134.760 ; 
                RECT 680.480 134.440 687.240 134.760 ; 
                RECT 2.880 135.800 102.120 136.120 ; 
                RECT 120.840 135.800 147.680 136.120 ; 
                RECT 153.480 135.800 202.760 136.120 ; 
                RECT 258.200 135.800 275.520 136.120 ; 
                RECT 680.480 135.800 687.240 136.120 ; 
                RECT 2.880 137.160 102.120 137.480 ; 
                RECT 120.840 137.160 126.600 137.480 ; 
                RECT 133.760 137.160 202.760 137.480 ; 
                RECT 258.200 137.160 275.520 137.480 ; 
                RECT 680.480 137.160 687.240 137.480 ; 
                RECT 2.880 138.520 102.120 138.840 ; 
                RECT 138.520 138.520 202.760 138.840 ; 
                RECT 258.200 138.520 275.520 138.840 ; 
                RECT 680.480 138.520 687.240 138.840 ; 
                RECT 2.880 139.880 102.120 140.200 ; 
                RECT 120.840 139.880 202.760 140.200 ; 
                RECT 680.480 139.880 687.240 140.200 ; 
                RECT 2.880 141.240 100.760 141.560 ; 
                RECT 133.760 141.240 146.320 141.560 ; 
                RECT 152.120 141.240 202.760 141.560 ; 
                RECT 258.200 141.240 275.520 141.560 ; 
                RECT 680.480 141.240 687.240 141.560 ; 
                RECT 2.880 142.600 126.600 142.920 ; 
                RECT 146.680 142.600 687.240 142.920 ; 
                RECT 2.880 143.960 31.400 144.280 ; 
                RECT 146.000 143.960 687.240 144.280 ; 
                RECT 2.880 145.320 272.800 145.640 ; 
                RECT 682.520 145.320 687.240 145.640 ; 
                RECT 2.880 146.680 272.800 147.000 ; 
                RECT 682.520 146.680 687.240 147.000 ; 
                RECT 2.880 148.040 26.640 148.360 ; 
                RECT 33.120 148.040 80.360 148.360 ; 
                RECT 682.520 148.040 687.240 148.360 ; 
                RECT 2.880 149.400 24.600 149.720 ; 
                RECT 46.720 149.400 80.360 149.720 ; 
                RECT 682.520 149.400 687.240 149.720 ; 
                RECT 2.880 150.760 24.600 151.080 ; 
                RECT 46.040 150.760 59.960 151.080 ; 
                RECT 69.840 150.760 80.360 151.080 ; 
                RECT 682.520 150.760 687.240 151.080 ; 
                RECT 2.880 152.120 38.200 152.440 ; 
                RECT 44.680 152.120 59.960 152.440 ; 
                RECT 69.840 152.120 80.360 152.440 ; 
                RECT 682.520 152.120 687.240 152.440 ; 
                RECT 2.880 153.480 24.600 153.800 ; 
                RECT 35.160 153.480 59.960 153.800 ; 
                RECT 69.840 153.480 80.360 153.800 ; 
                RECT 682.520 153.480 687.240 153.800 ; 
                RECT 2.880 154.840 24.600 155.160 ; 
                RECT 35.160 154.840 59.960 155.160 ; 
                RECT 69.840 154.840 80.360 155.160 ; 
                RECT 682.520 154.840 687.240 155.160 ; 
                RECT 2.880 156.200 24.600 156.520 ; 
                RECT 35.160 156.200 59.960 156.520 ; 
                RECT 69.840 156.200 80.360 156.520 ; 
                RECT 682.520 156.200 687.240 156.520 ; 
                RECT 2.880 157.560 24.600 157.880 ; 
                RECT 35.160 157.560 80.360 157.880 ; 
                RECT 682.520 157.560 687.240 157.880 ; 
                RECT 2.880 158.920 59.960 159.240 ; 
                RECT 69.840 158.920 80.360 159.240 ; 
                RECT 682.520 158.920 687.240 159.240 ; 
                RECT 2.880 160.280 59.960 160.600 ; 
                RECT 69.840 160.280 80.360 160.600 ; 
                RECT 682.520 160.280 687.240 160.600 ; 
                RECT 2.880 161.640 17.800 161.960 ; 
                RECT 20.200 161.640 59.960 161.960 ; 
                RECT 69.840 161.640 80.360 161.960 ; 
                RECT 682.520 161.640 687.240 161.960 ; 
                RECT 2.880 163.000 17.120 163.320 ; 
                RECT 20.200 163.000 59.960 163.320 ; 
                RECT 69.840 163.000 80.360 163.320 ; 
                RECT 682.520 163.000 687.240 163.320 ; 
                RECT 2.880 164.360 59.960 164.680 ; 
                RECT 67.120 164.360 80.360 164.680 ; 
                RECT 682.520 164.360 687.240 164.680 ; 
                RECT 2.880 165.720 16.440 166.040 ; 
                RECT 20.200 165.720 33.440 166.040 ; 
                RECT 37.200 165.720 64.040 166.040 ; 
                RECT 69.840 165.720 80.360 166.040 ; 
                RECT 682.520 165.720 687.240 166.040 ; 
                RECT 2.880 167.080 15.760 167.400 ; 
                RECT 20.200 167.080 33.440 167.400 ; 
                RECT 37.880 167.080 59.960 167.400 ; 
                RECT 69.840 167.080 80.360 167.400 ; 
                RECT 682.520 167.080 687.240 167.400 ; 
                RECT 2.880 168.440 59.960 168.760 ; 
                RECT 69.840 168.440 80.360 168.760 ; 
                RECT 682.520 168.440 687.240 168.760 ; 
                RECT 2.880 169.800 15.080 170.120 ; 
                RECT 20.200 169.800 33.440 170.120 ; 
                RECT 38.560 169.800 59.960 170.120 ; 
                RECT 69.840 169.800 80.360 170.120 ; 
                RECT 682.520 169.800 687.240 170.120 ; 
                RECT 2.880 171.160 14.400 171.480 ; 
                RECT 20.200 171.160 33.440 171.480 ; 
                RECT 39.240 171.160 59.960 171.480 ; 
                RECT 69.840 171.160 80.360 171.480 ; 
                RECT 682.520 171.160 687.240 171.480 ; 
                RECT 2.880 172.520 13.720 172.840 ; 
                RECT 20.200 172.520 33.440 172.840 ; 
                RECT 39.240 172.520 59.960 172.840 ; 
                RECT 67.800 172.520 80.360 172.840 ; 
                RECT 682.520 172.520 687.240 172.840 ; 
                RECT 2.880 173.880 13.040 174.200 ; 
                RECT 20.200 173.880 66.080 174.200 ; 
                RECT 69.840 173.880 80.360 174.200 ; 
                RECT 682.520 173.880 687.240 174.200 ; 
                RECT 2.880 175.240 59.960 175.560 ; 
                RECT 69.840 175.240 80.360 175.560 ; 
                RECT 682.520 175.240 687.240 175.560 ; 
                RECT 2.880 176.600 12.360 176.920 ; 
                RECT 20.200 176.600 59.960 176.920 ; 
                RECT 69.840 176.600 80.360 176.920 ; 
                RECT 682.520 176.600 687.240 176.920 ; 
                RECT 2.880 177.960 11.680 178.280 ; 
                RECT 20.200 177.960 59.960 178.280 ; 
                RECT 69.840 177.960 80.360 178.280 ; 
                RECT 682.520 177.960 687.240 178.280 ; 
                RECT 2.880 179.320 11.000 179.640 ; 
                RECT 20.200 179.320 59.960 179.640 ; 
                RECT 69.840 179.320 80.360 179.640 ; 
                RECT 682.520 179.320 687.240 179.640 ; 
                RECT 2.880 180.680 80.360 181.000 ; 
                RECT 682.520 180.680 687.240 181.000 ; 
                RECT 2.880 182.040 10.320 182.360 ; 
                RECT 20.200 182.040 33.440 182.360 ; 
                RECT 35.840 182.040 61.320 182.360 ; 
                RECT 69.840 182.040 80.360 182.360 ; 
                RECT 682.520 182.040 687.240 182.360 ; 
                RECT 2.880 183.400 64.720 183.720 ; 
                RECT 69.840 183.400 80.360 183.720 ; 
                RECT 682.520 183.400 687.240 183.720 ; 
                RECT 2.880 184.760 64.720 185.080 ; 
                RECT 69.840 184.760 80.360 185.080 ; 
                RECT 682.520 184.760 687.240 185.080 ; 
                RECT 2.880 186.120 61.320 186.440 ; 
                RECT 69.840 186.120 80.360 186.440 ; 
                RECT 682.520 186.120 687.240 186.440 ; 
                RECT 2.880 187.480 61.320 187.800 ; 
                RECT 69.840 187.480 80.360 187.800 ; 
                RECT 682.520 187.480 687.240 187.800 ; 
                RECT 2.880 188.840 37.520 189.160 ; 
                RECT 46.720 188.840 80.360 189.160 ; 
                RECT 682.520 188.840 687.240 189.160 ; 
                RECT 2.880 190.200 36.160 190.520 ; 
                RECT 46.040 190.200 61.320 190.520 ; 
                RECT 69.840 190.200 80.360 190.520 ; 
                RECT 682.520 190.200 687.240 190.520 ; 
                RECT 2.880 191.560 34.800 191.880 ; 
                RECT 44.680 191.560 59.960 191.880 ; 
                RECT 69.840 191.560 80.360 191.880 ; 
                RECT 682.520 191.560 687.240 191.880 ; 
                RECT 2.880 192.920 59.960 193.240 ; 
                RECT 69.840 192.920 80.360 193.240 ; 
                RECT 682.520 192.920 687.240 193.240 ; 
                RECT 2.880 194.280 59.960 194.600 ; 
                RECT 69.840 194.280 80.360 194.600 ; 
                RECT 682.520 194.280 687.240 194.600 ; 
                RECT 2.880 195.640 59.960 195.960 ; 
                RECT 69.840 195.640 80.360 195.960 ; 
                RECT 682.520 195.640 687.240 195.960 ; 
                RECT 2.880 197.000 80.360 197.320 ; 
                RECT 682.520 197.000 687.240 197.320 ; 
                RECT 2.880 198.360 59.960 198.680 ; 
                RECT 69.840 198.360 80.360 198.680 ; 
                RECT 682.520 198.360 687.240 198.680 ; 
                RECT 2.880 199.720 59.960 200.040 ; 
                RECT 69.840 199.720 80.360 200.040 ; 
                RECT 682.520 199.720 687.240 200.040 ; 
                RECT 2.880 201.080 59.960 201.400 ; 
                RECT 69.840 201.080 80.360 201.400 ; 
                RECT 682.520 201.080 687.240 201.400 ; 
                RECT 2.880 202.440 59.960 202.760 ; 
                RECT 69.840 202.440 80.360 202.760 ; 
                RECT 682.520 202.440 687.240 202.760 ; 
                RECT 2.880 203.800 59.960 204.120 ; 
                RECT 63.040 203.800 80.360 204.120 ; 
                RECT 682.520 203.800 687.240 204.120 ; 
                RECT 2.880 205.160 66.080 205.480 ; 
                RECT 69.840 205.160 80.360 205.480 ; 
                RECT 682.520 205.160 687.240 205.480 ; 
                RECT 2.880 206.520 59.960 206.840 ; 
                RECT 69.840 206.520 80.360 206.840 ; 
                RECT 682.520 206.520 687.240 206.840 ; 
                RECT 2.880 207.880 59.960 208.200 ; 
                RECT 69.840 207.880 80.360 208.200 ; 
                RECT 682.520 207.880 687.240 208.200 ; 
                RECT 2.880 209.240 59.960 209.560 ; 
                RECT 69.840 209.240 80.360 209.560 ; 
                RECT 682.520 209.240 687.240 209.560 ; 
                RECT 2.880 210.600 59.960 210.920 ; 
                RECT 69.840 210.600 80.360 210.920 ; 
                RECT 682.520 210.600 687.240 210.920 ; 
                RECT 2.880 211.960 59.960 212.280 ; 
                RECT 64.400 211.960 80.360 212.280 ; 
                RECT 682.520 211.960 687.240 212.280 ; 
                RECT 2.880 213.320 64.040 213.640 ; 
                RECT 69.840 213.320 80.360 213.640 ; 
                RECT 682.520 213.320 687.240 213.640 ; 
                RECT 2.880 214.680 59.960 215.000 ; 
                RECT 69.840 214.680 80.360 215.000 ; 
                RECT 682.520 214.680 687.240 215.000 ; 
                RECT 2.880 216.040 59.960 216.360 ; 
                RECT 69.840 216.040 80.360 216.360 ; 
                RECT 682.520 216.040 687.240 216.360 ; 
                RECT 2.880 217.400 59.960 217.720 ; 
                RECT 69.840 217.400 80.360 217.720 ; 
                RECT 682.520 217.400 687.240 217.720 ; 
                RECT 2.880 218.760 59.960 219.080 ; 
                RECT 69.840 218.760 80.360 219.080 ; 
                RECT 682.520 218.760 687.240 219.080 ; 
                RECT 2.880 220.120 80.360 220.440 ; 
                RECT 682.520 220.120 687.240 220.440 ; 
                RECT 2.880 221.480 62.000 221.800 ; 
                RECT 69.840 221.480 80.360 221.800 ; 
                RECT 682.520 221.480 687.240 221.800 ; 
                RECT 2.880 222.840 66.080 223.160 ; 
                RECT 69.840 222.840 80.360 223.160 ; 
                RECT 682.520 222.840 687.240 223.160 ; 
                RECT 2.880 224.200 62.000 224.520 ; 
                RECT 69.840 224.200 80.360 224.520 ; 
                RECT 682.520 224.200 687.240 224.520 ; 
                RECT 2.880 225.560 62.000 225.880 ; 
                RECT 69.840 225.560 80.360 225.880 ; 
                RECT 682.520 225.560 687.240 225.880 ; 
                RECT 2.880 226.920 62.000 227.240 ; 
                RECT 69.840 226.920 80.360 227.240 ; 
                RECT 682.520 226.920 687.240 227.240 ; 
                RECT 2.880 228.280 80.360 228.600 ; 
                RECT 682.520 228.280 687.240 228.600 ; 
                RECT 2.880 229.640 62.680 229.960 ; 
                RECT 69.840 229.640 80.360 229.960 ; 
                RECT 682.520 229.640 687.240 229.960 ; 
                RECT 2.880 231.000 62.680 231.320 ; 
                RECT 69.840 231.000 80.360 231.320 ; 
                RECT 682.520 231.000 687.240 231.320 ; 
                RECT 2.880 232.360 64.720 232.680 ; 
                RECT 69.840 232.360 80.360 232.680 ; 
                RECT 682.520 232.360 687.240 232.680 ; 
                RECT 2.880 233.720 65.400 234.040 ; 
                RECT 69.840 233.720 80.360 234.040 ; 
                RECT 682.520 233.720 687.240 234.040 ; 
                RECT 2.880 235.080 62.680 235.400 ; 
                RECT 69.840 235.080 80.360 235.400 ; 
                RECT 682.520 235.080 687.240 235.400 ; 
                RECT 2.880 236.440 80.360 236.760 ; 
                RECT 682.520 236.440 687.240 236.760 ; 
                RECT 2.880 237.800 62.680 238.120 ; 
                RECT 69.840 237.800 80.360 238.120 ; 
                RECT 682.520 237.800 687.240 238.120 ; 
                RECT 2.880 239.160 62.680 239.480 ; 
                RECT 69.840 239.160 80.360 239.480 ; 
                RECT 682.520 239.160 687.240 239.480 ; 
                RECT 2.880 240.520 62.680 240.840 ; 
                RECT 69.840 240.520 80.360 240.840 ; 
                RECT 682.520 240.520 687.240 240.840 ; 
                RECT 2.880 241.880 62.680 242.200 ; 
                RECT 69.840 241.880 80.360 242.200 ; 
                RECT 682.520 241.880 687.240 242.200 ; 
                RECT 2.880 243.240 80.360 243.560 ; 
                RECT 682.520 243.240 687.240 243.560 ; 
                RECT 2.880 244.600 64.040 244.920 ; 
                RECT 69.840 244.600 80.360 244.920 ; 
                RECT 682.520 244.600 687.240 244.920 ; 
                RECT 2.880 245.960 62.680 246.280 ; 
                RECT 69.840 245.960 80.360 246.280 ; 
                RECT 682.520 245.960 687.240 246.280 ; 
                RECT 2.880 247.320 62.680 247.640 ; 
                RECT 69.840 247.320 80.360 247.640 ; 
                RECT 682.520 247.320 687.240 247.640 ; 
                RECT 2.880 248.680 62.680 249.000 ; 
                RECT 69.840 248.680 80.360 249.000 ; 
                RECT 682.520 248.680 687.240 249.000 ; 
                RECT 2.880 250.040 62.680 250.360 ; 
                RECT 69.840 250.040 80.360 250.360 ; 
                RECT 682.520 250.040 687.240 250.360 ; 
                RECT 2.880 251.400 80.360 251.720 ; 
                RECT 682.520 251.400 687.240 251.720 ; 
                RECT 2.880 252.760 66.080 253.080 ; 
                RECT 69.840 252.760 80.360 253.080 ; 
                RECT 682.520 252.760 687.240 253.080 ; 
                RECT 2.880 254.120 62.680 254.440 ; 
                RECT 69.840 254.120 80.360 254.440 ; 
                RECT 682.520 254.120 687.240 254.440 ; 
                RECT 2.880 255.480 62.680 255.800 ; 
                RECT 69.840 255.480 80.360 255.800 ; 
                RECT 682.520 255.480 687.240 255.800 ; 
                RECT 2.880 256.840 62.680 257.160 ; 
                RECT 69.840 256.840 80.360 257.160 ; 
                RECT 682.520 256.840 687.240 257.160 ; 
                RECT 2.880 258.200 62.680 258.520 ; 
                RECT 69.840 258.200 80.360 258.520 ; 
                RECT 682.520 258.200 687.240 258.520 ; 
                RECT 2.880 259.560 80.360 259.880 ; 
                RECT 682.520 259.560 687.240 259.880 ; 
                RECT 2.880 260.920 63.360 261.240 ; 
                RECT 69.840 260.920 80.360 261.240 ; 
                RECT 682.520 260.920 687.240 261.240 ; 
                RECT 2.880 262.280 64.720 262.600 ; 
                RECT 69.840 262.280 80.360 262.600 ; 
                RECT 682.520 262.280 687.240 262.600 ; 
                RECT 2.880 263.640 63.360 263.960 ; 
                RECT 69.840 263.640 80.360 263.960 ; 
                RECT 682.520 263.640 687.240 263.960 ; 
                RECT 2.880 265.000 63.360 265.320 ; 
                RECT 69.840 265.000 80.360 265.320 ; 
                RECT 682.520 265.000 687.240 265.320 ; 
                RECT 2.880 266.360 63.360 266.680 ; 
                RECT 69.840 266.360 80.360 266.680 ; 
                RECT 682.520 266.360 687.240 266.680 ; 
                RECT 2.880 267.720 80.360 268.040 ; 
                RECT 682.520 267.720 687.240 268.040 ; 
                RECT 2.880 269.080 63.360 269.400 ; 
                RECT 69.840 269.080 80.360 269.400 ; 
                RECT 682.520 269.080 687.240 269.400 ; 
                RECT 2.880 270.440 63.360 270.760 ; 
                RECT 69.840 270.440 80.360 270.760 ; 
                RECT 682.520 270.440 687.240 270.760 ; 
                RECT 2.880 271.800 66.760 272.120 ; 
                RECT 69.840 271.800 80.360 272.120 ; 
                RECT 682.520 271.800 687.240 272.120 ; 
                RECT 2.880 273.160 63.360 273.480 ; 
                RECT 69.840 273.160 80.360 273.480 ; 
                RECT 682.520 273.160 687.240 273.480 ; 
                RECT 2.880 274.520 63.360 274.840 ; 
                RECT 69.840 274.520 80.360 274.840 ; 
                RECT 682.520 274.520 687.240 274.840 ; 
                RECT 2.880 275.880 80.360 276.200 ; 
                RECT 682.520 275.880 687.240 276.200 ; 
                RECT 2.880 277.240 272.800 277.560 ; 
                RECT 682.520 277.240 687.240 277.560 ; 
                RECT 2.880 278.600 272.800 278.920 ; 
                RECT 682.520 278.600 687.240 278.920 ; 
                RECT 2.880 279.960 272.800 280.280 ; 
                RECT 682.520 279.960 687.240 280.280 ; 
                RECT 2.880 281.320 687.240 281.640 ; 
                RECT 2.880 282.680 687.240 283.000 ; 
                RECT 2.880 284.040 687.240 284.360 ; 
                RECT 2.880 285.400 687.240 285.720 ; 
                RECT 2.880 2.880 687.240 4.240 ; 
                RECT 2.880 287.400 687.240 288.760 ; 
                RECT 276.940 29.630 282.740 30.750 ; 
                RECT 672.840 29.630 678.640 30.750 ; 
                RECT 276.940 35.495 282.740 36.265 ; 
                RECT 672.840 35.495 678.640 36.265 ; 
                RECT 276.940 41.530 282.740 42.230 ; 
                RECT 672.840 41.530 678.640 42.230 ; 
                RECT 276.940 47.120 282.740 47.820 ; 
                RECT 672.840 47.120 678.640 47.820 ; 
                RECT 276.940 78.350 678.640 79.150 ; 
                RECT 276.940 81.590 678.640 83.680 ; 
                RECT 276.940 61.400 678.640 63.200 ; 
                RECT 276.940 120.970 678.640 122.375 ; 
                RECT 276.940 70.450 678.640 71.250 ; 
                RECT 276.940 102.695 678.640 102.985 ; 
                RECT 276.940 73.460 678.640 74.260 ; 
                RECT 276.940 75.140 678.640 75.940 ; 
                RECT 276.940 20.260 678.640 22.060 ; 
                RECT 80.800 148.435 82.550 276.415 ; 
                RECT 94.785 148.435 96.705 276.415 ; 
                RECT 118.560 148.435 120.480 276.415 ; 
                RECT 122.400 148.435 124.320 276.415 ; 
                RECT 126.240 148.435 128.160 276.415 ; 
                RECT 168.810 148.435 170.730 276.415 ; 
                RECT 172.650 148.435 174.570 276.415 ; 
                RECT 176.490 148.435 178.410 276.415 ; 
                RECT 180.330 148.435 182.250 276.415 ; 
                RECT 184.170 148.435 186.090 276.415 ; 
                RECT 188.010 148.435 189.930 276.415 ; 
                RECT 191.850 148.435 193.770 276.415 ; 
                RECT 178.430 64.700 179.320 100.100 ; 
                RECT 185.190 64.700 186.080 100.100 ; 
                RECT 191.305 64.700 192.625 100.100 ; 
                RECT 201.635 64.700 203.555 100.100 ; 
                RECT 219.820 64.700 221.740 100.100 ; 
                RECT 223.660 64.700 225.580 100.100 ; 
                RECT 227.500 64.700 229.420 100.100 ; 
                RECT 203.455 118.840 204.565 141.800 ; 
                RECT 210.970 118.840 211.860 141.800 ; 
                RECT 217.730 118.840 218.620 141.800 ; 
                RECT 224.380 118.840 225.920 141.800 ; 
                RECT 237.185 118.840 239.105 141.800 ; 
                RECT 206.120 106.100 207.010 112.840 ; 
                RECT 212.770 106.100 214.310 112.840 ; 
                RECT 225.805 106.100 227.725 112.840 ; 
                RECT 229.645 106.100 231.565 112.840 ; 
                RECT 254.040 53.540 254.930 58.700 ; 
                RECT 25.030 149.500 34.190 149.870 ; 
                RECT 25.030 152.835 34.190 153.725 ; 
                RECT 102.600 135.860 119.840 136.530 ; 
                RECT 102.600 137.160 119.840 138.170 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 690.120 291.640 ; 
        LAYER met2 ;
            RECT 0.000 0.000 690.120 291.640 ; 
    END 
END sram22_256x64m4w8 
END LIBRARY 

