VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sramgen_sram_2048x32m8w8_replica_v1
  CLASS BLOCK ;
  ORIGIN 87.435 582.85 ;
  FOREIGN sramgen_sram_2048x32m8w8_replica_v1 -87.435 -582.85 ;
  SIZE 749.895 BY 594.565 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -81.8 -582.45 -81.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -80.2 -582.45 -79.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -78.6 -582.45 -78.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -77 -582.45 -76.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -75.4 -551.52 -75 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.8 -569.54 -73.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.8 -582.45 -73.4 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.2 -582.45 -71.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.6 -564.24 -70.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.6 -582.45 -70.2 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -69 -569.54 -68.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -569.54 -67 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -582.45 -67 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.8 -582.45 -65.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -564.24 -63.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -582.45 -63.8 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.6 -569.54 -62.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -61 -582.45 -60.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -562.12 -59 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -582.45 -59 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.8 -569.54 -57.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -569.54 -55.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -582.45 -55.8 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.6 -582.45 -54.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -561.06 -52.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -582.45 -52.6 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.4 -569.54 -51 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -569.54 -49.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -582.45 -49.4 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.2 -582.45 -47.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -561.06 -46.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -582.45 -46.2 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -569.54 -44.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -582.45 -44.6 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.4 -582.45 -43 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -558.94 -41.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -582.45 -41.4 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.2 -569.54 -39.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -569.54 -38.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -582.45 -38.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -37 -582.45 -36.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -557.88 -35 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -582.45 -35 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.8 -569.54 -33.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.2 -582.45 -31.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -557.88 -30.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -582.45 -30.2 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -557.88 -28.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -582.45 -28.6 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -569.54 -27 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -582.45 -27 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.8 -582.45 -25.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -556.82 -23.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -582.45 -23.8 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.6 -569.54 -22.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -569.54 -20.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -582.45 -20.6 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.4 -582.45 -19 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -555.76 -17.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -582.45 -17.4 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.2 -569.54 -15.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.6 -582.45 -14.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -554.7 -12.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -582.45 -12.6 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -554.7 -11 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -582.45 -11 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -413.72 -9.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -569.54 -9.4 -533.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -582.45 -9.4 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.2 -582.45 -7.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -550.46 -6.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -582.45 -6.2 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -5 -582.45 -4.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.4 -582.45 -3 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 2.86 -1.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 -582.45 -1.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 2.86 0.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 -582.45 0.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 2.86 1.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 -582.45 1.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 2.86 3.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 -582.45 3.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 2.86 5 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 -582.45 5 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 2.86 6.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -582.45 6.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 2.86 8.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -582.45 8.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 2.86 9.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -582.45 9.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 2.86 11.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -461.42 11.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -582.45 11.4 -531.8 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 2.86 13 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -424.32 13 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -497.46 13 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 2.86 14.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -434.92 14.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -582.45 14.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 2.86 16.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 -582.45 16.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 2.86 17.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 -582.45 17.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 2.86 19.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -582.45 19.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 2.86 21 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -582.45 21 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 2.86 22.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 -503.82 22.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 2.86 24.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 -502.76 24.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 2.86 25.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 -582.45 25.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 2.86 27.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 -582.45 27.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 2.86 29 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -582.45 29 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 2.86 30.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -582.45 30.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 2.86 32.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 -582.45 32.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 2.86 33.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -424.32 33.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -497.46 33.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 2.86 35.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -424.32 35.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -582.45 35.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 2.86 37 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -440.22 37 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -582.45 37 -521.2 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 2.86 38.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -582.45 38.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 2.86 40.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -582.45 40.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 2.86 41.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 -582.45 41.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 2.86 43.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 -582.45 43.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 2.86 45 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 -582.45 45 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 2.86 46.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 -582.45 46.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 2.86 48.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -582.45 48.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 2.86 49.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -582.45 49.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 2.86 51.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 -582.45 51.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 2.86 53 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -424.32 53 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -497.46 53 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 2.86 54.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -434.92 54.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -582.45 54.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 2.86 56.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 -582.45 56.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 2.86 57.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 -582.45 57.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 2.86 59.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -582.45 59.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 2.86 61 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -582.45 61 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 2.86 62.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 -503.82 62.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 2.86 64.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -502.76 64.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -582.45 64.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 2.86 65.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 -582.45 65.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 2.86 67.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 -582.45 67.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 2.86 69 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -582.45 69 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 2.86 70.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -582.45 70.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 2.86 72.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 -582.45 72.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 2.86 73.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -424.32 73.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -497.46 73.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 2.86 75.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -424.32 75.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -582.45 75.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 2.86 77 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 -582.45 77 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 2.86 78.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -582.45 78.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 2.86 80.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -582.45 80.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 2.86 81.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 -582.45 81.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 2.86 83.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 -582.45 83.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 2.86 85 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 -582.45 85 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 2.86 86.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 -582.45 86.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 2.86 88.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -582.45 88.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 2.86 89.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -582.45 89.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 2.86 91.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 -582.45 91.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 2.86 93 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -424.32 93 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -497.46 93 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 2.86 94.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -434.92 94.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -582.45 94.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 2.86 96.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 -582.45 96.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 2.86 97.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 -582.45 97.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 2.86 99.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -582.45 99.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 2.86 101 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -582.45 101 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 2.86 102.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 -503.82 102.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 2.86 104.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -502.76 104.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -582.45 104.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 2.86 105.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 -582.45 105.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 2.86 107.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 -582.45 107.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 2.86 109 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -582.45 109 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 2.86 110.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -582.45 110.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 2.86 112.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 -582.45 112.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 2.86 113.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -424.32 113.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -497.46 113.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 2.86 115.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -424.32 115.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -582.45 115.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 2.86 117 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 -582.45 117 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 2.86 118.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -582.45 118.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 2.86 120.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -582.45 120.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 2.86 121.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 -582.45 121.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 2.86 123.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 -582.45 123.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 2.86 125 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 -582.45 125 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 2.86 126.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 -582.45 126.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 2.86 128.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -582.45 128.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 2.86 129.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -582.45 129.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 2.86 131.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 -582.45 131.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 2.86 133 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -424.32 133 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -497.46 133 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 2.86 134.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -434.92 134.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -582.45 134.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 2.86 136.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 -582.45 136.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 2.86 137.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 -582.45 137.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 2.86 139.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -582.45 139.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 2.86 141 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -582.45 141 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 2.86 142.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 -503.82 142.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 2.86 144.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -502.76 144.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -582.45 144.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 2.86 145.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 -582.45 145.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 2.86 147.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 -582.45 147.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 2.86 149 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -582.45 149 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 2.86 150.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -582.45 150.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 2.86 152.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 -582.45 152.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 2.86 153.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -424.32 153.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -497.46 153.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 2.86 155.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -424.32 155.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -582.45 155.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 2.86 157 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 -582.45 157 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 2.86 158.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -582.45 158.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 2.86 160.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -582.45 160.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 2.86 161.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 -582.45 161.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 2.86 163.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 -582.45 163.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 2.86 165 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 -582.45 165 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 2.86 166.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 -582.45 166.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 2.86 168.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -582.45 168.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 2.86 169.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -582.45 169.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 2.86 171.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 -582.45 171.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 2.86 173 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -424.32 173 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -497.46 173 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 2.86 174.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -434.92 174.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -582.45 174.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 2.86 176.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 -582.45 176.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 2.86 177.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 -582.45 177.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 2.86 179.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 -582.45 179.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 2.86 181 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 -582.45 181 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 2.86 182.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 -503.82 182.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 2.86 184.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 -502.76 184.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 2.86 185.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 -582.45 185.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 2.86 187.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 -582.45 187.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 2.86 189 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 -582.45 189 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 2.86 190.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 -582.45 190.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 2.86 192.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 -582.45 192.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 2.86 193.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -424.32 193.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -497.46 193.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 2.86 195.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -424.32 195.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -582.45 195.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 2.86 197 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 -440.22 197 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 -582.45 197 -521.2 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 2.86 198.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 -582.45 198.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 2.86 200.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 -582.45 200.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 2.86 201.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 -582.45 201.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 2.86 203.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 -582.45 203.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 2.86 205 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 -582.45 205 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 2.86 206.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 -582.45 206.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 2.86 208.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 -582.45 208.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 2.86 209.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 -582.45 209.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 2.86 211.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 -582.45 211.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 2.86 213 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 -424.32 213 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 -497.46 213 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 2.86 214.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 -434.92 214.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 -582.45 214.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 2.86 216.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 -582.45 216.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 2.86 217.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 -582.45 217.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 2.86 219.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 -582.45 219.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 2.86 221 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 -582.45 221 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 2.86 222.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 -503.82 222.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 2.86 224.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 -502.76 224.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 -582.45 224.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 2.86 225.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 -582.45 225.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 2.86 227.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 -582.45 227.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 2.86 229 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 -582.45 229 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 2.86 230.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 -582.45 230.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 2.86 232.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 -582.45 232.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 2.86 233.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -424.32 233.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -497.46 233.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 2.86 235.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 -424.32 235.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 -582.45 235.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 2.86 237 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 -582.45 237 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 2.86 238.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 -582.45 238.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 2.86 240.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 -582.45 240.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 2.86 241.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 -582.45 241.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 2.86 243.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 -582.45 243.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 2.86 245 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 -582.45 245 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 2.86 246.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 -582.45 246.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 2.86 248.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 -582.45 248.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 2.86 249.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -582.45 249.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 2.86 251.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 -582.45 251.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 2.86 253 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 -424.32 253 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 -497.46 253 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 2.86 254.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 -434.92 254.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 -582.45 254.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 2.86 256.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 -582.45 256.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 2.86 257.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 -582.45 257.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 2.86 259.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 -582.45 259.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 2.86 261 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 -582.45 261 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 2.86 262.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 -503.82 262.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 2.86 264.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 -502.76 264.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 -582.45 264.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 2.86 265.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 -582.45 265.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 2.86 267.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 -582.45 267.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 2.86 269 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 -582.45 269 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 2.86 270.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 -582.45 270.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 2.86 272.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 -582.45 272.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 2.86 273.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -424.32 273.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -497.46 273.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 2.86 275.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 -424.32 275.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 -582.45 275.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 2.86 277 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 -582.45 277 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 2.86 278.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 -582.45 278.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 2.86 280.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 -582.45 280.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 2.86 281.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 -582.45 281.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 2.86 283.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 -582.45 283.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 2.86 285 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 -582.45 285 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 2.86 286.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 -582.45 286.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 2.86 288.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 -582.45 288.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 2.86 289.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 -582.45 289.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 2.86 291.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 -582.45 291.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 2.86 293 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 -424.32 293 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 -497.46 293 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 2.86 294.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 -434.92 294.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 -582.45 294.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 2.86 296.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 -582.45 296.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 2.86 297.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 -582.45 297.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 2.86 299.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 -582.45 299.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 2.86 301 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 -582.45 301 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 2.86 302.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 -503.82 302.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 2.86 304.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 -502.76 304.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 -582.45 304.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 2.86 305.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 -582.45 305.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 2.86 307.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 -582.45 307.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 2.86 309 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 -582.45 309 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 2.86 310.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 -582.45 310.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 2.86 312.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 -582.45 312.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 2.86 313.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -424.32 313.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -497.46 313.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 2.86 315.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 -424.32 315.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 -582.45 315.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 2.86 317 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 -582.45 317 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 2.86 318.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 -582.45 318.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 2.86 320.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 -582.45 320.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 2.86 321.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 -582.45 321.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 2.86 323.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 -582.45 323.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 2.86 325 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 -582.45 325 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 2.86 326.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 -582.45 326.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 2.86 328.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 -582.45 328.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 2.86 329.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 -582.45 329.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 331 2.86 331.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 331 -582.45 331.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 2.86 333 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 -424.32 333 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 -497.46 333 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 2.86 334.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 -434.92 334.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 -582.45 334.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.8 2.86 336.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.8 -582.45 336.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.4 2.86 337.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.4 -582.45 337.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 339 2.86 339.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 339 -582.45 339.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.6 2.86 341 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.6 -582.45 341 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.2 2.86 342.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.2 -503.82 342.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.8 2.86 344.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.8 -502.76 344.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.4 2.86 345.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.4 -582.45 345.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 347 2.86 347.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 347 -582.45 347.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.6 2.86 349 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.6 -582.45 349 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.2 2.86 350.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.2 -582.45 350.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.8 2.86 352.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.8 -582.45 352.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 2.86 353.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 -424.32 353.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 -497.46 353.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 2.86 355.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 -424.32 355.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 -582.45 355.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 2.86 357 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 -440.22 357 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 -582.45 357 -521.2 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.2 2.86 358.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.2 -582.45 358.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.8 2.86 360.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.8 -582.45 360.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.4 2.86 361.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.4 -582.45 361.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 363 2.86 363.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 363 -582.45 363.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.6 2.86 365 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.6 -582.45 365 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.2 2.86 366.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.2 -582.45 366.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.8 2.86 368.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.8 -582.45 368.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.4 2.86 369.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.4 -582.45 369.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 371 2.86 371.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 371 -582.45 371.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 2.86 373 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 -424.32 373 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 -497.46 373 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 2.86 374.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 -434.92 374.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 -582.45 374.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.8 2.86 376.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.8 -582.45 376.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.4 2.86 377.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.4 -582.45 377.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 379 2.86 379.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 379 -582.45 379.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.6 2.86 381 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.6 -582.45 381 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.2 2.86 382.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.2 -503.82 382.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 2.86 384.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 -502.76 384.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 -582.45 384.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.4 2.86 385.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.4 -582.45 385.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 387 2.86 387.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 387 -582.45 387.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.6 2.86 389 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.6 -582.45 389 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.2 2.86 390.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.2 -582.45 390.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.8 2.86 392.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.8 -582.45 392.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 2.86 393.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 -424.32 393.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 -497.46 393.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 2.86 395.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 -424.32 395.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 -582.45 395.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.6 2.86 397 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.6 -582.45 397 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.2 2.86 398.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.2 -582.45 398.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.8 2.86 400.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.8 -582.45 400.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.4 2.86 401.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.4 -582.45 401.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 403 2.86 403.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 403 -582.45 403.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.6 2.86 405 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.6 -582.45 405 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.2 2.86 406.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.2 -582.45 406.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.8 2.86 408.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.8 -582.45 408.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.4 2.86 409.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.4 -582.45 409.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 411 2.86 411.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 411 -582.45 411.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 2.86 413 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 -424.32 413 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 -497.46 413 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 2.86 414.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 -434.92 414.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 -582.45 414.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.8 2.86 416.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.8 -582.45 416.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.4 2.86 417.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.4 -582.45 417.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 419 2.86 419.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 419 -582.45 419.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.6 2.86 421 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.6 -582.45 421 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.2 2.86 422.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.2 -503.82 422.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 2.86 424.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 -502.76 424.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 -582.45 424.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.4 2.86 425.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.4 -582.45 425.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 427 2.86 427.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 427 -582.45 427.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.6 2.86 429 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.6 -582.45 429 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.2 2.86 430.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.2 -582.45 430.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.8 2.86 432.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.8 -582.45 432.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 2.86 433.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 -424.32 433.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 -497.46 433.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 2.86 435.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 -424.32 435.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 -582.45 435.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.6 2.86 437 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.6 -582.45 437 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.2 2.86 438.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.2 -582.45 438.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.8 2.86 440.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.8 -582.45 440.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.4 2.86 441.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.4 -582.45 441.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 443 2.86 443.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 443 -582.45 443.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.6 2.86 445 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.6 -582.45 445 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.2 2.86 446.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.2 -582.45 446.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.8 2.86 448.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.8 -582.45 448.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.4 2.86 449.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.4 -582.45 449.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 451 2.86 451.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 451 -582.45 451.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 2.86 453 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 -424.32 453 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 -497.46 453 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 2.86 454.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 -434.92 454.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 -582.45 454.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.8 2.86 456.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.8 -582.45 456.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.4 2.86 457.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.4 -582.45 457.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 459 2.86 459.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 459 -582.45 459.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.6 2.86 461 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.6 -582.45 461 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.2 2.86 462.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.2 -503.82 462.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 2.86 464.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 -502.76 464.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 -582.45 464.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.4 2.86 465.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.4 -582.45 465.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 467 2.86 467.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 467 -582.45 467.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.6 2.86 469 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.6 -582.45 469 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.2 2.86 470.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.2 -582.45 470.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.8 2.86 472.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.8 -582.45 472.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 2.86 473.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 -424.32 473.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 -497.46 473.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 2.86 475.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 -424.32 475.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 -582.45 475.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.6 2.86 477 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.6 -582.45 477 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.2 2.86 478.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.2 -582.45 478.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.8 2.86 480.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.8 -582.45 480.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.4 2.86 481.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.4 -582.45 481.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 483 2.86 483.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 483 -582.45 483.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.6 2.86 485 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.6 -582.45 485 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.2 2.86 486.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.2 -582.45 486.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.8 2.86 488.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.8 -582.45 488.2 -414.14 ;
        RECT 487.75 -500.595 488.2 -500.265 ;
        RECT 487.75 -514.735 488.2 -514.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.4 2.86 489.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.4 -582.45 489.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 491 2.86 491.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 491 -582.45 491.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 2.86 493 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 -424.32 493 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 -497.46 493 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 2.86 494.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 -434.92 494.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 -582.45 494.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.8 2.86 496.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.8 -582.45 496.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.4 2.86 497.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.4 -582.45 497.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 499 2.86 499.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 499 -582.45 499.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.6 2.86 501 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.6 -582.45 501 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.2 2.86 502.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.2 -503.82 502.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.8 2.86 504.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.8 -502.76 504.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.4 2.86 505.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.4 -582.45 505.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 507 2.86 507.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 507 -582.45 507.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.6 2.86 509 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.6 -582.45 509 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.2 2.86 510.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.2 -582.45 510.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.8 2.86 512.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.8 -582.45 512.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 2.86 513.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 -424.32 513.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 -497.46 513.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 2.86 515.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 -424.32 515.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 -582.45 515.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 2.86 517 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 -440.22 517 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 -582.45 517 -521.2 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.2 2.86 518.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.2 -582.45 518.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.8 2.86 520.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.8 -582.45 520.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.4 2.86 521.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.4 -582.45 521.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 523 2.86 523.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 523 -582.45 523.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.6 2.86 525 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.6 -582.45 525 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.2 2.86 526.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.2 -582.45 526.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.8 2.86 528.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.8 -582.45 528.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.4 2.86 529.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.4 -582.45 529.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 531 2.86 531.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 531 -582.45 531.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 2.86 533 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 -424.32 533 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 -497.46 533 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 2.86 534.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 -434.92 534.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 -582.45 534.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.8 2.86 536.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.8 -582.45 536.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.4 2.86 537.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.4 -582.45 537.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 539 2.86 539.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 539 -582.45 539.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.6 2.86 541 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.6 -582.45 541 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.2 2.86 542.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.2 -503.82 542.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 2.86 544.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 -502.76 544.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 -582.45 544.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.4 2.86 545.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.4 -582.45 545.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 547 2.86 547.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 547 -582.45 547.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.6 2.86 549 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.6 -582.45 549 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.2 2.86 550.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.2 -582.45 550.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.8 2.86 552.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.8 -582.45 552.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 2.86 553.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 -424.32 553.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 -497.46 553.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 2.86 555.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 -424.32 555.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 -582.45 555.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.6 2.86 557 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.6 -582.45 557 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.2 2.86 558.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.2 -582.45 558.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.8 2.86 560.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.8 -582.45 560.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.4 2.86 561.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.4 -582.45 561.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 563 2.86 563.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 563 -582.45 563.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.6 2.86 565 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.6 -582.45 565 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.2 2.86 566.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.2 -582.45 566.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.8 2.86 568.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.8 -582.45 568.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.4 2.86 569.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.4 -582.45 569.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 571 2.86 571.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 571 -582.45 571.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 2.86 573 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 -424.32 573 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 -497.46 573 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 2.86 574.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 -434.92 574.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 -582.45 574.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.8 2.86 576.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.8 -582.45 576.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.4 2.86 577.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.4 -582.45 577.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 579 2.86 579.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 579 -582.45 579.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.6 2.86 581 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.6 -582.45 581 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.2 2.86 582.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.2 -503.82 582.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 2.86 584.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 -502.76 584.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 -582.45 584.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.4 2.86 585.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.4 -582.45 585.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 587 2.86 587.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 587 -582.45 587.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.6 2.86 589 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.6 -582.45 589 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.2 2.86 590.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.2 -582.45 590.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.8 2.86 592.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.8 -582.45 592.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 2.86 593.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 -424.32 593.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 -497.46 593.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 2.86 595.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 -424.32 595.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 -582.45 595.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.6 2.86 597 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.6 -582.45 597 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.2 2.86 598.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.2 -582.45 598.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.8 2.86 600.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.8 -582.45 600.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.4 2.86 601.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.4 -582.45 601.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 603 2.86 603.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 603 -582.45 603.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.6 2.86 605 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.6 -582.45 605 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.2 2.86 606.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.2 -582.45 606.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.8 2.86 608.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.8 -582.45 608.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.4 2.86 609.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.4 -582.45 609.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 611 2.86 611.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 611 -582.45 611.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 2.86 613 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 -424.32 613 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 -497.46 613 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 2.86 614.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 -434.92 614.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 -582.45 614.6 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.8 2.86 616.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.8 -582.45 616.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.4 2.86 617.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.4 -582.45 617.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 619 2.86 619.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 619 -582.45 619.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.6 2.86 621 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.6 -582.45 621 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.2 2.86 622.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.2 -503.82 622.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 2.86 624.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 -502.76 624.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 -582.45 624.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.4 2.86 625.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.4 -582.45 625.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 627 2.86 627.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 627 -582.45 627.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.6 2.86 629 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.6 -582.45 629 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.2 2.86 630.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.2 -582.45 630.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.8 2.86 632.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.8 -582.45 632.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 2.86 633.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 -424.32 633.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 -497.46 633.8 -488.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 2.86 635.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 -424.32 635.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 -582.45 635.4 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.6 2.86 637 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.6 -582.45 637 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.2 2.86 638.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.2 -582.45 638.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.8 2.86 640.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.8 -582.45 640.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.4 2.86 641.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.4 -582.45 641.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 643 2.86 643.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 643 -582.45 643.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.6 2.86 645 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.6 -582.45 645 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.2 2.86 646.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.2 -582.45 646.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.8 2.86 648.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.8 -582.45 648.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.4 2.86 649.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.4 -582.45 649.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 651 -582.45 651.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 652.6 -582.45 653 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 654.2 -582.45 654.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 655.8 -582.45 656.2 11.315 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -81 -580.91 -80.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.4 -580.91 -79 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -77.8 -580.91 -77.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -76.2 -551.52 -75.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.6 -569.54 -74.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -73 -580.91 -72.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.4 -564.24 -71 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.4 -580.91 -71 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.8 -565.3 -69.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.8 -580.91 -69.4 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -569.54 -67.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -580.91 -67.8 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.6 -580.91 -66.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -563.18 -64.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -580.91 -64.6 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.4 -569.54 -63 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -569.54 -61.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -580.91 -61.4 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.2 -580.91 -59.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -562.12 -58.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -580.91 -58.2 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -57 -569.54 -56.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.4 -580.91 -55 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -561.06 -53.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -580.91 -53.4 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.2 -562.12 -51.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -569.54 -50.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -580.91 -50.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -49 -580.91 -48.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -560 -47 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -580.91 -47 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.8 -569.54 -45.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -569.54 -43.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -580.91 -43.8 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.6 -580.91 -42.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -558.94 -40.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -580.91 -40.6 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.4 -569.54 -39 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.8 -580.91 -37.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -557.88 -35.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -580.91 -35.8 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.6 -558.94 -34.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -569.54 -32.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -580.91 -32.6 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.4 -580.91 -31 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -557.88 -29.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -580.91 -29.4 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.2 -569.54 -27.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -569.54 -26.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -580.91 -26.2 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -25 -580.91 -24.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -556.82 -23 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -580.91 -23 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.8 -569.54 -21.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.2 -580.91 -19.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -555.76 -18.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -580.91 -18.2 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -17 -555.76 -16.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -569.54 -15 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -580.91 -15 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.8 -580.91 -13.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -554.7 -11.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -580.91 -11.8 -572.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -413.72 -10.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -569.54 -10.2 -533.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -569.54 -8.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -580.91 -8.6 -575.26 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.4 -580.91 -7 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -550.46 -5.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -580.91 -5.4 -572.08 ;
        RECT -5.805 -573.905 -5.4 -573.575 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.2 -580.91 -3.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.6 -580.91 -2.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 2.86 -0.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 -580.91 -0.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 2.86 1 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 -580.91 1 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 2.86 2.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 -580.91 2.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 2.86 4.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 -580.91 4.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 2.86 5.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -580.91 5.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 2.86 7.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 -580.91 7.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 2.86 9 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -580.91 9 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 2.86 10.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -580.91 10.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 2.86 12.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 -580.91 12.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 2.86 13.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -424.32 13.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -497.46 13.8 -488.34 ;
        RECT 13.435 -497.46 13.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 2.86 15.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -424.32 15.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -580.91 15.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 2.86 17 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 -580.91 17 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 2.86 18.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -580.91 18.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 2.86 20.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -580.91 20.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 2.86 21.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -503.82 21.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 2.86 23.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 -502.76 23.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 2.86 25 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 -519.72 25 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 2.86 26.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 -580.91 26.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 2.86 28.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -580.91 28.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 2.86 29.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -580.91 29.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 2.86 31.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 -580.91 31.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 2.86 33 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -424.32 33 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -497.46 33 -488.34 ;
        RECT 32.635 -497.46 32.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 2.86 34.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -434.92 34.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -580.91 34.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 2.86 36.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -440.22 36.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -580.91 36.2 -521.2 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 2.86 37.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 -580.91 37.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 2.86 39.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -580.91 39.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 2.86 41 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -580.91 41 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 2.86 42.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 -580.91 42.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 2.86 44.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 -580.91 44.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 2.86 45.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 -580.91 45.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 2.86 47.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 -580.91 47.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 2.86 49 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -580.91 49 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 2.86 50.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -580.91 50.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 2.86 52.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 -580.91 52.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 2.86 53.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -424.32 53.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -497.46 53.8 -488.34 ;
        RECT 53.435 -497.46 53.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 2.86 55.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -424.32 55.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -580.91 55.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 2.86 57 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 -580.91 57 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 2.86 58.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -580.91 58.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 2.86 60.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -580.91 60.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 2.86 61.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 -503.82 61.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 2.86 63.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 -502.76 63.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 2.86 65 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 -580.91 65 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 2.86 66.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 -580.91 66.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 2.86 68.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -580.91 68.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 2.86 69.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -580.91 69.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 2.86 71.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 -580.91 71.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 2.86 73 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -424.32 73 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -497.46 73 -488.34 ;
        RECT 72.635 -497.46 72.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 2.86 74.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -434.92 74.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -580.91 74.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 2.86 76.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 -580.91 76.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 2.86 77.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 -580.91 77.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 2.86 79.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -580.91 79.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 2.86 81 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -580.91 81 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 2.86 82.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 -580.91 82.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 2.86 84.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 -580.91 84.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 2.86 85.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 -580.91 85.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 2.86 87.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 -580.91 87.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 2.86 89 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -580.91 89 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 2.86 90.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -580.91 90.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 2.86 92.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 -580.91 92.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 2.86 93.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -424.32 93.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -497.46 93.8 -488.34 ;
        RECT 93.435 -497.46 93.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 2.86 95.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -424.32 95.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -580.91 95.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 2.86 97 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 -580.91 97 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 2.86 98.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -580.91 98.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 2.86 100.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -580.91 100.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 2.86 101.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -503.82 101.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 2.86 103.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 -502.76 103.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 2.86 105 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 -580.91 105 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 2.86 106.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 -580.91 106.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 2.86 108.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -580.91 108.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 2.86 109.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -580.91 109.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 2.86 111.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 -580.91 111.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 2.86 113 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -424.32 113 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -497.46 113 -488.34 ;
        RECT 112.635 -497.46 112.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 2.86 114.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -434.92 114.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -580.91 114.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 2.86 116.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 -580.91 116.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 2.86 117.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 -580.91 117.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 2.86 119.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -580.91 119.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 2.86 121 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -580.91 121 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 2.86 122.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 -580.91 122.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 2.86 124.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 -580.91 124.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 2.86 125.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 -580.91 125.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 2.86 127.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 -580.91 127.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 2.86 129 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -580.91 129 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 2.86 130.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -580.91 130.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 2.86 132.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 -580.91 132.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 2.86 133.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -424.32 133.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -497.46 133.8 -488.34 ;
        RECT 133.435 -497.46 133.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 2.86 135.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -424.32 135.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -580.91 135.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 2.86 137 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 -580.91 137 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 2.86 138.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -580.91 138.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 2.86 140.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -580.91 140.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 2.86 141.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 -503.82 141.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 2.86 143.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 -502.76 143.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 2.86 145 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 -580.91 145 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 2.86 146.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 -580.91 146.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 2.86 148.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -580.91 148.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 2.86 149.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -580.91 149.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 2.86 151.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 -580.91 151.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 2.86 153 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -424.32 153 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -497.46 153 -488.34 ;
        RECT 152.635 -497.46 152.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 2.86 154.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -434.92 154.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -580.91 154.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 2.86 156.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 -580.91 156.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 2.86 157.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 -580.91 157.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 2.86 159.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -580.91 159.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 2.86 161 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -580.91 161 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 2.86 162.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 -580.91 162.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 2.86 164.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 -580.91 164.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 2.86 165.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 -580.91 165.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 2.86 167.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 -580.91 167.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 2.86 169 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -580.91 169 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 2.86 170.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -580.91 170.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 2.86 172.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 -580.91 172.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 2.86 173.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -424.32 173.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -497.46 173.8 -488.34 ;
        RECT 173.435 -497.46 173.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 2.86 175.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -424.32 175.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -580.91 175.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 2.86 177 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 -580.91 177 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 2.86 178.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 -580.91 178.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 2.86 180.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 -580.91 180.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 2.86 181.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 -503.82 181.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 2.86 183.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 -502.76 183.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 2.86 185 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 -519.72 185 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 2.86 186.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 -580.91 186.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 2.86 188.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 -580.91 188.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 2.86 189.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 -580.91 189.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 2.86 191.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 -580.91 191.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 2.86 193 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 -424.32 193 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 -497.46 193 -488.34 ;
        RECT 192.635 -497.46 192.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 2.86 194.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 -434.92 194.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 -580.91 194.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 2.86 196.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 -440.22 196.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 -580.91 196.2 -521.2 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 2.86 197.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 -580.91 197.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 2.86 199.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 -580.91 199.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 2.86 201 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 -580.91 201 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 2.86 202.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 -580.91 202.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 2.86 204.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 -580.91 204.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 2.86 205.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 -580.91 205.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 2.86 207.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 -580.91 207.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 2.86 209 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 -580.91 209 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 2.86 210.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 -580.91 210.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 2.86 212.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 -580.91 212.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 2.86 213.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -424.32 213.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -497.46 213.8 -488.34 ;
        RECT 213.435 -497.46 213.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 2.86 215.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 -424.32 215.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 -580.91 215.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 2.86 217 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 -580.91 217 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 2.86 218.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 -580.91 218.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 2.86 220.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 -580.91 220.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 2.86 221.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 -503.82 221.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 2.86 223.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 -502.76 223.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 2.86 225 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 -580.91 225 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 2.86 226.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 -580.91 226.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 2.86 228.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 -580.91 228.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 2.86 229.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 -580.91 229.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 2.86 231.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 -580.91 231.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 2.86 233 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 -424.32 233 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 -497.46 233 -488.34 ;
        RECT 232.635 -497.46 232.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 2.86 234.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 -434.92 234.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 -580.91 234.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 2.86 236.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 -580.91 236.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 2.86 237.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 -580.91 237.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 2.86 239.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 -580.91 239.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 2.86 241 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 -580.91 241 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 2.86 242.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 -580.91 242.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 2.86 244.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 -580.91 244.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 2.86 245.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 -580.91 245.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 2.86 247.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 -580.91 247.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 2.86 249 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 -580.91 249 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 2.86 250.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 -580.91 250.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 2.86 252.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 -580.91 252.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 2.86 253.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -424.32 253.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -497.46 253.8 -488.34 ;
        RECT 253.435 -497.46 253.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 2.86 255.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 -424.32 255.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 -580.91 255.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 2.86 257 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 -580.91 257 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 2.86 258.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 -580.91 258.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 2.86 260.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 -580.91 260.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 2.86 261.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 -503.82 261.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 2.86 263.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 -502.76 263.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 2.86 265 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 -580.91 265 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 2.86 266.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 -580.91 266.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 2.86 268.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 -580.91 268.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 2.86 269.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 -580.91 269.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 2.86 271.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 -580.91 271.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 2.86 273 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 -424.32 273 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 -497.46 273 -488.34 ;
        RECT 272.635 -497.46 272.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 2.86 274.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 -434.92 274.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 -580.91 274.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 2.86 276.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 -580.91 276.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 2.86 277.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 -580.91 277.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 2.86 279.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 -580.91 279.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 2.86 281 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 -580.91 281 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 2.86 282.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 -580.91 282.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 2.86 284.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 -580.91 284.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 2.86 285.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 -580.91 285.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 2.86 287.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 -580.91 287.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 2.86 289 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 -580.91 289 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 2.86 290.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -580.91 290.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 2.86 292.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 -580.91 292.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 2.86 293.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -424.32 293.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -497.46 293.8 -488.34 ;
        RECT 293.435 -497.46 293.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 2.86 295.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 -424.32 295.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 -580.91 295.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 2.86 297 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 -580.91 297 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 2.86 298.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 -580.91 298.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 2.86 300.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 -580.91 300.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 2.86 301.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 -503.82 301.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 2.86 303.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 -502.76 303.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 2.86 305 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 -580.91 305 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 2.86 306.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 -580.91 306.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 2.86 308.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 -580.91 308.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 2.86 309.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 -580.91 309.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 2.86 311.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 -580.91 311.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 2.86 313 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 -424.32 313 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 -497.46 313 -488.34 ;
        RECT 312.635 -497.46 312.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 2.86 314.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 -434.92 314.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 -580.91 314.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 2.86 316.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 -580.91 316.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 2.86 317.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 -580.91 317.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 2.86 319.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 -580.91 319.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 2.86 321 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 -580.91 321 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 2.86 322.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 -580.91 322.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 2.86 324.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 -580.91 324.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 2.86 325.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 -580.91 325.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 2.86 327.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 -580.91 327.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 2.86 329 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 -580.91 329 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 2.86 330.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 -580.91 330.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.8 2.86 332.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.8 -580.91 332.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 2.86 333.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 -424.32 333.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 -497.46 333.8 -488.34 ;
        RECT 333.435 -497.46 333.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 2.86 335.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 -424.32 335.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 -580.91 335.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.6 2.86 337 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.6 -580.91 337 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.2 2.86 338.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.2 -580.91 338.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.8 2.86 340.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.8 -580.91 340.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.4 2.86 341.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.4 -503.82 341.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 343 2.86 343.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 343 -502.76 343.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.6 2.86 345 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.6 -519.72 345 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.2 2.86 346.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.2 -580.91 346.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.8 2.86 348.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.8 -580.91 348.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.4 2.86 349.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.4 -580.91 349.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 351 2.86 351.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 351 -580.91 351.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 2.86 353 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 -424.32 353 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 -497.46 353 -488.34 ;
        RECT 352.635 -497.46 352.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 2.86 354.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 -434.92 354.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 -580.91 354.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 2.86 356.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 -440.22 356.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 -580.91 356.2 -521.2 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.4 2.86 357.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.4 -580.91 357.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 359 2.86 359.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 359 -580.91 359.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.6 2.86 361 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.6 -580.91 361 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.2 2.86 362.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.2 -580.91 362.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.8 2.86 364.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.8 -580.91 364.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.4 2.86 365.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.4 -580.91 365.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 367 2.86 367.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 367 -580.91 367.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.6 2.86 369 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.6 -580.91 369 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.2 2.86 370.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.2 -580.91 370.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.8 2.86 372.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.8 -580.91 372.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 2.86 373.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 -424.32 373.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 -497.46 373.8 -488.34 ;
        RECT 373.435 -497.46 373.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 2.86 375.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 -424.32 375.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 -580.91 375.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.6 2.86 377 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.6 -580.91 377 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.2 2.86 378.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.2 -580.91 378.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.8 2.86 380.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.8 -580.91 380.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.4 2.86 381.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.4 -503.82 381.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 383 2.86 383.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 383 -502.76 383.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.6 2.86 385 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.6 -580.91 385 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.2 2.86 386.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.2 -580.91 386.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.8 2.86 388.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.8 -580.91 388.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.4 2.86 389.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.4 -580.91 389.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 391 2.86 391.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 391 -580.91 391.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 2.86 393 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 -424.32 393 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 -497.46 393 -488.34 ;
        RECT 392.635 -497.46 392.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 2.86 394.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 -434.92 394.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 -580.91 394.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.8 2.86 396.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.8 -580.91 396.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.4 2.86 397.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.4 -580.91 397.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 399 2.86 399.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 399 -580.91 399.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.6 2.86 401 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.6 -580.91 401 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.2 2.86 402.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.2 -580.91 402.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.8 2.86 404.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.8 -580.91 404.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.4 2.86 405.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.4 -580.91 405.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 407 2.86 407.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 407 -580.91 407.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.6 2.86 409 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.6 -580.91 409 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.2 2.86 410.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.2 -580.91 410.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.8 2.86 412.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.8 -580.91 412.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 2.86 413.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 -424.32 413.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 -497.46 413.8 -488.34 ;
        RECT 413.435 -497.46 413.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 2.86 415.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 -424.32 415.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 -580.91 415.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.6 2.86 417 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.6 -580.91 417 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.2 2.86 418.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.2 -580.91 418.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.8 2.86 420.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.8 -580.91 420.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.4 2.86 421.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.4 -503.82 421.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 423 2.86 423.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 423 -502.76 423.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.6 2.86 425 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.6 -580.91 425 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.2 2.86 426.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.2 -580.91 426.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.8 2.86 428.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.8 -580.91 428.2 -414.14 ;
        RECT 427.75 -523.605 428.2 -523.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.4 2.86 429.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.4 -580.91 429.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 431 2.86 431.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 431 -580.91 431.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 2.86 433 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 -424.32 433 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 -497.46 433 -488.34 ;
        RECT 432.635 -497.46 432.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 2.86 434.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 -434.92 434.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 -580.91 434.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.8 2.86 436.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.8 -580.91 436.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.4 2.86 437.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.4 -580.91 437.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 439 2.86 439.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 439 -580.91 439.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.6 2.86 441 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.6 -580.91 441 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.2 2.86 442.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.2 -580.91 442.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.8 2.86 444.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.8 -580.91 444.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.4 2.86 445.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.4 -580.91 445.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 447 2.86 447.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 447 -580.91 447.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.6 2.86 449 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.6 -580.91 449 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.2 2.86 450.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.2 -580.91 450.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.8 2.86 452.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.8 -580.91 452.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 2.86 453.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 -424.32 453.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 -497.46 453.8 -488.34 ;
        RECT 453.435 -497.46 453.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 2.86 455.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 -424.32 455.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 -580.91 455.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.6 2.86 457 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.6 -580.91 457 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.2 2.86 458.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.2 -580.91 458.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.8 2.86 460.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.8 -580.91 460.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.4 2.86 461.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.4 -503.82 461.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 463 2.86 463.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 463 -502.76 463.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.6 2.86 465 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.6 -580.91 465 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.2 2.86 466.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.2 -580.91 466.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.8 2.86 468.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.8 -580.91 468.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.4 2.86 469.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.4 -580.91 469.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 471 2.86 471.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 471 -580.91 471.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 2.86 473 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 -424.32 473 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 -497.46 473 -488.34 ;
        RECT 472.635 -497.46 472.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 2.86 474.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 -434.92 474.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 -580.91 474.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.8 2.86 476.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.8 -580.91 476.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.4 2.86 477.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.4 -580.91 477.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 479 2.86 479.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 479 -580.91 479.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.6 2.86 481 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.6 -580.91 481 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.2 2.86 482.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.2 -580.91 482.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.8 2.86 484.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.8 -580.91 484.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.4 2.86 485.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.4 -580.91 485.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 487 2.86 487.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 487 -580.91 487.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.6 2.86 489 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.6 -580.91 489 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.2 2.86 490.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.2 -580.91 490.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.8 2.86 492.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.8 -580.91 492.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 2.86 493.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 -424.32 493.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 -497.46 493.8 -488.34 ;
        RECT 493.435 -497.46 493.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 2.86 495.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 -424.32 495.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 -580.91 495.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.6 2.86 497 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.6 -580.91 497 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.2 2.86 498.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.2 -580.91 498.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.8 2.86 500.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.8 -580.91 500.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.4 2.86 501.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.4 -503.82 501.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 503 2.86 503.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 503 -502.76 503.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.6 2.86 505 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.6 -519.72 505 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.2 2.86 506.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.2 -580.91 506.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.8 2.86 508.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.8 -580.91 508.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.4 2.86 509.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.4 -580.91 509.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 511 2.86 511.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 511 -580.91 511.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 2.86 513 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 -424.32 513 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 -497.46 513 -488.34 ;
        RECT 512.635 -497.46 512.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 2.86 514.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 -434.92 514.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 -580.91 514.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 2.86 516.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 -440.22 516.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 -580.91 516.2 -521.2 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.4 2.86 517.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.4 -580.91 517.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 519 2.86 519.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 519 -580.91 519.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.6 2.86 521 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.6 -580.91 521 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.2 2.86 522.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.2 -580.91 522.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.8 2.86 524.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.8 -580.91 524.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.4 2.86 525.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.4 -580.91 525.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 527 2.86 527.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 527 -580.91 527.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.6 2.86 529 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.6 -580.91 529 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.2 2.86 530.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.2 -580.91 530.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.8 2.86 532.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.8 -580.91 532.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 2.86 533.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 -424.32 533.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 -497.46 533.8 -488.34 ;
        RECT 533.435 -497.46 533.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 2.86 535.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 -424.32 535.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 -580.91 535.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.6 2.86 537 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.6 -580.91 537 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.2 2.86 538.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.2 -580.91 538.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.8 2.86 540.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.8 -580.91 540.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.4 2.86 541.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.4 -503.82 541.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 543 2.86 543.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 543 -502.76 543.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.6 2.86 545 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.6 -580.91 545 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.2 2.86 546.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.2 -580.91 546.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.8 2.86 548.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.8 -580.91 548.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.4 2.86 549.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.4 -580.91 549.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 551 2.86 551.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 551 -580.91 551.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 2.86 553 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 -424.32 553 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 -497.46 553 -488.34 ;
        RECT 552.635 -497.46 552.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 2.86 554.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 -434.92 554.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 -580.91 554.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.8 2.86 556.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.8 -580.91 556.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 557.4 2.86 557.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 557.4 -580.91 557.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 559 2.86 559.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 559 -580.91 559.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.6 2.86 561 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.6 -580.91 561 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 2.86 562.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 -580.91 562.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.8 2.86 564.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.8 -580.91 564.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.4 2.86 565.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.4 -580.91 565.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 567 2.86 567.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 567 -580.91 567.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.6 2.86 569 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.6 -580.91 569 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.2 2.86 570.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.2 -580.91 570.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.8 2.86 572.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.8 -580.91 572.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 2.86 573.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 -424.32 573.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 -497.46 573.8 -488.34 ;
        RECT 573.435 -497.46 573.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 2.86 575.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 -424.32 575.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 -580.91 575.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.6 2.86 577 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.6 -580.91 577 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.2 2.86 578.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.2 -580.91 578.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.8 2.86 580.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.8 -580.91 580.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.4 2.86 581.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.4 -503.82 581.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 583 2.86 583.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 583 -502.76 583.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.6 2.86 585 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.6 -580.91 585 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.2 2.86 586.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.2 -580.91 586.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.8 2.86 588.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.8 -580.91 588.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.4 2.86 589.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.4 -580.91 589.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 591 2.86 591.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 591 -580.91 591.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 2.86 593 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 -424.32 593 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 -497.46 593 -488.34 ;
        RECT 592.635 -497.46 592.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 2.86 594.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 -434.92 594.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 -580.91 594.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.8 2.86 596.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.8 -580.91 596.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.4 2.86 597.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.4 -580.91 597.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 599 2.86 599.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 599 -580.91 599.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.6 2.86 601 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.6 -580.91 601 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.2 2.86 602.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.2 -580.91 602.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.8 2.86 604.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.8 -580.91 604.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.4 2.86 605.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.4 -580.91 605.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 607 2.86 607.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 607 -580.91 607.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.6 2.86 609 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.6 -580.91 609 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.2 2.86 610.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.2 -580.91 610.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.8 2.86 612.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.8 -580.91 612.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 2.86 613.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 -424.32 613.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 -497.46 613.8 -488.34 ;
        RECT 613.435 -497.46 613.765 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 2.86 615.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 -424.32 615.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 -580.91 615.4 -504.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.6 2.86 617 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.6 -580.91 617 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.2 2.86 618.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.2 -580.91 618.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.8 2.86 620.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.8 -580.91 620.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.4 2.86 621.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.4 -503.82 621.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 623 2.86 623.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 623 -502.76 623.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.6 2.86 625 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.6 -580.91 625 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.2 2.86 626.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.2 -580.91 626.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.8 2.86 628.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.8 -580.91 628.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.4 2.86 629.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.4 -580.91 629.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 631 2.86 631.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 631 -580.91 631.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 2.86 633 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 -424.32 633 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 -497.46 633 -488.34 ;
        RECT 632.635 -497.46 632.965 -488.25 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 2.86 634.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 -434.92 634.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 -580.91 634.6 -512.72 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.8 2.86 636.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.8 -580.91 636.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.4 2.86 637.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.4 -580.91 637.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 639 2.86 639.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 639 -580.91 639.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.6 2.86 641 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.6 -580.91 641 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.2 2.86 642.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.2 -580.91 642.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.8 2.86 644.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.8 -580.91 644.2 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.4 2.86 645.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.4 -580.91 645.8 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 647 2.86 647.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 647 -580.91 647.4 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.6 2.86 649 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.6 -580.91 649 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.2 2.86 650.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.2 -580.91 650.6 -414.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.8 -580.91 652.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.4 -580.91 653.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 655 -580.91 655.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.6 -580.91 657 9.775 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -16.46 -582.85 -16.16 -582.55 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -74.86 -582.85 -74.56 -582.55 ;
    END
  END addr[10]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -22.3 -582.85 -22 -582.55 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.14 -582.85 -27.84 -582.55 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -33.98 -582.85 -33.68 -582.55 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -39.82 -582.85 -39.52 -582.55 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -45.66 -582.85 -45.36 -582.55 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -51.5 -582.85 -51.2 -582.55 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -57.34 -582.85 -57.04 -582.55 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -63.18 -582.85 -62.88 -582.55 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -69.02 -582.85 -68.72 -582.55 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -75.88 -582.85 -75.46 -582.43 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.015 -582.85 22.315 -582.55 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.015 -582.85 222.315 -582.55 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.63 -582.85 222.93 -582.55 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.015 -582.85 262.315 -582.55 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.63 -582.85 262.93 -582.55 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 302.015 -582.85 302.315 -582.55 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 302.63 -582.85 302.93 -582.55 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 342.015 -582.85 342.315 -582.55 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 342.63 -582.85 342.93 -582.55 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 382.015 -582.85 382.315 -582.55 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 382.63 -582.85 382.93 -582.55 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.63 -582.85 22.93 -582.55 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 422.015 -582.85 422.315 -582.55 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 422.63 -582.85 422.93 -582.55 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 462.015 -582.85 462.315 -582.55 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 462.63 -582.85 462.93 -582.55 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 502.015 -582.85 502.315 -582.55 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 502.63 -582.85 502.93 -582.55 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 542.015 -582.85 542.315 -582.55 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 542.63 -582.85 542.93 -582.55 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.015 -582.85 582.315 -582.55 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.63 -582.85 582.93 -582.55 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.015 -582.85 62.315 -582.55 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 622.015 -582.85 622.315 -582.55 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 622.63 -582.85 622.93 -582.55 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.63 -582.85 62.93 -582.55 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.015 -582.85 102.315 -582.55 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.63 -582.85 102.93 -582.55 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.015 -582.85 142.315 -582.55 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.63 -582.85 142.93 -582.55 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.015 -582.85 182.315 -582.55 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.63 -582.85 182.93 -582.55 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 13.285 -582.85 13.585 -582.55 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.285 -582.85 213.585 -582.55 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.285 -582.85 233.585 -582.55 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 253.285 -582.85 253.585 -582.55 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.285 -582.85 273.585 -582.55 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 293.285 -582.85 293.585 -582.55 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.285 -582.85 313.585 -582.55 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 333.285 -582.85 333.585 -582.55 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 353.285 -582.85 353.585 -582.55 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 373.285 -582.85 373.585 -582.55 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.285 -582.85 393.585 -582.55 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 33.285 -582.85 33.585 -582.55 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 413.285 -582.85 413.585 -582.55 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 433.285 -582.85 433.585 -582.55 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 453.285 -582.85 453.585 -582.55 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.285 -582.85 473.585 -582.55 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.285 -582.85 493.585 -582.55 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 513.285 -582.85 513.585 -582.55 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 533.285 -582.85 533.585 -582.55 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 553.285 -582.85 553.585 -582.55 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 573.285 -582.85 573.585 -582.55 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 593.285 -582.85 593.585 -582.55 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.285 -582.85 53.585 -582.55 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.285 -582.85 613.585 -582.55 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 633.285 -582.85 633.585 -582.55 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 73.285 -582.85 73.585 -582.55 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 93.285 -582.85 93.585 -582.55 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.285 -582.85 113.585 -582.55 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.285 -582.85 133.585 -582.55 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 153.285 -582.85 153.585 -582.55 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.285 -582.85 173.585 -582.55 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.285 -582.85 193.585 -582.55 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -10.62 -582.85 -10.32 -582.55 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.125 -582.85 24.425 -582.55 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 184.125 -582.85 184.425 -582.55 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 344.125 -582.85 344.425 -582.55 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 504.125 -582.85 504.425 -582.55 ;
    END
  END wmask[3]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -87.435 -582.85 662.46 11.715 ;
    LAYER met2 SPACING 0.14 ;
      RECT -87.435 -582.85 662.46 11.715 ;
    LAYER met3 SPACING 0.3 ;
      RECT 635.115 -472.25 635.445 -471.92 ;
      RECT 635.13 -487.68 635.43 -471.92 ;
      RECT 635.115 -487.68 635.445 -487.35 ;
      RECT 635.13 -468.465 635.43 -424.72 ;
      RECT 635.115 -426.695 635.445 -426.365 ;
      RECT 635.115 -468.055 635.445 -467.725 ;
      RECT 634.515 -511.57 634.815 -435.98 ;
      RECT 634.5 -436.355 634.83 -436.025 ;
      RECT 634.5 -455.835 634.83 -455.505 ;
      RECT 634.5 -511.57 634.83 -511.24 ;
      RECT 633.9 -451.175 634.2 -436.61 ;
      RECT 633.885 -436.985 634.215 -436.655 ;
      RECT 633.885 -451.175 634.215 -450.845 ;
      RECT 633.27 -498.655 633.6 -498.325 ;
      RECT 633.285 -582.06 633.585 -498.325 ;
      RECT 633.27 -472.71 633.6 -472.38 ;
      RECT 633.285 -487.68 633.585 -472.38 ;
      RECT 633.27 -487.68 633.6 -487.35 ;
      RECT 633.285 -468.485 633.585 -424.72 ;
      RECT 633.27 -425.095 633.6 -424.765 ;
      RECT 633.27 -468.485 633.6 -468.155 ;
      RECT 623.245 -504.045 623.575 -503.715 ;
      RECT 623.26 -574.79 623.56 -503.715 ;
      RECT 623.245 -511.285 623.575 -510.955 ;
      RECT 623.245 -574.745 623.575 -574.415 ;
      RECT 622.615 -510.485 622.945 -510.155 ;
      RECT 622.63 -582.06 622.93 -510.155 ;
      RECT 622 -504.845 622.33 -504.515 ;
      RECT 622.015 -582.06 622.315 -504.515 ;
      RECT 615.115 -472.25 615.445 -471.92 ;
      RECT 615.13 -487.68 615.43 -471.92 ;
      RECT 615.115 -487.68 615.445 -487.35 ;
      RECT 615.13 -468.465 615.43 -424.72 ;
      RECT 615.115 -426.695 615.445 -426.365 ;
      RECT 615.115 -468.055 615.445 -467.725 ;
      RECT 614.515 -503.56 614.815 -435.98 ;
      RECT 614.5 -436.355 614.83 -436.025 ;
      RECT 614.5 -455.835 614.83 -455.505 ;
      RECT 614.5 -503.56 614.83 -503.23 ;
      RECT 613.9 -451.175 614.2 -436.61 ;
      RECT 613.885 -436.985 614.215 -436.655 ;
      RECT 613.885 -451.175 614.215 -450.845 ;
      RECT 613.27 -498.655 613.6 -498.325 ;
      RECT 613.285 -582.06 613.585 -498.325 ;
      RECT 613.27 -472.71 613.6 -472.38 ;
      RECT 613.285 -487.68 613.585 -472.38 ;
      RECT 613.27 -487.68 613.6 -487.35 ;
      RECT 613.285 -468.485 613.585 -424.72 ;
      RECT 613.27 -425.095 613.6 -424.765 ;
      RECT 613.27 -468.485 613.6 -468.155 ;
      RECT 595.115 -472.25 595.445 -471.92 ;
      RECT 595.13 -487.68 595.43 -471.92 ;
      RECT 595.115 -487.68 595.445 -487.35 ;
      RECT 595.13 -468.465 595.43 -424.72 ;
      RECT 595.115 -426.695 595.445 -426.365 ;
      RECT 595.115 -468.055 595.445 -467.725 ;
      RECT 594.515 -511.57 594.815 -435.98 ;
      RECT 594.5 -436.355 594.83 -436.025 ;
      RECT 594.5 -455.835 594.83 -455.505 ;
      RECT 594.5 -511.57 594.83 -511.24 ;
      RECT 593.9 -451.175 594.2 -436.61 ;
      RECT 593.885 -436.985 594.215 -436.655 ;
      RECT 593.885 -451.175 594.215 -450.845 ;
      RECT 593.27 -498.655 593.6 -498.325 ;
      RECT 593.285 -582.06 593.585 -498.325 ;
      RECT 593.27 -472.71 593.6 -472.38 ;
      RECT 593.285 -487.68 593.585 -472.38 ;
      RECT 593.27 -487.68 593.6 -487.35 ;
      RECT 593.285 -468.485 593.585 -424.72 ;
      RECT 593.27 -425.095 593.6 -424.765 ;
      RECT 593.27 -468.485 593.6 -468.155 ;
      RECT 583.245 -504.045 583.575 -503.715 ;
      RECT 583.26 -574.79 583.56 -503.715 ;
      RECT 583.245 -511.285 583.575 -510.955 ;
      RECT 583.245 -574.745 583.575 -574.415 ;
      RECT 582.615 -510.485 582.945 -510.155 ;
      RECT 582.63 -582.06 582.93 -510.155 ;
      RECT 582 -504.845 582.33 -504.515 ;
      RECT 582.015 -582.06 582.315 -504.515 ;
      RECT 575.115 -472.25 575.445 -471.92 ;
      RECT 575.13 -487.68 575.43 -471.92 ;
      RECT 575.115 -487.68 575.445 -487.35 ;
      RECT 575.13 -468.465 575.43 -424.72 ;
      RECT 575.115 -426.695 575.445 -426.365 ;
      RECT 575.115 -468.055 575.445 -467.725 ;
      RECT 574.515 -503.56 574.815 -435.98 ;
      RECT 574.5 -436.355 574.83 -436.025 ;
      RECT 574.5 -455.835 574.83 -455.505 ;
      RECT 574.5 -503.56 574.83 -503.23 ;
      RECT 573.9 -451.175 574.2 -436.61 ;
      RECT 573.885 -436.985 574.215 -436.655 ;
      RECT 573.885 -451.175 574.215 -450.845 ;
      RECT 573.27 -498.655 573.6 -498.325 ;
      RECT 573.285 -582.06 573.585 -498.325 ;
      RECT 573.27 -472.71 573.6 -472.38 ;
      RECT 573.285 -487.68 573.585 -472.38 ;
      RECT 573.27 -487.68 573.6 -487.35 ;
      RECT 573.285 -468.485 573.585 -424.72 ;
      RECT 573.27 -425.095 573.6 -424.765 ;
      RECT 573.27 -468.485 573.6 -468.155 ;
      RECT 555.115 -472.25 555.445 -471.92 ;
      RECT 555.13 -487.68 555.43 -471.92 ;
      RECT 555.115 -487.68 555.445 -487.35 ;
      RECT 555.13 -468.465 555.43 -424.72 ;
      RECT 555.115 -426.695 555.445 -426.365 ;
      RECT 555.115 -468.055 555.445 -467.725 ;
      RECT 554.515 -511.57 554.815 -435.98 ;
      RECT 554.5 -436.355 554.83 -436.025 ;
      RECT 554.5 -455.835 554.83 -455.505 ;
      RECT 554.5 -511.57 554.83 -511.24 ;
      RECT 553.9 -451.175 554.2 -436.61 ;
      RECT 553.885 -436.985 554.215 -436.655 ;
      RECT 553.885 -451.175 554.215 -450.845 ;
      RECT 553.27 -498.655 553.6 -498.325 ;
      RECT 553.285 -582.06 553.585 -498.325 ;
      RECT 553.27 -472.71 553.6 -472.38 ;
      RECT 553.285 -487.68 553.585 -472.38 ;
      RECT 553.27 -487.68 553.6 -487.35 ;
      RECT 553.285 -468.485 553.585 -424.72 ;
      RECT 553.27 -425.095 553.6 -424.765 ;
      RECT 553.27 -468.485 553.6 -468.155 ;
      RECT 543.245 -504.045 543.575 -503.715 ;
      RECT 543.26 -574.79 543.56 -503.715 ;
      RECT 543.245 -511.285 543.575 -510.955 ;
      RECT 543.245 -574.745 543.575 -574.415 ;
      RECT 542.615 -510.485 542.945 -510.155 ;
      RECT 542.63 -582.06 542.93 -510.155 ;
      RECT 542 -504.845 542.33 -504.515 ;
      RECT 542.015 -582.06 542.315 -504.515 ;
      RECT 535.115 -472.25 535.445 -471.92 ;
      RECT 535.13 -487.68 535.43 -471.92 ;
      RECT 535.115 -487.68 535.445 -487.35 ;
      RECT 535.13 -468.465 535.43 -424.72 ;
      RECT 535.115 -426.695 535.445 -426.365 ;
      RECT 535.115 -468.055 535.445 -467.725 ;
      RECT 534.515 -503.56 534.815 -435.98 ;
      RECT 534.5 -436.355 534.83 -436.025 ;
      RECT 534.5 -455.835 534.83 -455.505 ;
      RECT 534.5 -503.56 534.83 -503.23 ;
      RECT 533.9 -451.175 534.2 -436.61 ;
      RECT 533.885 -436.985 534.215 -436.655 ;
      RECT 533.885 -451.175 534.215 -450.845 ;
      RECT 533.27 -498.655 533.6 -498.325 ;
      RECT 533.285 -582.06 533.585 -498.325 ;
      RECT 533.27 -472.71 533.6 -472.38 ;
      RECT 533.285 -487.68 533.585 -472.38 ;
      RECT 533.27 -487.68 533.6 -487.35 ;
      RECT 533.285 -468.485 533.585 -424.72 ;
      RECT 533.27 -425.095 533.6 -424.765 ;
      RECT 533.27 -468.485 533.6 -468.155 ;
      RECT 516.3 -520.41 516.6 -440.705 ;
      RECT 516.285 -441.08 516.615 -440.75 ;
      RECT 516.285 -520.41 516.615 -520.08 ;
      RECT 515.115 -472.25 515.445 -471.92 ;
      RECT 515.13 -487.68 515.43 -471.92 ;
      RECT 515.115 -487.68 515.445 -487.35 ;
      RECT 515.13 -468.465 515.43 -424.72 ;
      RECT 515.115 -426.695 515.445 -426.365 ;
      RECT 515.115 -468.055 515.445 -467.725 ;
      RECT 514.515 -511.57 514.815 -435.98 ;
      RECT 514.5 -436.355 514.83 -436.025 ;
      RECT 514.5 -455.835 514.83 -455.505 ;
      RECT 514.5 -511.57 514.83 -511.24 ;
      RECT 513.9 -451.175 514.2 -436.61 ;
      RECT 513.885 -436.985 514.215 -436.655 ;
      RECT 513.885 -451.175 514.215 -450.845 ;
      RECT 513.27 -498.655 513.6 -498.325 ;
      RECT 513.285 -582.06 513.585 -498.325 ;
      RECT 513.27 -472.71 513.6 -472.38 ;
      RECT 513.285 -487.68 513.585 -472.38 ;
      RECT 513.27 -487.68 513.6 -487.35 ;
      RECT 513.285 -468.485 513.585 -424.72 ;
      RECT 513.27 -425.095 513.6 -424.765 ;
      RECT 513.27 -468.485 513.6 -468.155 ;
      RECT 504.11 -520.785 504.44 -520.455 ;
      RECT 504.125 -582.06 504.425 -520.455 ;
      RECT 503.245 -504.045 503.575 -503.715 ;
      RECT 503.26 -574.79 503.56 -503.715 ;
      RECT 503.245 -511.285 503.575 -510.955 ;
      RECT 503.245 -519.985 503.575 -519.655 ;
      RECT 503.245 -574.745 503.575 -574.415 ;
      RECT 502.615 -510.485 502.945 -510.155 ;
      RECT 502.63 -582.06 502.93 -510.155 ;
      RECT 502 -504.845 502.33 -504.515 ;
      RECT 502.015 -582.06 502.315 -504.515 ;
      RECT 495.115 -472.25 495.445 -471.92 ;
      RECT 495.13 -487.68 495.43 -471.92 ;
      RECT 495.115 -487.68 495.445 -487.35 ;
      RECT 495.13 -468.465 495.43 -424.72 ;
      RECT 495.115 -426.695 495.445 -426.365 ;
      RECT 495.115 -468.055 495.445 -467.725 ;
      RECT 494.515 -503.56 494.815 -435.98 ;
      RECT 494.5 -436.355 494.83 -436.025 ;
      RECT 494.5 -455.835 494.83 -455.505 ;
      RECT 494.5 -503.56 494.83 -503.23 ;
      RECT 493.9 -451.175 494.2 -436.61 ;
      RECT 493.885 -436.985 494.215 -436.655 ;
      RECT 493.885 -451.175 494.215 -450.845 ;
      RECT 493.27 -498.655 493.6 -498.325 ;
      RECT 493.285 -582.06 493.585 -498.325 ;
      RECT 493.27 -472.71 493.6 -472.38 ;
      RECT 493.285 -487.68 493.585 -472.38 ;
      RECT 493.27 -487.68 493.6 -487.35 ;
      RECT 493.285 -468.485 493.585 -424.72 ;
      RECT 493.27 -425.095 493.6 -424.765 ;
      RECT 493.27 -468.485 493.6 -468.155 ;
      RECT 475.115 -472.25 475.445 -471.92 ;
      RECT 475.13 -487.68 475.43 -471.92 ;
      RECT 475.115 -487.68 475.445 -487.35 ;
      RECT 475.13 -468.465 475.43 -424.72 ;
      RECT 475.115 -426.695 475.445 -426.365 ;
      RECT 475.115 -468.055 475.445 -467.725 ;
      RECT 474.515 -511.57 474.815 -435.98 ;
      RECT 474.5 -436.355 474.83 -436.025 ;
      RECT 474.5 -455.835 474.83 -455.505 ;
      RECT 474.5 -511.57 474.83 -511.24 ;
      RECT 473.9 -451.175 474.2 -436.61 ;
      RECT 473.885 -436.985 474.215 -436.655 ;
      RECT 473.885 -451.175 474.215 -450.845 ;
      RECT 473.27 -498.655 473.6 -498.325 ;
      RECT 473.285 -582.06 473.585 -498.325 ;
      RECT 473.27 -472.71 473.6 -472.38 ;
      RECT 473.285 -487.68 473.585 -472.38 ;
      RECT 473.27 -487.68 473.6 -487.35 ;
      RECT 473.285 -468.485 473.585 -424.72 ;
      RECT 473.27 -425.095 473.6 -424.765 ;
      RECT 473.27 -468.485 473.6 -468.155 ;
      RECT 463.245 -504.045 463.575 -503.715 ;
      RECT 463.26 -574.79 463.56 -503.715 ;
      RECT 463.245 -511.285 463.575 -510.955 ;
      RECT 463.245 -574.745 463.575 -574.415 ;
      RECT 462.615 -510.485 462.945 -510.155 ;
      RECT 462.63 -582.06 462.93 -510.155 ;
      RECT 462 -504.845 462.33 -504.515 ;
      RECT 462.015 -582.06 462.315 -504.515 ;
      RECT 455.115 -472.25 455.445 -471.92 ;
      RECT 455.13 -487.68 455.43 -471.92 ;
      RECT 455.115 -487.68 455.445 -487.35 ;
      RECT 455.13 -468.465 455.43 -424.72 ;
      RECT 455.115 -426.695 455.445 -426.365 ;
      RECT 455.115 -468.055 455.445 -467.725 ;
      RECT 454.515 -503.56 454.815 -435.98 ;
      RECT 454.5 -436.355 454.83 -436.025 ;
      RECT 454.5 -455.835 454.83 -455.505 ;
      RECT 454.5 -503.56 454.83 -503.23 ;
      RECT 453.9 -451.175 454.2 -436.61 ;
      RECT 453.885 -436.985 454.215 -436.655 ;
      RECT 453.885 -451.175 454.215 -450.845 ;
      RECT 453.27 -498.655 453.6 -498.325 ;
      RECT 453.285 -582.06 453.585 -498.325 ;
      RECT 453.27 -472.71 453.6 -472.38 ;
      RECT 453.285 -487.68 453.585 -472.38 ;
      RECT 453.27 -487.68 453.6 -487.35 ;
      RECT 453.285 -468.485 453.585 -424.72 ;
      RECT 453.27 -425.095 453.6 -424.765 ;
      RECT 453.27 -468.485 453.6 -468.155 ;
      RECT 435.115 -472.25 435.445 -471.92 ;
      RECT 435.13 -487.68 435.43 -471.92 ;
      RECT 435.115 -487.68 435.445 -487.35 ;
      RECT 435.13 -468.465 435.43 -424.72 ;
      RECT 435.115 -426.695 435.445 -426.365 ;
      RECT 435.115 -468.055 435.445 -467.725 ;
      RECT 434.515 -511.57 434.815 -435.98 ;
      RECT 434.5 -436.355 434.83 -436.025 ;
      RECT 434.5 -455.835 434.83 -455.505 ;
      RECT 434.5 -511.57 434.83 -511.24 ;
      RECT 433.9 -451.175 434.2 -436.61 ;
      RECT 433.885 -436.985 434.215 -436.655 ;
      RECT 433.885 -451.175 434.215 -450.845 ;
      RECT 433.27 -498.655 433.6 -498.325 ;
      RECT 433.285 -582.06 433.585 -498.325 ;
      RECT 433.27 -472.71 433.6 -472.38 ;
      RECT 433.285 -487.68 433.585 -472.38 ;
      RECT 433.27 -487.68 433.6 -487.35 ;
      RECT 433.285 -468.485 433.585 -424.72 ;
      RECT 433.27 -425.095 433.6 -424.765 ;
      RECT 433.27 -468.485 433.6 -468.155 ;
      RECT 423.245 -504.045 423.575 -503.715 ;
      RECT 423.26 -574.79 423.56 -503.715 ;
      RECT 423.245 -511.285 423.575 -510.955 ;
      RECT 423.245 -574.745 423.575 -574.415 ;
      RECT 422.615 -510.485 422.945 -510.155 ;
      RECT 422.63 -582.06 422.93 -510.155 ;
      RECT 422 -504.845 422.33 -504.515 ;
      RECT 422.015 -582.06 422.315 -504.515 ;
      RECT 415.115 -472.25 415.445 -471.92 ;
      RECT 415.13 -487.68 415.43 -471.92 ;
      RECT 415.115 -487.68 415.445 -487.35 ;
      RECT 415.13 -468.465 415.43 -424.72 ;
      RECT 415.115 -426.695 415.445 -426.365 ;
      RECT 415.115 -468.055 415.445 -467.725 ;
      RECT 414.515 -503.56 414.815 -435.98 ;
      RECT 414.5 -436.355 414.83 -436.025 ;
      RECT 414.5 -455.835 414.83 -455.505 ;
      RECT 414.5 -503.56 414.83 -503.23 ;
      RECT 413.9 -451.175 414.2 -436.61 ;
      RECT 413.885 -436.985 414.215 -436.655 ;
      RECT 413.885 -451.175 414.215 -450.845 ;
      RECT 413.27 -498.655 413.6 -498.325 ;
      RECT 413.285 -582.06 413.585 -498.325 ;
      RECT 413.27 -472.71 413.6 -472.38 ;
      RECT 413.285 -487.68 413.585 -472.38 ;
      RECT 413.27 -487.68 413.6 -487.35 ;
      RECT 413.285 -468.485 413.585 -424.72 ;
      RECT 413.27 -425.095 413.6 -424.765 ;
      RECT 413.27 -468.485 413.6 -468.155 ;
      RECT 395.115 -472.25 395.445 -471.92 ;
      RECT 395.13 -487.68 395.43 -471.92 ;
      RECT 395.115 -487.68 395.445 -487.35 ;
      RECT 395.13 -468.465 395.43 -424.72 ;
      RECT 395.115 -426.695 395.445 -426.365 ;
      RECT 395.115 -468.055 395.445 -467.725 ;
      RECT 394.515 -511.57 394.815 -435.98 ;
      RECT 394.5 -436.355 394.83 -436.025 ;
      RECT 394.5 -455.835 394.83 -455.505 ;
      RECT 394.5 -511.57 394.83 -511.24 ;
      RECT 393.9 -451.175 394.2 -436.61 ;
      RECT 393.885 -436.985 394.215 -436.655 ;
      RECT 393.885 -451.175 394.215 -450.845 ;
      RECT 393.27 -498.655 393.6 -498.325 ;
      RECT 393.285 -582.06 393.585 -498.325 ;
      RECT 393.27 -472.71 393.6 -472.38 ;
      RECT 393.285 -487.68 393.585 -472.38 ;
      RECT 393.27 -487.68 393.6 -487.35 ;
      RECT 393.285 -468.485 393.585 -424.72 ;
      RECT 393.27 -425.095 393.6 -424.765 ;
      RECT 393.27 -468.485 393.6 -468.155 ;
      RECT 383.245 -504.045 383.575 -503.715 ;
      RECT 383.26 -574.79 383.56 -503.715 ;
      RECT 383.245 -511.285 383.575 -510.955 ;
      RECT 383.245 -574.745 383.575 -574.415 ;
      RECT 382.615 -510.485 382.945 -510.155 ;
      RECT 382.63 -582.06 382.93 -510.155 ;
      RECT 382 -504.845 382.33 -504.515 ;
      RECT 382.015 -582.06 382.315 -504.515 ;
      RECT 375.115 -472.25 375.445 -471.92 ;
      RECT 375.13 -487.68 375.43 -471.92 ;
      RECT 375.115 -487.68 375.445 -487.35 ;
      RECT 375.13 -468.465 375.43 -424.72 ;
      RECT 375.115 -426.695 375.445 -426.365 ;
      RECT 375.115 -468.055 375.445 -467.725 ;
      RECT 374.515 -503.56 374.815 -435.98 ;
      RECT 374.5 -436.355 374.83 -436.025 ;
      RECT 374.5 -455.835 374.83 -455.505 ;
      RECT 374.5 -503.56 374.83 -503.23 ;
      RECT 373.9 -451.175 374.2 -436.61 ;
      RECT 373.885 -436.985 374.215 -436.655 ;
      RECT 373.885 -451.175 374.215 -450.845 ;
      RECT 373.27 -498.655 373.6 -498.325 ;
      RECT 373.285 -582.06 373.585 -498.325 ;
      RECT 373.27 -472.71 373.6 -472.38 ;
      RECT 373.285 -487.68 373.585 -472.38 ;
      RECT 373.27 -487.68 373.6 -487.35 ;
      RECT 373.285 -468.485 373.585 -424.72 ;
      RECT 373.27 -425.095 373.6 -424.765 ;
      RECT 373.27 -468.485 373.6 -468.155 ;
      RECT 356.3 -520.41 356.6 -440.705 ;
      RECT 356.285 -441.08 356.615 -440.75 ;
      RECT 356.285 -520.41 356.615 -520.08 ;
      RECT 355.115 -472.25 355.445 -471.92 ;
      RECT 355.13 -487.68 355.43 -471.92 ;
      RECT 355.115 -487.68 355.445 -487.35 ;
      RECT 355.13 -468.465 355.43 -424.72 ;
      RECT 355.115 -426.695 355.445 -426.365 ;
      RECT 355.115 -468.055 355.445 -467.725 ;
      RECT 354.515 -511.57 354.815 -435.98 ;
      RECT 354.5 -436.355 354.83 -436.025 ;
      RECT 354.5 -455.835 354.83 -455.505 ;
      RECT 354.5 -511.57 354.83 -511.24 ;
      RECT 353.9 -451.175 354.2 -436.61 ;
      RECT 353.885 -436.985 354.215 -436.655 ;
      RECT 353.885 -451.175 354.215 -450.845 ;
      RECT 353.27 -498.655 353.6 -498.325 ;
      RECT 353.285 -582.06 353.585 -498.325 ;
      RECT 353.27 -472.71 353.6 -472.38 ;
      RECT 353.285 -487.68 353.585 -472.38 ;
      RECT 353.27 -487.68 353.6 -487.35 ;
      RECT 353.285 -468.485 353.585 -424.72 ;
      RECT 353.27 -425.095 353.6 -424.765 ;
      RECT 353.27 -468.485 353.6 -468.155 ;
      RECT 344.11 -520.785 344.44 -520.455 ;
      RECT 344.125 -582.06 344.425 -520.455 ;
      RECT 343.245 -504.045 343.575 -503.715 ;
      RECT 343.26 -574.79 343.56 -503.715 ;
      RECT 343.245 -511.285 343.575 -510.955 ;
      RECT 343.245 -519.985 343.575 -519.655 ;
      RECT 343.245 -574.745 343.575 -574.415 ;
      RECT 342.615 -510.485 342.945 -510.155 ;
      RECT 342.63 -582.06 342.93 -510.155 ;
      RECT 342 -504.845 342.33 -504.515 ;
      RECT 342.015 -582.06 342.315 -504.515 ;
      RECT 335.115 -472.25 335.445 -471.92 ;
      RECT 335.13 -487.68 335.43 -471.92 ;
      RECT 335.115 -487.68 335.445 -487.35 ;
      RECT 335.13 -468.465 335.43 -424.72 ;
      RECT 335.115 -426.695 335.445 -426.365 ;
      RECT 335.115 -468.055 335.445 -467.725 ;
      RECT 334.515 -503.56 334.815 -435.98 ;
      RECT 334.5 -436.355 334.83 -436.025 ;
      RECT 334.5 -455.835 334.83 -455.505 ;
      RECT 334.5 -503.56 334.83 -503.23 ;
      RECT 333.9 -451.175 334.2 -436.61 ;
      RECT 333.885 -436.985 334.215 -436.655 ;
      RECT 333.885 -451.175 334.215 -450.845 ;
      RECT 333.27 -498.655 333.6 -498.325 ;
      RECT 333.285 -582.06 333.585 -498.325 ;
      RECT 333.27 -472.71 333.6 -472.38 ;
      RECT 333.285 -487.68 333.585 -472.38 ;
      RECT 333.27 -487.68 333.6 -487.35 ;
      RECT 333.285 -468.485 333.585 -424.72 ;
      RECT 333.27 -425.095 333.6 -424.765 ;
      RECT 333.27 -468.485 333.6 -468.155 ;
      RECT 315.115 -472.25 315.445 -471.92 ;
      RECT 315.13 -487.68 315.43 -471.92 ;
      RECT 315.115 -487.68 315.445 -487.35 ;
      RECT 315.13 -468.465 315.43 -424.72 ;
      RECT 315.115 -426.695 315.445 -426.365 ;
      RECT 315.115 -468.055 315.445 -467.725 ;
      RECT 314.515 -511.57 314.815 -435.98 ;
      RECT 314.5 -436.355 314.83 -436.025 ;
      RECT 314.5 -455.835 314.83 -455.505 ;
      RECT 314.5 -511.57 314.83 -511.24 ;
      RECT 313.9 -451.175 314.2 -436.61 ;
      RECT 313.885 -436.985 314.215 -436.655 ;
      RECT 313.885 -451.175 314.215 -450.845 ;
      RECT 313.27 -498.655 313.6 -498.325 ;
      RECT 313.285 -582.06 313.585 -498.325 ;
      RECT 313.27 -472.71 313.6 -472.38 ;
      RECT 313.285 -487.68 313.585 -472.38 ;
      RECT 313.27 -487.68 313.6 -487.35 ;
      RECT 313.285 -468.485 313.585 -424.72 ;
      RECT 313.27 -425.095 313.6 -424.765 ;
      RECT 313.27 -468.485 313.6 -468.155 ;
      RECT 303.245 -504.045 303.575 -503.715 ;
      RECT 303.26 -574.79 303.56 -503.715 ;
      RECT 303.245 -511.285 303.575 -510.955 ;
      RECT 303.245 -574.745 303.575 -574.415 ;
      RECT 302.615 -510.485 302.945 -510.155 ;
      RECT 302.63 -582.06 302.93 -510.155 ;
      RECT 302 -504.845 302.33 -504.515 ;
      RECT 302.015 -582.06 302.315 -504.515 ;
      RECT 295.115 -472.25 295.445 -471.92 ;
      RECT 295.13 -487.68 295.43 -471.92 ;
      RECT 295.115 -487.68 295.445 -487.35 ;
      RECT 295.13 -468.465 295.43 -424.72 ;
      RECT 295.115 -426.695 295.445 -426.365 ;
      RECT 295.115 -468.055 295.445 -467.725 ;
      RECT 294.515 -503.56 294.815 -435.98 ;
      RECT 294.5 -436.355 294.83 -436.025 ;
      RECT 294.5 -455.835 294.83 -455.505 ;
      RECT 294.5 -503.56 294.83 -503.23 ;
      RECT 293.9 -451.175 294.2 -436.61 ;
      RECT 293.885 -436.985 294.215 -436.655 ;
      RECT 293.885 -451.175 294.215 -450.845 ;
      RECT 293.27 -498.655 293.6 -498.325 ;
      RECT 293.285 -582.06 293.585 -498.325 ;
      RECT 293.27 -472.71 293.6 -472.38 ;
      RECT 293.285 -487.68 293.585 -472.38 ;
      RECT 293.27 -487.68 293.6 -487.35 ;
      RECT 293.285 -468.485 293.585 -424.72 ;
      RECT 293.27 -425.095 293.6 -424.765 ;
      RECT 293.27 -468.485 293.6 -468.155 ;
      RECT 275.115 -472.25 275.445 -471.92 ;
      RECT 275.13 -487.68 275.43 -471.92 ;
      RECT 275.115 -487.68 275.445 -487.35 ;
      RECT 275.13 -468.465 275.43 -424.72 ;
      RECT 275.115 -426.695 275.445 -426.365 ;
      RECT 275.115 -468.055 275.445 -467.725 ;
      RECT 274.515 -511.57 274.815 -435.98 ;
      RECT 274.5 -436.355 274.83 -436.025 ;
      RECT 274.5 -455.835 274.83 -455.505 ;
      RECT 274.5 -511.57 274.83 -511.24 ;
      RECT 273.9 -451.175 274.2 -436.61 ;
      RECT 273.885 -436.985 274.215 -436.655 ;
      RECT 273.885 -451.175 274.215 -450.845 ;
      RECT 273.27 -498.655 273.6 -498.325 ;
      RECT 273.285 -582.06 273.585 -498.325 ;
      RECT 273.27 -472.71 273.6 -472.38 ;
      RECT 273.285 -487.68 273.585 -472.38 ;
      RECT 273.27 -487.68 273.6 -487.35 ;
      RECT 273.285 -468.485 273.585 -424.72 ;
      RECT 273.27 -425.095 273.6 -424.765 ;
      RECT 273.27 -468.485 273.6 -468.155 ;
      RECT 263.245 -504.045 263.575 -503.715 ;
      RECT 263.26 -574.79 263.56 -503.715 ;
      RECT 263.245 -511.285 263.575 -510.955 ;
      RECT 263.245 -574.745 263.575 -574.415 ;
      RECT 262.615 -510.485 262.945 -510.155 ;
      RECT 262.63 -582.06 262.93 -510.155 ;
      RECT 262 -504.845 262.33 -504.515 ;
      RECT 262.015 -582.06 262.315 -504.515 ;
      RECT 255.115 -472.25 255.445 -471.92 ;
      RECT 255.13 -487.68 255.43 -471.92 ;
      RECT 255.115 -487.68 255.445 -487.35 ;
      RECT 255.13 -468.465 255.43 -424.72 ;
      RECT 255.115 -426.695 255.445 -426.365 ;
      RECT 255.115 -468.055 255.445 -467.725 ;
      RECT 254.515 -503.56 254.815 -435.98 ;
      RECT 254.5 -436.355 254.83 -436.025 ;
      RECT 254.5 -455.835 254.83 -455.505 ;
      RECT 254.5 -503.56 254.83 -503.23 ;
      RECT 253.9 -451.175 254.2 -436.61 ;
      RECT 253.885 -436.985 254.215 -436.655 ;
      RECT 253.885 -451.175 254.215 -450.845 ;
      RECT 253.27 -498.655 253.6 -498.325 ;
      RECT 253.285 -582.06 253.585 -498.325 ;
      RECT 253.27 -472.71 253.6 -472.38 ;
      RECT 253.285 -487.68 253.585 -472.38 ;
      RECT 253.27 -487.68 253.6 -487.35 ;
      RECT 253.285 -468.485 253.585 -424.72 ;
      RECT 253.27 -425.095 253.6 -424.765 ;
      RECT 253.27 -468.485 253.6 -468.155 ;
      RECT 235.115 -472.25 235.445 -471.92 ;
      RECT 235.13 -487.68 235.43 -471.92 ;
      RECT 235.115 -487.68 235.445 -487.35 ;
      RECT 235.13 -468.465 235.43 -424.72 ;
      RECT 235.115 -426.695 235.445 -426.365 ;
      RECT 235.115 -468.055 235.445 -467.725 ;
      RECT 234.515 -511.57 234.815 -435.98 ;
      RECT 234.5 -436.355 234.83 -436.025 ;
      RECT 234.5 -455.835 234.83 -455.505 ;
      RECT 234.5 -511.57 234.83 -511.24 ;
      RECT 233.9 -451.175 234.2 -436.61 ;
      RECT 233.885 -436.985 234.215 -436.655 ;
      RECT 233.885 -451.175 234.215 -450.845 ;
      RECT 233.27 -498.655 233.6 -498.325 ;
      RECT 233.285 -582.06 233.585 -498.325 ;
      RECT 233.27 -472.71 233.6 -472.38 ;
      RECT 233.285 -487.68 233.585 -472.38 ;
      RECT 233.27 -487.68 233.6 -487.35 ;
      RECT 233.285 -468.485 233.585 -424.72 ;
      RECT 233.27 -425.095 233.6 -424.765 ;
      RECT 233.27 -468.485 233.6 -468.155 ;
      RECT 223.245 -504.045 223.575 -503.715 ;
      RECT 223.26 -574.79 223.56 -503.715 ;
      RECT 223.245 -511.285 223.575 -510.955 ;
      RECT 223.245 -574.745 223.575 -574.415 ;
      RECT 222.615 -510.485 222.945 -510.155 ;
      RECT 222.63 -582.06 222.93 -510.155 ;
      RECT 222 -504.845 222.33 -504.515 ;
      RECT 222.015 -582.06 222.315 -504.515 ;
      RECT 215.115 -472.25 215.445 -471.92 ;
      RECT 215.13 -487.68 215.43 -471.92 ;
      RECT 215.115 -487.68 215.445 -487.35 ;
      RECT 215.13 -468.465 215.43 -424.72 ;
      RECT 215.115 -426.695 215.445 -426.365 ;
      RECT 215.115 -468.055 215.445 -467.725 ;
      RECT 214.515 -503.56 214.815 -435.98 ;
      RECT 214.5 -436.355 214.83 -436.025 ;
      RECT 214.5 -455.835 214.83 -455.505 ;
      RECT 214.5 -503.56 214.83 -503.23 ;
      RECT 213.9 -451.175 214.2 -436.61 ;
      RECT 213.885 -436.985 214.215 -436.655 ;
      RECT 213.885 -451.175 214.215 -450.845 ;
      RECT 213.27 -498.655 213.6 -498.325 ;
      RECT 213.285 -582.06 213.585 -498.325 ;
      RECT 213.27 -472.71 213.6 -472.38 ;
      RECT 213.285 -487.68 213.585 -472.38 ;
      RECT 213.27 -487.68 213.6 -487.35 ;
      RECT 213.285 -468.485 213.585 -424.72 ;
      RECT 213.27 -425.095 213.6 -424.765 ;
      RECT 213.27 -468.485 213.6 -468.155 ;
      RECT 196.3 -520.41 196.6 -440.705 ;
      RECT 196.285 -441.08 196.615 -440.75 ;
      RECT 196.285 -520.41 196.615 -520.08 ;
      RECT 195.115 -472.25 195.445 -471.92 ;
      RECT 195.13 -487.68 195.43 -471.92 ;
      RECT 195.115 -487.68 195.445 -487.35 ;
      RECT 195.13 -468.465 195.43 -424.72 ;
      RECT 195.115 -426.695 195.445 -426.365 ;
      RECT 195.115 -468.055 195.445 -467.725 ;
      RECT 194.515 -511.57 194.815 -435.98 ;
      RECT 194.5 -436.355 194.83 -436.025 ;
      RECT 194.5 -455.835 194.83 -455.505 ;
      RECT 194.5 -511.57 194.83 -511.24 ;
      RECT 193.9 -451.175 194.2 -436.61 ;
      RECT 193.885 -436.985 194.215 -436.655 ;
      RECT 193.885 -451.175 194.215 -450.845 ;
      RECT 193.27 -498.655 193.6 -498.325 ;
      RECT 193.285 -582.06 193.585 -498.325 ;
      RECT 193.27 -472.71 193.6 -472.38 ;
      RECT 193.285 -487.68 193.585 -472.38 ;
      RECT 193.27 -487.68 193.6 -487.35 ;
      RECT 193.285 -468.485 193.585 -424.72 ;
      RECT 193.27 -425.095 193.6 -424.765 ;
      RECT 193.27 -468.485 193.6 -468.155 ;
      RECT 184.11 -520.785 184.44 -520.455 ;
      RECT 184.125 -582.06 184.425 -520.455 ;
      RECT 183.245 -504.045 183.575 -503.715 ;
      RECT 183.26 -574.79 183.56 -503.715 ;
      RECT 183.245 -511.285 183.575 -510.955 ;
      RECT 183.245 -519.985 183.575 -519.655 ;
      RECT 183.245 -574.745 183.575 -574.415 ;
      RECT 182.615 -510.485 182.945 -510.155 ;
      RECT 182.63 -582.06 182.93 -510.155 ;
      RECT 182 -504.845 182.33 -504.515 ;
      RECT 182.015 -582.06 182.315 -504.515 ;
      RECT 175.115 -472.25 175.445 -471.92 ;
      RECT 175.13 -487.68 175.43 -471.92 ;
      RECT 175.115 -487.68 175.445 -487.35 ;
      RECT 175.13 -468.465 175.43 -424.72 ;
      RECT 175.115 -426.695 175.445 -426.365 ;
      RECT 175.115 -468.055 175.445 -467.725 ;
      RECT 174.515 -503.56 174.815 -435.98 ;
      RECT 174.5 -436.355 174.83 -436.025 ;
      RECT 174.5 -455.835 174.83 -455.505 ;
      RECT 174.5 -503.56 174.83 -503.23 ;
      RECT 173.9 -451.175 174.2 -436.61 ;
      RECT 173.885 -436.985 174.215 -436.655 ;
      RECT 173.885 -451.175 174.215 -450.845 ;
      RECT 173.27 -498.655 173.6 -498.325 ;
      RECT 173.285 -582.06 173.585 -498.325 ;
      RECT 173.27 -472.71 173.6 -472.38 ;
      RECT 173.285 -487.68 173.585 -472.38 ;
      RECT 173.27 -487.68 173.6 -487.35 ;
      RECT 173.285 -468.485 173.585 -424.72 ;
      RECT 173.27 -425.095 173.6 -424.765 ;
      RECT 173.27 -468.485 173.6 -468.155 ;
      RECT 155.115 -472.25 155.445 -471.92 ;
      RECT 155.13 -487.68 155.43 -471.92 ;
      RECT 155.115 -487.68 155.445 -487.35 ;
      RECT 155.13 -468.465 155.43 -424.72 ;
      RECT 155.115 -426.695 155.445 -426.365 ;
      RECT 155.115 -468.055 155.445 -467.725 ;
      RECT 154.515 -511.57 154.815 -435.98 ;
      RECT 154.5 -436.355 154.83 -436.025 ;
      RECT 154.5 -455.835 154.83 -455.505 ;
      RECT 154.5 -511.57 154.83 -511.24 ;
      RECT 153.9 -451.175 154.2 -436.61 ;
      RECT 153.885 -436.985 154.215 -436.655 ;
      RECT 153.885 -451.175 154.215 -450.845 ;
      RECT 153.27 -498.655 153.6 -498.325 ;
      RECT 153.285 -582.06 153.585 -498.325 ;
      RECT 153.27 -472.71 153.6 -472.38 ;
      RECT 153.285 -487.68 153.585 -472.38 ;
      RECT 153.27 -487.68 153.6 -487.35 ;
      RECT 153.285 -468.485 153.585 -424.72 ;
      RECT 153.27 -425.095 153.6 -424.765 ;
      RECT 153.27 -468.485 153.6 -468.155 ;
      RECT 143.245 -504.045 143.575 -503.715 ;
      RECT 143.26 -574.79 143.56 -503.715 ;
      RECT 143.245 -511.285 143.575 -510.955 ;
      RECT 143.245 -574.745 143.575 -574.415 ;
      RECT 142.615 -510.485 142.945 -510.155 ;
      RECT 142.63 -582.06 142.93 -510.155 ;
      RECT 142 -504.845 142.33 -504.515 ;
      RECT 142.015 -582.06 142.315 -504.515 ;
      RECT 135.115 -472.25 135.445 -471.92 ;
      RECT 135.13 -487.68 135.43 -471.92 ;
      RECT 135.115 -487.68 135.445 -487.35 ;
      RECT 135.13 -468.465 135.43 -424.72 ;
      RECT 135.115 -426.695 135.445 -426.365 ;
      RECT 135.115 -468.055 135.445 -467.725 ;
      RECT 134.515 -503.56 134.815 -435.98 ;
      RECT 134.5 -436.355 134.83 -436.025 ;
      RECT 134.5 -455.835 134.83 -455.505 ;
      RECT 134.5 -503.56 134.83 -503.23 ;
      RECT 133.9 -451.175 134.2 -436.61 ;
      RECT 133.885 -436.985 134.215 -436.655 ;
      RECT 133.885 -451.175 134.215 -450.845 ;
      RECT 133.27 -498.655 133.6 -498.325 ;
      RECT 133.285 -582.06 133.585 -498.325 ;
      RECT 133.27 -472.71 133.6 -472.38 ;
      RECT 133.285 -487.68 133.585 -472.38 ;
      RECT 133.27 -487.68 133.6 -487.35 ;
      RECT 133.285 -468.485 133.585 -424.72 ;
      RECT 133.27 -425.095 133.6 -424.765 ;
      RECT 133.27 -468.485 133.6 -468.155 ;
      RECT 115.115 -472.25 115.445 -471.92 ;
      RECT 115.13 -487.68 115.43 -471.92 ;
      RECT 115.115 -487.68 115.445 -487.35 ;
      RECT 115.13 -468.465 115.43 -424.72 ;
      RECT 115.115 -426.695 115.445 -426.365 ;
      RECT 115.115 -468.055 115.445 -467.725 ;
      RECT 114.515 -511.57 114.815 -435.98 ;
      RECT 114.5 -436.355 114.83 -436.025 ;
      RECT 114.5 -455.835 114.83 -455.505 ;
      RECT 114.5 -511.57 114.83 -511.24 ;
      RECT 113.9 -451.175 114.2 -436.61 ;
      RECT 113.885 -436.985 114.215 -436.655 ;
      RECT 113.885 -451.175 114.215 -450.845 ;
      RECT 113.27 -498.655 113.6 -498.325 ;
      RECT 113.285 -582.06 113.585 -498.325 ;
      RECT 113.27 -472.71 113.6 -472.38 ;
      RECT 113.285 -487.68 113.585 -472.38 ;
      RECT 113.27 -487.68 113.6 -487.35 ;
      RECT 113.285 -468.485 113.585 -424.72 ;
      RECT 113.27 -425.095 113.6 -424.765 ;
      RECT 113.27 -468.485 113.6 -468.155 ;
      RECT 103.245 -504.045 103.575 -503.715 ;
      RECT 103.26 -574.79 103.56 -503.715 ;
      RECT 103.245 -511.285 103.575 -510.955 ;
      RECT 103.245 -574.745 103.575 -574.415 ;
      RECT 102.615 -510.485 102.945 -510.155 ;
      RECT 102.63 -582.06 102.93 -510.155 ;
      RECT 102 -504.845 102.33 -504.515 ;
      RECT 102.015 -582.06 102.315 -504.515 ;
      RECT 95.115 -472.25 95.445 -471.92 ;
      RECT 95.13 -487.68 95.43 -471.92 ;
      RECT 95.115 -487.68 95.445 -487.35 ;
      RECT 95.13 -468.465 95.43 -424.72 ;
      RECT 95.115 -426.695 95.445 -426.365 ;
      RECT 95.115 -468.055 95.445 -467.725 ;
      RECT 94.515 -503.56 94.815 -435.98 ;
      RECT 94.5 -436.355 94.83 -436.025 ;
      RECT 94.5 -455.835 94.83 -455.505 ;
      RECT 94.5 -503.56 94.83 -503.23 ;
      RECT 93.9 -451.175 94.2 -436.61 ;
      RECT 93.885 -436.985 94.215 -436.655 ;
      RECT 93.885 -451.175 94.215 -450.845 ;
      RECT 93.27 -498.655 93.6 -498.325 ;
      RECT 93.285 -582.06 93.585 -498.325 ;
      RECT 93.27 -472.71 93.6 -472.38 ;
      RECT 93.285 -487.68 93.585 -472.38 ;
      RECT 93.27 -487.68 93.6 -487.35 ;
      RECT 93.285 -468.485 93.585 -424.72 ;
      RECT 93.27 -425.095 93.6 -424.765 ;
      RECT 93.27 -468.485 93.6 -468.155 ;
      RECT 75.115 -472.25 75.445 -471.92 ;
      RECT 75.13 -487.68 75.43 -471.92 ;
      RECT 75.115 -487.68 75.445 -487.35 ;
      RECT 75.13 -468.465 75.43 -424.72 ;
      RECT 75.115 -426.695 75.445 -426.365 ;
      RECT 75.115 -468.055 75.445 -467.725 ;
      RECT 74.515 -511.57 74.815 -435.98 ;
      RECT 74.5 -436.355 74.83 -436.025 ;
      RECT 74.5 -455.835 74.83 -455.505 ;
      RECT 74.5 -511.57 74.83 -511.24 ;
      RECT 73.9 -451.175 74.2 -436.61 ;
      RECT 73.885 -436.985 74.215 -436.655 ;
      RECT 73.885 -451.175 74.215 -450.845 ;
      RECT 73.27 -498.655 73.6 -498.325 ;
      RECT 73.285 -582.06 73.585 -498.325 ;
      RECT 73.27 -472.71 73.6 -472.38 ;
      RECT 73.285 -487.68 73.585 -472.38 ;
      RECT 73.27 -487.68 73.6 -487.35 ;
      RECT 73.285 -468.485 73.585 -424.72 ;
      RECT 73.27 -425.095 73.6 -424.765 ;
      RECT 73.27 -468.485 73.6 -468.155 ;
      RECT 63.245 -504.045 63.575 -503.715 ;
      RECT 63.26 -574.79 63.56 -503.715 ;
      RECT 63.245 -511.285 63.575 -510.955 ;
      RECT 63.245 -574.745 63.575 -574.415 ;
      RECT 62.615 -510.485 62.945 -510.155 ;
      RECT 62.63 -582.06 62.93 -510.155 ;
      RECT 62 -504.845 62.33 -504.515 ;
      RECT 62.015 -582.06 62.315 -504.515 ;
      RECT 55.115 -472.25 55.445 -471.92 ;
      RECT 55.13 -487.68 55.43 -471.92 ;
      RECT 55.115 -487.68 55.445 -487.35 ;
      RECT 55.13 -468.465 55.43 -424.72 ;
      RECT 55.115 -426.695 55.445 -426.365 ;
      RECT 55.115 -468.055 55.445 -467.725 ;
      RECT 54.515 -503.56 54.815 -435.98 ;
      RECT 54.5 -436.355 54.83 -436.025 ;
      RECT 54.5 -455.835 54.83 -455.505 ;
      RECT 54.5 -503.56 54.83 -503.23 ;
      RECT 53.9 -451.175 54.2 -436.61 ;
      RECT 53.885 -436.985 54.215 -436.655 ;
      RECT 53.885 -451.175 54.215 -450.845 ;
      RECT 53.27 -498.655 53.6 -498.325 ;
      RECT 53.285 -582.06 53.585 -498.325 ;
      RECT 53.27 -472.71 53.6 -472.38 ;
      RECT 53.285 -487.68 53.585 -472.38 ;
      RECT 53.27 -487.68 53.6 -487.35 ;
      RECT 53.285 -468.485 53.585 -424.72 ;
      RECT 53.27 -425.095 53.6 -424.765 ;
      RECT 53.27 -468.485 53.6 -468.155 ;
      RECT 36.3 -520.41 36.6 -440.705 ;
      RECT 36.285 -441.08 36.615 -440.75 ;
      RECT 36.285 -520.41 36.615 -520.08 ;
      RECT 35.115 -472.25 35.445 -471.92 ;
      RECT 35.13 -487.68 35.43 -471.92 ;
      RECT 35.115 -487.68 35.445 -487.35 ;
      RECT 35.13 -468.465 35.43 -424.72 ;
      RECT 35.115 -426.695 35.445 -426.365 ;
      RECT 35.115 -468.055 35.445 -467.725 ;
      RECT 34.515 -511.57 34.815 -435.98 ;
      RECT 34.5 -436.355 34.83 -436.025 ;
      RECT 34.5 -455.835 34.83 -455.505 ;
      RECT 34.5 -511.57 34.83 -511.24 ;
      RECT 33.9 -451.175 34.2 -436.61 ;
      RECT 33.885 -436.985 34.215 -436.655 ;
      RECT 33.885 -451.175 34.215 -450.845 ;
      RECT 33.27 -498.655 33.6 -498.325 ;
      RECT 33.285 -582.06 33.585 -498.325 ;
      RECT 33.27 -472.71 33.6 -472.38 ;
      RECT 33.285 -487.68 33.585 -472.38 ;
      RECT 33.27 -487.68 33.6 -487.35 ;
      RECT 33.285 -468.485 33.585 -424.72 ;
      RECT 33.27 -425.095 33.6 -424.765 ;
      RECT 33.27 -468.485 33.6 -468.155 ;
      RECT 24.11 -520.785 24.44 -520.455 ;
      RECT 24.125 -582.06 24.425 -520.455 ;
      RECT 23.245 -504.045 23.575 -503.715 ;
      RECT 23.26 -574.79 23.56 -503.715 ;
      RECT 23.245 -511.285 23.575 -510.955 ;
      RECT 23.245 -519.985 23.575 -519.655 ;
      RECT 23.245 -574.745 23.575 -574.415 ;
      RECT 22.615 -510.485 22.945 -510.155 ;
      RECT 22.63 -582.06 22.93 -510.155 ;
      RECT 22 -504.845 22.33 -504.515 ;
      RECT 22.015 -582.06 22.315 -504.515 ;
      RECT 15.115 -472.25 15.445 -471.92 ;
      RECT 15.13 -487.68 15.43 -471.92 ;
      RECT 15.115 -487.68 15.445 -487.35 ;
      RECT 15.13 -468.465 15.43 -424.72 ;
      RECT 15.115 -426.695 15.445 -426.365 ;
      RECT 15.115 -468.055 15.445 -467.725 ;
      RECT 14.515 -503.56 14.815 -435.98 ;
      RECT 14.5 -436.355 14.83 -436.025 ;
      RECT 14.5 -455.835 14.83 -455.505 ;
      RECT 14.5 -503.56 14.83 -503.23 ;
      RECT 13.9 -451.175 14.2 -436.61 ;
      RECT 13.885 -436.985 14.215 -436.655 ;
      RECT 13.885 -451.175 14.215 -450.845 ;
      RECT 13.27 -498.655 13.6 -498.325 ;
      RECT 13.285 -582.06 13.585 -498.325 ;
      RECT 13.27 -472.71 13.6 -472.38 ;
      RECT 13.285 -487.68 13.585 -472.38 ;
      RECT 13.27 -487.68 13.6 -487.35 ;
      RECT 13.285 -468.485 13.585 -424.72 ;
      RECT 13.27 -425.095 13.6 -424.765 ;
      RECT 13.27 -468.485 13.6 -468.155 ;
      RECT 11.005 -462.47 11.335 -462.14 ;
      RECT 11.02 -530.86 11.32 -462.14 ;
      RECT 11.005 -530.86 11.335 -530.53 ;
      RECT -5.91 -551.295 -5.58 -550.965 ;
      RECT -5.895 -570.73 -5.595 -550.965 ;
      RECT -5.91 -570.73 -5.58 -570.4 ;
      RECT -9.505 -570.285 -9.175 -569.955 ;
      RECT -9.49 -574.79 -9.19 -569.955 ;
      RECT -9.505 -574.745 -9.175 -574.415 ;
      RECT -10.34 -415.26 -10.01 -414.93 ;
      RECT -10.325 -532.65 -10.025 -414.93 ;
      RECT -10.34 -532.65 -10.01 -532.32 ;
      RECT -10.635 -571.085 -10.305 -570.755 ;
      RECT -10.62 -582.06 -10.32 -570.755 ;
      RECT -11.75 -556.06 -11.42 -555.73 ;
      RECT -11.735 -570.73 -11.435 -555.73 ;
      RECT -11.75 -570.73 -11.42 -570.4 ;
      RECT -12.385 -555.56 -12.055 -555.23 ;
      RECT -12.37 -571.485 -12.07 -555.23 ;
      RECT -12.385 -571.485 -12.055 -571.155 ;
      RECT -15.345 -570.285 -15.015 -569.955 ;
      RECT -15.33 -574.79 -15.03 -569.955 ;
      RECT -15.345 -574.745 -15.015 -574.415 ;
      RECT -16.475 -571.085 -16.145 -570.755 ;
      RECT -16.46 -582.06 -16.16 -570.755 ;
      RECT -17.59 -557.06 -17.26 -556.73 ;
      RECT -17.575 -570.73 -17.275 -556.73 ;
      RECT -17.59 -570.73 -17.26 -570.4 ;
      RECT -18.225 -556.56 -17.895 -556.23 ;
      RECT -18.21 -571.485 -17.91 -556.23 ;
      RECT -18.225 -571.485 -17.895 -571.155 ;
      RECT -21.185 -570.285 -20.855 -569.955 ;
      RECT -21.17 -574.79 -20.87 -569.955 ;
      RECT -21.185 -574.745 -20.855 -574.415 ;
      RECT -22.315 -571.085 -21.985 -570.755 ;
      RECT -22.3 -582.06 -22 -570.755 ;
      RECT -23.43 -558.06 -23.1 -557.73 ;
      RECT -23.415 -570.73 -23.115 -557.73 ;
      RECT -23.43 -570.73 -23.1 -570.4 ;
      RECT -24.065 -557.56 -23.735 -557.23 ;
      RECT -24.05 -571.485 -23.75 -557.23 ;
      RECT -24.065 -571.485 -23.735 -571.155 ;
      RECT -27.025 -570.285 -26.695 -569.955 ;
      RECT -27.01 -574.79 -26.71 -569.955 ;
      RECT -27.025 -574.745 -26.695 -574.415 ;
      RECT -28.155 -571.085 -27.825 -570.755 ;
      RECT -28.14 -582.06 -27.84 -570.755 ;
      RECT -29.27 -559.06 -28.94 -558.73 ;
      RECT -29.255 -570.73 -28.955 -558.73 ;
      RECT -29.27 -570.73 -28.94 -570.4 ;
      RECT -29.905 -558.56 -29.575 -558.23 ;
      RECT -29.89 -571.485 -29.59 -558.23 ;
      RECT -29.905 -571.485 -29.575 -571.155 ;
      RECT -32.865 -570.285 -32.535 -569.955 ;
      RECT -32.85 -574.79 -32.55 -569.955 ;
      RECT -32.865 -574.745 -32.535 -574.415 ;
      RECT -33.995 -571.085 -33.665 -570.755 ;
      RECT -33.98 -582.06 -33.68 -570.755 ;
      RECT -35.11 -560.06 -34.78 -559.73 ;
      RECT -35.095 -570.73 -34.795 -559.73 ;
      RECT -35.11 -570.73 -34.78 -570.4 ;
      RECT -35.745 -559.56 -35.415 -559.23 ;
      RECT -35.73 -571.485 -35.43 -559.23 ;
      RECT -35.745 -571.485 -35.415 -571.155 ;
      RECT -38.705 -570.285 -38.375 -569.955 ;
      RECT -38.69 -574.79 -38.39 -569.955 ;
      RECT -38.705 -574.745 -38.375 -574.415 ;
      RECT -39.835 -571.085 -39.505 -570.755 ;
      RECT -39.82 -582.06 -39.52 -570.755 ;
      RECT -40.95 -561.06 -40.62 -560.73 ;
      RECT -40.935 -570.73 -40.635 -560.73 ;
      RECT -40.95 -570.73 -40.62 -570.4 ;
      RECT -41.585 -560.56 -41.255 -560.23 ;
      RECT -41.57 -571.485 -41.27 -560.23 ;
      RECT -41.585 -571.485 -41.255 -571.155 ;
      RECT -44.545 -570.285 -44.215 -569.955 ;
      RECT -44.53 -574.79 -44.23 -569.955 ;
      RECT -44.545 -574.745 -44.215 -574.415 ;
      RECT -45.675 -571.085 -45.345 -570.755 ;
      RECT -45.66 -582.06 -45.36 -570.755 ;
      RECT -46.79 -562.06 -46.46 -561.73 ;
      RECT -46.775 -570.73 -46.475 -561.73 ;
      RECT -46.79 -570.73 -46.46 -570.4 ;
      RECT -47.425 -561.56 -47.095 -561.23 ;
      RECT -47.41 -571.485 -47.11 -561.23 ;
      RECT -47.425 -571.485 -47.095 -571.155 ;
      RECT -50.385 -570.285 -50.055 -569.955 ;
      RECT -50.37 -574.79 -50.07 -569.955 ;
      RECT -50.385 -574.745 -50.055 -574.415 ;
      RECT -51.515 -571.085 -51.185 -570.755 ;
      RECT -51.5 -582.06 -51.2 -570.755 ;
      RECT -52.63 -563.06 -52.3 -562.73 ;
      RECT -52.615 -570.73 -52.315 -562.73 ;
      RECT -52.63 -570.73 -52.3 -570.4 ;
      RECT -53.265 -562.56 -52.935 -562.23 ;
      RECT -53.25 -571.485 -52.95 -562.23 ;
      RECT -53.265 -571.485 -52.935 -571.155 ;
      RECT -56.225 -570.285 -55.895 -569.955 ;
      RECT -56.21 -574.79 -55.91 -569.955 ;
      RECT -56.225 -574.745 -55.895 -574.415 ;
      RECT -57.355 -571.085 -57.025 -570.755 ;
      RECT -57.34 -582.06 -57.04 -570.755 ;
      RECT -58.47 -564.06 -58.14 -563.73 ;
      RECT -58.455 -570.73 -58.155 -563.73 ;
      RECT -58.47 -570.73 -58.14 -570.4 ;
      RECT -59.105 -563.56 -58.775 -563.23 ;
      RECT -59.09 -571.485 -58.79 -563.23 ;
      RECT -59.105 -571.485 -58.775 -571.155 ;
      RECT -62.065 -570.285 -61.735 -569.955 ;
      RECT -62.05 -574.79 -61.75 -569.955 ;
      RECT -62.065 -574.745 -61.735 -574.415 ;
      RECT -63.195 -571.085 -62.865 -570.755 ;
      RECT -63.18 -582.06 -62.88 -570.755 ;
      RECT -64.31 -565.06 -63.98 -564.73 ;
      RECT -64.295 -570.73 -63.995 -564.73 ;
      RECT -64.31 -570.73 -63.98 -570.4 ;
      RECT -64.945 -564.56 -64.615 -564.23 ;
      RECT -64.93 -571.485 -64.63 -564.23 ;
      RECT -64.945 -571.485 -64.615 -571.155 ;
      RECT -67.905 -570.285 -67.575 -569.955 ;
      RECT -67.89 -574.79 -67.59 -569.955 ;
      RECT -67.905 -574.745 -67.575 -574.415 ;
      RECT -69.035 -571.085 -68.705 -570.755 ;
      RECT -69.02 -582.06 -68.72 -570.755 ;
      RECT -70.15 -566.06 -69.82 -565.73 ;
      RECT -70.135 -570.73 -69.835 -565.73 ;
      RECT -70.15 -570.73 -69.82 -570.4 ;
      RECT -70.785 -565.56 -70.455 -565.23 ;
      RECT -70.77 -571.485 -70.47 -565.23 ;
      RECT -70.785 -571.485 -70.455 -571.155 ;
      RECT -73.745 -570.285 -73.415 -569.955 ;
      RECT -73.73 -574.79 -73.43 -569.955 ;
      RECT -73.745 -574.745 -73.415 -574.415 ;
      RECT -74.875 -571.085 -74.545 -570.755 ;
      RECT -74.86 -582.06 -74.56 -570.755 ;
      RECT -75.74 -574.79 -75.34 -552.605 ;
      RECT -75.88 -581.94 -75.46 -574.37 ;
  END
END sramgen_sram_2048x32m8w8_replica_v1

END LIBRARY
