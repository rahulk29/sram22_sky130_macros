VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_1024x8m8w1
    CLASS BLOCK  ;
    FOREIGN sram22_1024x8m8w1   ;
    SIZE 293.000 BY 452.800 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.496400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 195.270 0.000 195.410 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.496400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 206.170 0.000 206.310 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.496400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 217.070 0.000 217.210 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.496400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 227.970 0.000 228.110 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.496400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 238.870 0.000 239.010 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.496400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 249.770 0.000 249.910 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.496400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 260.670 0.000 260.810 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.496400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 271.570 0.000 271.710 0.140 ; 
        END 
    END dout[7] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.220700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.218000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.850 0.000 194.990 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.220700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.218000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 205.750 0.000 205.890 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.220700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.218000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 216.650 0.000 216.790 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.220700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.218000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 227.550 0.000 227.690 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.220700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.218000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 238.450 0.000 238.590 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.220700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.218000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 249.350 0.000 249.490 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.220700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.218000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 260.250 0.000 260.390 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.220700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.218000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 271.150 0.000 271.290 0.140 ; 
        END 
    END din[7] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.031100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.500 0.000 194.640 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.031100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 205.400 0.000 205.540 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.031100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 216.300 0.000 216.440 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.031100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 227.200 0.000 227.340 0.140 ; 
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.031100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 238.100 0.000 238.240 0.140 ; 
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.031100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 249.000 0.000 249.140 0.140 ; 
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.031100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 259.900 0.000 260.040 0.140 ; 
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.031100 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 270.800 0.000 270.940 0.140 ; 
        END 
    END wmask[7] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 139.200 0.000 139.520 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 133.080 0.000 133.400 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 126.960 0.000 127.280 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 120.840 0.000 121.160 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 115.400 0.000 115.720 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 109.280 0.000 109.600 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 103.160 0.000 103.480 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 97.040 0.000 97.360 0.320 ; 
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 90.920 0.000 91.240 0.320 ; 
        END 
    END addr[8] 
    PIN addr[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 84.800 0.000 85.120 0.320 ; 
        END 
    END addr[9] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 151.440 0.000 151.760 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.768700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 145.320 0.000 145.640 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 10.602000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 154.840 0.000 155.160 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 14.508000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 155.520 0.000 155.840 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 194.600 6.240 ; 
                RECT 196.320 5.920 205.480 6.240 ; 
                RECT 207.200 5.920 216.360 6.240 ; 
                RECT 218.080 5.920 227.240 6.240 ; 
                RECT 228.960 5.920 238.120 6.240 ; 
                RECT 239.840 5.920 249.000 6.240 ; 
                RECT 250.720 5.920 259.880 6.240 ; 
                RECT 261.600 5.920 270.760 6.240 ; 
                RECT 272.480 5.920 292.840 6.240 ; 
                RECT 0.160 7.280 292.840 7.600 ; 
                RECT 0.160 8.640 292.840 8.960 ; 
                RECT 0.160 10.000 154.480 10.320 ; 
                RECT 188.160 10.000 292.840 10.320 ; 
                RECT 0.160 11.360 292.840 11.680 ; 
                RECT 0.160 12.720 80.360 13.040 ; 
                RECT 156.200 12.720 193.920 13.040 ; 
                RECT 271.800 12.720 292.840 13.040 ; 
                RECT 0.160 14.080 181.680 14.400 ; 
                RECT 283.360 14.080 292.840 14.400 ; 
                RECT 0.160 15.440 181.680 15.760 ; 
                RECT 283.360 15.440 292.840 15.760 ; 
                RECT 0.160 16.800 181.680 17.120 ; 
                RECT 283.360 16.800 292.840 17.120 ; 
                RECT 0.160 18.160 80.360 18.480 ; 
                RECT 155.520 18.160 181.680 18.480 ; 
                RECT 283.360 18.160 292.840 18.480 ; 
                RECT 0.160 19.520 181.680 19.840 ; 
                RECT 283.360 19.520 292.840 19.840 ; 
                RECT 0.160 20.880 181.680 21.200 ; 
                RECT 283.360 20.880 292.840 21.200 ; 
                RECT 0.160 22.240 181.680 22.560 ; 
                RECT 283.360 22.240 292.840 22.560 ; 
                RECT 0.160 23.600 181.680 23.920 ; 
                RECT 283.360 23.600 292.840 23.920 ; 
                RECT 0.160 24.960 181.680 25.280 ; 
                RECT 283.360 24.960 292.840 25.280 ; 
                RECT 0.160 26.320 181.680 26.640 ; 
                RECT 283.360 26.320 292.840 26.640 ; 
                RECT 0.160 27.680 181.680 28.000 ; 
                RECT 283.360 27.680 292.840 28.000 ; 
                RECT 0.160 29.040 181.680 29.360 ; 
                RECT 283.360 29.040 292.840 29.360 ; 
                RECT 0.160 30.400 181.000 30.720 ; 
                RECT 283.360 30.400 292.840 30.720 ; 
                RECT 0.160 31.760 181.680 32.080 ; 
                RECT 283.360 31.760 292.840 32.080 ; 
                RECT 0.160 33.120 181.680 33.440 ; 
                RECT 283.360 33.120 292.840 33.440 ; 
                RECT 0.160 34.480 115.040 34.800 ; 
                RECT 128.320 34.480 181.680 34.800 ; 
                RECT 283.360 34.480 292.840 34.800 ; 
                RECT 0.160 35.840 113.680 36.160 ; 
                RECT 134.440 35.840 181.680 36.160 ; 
                RECT 283.360 35.840 292.840 36.160 ; 
                RECT 0.160 37.200 112.320 37.520 ; 
                RECT 140.560 37.200 181.680 37.520 ; 
                RECT 283.360 37.200 292.840 37.520 ; 
                RECT 0.160 38.560 89.880 38.880 ; 
                RECT 155.520 38.560 181.680 38.880 ; 
                RECT 283.360 38.560 292.840 38.880 ; 
                RECT 0.160 39.920 90.560 40.240 ; 
                RECT 146.000 39.920 181.680 40.240 ; 
                RECT 283.360 39.920 292.840 40.240 ; 
                RECT 0.160 41.280 181.680 41.600 ; 
                RECT 283.360 41.280 292.840 41.600 ; 
                RECT 0.160 42.640 181.680 42.960 ; 
                RECT 283.360 42.640 292.840 42.960 ; 
                RECT 0.160 44.000 148.360 44.320 ; 
                RECT 154.160 44.000 181.680 44.320 ; 
                RECT 283.360 44.000 292.840 44.320 ; 
                RECT 0.160 45.360 148.360 45.680 ; 
                RECT 154.160 45.360 181.680 45.680 ; 
                RECT 283.360 45.360 292.840 45.680 ; 
                RECT 0.160 46.720 148.360 47.040 ; 
                RECT 283.360 46.720 292.840 47.040 ; 
                RECT 0.160 48.080 148.360 48.400 ; 
                RECT 283.360 48.080 292.840 48.400 ; 
                RECT 0.160 49.440 148.360 49.760 ; 
                RECT 154.160 49.440 181.680 49.760 ; 
                RECT 283.360 49.440 292.840 49.760 ; 
                RECT 0.160 50.800 181.680 51.120 ; 
                RECT 283.360 50.800 292.840 51.120 ; 
                RECT 0.160 52.160 181.680 52.480 ; 
                RECT 283.360 52.160 292.840 52.480 ; 
                RECT 0.160 53.520 181.680 53.840 ; 
                RECT 283.360 53.520 292.840 53.840 ; 
                RECT 0.160 54.880 181.680 55.200 ; 
                RECT 283.360 54.880 292.840 55.200 ; 
                RECT 0.160 56.240 111.640 56.560 ; 
                RECT 120.160 56.240 126.600 56.560 ; 
                RECT 153.480 56.240 181.680 56.560 ; 
                RECT 283.360 56.240 292.840 56.560 ; 
                RECT 0.160 57.600 113.000 57.920 ; 
                RECT 119.480 57.600 126.600 57.920 ; 
                RECT 163.000 57.600 181.680 57.920 ; 
                RECT 283.360 57.600 292.840 57.920 ; 
                RECT 0.160 58.960 114.360 59.280 ; 
                RECT 118.120 58.960 126.600 59.280 ; 
                RECT 163.000 58.960 181.680 59.280 ; 
                RECT 283.360 58.960 292.840 59.280 ; 
                RECT 0.160 60.320 126.600 60.640 ; 
                RECT 161.640 60.320 181.680 60.640 ; 
                RECT 283.360 60.320 292.840 60.640 ; 
                RECT 0.160 61.680 126.600 62.000 ; 
                RECT 163.000 61.680 181.680 62.000 ; 
                RECT 283.360 61.680 292.840 62.000 ; 
                RECT 0.160 63.040 126.600 63.360 ; 
                RECT 165.720 63.040 181.680 63.360 ; 
                RECT 283.360 63.040 292.840 63.360 ; 
                RECT 0.160 64.400 126.600 64.720 ; 
                RECT 153.480 64.400 181.680 64.720 ; 
                RECT 283.360 64.400 292.840 64.720 ; 
                RECT 0.160 65.760 126.600 66.080 ; 
                RECT 165.720 65.760 181.680 66.080 ; 
                RECT 283.360 65.760 292.840 66.080 ; 
                RECT 0.160 67.120 126.600 67.440 ; 
                RECT 164.360 67.120 181.680 67.440 ; 
                RECT 283.360 67.120 292.840 67.440 ; 
                RECT 0.160 68.480 126.600 68.800 ; 
                RECT 165.720 68.480 181.680 68.800 ; 
                RECT 283.360 68.480 292.840 68.800 ; 
                RECT 0.160 69.840 126.600 70.160 ; 
                RECT 168.440 69.840 181.680 70.160 ; 
                RECT 283.360 69.840 292.840 70.160 ; 
                RECT 0.160 71.200 126.600 71.520 ; 
                RECT 168.440 71.200 181.680 71.520 ; 
                RECT 283.360 71.200 292.840 71.520 ; 
                RECT 0.160 72.560 126.600 72.880 ; 
                RECT 167.080 72.560 181.680 72.880 ; 
                RECT 283.360 72.560 292.840 72.880 ; 
                RECT 0.160 73.920 126.600 74.240 ; 
                RECT 153.480 73.920 181.680 74.240 ; 
                RECT 283.360 73.920 292.840 74.240 ; 
                RECT 0.160 75.280 126.600 75.600 ; 
                RECT 167.080 75.280 181.680 75.600 ; 
                RECT 283.360 75.280 292.840 75.600 ; 
                RECT 0.160 76.640 126.600 76.960 ; 
                RECT 171.160 76.640 181.680 76.960 ; 
                RECT 283.360 76.640 292.840 76.960 ; 
                RECT 0.160 78.000 126.600 78.320 ; 
                RECT 171.160 78.000 181.680 78.320 ; 
                RECT 283.360 78.000 292.840 78.320 ; 
                RECT 0.160 79.360 126.600 79.680 ; 
                RECT 169.800 79.360 181.680 79.680 ; 
                RECT 283.360 79.360 292.840 79.680 ; 
                RECT 0.160 80.720 126.600 81.040 ; 
                RECT 171.160 80.720 181.680 81.040 ; 
                RECT 283.360 80.720 292.840 81.040 ; 
                RECT 0.160 82.080 87.840 82.400 ; 
                RECT 99.080 82.080 126.600 82.400 ; 
                RECT 153.480 82.080 181.680 82.400 ; 
                RECT 283.360 82.080 292.840 82.400 ; 
                RECT 0.160 83.440 89.200 83.760 ; 
                RECT 91.600 83.440 126.600 83.760 ; 
                RECT 173.880 83.440 181.680 83.760 ; 
                RECT 283.360 83.440 292.840 83.760 ; 
                RECT 0.160 84.800 90.560 85.120 ; 
                RECT 95.000 84.800 102.800 85.120 ; 
                RECT 105.200 84.800 126.600 85.120 ; 
                RECT 173.880 84.800 181.680 85.120 ; 
                RECT 283.360 84.800 292.840 85.120 ; 
                RECT 0.160 86.160 90.560 86.480 ; 
                RECT 94.320 86.160 126.600 86.480 ; 
                RECT 172.520 86.160 181.680 86.480 ; 
                RECT 283.360 86.160 292.840 86.480 ; 
                RECT 0.160 87.520 97.360 87.840 ; 
                RECT 105.880 87.520 126.600 87.840 ; 
                RECT 173.880 87.520 181.680 87.840 ; 
                RECT 283.360 87.520 292.840 87.840 ; 
                RECT 0.160 88.880 92.600 89.200 ; 
                RECT 99.080 88.880 126.600 89.200 ; 
                RECT 176.600 88.880 181.680 89.200 ; 
                RECT 283.360 88.880 292.840 89.200 ; 
                RECT 0.160 90.240 89.880 90.560 ; 
                RECT 99.080 90.240 126.600 90.560 ; 
                RECT 153.480 90.240 181.680 90.560 ; 
                RECT 283.360 90.240 292.840 90.560 ; 
                RECT 0.160 91.600 126.600 91.920 ; 
                RECT 176.600 91.600 181.680 91.920 ; 
                RECT 283.360 91.600 292.840 91.920 ; 
                RECT 0.160 92.960 87.160 93.280 ; 
                RECT 99.080 92.960 126.600 93.280 ; 
                RECT 175.240 92.960 181.680 93.280 ; 
                RECT 283.360 92.960 292.840 93.280 ; 
                RECT 0.160 94.320 97.360 94.640 ; 
                RECT 104.520 94.320 126.600 94.640 ; 
                RECT 176.600 94.320 181.680 94.640 ; 
                RECT 283.360 94.320 292.840 94.640 ; 
                RECT 0.160 95.680 96.000 96.000 ; 
                RECT 99.080 95.680 126.600 96.000 ; 
                RECT 179.320 95.680 181.680 96.000 ; 
                RECT 283.360 95.680 292.840 96.000 ; 
                RECT 0.160 97.040 126.600 97.360 ; 
                RECT 179.320 97.040 181.680 97.360 ; 
                RECT 283.360 97.040 292.840 97.360 ; 
                RECT 0.160 98.400 97.360 98.720 ; 
                RECT 105.200 98.400 126.600 98.720 ; 
                RECT 177.960 98.400 181.680 98.720 ; 
                RECT 283.360 98.400 292.840 98.720 ; 
                RECT 0.160 99.760 93.960 100.080 ; 
                RECT 99.080 99.760 126.600 100.080 ; 
                RECT 179.320 99.760 181.680 100.080 ; 
                RECT 283.360 99.760 292.840 100.080 ; 
                RECT 0.160 101.120 96.000 101.440 ; 
                RECT 99.080 101.120 126.600 101.440 ; 
                RECT 177.960 101.120 181.680 101.440 ; 
                RECT 283.360 101.120 292.840 101.440 ; 
                RECT 0.160 102.480 126.600 102.800 ; 
                RECT 283.360 102.480 292.840 102.800 ; 
                RECT 0.160 103.840 87.160 104.160 ; 
                RECT 109.960 103.840 126.600 104.160 ; 
                RECT 283.360 103.840 292.840 104.160 ; 
                RECT 0.160 105.200 104.160 105.520 ; 
                RECT 111.320 105.200 126.600 105.520 ; 
                RECT 283.360 105.200 292.840 105.520 ; 
                RECT 0.160 106.560 96.000 106.880 ; 
                RECT 99.080 106.560 108.240 106.880 ; 
                RECT 112.000 106.560 126.600 106.880 ; 
                RECT 283.360 106.560 292.840 106.880 ; 
                RECT 0.160 107.920 87.840 108.240 ; 
                RECT 101.800 107.920 126.600 108.240 ; 
                RECT 153.480 107.920 181.680 108.240 ; 
                RECT 283.360 107.920 292.840 108.240 ; 
                RECT 0.160 109.280 96.680 109.600 ; 
                RECT 105.200 109.280 181.680 109.600 ; 
                RECT 283.360 109.280 292.840 109.600 ; 
                RECT 0.160 110.640 93.960 110.960 ; 
                RECT 105.880 110.640 157.200 110.960 ; 
                RECT 283.360 110.640 292.840 110.960 ; 
                RECT 0.160 112.000 178.960 112.320 ; 
                RECT 283.360 112.000 292.840 112.320 ; 
                RECT 0.160 113.360 176.240 113.680 ; 
                RECT 283.360 113.360 292.840 113.680 ; 
                RECT 0.160 114.720 89.880 115.040 ; 
                RECT 99.080 114.720 173.520 115.040 ; 
                RECT 283.360 114.720 292.840 115.040 ; 
                RECT 0.160 116.080 89.880 116.400 ; 
                RECT 95.680 116.080 170.800 116.400 ; 
                RECT 283.360 116.080 292.840 116.400 ; 
                RECT 0.160 117.440 168.080 117.760 ; 
                RECT 283.360 117.440 292.840 117.760 ; 
                RECT 0.160 118.800 96.000 119.120 ; 
                RECT 98.400 118.800 165.360 119.120 ; 
                RECT 283.360 118.800 292.840 119.120 ; 
                RECT 0.160 120.160 89.200 120.480 ; 
                RECT 104.520 120.160 162.640 120.480 ; 
                RECT 283.360 120.160 292.840 120.480 ; 
                RECT 0.160 121.520 159.920 121.840 ; 
                RECT 283.360 121.520 292.840 121.840 ; 
                RECT 0.160 122.880 96.000 123.200 ; 
                RECT 98.400 122.880 181.680 123.200 ; 
                RECT 283.360 122.880 292.840 123.200 ; 
                RECT 0.160 124.240 91.240 124.560 ; 
                RECT 99.080 124.240 181.680 124.560 ; 
                RECT 283.360 124.240 292.840 124.560 ; 
                RECT 0.160 125.600 66.080 125.920 ; 
                RECT 84.800 125.600 87.840 125.920 ; 
                RECT 95.000 125.600 96.680 125.920 ; 
                RECT 99.080 125.600 181.680 125.920 ; 
                RECT 283.360 125.600 292.840 125.920 ; 
                RECT 0.160 126.960 66.080 127.280 ; 
                RECT 84.800 126.960 181.680 127.280 ; 
                RECT 283.360 126.960 292.840 127.280 ; 
                RECT 0.160 128.320 66.080 128.640 ; 
                RECT 84.800 128.320 87.160 128.640 ; 
                RECT 105.200 128.320 181.680 128.640 ; 
                RECT 283.360 128.320 292.840 128.640 ; 
                RECT 0.160 129.680 66.080 130.000 ; 
                RECT 97.720 129.680 181.680 130.000 ; 
                RECT 283.360 129.680 292.840 130.000 ; 
                RECT 0.160 131.040 66.080 131.360 ; 
                RECT 84.800 131.040 87.840 131.360 ; 
                RECT 101.800 131.040 181.680 131.360 ; 
                RECT 283.360 131.040 292.840 131.360 ; 
                RECT 0.160 132.400 66.080 132.720 ; 
                RECT 84.800 132.400 181.680 132.720 ; 
                RECT 283.360 132.400 292.840 132.720 ; 
                RECT 0.160 133.760 66.080 134.080 ; 
                RECT 84.800 133.760 181.680 134.080 ; 
                RECT 283.360 133.760 292.840 134.080 ; 
                RECT 0.160 135.120 66.080 135.440 ; 
                RECT 84.800 135.120 100.080 135.440 ; 
                RECT 105.880 135.120 181.680 135.440 ; 
                RECT 283.360 135.120 292.840 135.440 ; 
                RECT 0.160 136.480 66.080 136.800 ; 
                RECT 84.800 136.480 102.800 136.800 ; 
                RECT 105.200 136.480 181.680 136.800 ; 
                RECT 283.360 136.480 292.840 136.800 ; 
                RECT 0.160 137.840 66.080 138.160 ; 
                RECT 84.800 137.840 181.680 138.160 ; 
                RECT 283.360 137.840 292.840 138.160 ; 
                RECT 0.160 139.200 66.080 139.520 ; 
                RECT 84.800 139.200 89.880 139.520 ; 
                RECT 92.960 139.200 147.680 139.520 ; 
                RECT 153.480 139.200 181.680 139.520 ; 
                RECT 283.360 139.200 292.840 139.520 ; 
                RECT 0.160 140.560 66.080 140.880 ; 
                RECT 84.800 140.560 87.160 140.880 ; 
                RECT 91.600 140.560 147.680 140.880 ; 
                RECT 153.480 140.560 181.680 140.880 ; 
                RECT 283.360 140.560 292.840 140.880 ; 
                RECT 0.160 141.920 66.080 142.240 ; 
                RECT 84.800 141.920 147.680 142.240 ; 
                RECT 153.480 141.920 181.680 142.240 ; 
                RECT 283.360 141.920 292.840 142.240 ; 
                RECT 0.160 143.280 66.080 143.600 ; 
                RECT 85.480 143.280 147.680 143.600 ; 
                RECT 153.480 143.280 181.680 143.600 ; 
                RECT 283.360 143.280 292.840 143.600 ; 
                RECT 0.160 144.640 66.080 144.960 ; 
                RECT 84.800 144.640 147.680 144.960 ; 
                RECT 153.480 144.640 181.680 144.960 ; 
                RECT 283.360 144.640 292.840 144.960 ; 
                RECT 0.160 146.000 66.080 146.320 ; 
                RECT 84.800 146.000 181.680 146.320 ; 
                RECT 283.360 146.000 292.840 146.320 ; 
                RECT 0.160 147.360 66.080 147.680 ; 
                RECT 84.800 147.360 92.600 147.680 ; 
                RECT 105.200 147.360 181.680 147.680 ; 
                RECT 283.360 147.360 292.840 147.680 ; 
                RECT 0.160 148.720 66.080 149.040 ; 
                RECT 84.800 148.720 89.880 149.040 ; 
                RECT 94.320 148.720 161.280 149.040 ; 
                RECT 283.360 148.720 292.840 149.040 ; 
                RECT 0.160 150.080 66.080 150.400 ; 
                RECT 84.800 150.080 164.000 150.400 ; 
                RECT 283.360 150.080 292.840 150.400 ; 
                RECT 0.160 151.440 66.080 151.760 ; 
                RECT 84.800 151.440 132.720 151.760 ; 
                RECT 152.800 151.440 166.720 151.760 ; 
                RECT 283.360 151.440 292.840 151.760 ; 
                RECT 0.160 152.800 66.080 153.120 ; 
                RECT 84.800 152.800 132.720 153.120 ; 
                RECT 152.800 152.800 169.440 153.120 ; 
                RECT 283.360 152.800 292.840 153.120 ; 
                RECT 0.160 154.160 66.080 154.480 ; 
                RECT 84.800 154.160 92.600 154.480 ; 
                RECT 95.000 154.160 132.720 154.480 ; 
                RECT 152.800 154.160 172.160 154.480 ; 
                RECT 283.360 154.160 292.840 154.480 ; 
                RECT 0.160 155.520 66.080 155.840 ; 
                RECT 84.800 155.520 89.200 155.840 ; 
                RECT 92.280 155.520 102.800 155.840 ; 
                RECT 105.880 155.520 132.720 155.840 ; 
                RECT 152.800 155.520 174.880 155.840 ; 
                RECT 283.360 155.520 292.840 155.840 ; 
                RECT 0.160 156.880 66.080 157.200 ; 
                RECT 84.800 156.880 132.720 157.200 ; 
                RECT 152.800 156.880 177.600 157.200 ; 
                RECT 283.360 156.880 292.840 157.200 ; 
                RECT 0.160 158.240 66.080 158.560 ; 
                RECT 84.800 158.240 132.720 158.560 ; 
                RECT 283.360 158.240 292.840 158.560 ; 
                RECT 0.160 159.600 66.080 159.920 ; 
                RECT 84.800 159.600 132.720 159.920 ; 
                RECT 283.360 159.600 292.840 159.920 ; 
                RECT 0.160 160.960 66.080 161.280 ; 
                RECT 84.800 160.960 132.720 161.280 ; 
                RECT 152.800 160.960 181.680 161.280 ; 
                RECT 283.360 160.960 292.840 161.280 ; 
                RECT 0.160 162.320 66.080 162.640 ; 
                RECT 84.800 162.320 132.720 162.640 ; 
                RECT 152.800 162.320 181.680 162.640 ; 
                RECT 283.360 162.320 292.840 162.640 ; 
                RECT 0.160 163.680 66.080 164.000 ; 
                RECT 84.800 163.680 132.720 164.000 ; 
                RECT 152.800 163.680 181.680 164.000 ; 
                RECT 283.360 163.680 292.840 164.000 ; 
                RECT 0.160 165.040 91.240 165.360 ; 
                RECT 104.520 165.040 132.720 165.360 ; 
                RECT 152.800 165.040 181.680 165.360 ; 
                RECT 283.360 165.040 292.840 165.360 ; 
                RECT 0.160 166.400 132.720 166.720 ; 
                RECT 152.800 166.400 181.680 166.720 ; 
                RECT 283.360 166.400 292.840 166.720 ; 
                RECT 0.160 167.760 132.720 168.080 ; 
                RECT 152.800 167.760 181.680 168.080 ; 
                RECT 283.360 167.760 292.840 168.080 ; 
                RECT 0.160 169.120 45.000 169.440 ; 
                RECT 65.760 169.120 132.720 169.440 ; 
                RECT 152.800 169.120 181.680 169.440 ; 
                RECT 283.360 169.120 292.840 169.440 ; 
                RECT 0.160 170.480 45.000 170.800 ; 
                RECT 65.760 170.480 93.280 170.800 ; 
                RECT 99.080 170.480 132.720 170.800 ; 
                RECT 152.800 170.480 181.680 170.800 ; 
                RECT 283.360 170.480 292.840 170.800 ; 
                RECT 0.160 171.840 45.000 172.160 ; 
                RECT 65.760 171.840 72.200 172.160 ; 
                RECT 79.360 171.840 132.720 172.160 ; 
                RECT 152.800 171.840 181.680 172.160 ; 
                RECT 283.360 171.840 292.840 172.160 ; 
                RECT 0.160 173.200 45.000 173.520 ; 
                RECT 65.760 173.200 66.760 173.520 ; 
                RECT 84.120 173.200 132.720 173.520 ; 
                RECT 152.800 173.200 181.680 173.520 ; 
                RECT 283.360 173.200 292.840 173.520 ; 
                RECT 0.160 174.560 45.000 174.880 ; 
                RECT 65.760 174.560 132.720 174.880 ; 
                RECT 283.360 174.560 292.840 174.880 ; 
                RECT 0.160 175.920 32.760 176.240 ; 
                RECT 79.360 175.920 87.840 176.240 ; 
                RECT 97.720 175.920 132.720 176.240 ; 
                RECT 152.800 175.920 181.680 176.240 ; 
                RECT 283.360 175.920 292.840 176.240 ; 
                RECT 0.160 177.280 72.200 177.600 ; 
                RECT 92.280 177.280 292.840 177.600 ; 
                RECT 0.160 178.640 32.760 178.960 ; 
                RECT 91.600 178.640 292.840 178.960 ; 
                RECT 0.160 180.000 178.960 180.320 ; 
                RECT 286.080 180.000 292.840 180.320 ; 
                RECT 0.160 181.360 178.960 181.680 ; 
                RECT 286.080 181.360 292.840 181.680 ; 
                RECT 0.160 182.720 28.000 183.040 ; 
                RECT 34.480 182.720 99.400 183.040 ; 
                RECT 286.080 182.720 292.840 183.040 ; 
                RECT 0.160 184.080 25.960 184.400 ; 
                RECT 48.760 184.080 99.400 184.400 ; 
                RECT 286.080 184.080 292.840 184.400 ; 
                RECT 0.160 185.440 25.960 185.760 ; 
                RECT 48.080 185.440 59.960 185.760 ; 
                RECT 61.680 185.440 76.280 185.760 ; 
                RECT 90.240 185.440 99.400 185.760 ; 
                RECT 286.080 185.440 292.840 185.760 ; 
                RECT 0.160 186.800 59.960 187.120 ; 
                RECT 61.680 186.800 76.280 187.120 ; 
                RECT 90.240 186.800 99.400 187.120 ; 
                RECT 286.080 186.800 292.840 187.120 ; 
                RECT 0.160 188.160 25.960 188.480 ; 
                RECT 36.520 188.160 59.960 188.480 ; 
                RECT 64.400 188.160 76.280 188.480 ; 
                RECT 90.240 188.160 99.400 188.480 ; 
                RECT 286.080 188.160 292.840 188.480 ; 
                RECT 0.160 189.520 59.960 189.840 ; 
                RECT 65.080 189.520 76.280 189.840 ; 
                RECT 90.240 189.520 99.400 189.840 ; 
                RECT 286.080 189.520 292.840 189.840 ; 
                RECT 0.160 190.880 25.960 191.200 ; 
                RECT 36.520 190.880 59.960 191.200 ; 
                RECT 65.080 190.880 76.280 191.200 ; 
                RECT 90.240 190.880 99.400 191.200 ; 
                RECT 286.080 190.880 292.840 191.200 ; 
                RECT 0.160 192.240 25.960 192.560 ; 
                RECT 36.520 192.240 99.400 192.560 ; 
                RECT 286.080 192.240 292.840 192.560 ; 
                RECT 0.160 193.600 76.280 193.920 ; 
                RECT 90.240 193.600 99.400 193.920 ; 
                RECT 286.080 193.600 292.840 193.920 ; 
                RECT 0.160 194.960 76.280 195.280 ; 
                RECT 90.240 194.960 99.400 195.280 ; 
                RECT 286.080 194.960 292.840 195.280 ; 
                RECT 0.160 196.320 76.280 196.640 ; 
                RECT 90.240 196.320 99.400 196.640 ; 
                RECT 286.080 196.320 292.840 196.640 ; 
                RECT 0.160 197.680 19.160 198.000 ; 
                RECT 21.560 197.680 34.800 198.000 ; 
                RECT 37.200 197.680 76.280 198.000 ; 
                RECT 90.240 197.680 99.400 198.000 ; 
                RECT 286.080 197.680 292.840 198.000 ; 
                RECT 0.160 199.040 18.480 199.360 ; 
                RECT 21.560 199.040 38.880 199.360 ; 
                RECT 49.440 199.040 76.280 199.360 ; 
                RECT 83.440 199.040 99.400 199.360 ; 
                RECT 286.080 199.040 292.840 199.360 ; 
                RECT 0.160 200.400 17.800 200.720 ; 
                RECT 21.560 200.400 40.240 200.720 ; 
                RECT 48.080 200.400 84.440 200.720 ; 
                RECT 90.240 200.400 99.400 200.720 ; 
                RECT 286.080 200.400 292.840 200.720 ; 
                RECT 0.160 201.760 17.120 202.080 ; 
                RECT 21.560 201.760 59.960 202.080 ; 
                RECT 61.680 201.760 76.280 202.080 ; 
                RECT 90.240 201.760 99.400 202.080 ; 
                RECT 286.080 201.760 292.840 202.080 ; 
                RECT 0.160 203.120 59.960 203.440 ; 
                RECT 62.360 203.120 76.280 203.440 ; 
                RECT 90.240 203.120 99.400 203.440 ; 
                RECT 286.080 203.120 292.840 203.440 ; 
                RECT 0.160 204.480 16.440 204.800 ; 
                RECT 21.560 204.480 59.960 204.800 ; 
                RECT 63.040 204.480 76.280 204.800 ; 
                RECT 90.240 204.480 99.400 204.800 ; 
                RECT 286.080 204.480 292.840 204.800 ; 
                RECT 0.160 205.840 15.760 206.160 ; 
                RECT 21.560 205.840 59.960 206.160 ; 
                RECT 61.680 205.840 76.280 206.160 ; 
                RECT 90.240 205.840 99.400 206.160 ; 
                RECT 286.080 205.840 292.840 206.160 ; 
                RECT 0.160 207.200 59.960 207.520 ; 
                RECT 63.040 207.200 76.280 207.520 ; 
                RECT 84.800 207.200 99.400 207.520 ; 
                RECT 286.080 207.200 292.840 207.520 ; 
                RECT 0.160 208.560 15.080 208.880 ; 
                RECT 21.560 208.560 34.800 208.880 ; 
                RECT 41.280 208.560 76.280 208.880 ; 
                RECT 90.240 208.560 99.400 208.880 ; 
                RECT 286.080 208.560 292.840 208.880 ; 
                RECT 0.160 209.920 14.400 210.240 ; 
                RECT 21.560 209.920 34.800 210.240 ; 
                RECT 41.960 209.920 76.280 210.240 ; 
                RECT 90.240 209.920 99.400 210.240 ; 
                RECT 286.080 209.920 292.840 210.240 ; 
                RECT 0.160 211.280 76.280 211.600 ; 
                RECT 90.240 211.280 99.400 211.600 ; 
                RECT 286.080 211.280 292.840 211.600 ; 
                RECT 0.160 212.640 13.720 212.960 ; 
                RECT 21.560 212.640 34.800 212.960 ; 
                RECT 40.600 212.640 76.280 212.960 ; 
                RECT 90.240 212.640 99.400 212.960 ; 
                RECT 286.080 212.640 292.840 212.960 ; 
                RECT 0.160 214.000 13.040 214.320 ; 
                RECT 21.560 214.000 34.800 214.320 ; 
                RECT 39.920 214.000 76.280 214.320 ; 
                RECT 90.240 214.000 99.400 214.320 ; 
                RECT 286.080 214.000 292.840 214.320 ; 
                RECT 0.160 215.360 12.360 215.680 ; 
                RECT 21.560 215.360 99.400 215.680 ; 
                RECT 286.080 215.360 292.840 215.680 ; 
                RECT 0.160 216.720 11.680 217.040 ; 
                RECT 21.560 216.720 76.280 217.040 ; 
                RECT 90.240 216.720 99.400 217.040 ; 
                RECT 286.080 216.720 292.840 217.040 ; 
                RECT 0.160 218.080 76.280 218.400 ; 
                RECT 90.240 218.080 99.400 218.400 ; 
                RECT 286.080 218.080 292.840 218.400 ; 
                RECT 0.160 219.440 11.000 219.760 ; 
                RECT 21.560 219.440 76.280 219.760 ; 
                RECT 90.240 219.440 99.400 219.760 ; 
                RECT 286.080 219.440 292.840 219.760 ; 
                RECT 0.160 220.800 10.320 221.120 ; 
                RECT 21.560 220.800 76.280 221.120 ; 
                RECT 90.240 220.800 99.400 221.120 ; 
                RECT 286.080 220.800 292.840 221.120 ; 
                RECT 0.160 222.160 76.280 222.480 ; 
                RECT 90.240 222.160 99.400 222.480 ; 
                RECT 286.080 222.160 292.840 222.480 ; 
                RECT 0.160 223.520 99.400 223.840 ; 
                RECT 286.080 223.520 292.840 223.840 ; 
                RECT 0.160 224.880 76.280 225.200 ; 
                RECT 90.240 224.880 99.400 225.200 ; 
                RECT 286.080 224.880 292.840 225.200 ; 
                RECT 0.160 226.240 76.280 226.560 ; 
                RECT 90.240 226.240 99.400 226.560 ; 
                RECT 286.080 226.240 292.840 226.560 ; 
                RECT 0.160 227.600 76.280 227.920 ; 
                RECT 90.240 227.600 99.400 227.920 ; 
                RECT 286.080 227.600 292.840 227.920 ; 
                RECT 0.160 228.960 76.280 229.280 ; 
                RECT 90.240 228.960 99.400 229.280 ; 
                RECT 286.080 228.960 292.840 229.280 ; 
                RECT 0.160 230.320 76.280 230.640 ; 
                RECT 90.240 230.320 99.400 230.640 ; 
                RECT 286.080 230.320 292.840 230.640 ; 
                RECT 0.160 231.680 99.400 232.000 ; 
                RECT 286.080 231.680 292.840 232.000 ; 
                RECT 0.160 233.040 76.280 233.360 ; 
                RECT 90.240 233.040 99.400 233.360 ; 
                RECT 286.080 233.040 292.840 233.360 ; 
                RECT 0.160 234.400 76.280 234.720 ; 
                RECT 90.240 234.400 99.400 234.720 ; 
                RECT 286.080 234.400 292.840 234.720 ; 
                RECT 0.160 235.760 76.280 236.080 ; 
                RECT 90.240 235.760 99.400 236.080 ; 
                RECT 286.080 235.760 292.840 236.080 ; 
                RECT 0.160 237.120 76.280 237.440 ; 
                RECT 90.240 237.120 99.400 237.440 ; 
                RECT 286.080 237.120 292.840 237.440 ; 
                RECT 0.160 238.480 76.280 238.800 ; 
                RECT 88.200 238.480 99.400 238.800 ; 
                RECT 286.080 238.480 292.840 238.800 ; 
                RECT 0.160 239.840 86.480 240.160 ; 
                RECT 90.240 239.840 99.400 240.160 ; 
                RECT 286.080 239.840 292.840 240.160 ; 
                RECT 0.160 241.200 76.280 241.520 ; 
                RECT 90.240 241.200 99.400 241.520 ; 
                RECT 286.080 241.200 292.840 241.520 ; 
                RECT 0.160 242.560 76.280 242.880 ; 
                RECT 90.240 242.560 99.400 242.880 ; 
                RECT 286.080 242.560 292.840 242.880 ; 
                RECT 0.160 243.920 76.280 244.240 ; 
                RECT 90.240 243.920 99.400 244.240 ; 
                RECT 286.080 243.920 292.840 244.240 ; 
                RECT 0.160 245.280 76.280 245.600 ; 
                RECT 90.240 245.280 99.400 245.600 ; 
                RECT 286.080 245.280 292.840 245.600 ; 
                RECT 0.160 246.640 76.280 246.960 ; 
                RECT 89.560 246.640 99.400 246.960 ; 
                RECT 286.080 246.640 292.840 246.960 ; 
                RECT 0.160 248.000 80.360 248.320 ; 
                RECT 90.240 248.000 99.400 248.320 ; 
                RECT 286.080 248.000 292.840 248.320 ; 
                RECT 0.160 249.360 77.640 249.680 ; 
                RECT 90.240 249.360 99.400 249.680 ; 
                RECT 286.080 249.360 292.840 249.680 ; 
                RECT 0.160 250.720 77.640 251.040 ; 
                RECT 90.240 250.720 99.400 251.040 ; 
                RECT 286.080 250.720 292.840 251.040 ; 
                RECT 0.160 252.080 77.640 252.400 ; 
                RECT 90.240 252.080 99.400 252.400 ; 
                RECT 286.080 252.080 292.840 252.400 ; 
                RECT 0.160 253.440 77.640 253.760 ; 
                RECT 90.240 253.440 99.400 253.760 ; 
                RECT 286.080 253.440 292.840 253.760 ; 
                RECT 0.160 254.800 39.560 255.120 ; 
                RECT 65.760 254.800 99.400 255.120 ; 
                RECT 286.080 254.800 292.840 255.120 ; 
                RECT 0.160 256.160 38.200 256.480 ; 
                RECT 64.400 256.160 77.640 256.480 ; 
                RECT 90.240 256.160 99.400 256.480 ; 
                RECT 286.080 256.160 292.840 256.480 ; 
                RECT 0.160 257.520 36.840 257.840 ; 
                RECT 63.720 257.520 76.280 257.840 ; 
                RECT 90.240 257.520 99.400 257.840 ; 
                RECT 286.080 257.520 292.840 257.840 ; 
                RECT 0.160 258.880 76.280 259.200 ; 
                RECT 90.240 258.880 99.400 259.200 ; 
                RECT 286.080 258.880 292.840 259.200 ; 
                RECT 0.160 260.240 76.280 260.560 ; 
                RECT 90.240 260.240 99.400 260.560 ; 
                RECT 286.080 260.240 292.840 260.560 ; 
                RECT 0.160 261.600 76.280 261.920 ; 
                RECT 90.240 261.600 99.400 261.920 ; 
                RECT 286.080 261.600 292.840 261.920 ; 
                RECT 0.160 262.960 99.400 263.280 ; 
                RECT 286.080 262.960 292.840 263.280 ; 
                RECT 0.160 264.320 77.640 264.640 ; 
                RECT 90.240 264.320 99.400 264.640 ; 
                RECT 286.080 264.320 292.840 264.640 ; 
                RECT 0.160 265.680 76.280 266.000 ; 
                RECT 90.240 265.680 99.400 266.000 ; 
                RECT 286.080 265.680 292.840 266.000 ; 
                RECT 0.160 267.040 76.280 267.360 ; 
                RECT 90.240 267.040 99.400 267.360 ; 
                RECT 286.080 267.040 292.840 267.360 ; 
                RECT 0.160 268.400 76.280 268.720 ; 
                RECT 90.240 268.400 99.400 268.720 ; 
                RECT 286.080 268.400 292.840 268.720 ; 
                RECT 0.160 269.760 76.280 270.080 ; 
                RECT 90.240 269.760 99.400 270.080 ; 
                RECT 286.080 269.760 292.840 270.080 ; 
                RECT 0.160 271.120 99.400 271.440 ; 
                RECT 286.080 271.120 292.840 271.440 ; 
                RECT 0.160 272.480 76.280 272.800 ; 
                RECT 90.240 272.480 99.400 272.800 ; 
                RECT 286.080 272.480 292.840 272.800 ; 
                RECT 0.160 273.840 76.280 274.160 ; 
                RECT 90.240 273.840 99.400 274.160 ; 
                RECT 286.080 273.840 292.840 274.160 ; 
                RECT 0.160 275.200 76.280 275.520 ; 
                RECT 90.240 275.200 99.400 275.520 ; 
                RECT 286.080 275.200 292.840 275.520 ; 
                RECT 0.160 276.560 76.280 276.880 ; 
                RECT 90.240 276.560 99.400 276.880 ; 
                RECT 286.080 276.560 292.840 276.880 ; 
                RECT 0.160 277.920 76.280 278.240 ; 
                RECT 79.360 277.920 99.400 278.240 ; 
                RECT 286.080 277.920 292.840 278.240 ; 
                RECT 0.160 279.280 80.360 279.600 ; 
                RECT 90.240 279.280 99.400 279.600 ; 
                RECT 286.080 279.280 292.840 279.600 ; 
                RECT 0.160 280.640 76.280 280.960 ; 
                RECT 90.240 280.640 99.400 280.960 ; 
                RECT 286.080 280.640 292.840 280.960 ; 
                RECT 0.160 282.000 76.280 282.320 ; 
                RECT 90.240 282.000 99.400 282.320 ; 
                RECT 286.080 282.000 292.840 282.320 ; 
                RECT 0.160 283.360 78.320 283.680 ; 
                RECT 90.240 283.360 99.400 283.680 ; 
                RECT 286.080 283.360 292.840 283.680 ; 
                RECT 0.160 284.720 76.280 285.040 ; 
                RECT 90.240 284.720 99.400 285.040 ; 
                RECT 286.080 284.720 292.840 285.040 ; 
                RECT 0.160 286.080 76.280 286.400 ; 
                RECT 80.040 286.080 99.400 286.400 ; 
                RECT 286.080 286.080 292.840 286.400 ; 
                RECT 0.160 287.440 82.400 287.760 ; 
                RECT 90.240 287.440 99.400 287.760 ; 
                RECT 286.080 287.440 292.840 287.760 ; 
                RECT 0.160 288.800 76.280 289.120 ; 
                RECT 90.240 288.800 99.400 289.120 ; 
                RECT 286.080 288.800 292.840 289.120 ; 
                RECT 0.160 290.160 76.280 290.480 ; 
                RECT 90.240 290.160 99.400 290.480 ; 
                RECT 286.080 290.160 292.840 290.480 ; 
                RECT 0.160 291.520 76.280 291.840 ; 
                RECT 90.240 291.520 99.400 291.840 ; 
                RECT 286.080 291.520 292.840 291.840 ; 
                RECT 0.160 292.880 76.280 293.200 ; 
                RECT 90.240 292.880 99.400 293.200 ; 
                RECT 286.080 292.880 292.840 293.200 ; 
                RECT 0.160 294.240 99.400 294.560 ; 
                RECT 286.080 294.240 292.840 294.560 ; 
                RECT 0.160 295.600 78.320 295.920 ; 
                RECT 90.240 295.600 99.400 295.920 ; 
                RECT 286.080 295.600 292.840 295.920 ; 
                RECT 0.160 296.960 76.280 297.280 ; 
                RECT 90.240 296.960 99.400 297.280 ; 
                RECT 286.080 296.960 292.840 297.280 ; 
                RECT 0.160 298.320 76.280 298.640 ; 
                RECT 90.240 298.320 99.400 298.640 ; 
                RECT 286.080 298.320 292.840 298.640 ; 
                RECT 0.160 299.680 76.280 300.000 ; 
                RECT 90.240 299.680 99.400 300.000 ; 
                RECT 286.080 299.680 292.840 300.000 ; 
                RECT 0.160 301.040 76.280 301.360 ; 
                RECT 90.240 301.040 99.400 301.360 ; 
                RECT 286.080 301.040 292.840 301.360 ; 
                RECT 0.160 302.400 99.400 302.720 ; 
                RECT 286.080 302.400 292.840 302.720 ; 
                RECT 0.160 303.760 78.320 304.080 ; 
                RECT 90.240 303.760 99.400 304.080 ; 
                RECT 286.080 303.760 292.840 304.080 ; 
                RECT 0.160 305.120 76.280 305.440 ; 
                RECT 90.240 305.120 99.400 305.440 ; 
                RECT 286.080 305.120 292.840 305.440 ; 
                RECT 0.160 306.480 76.280 306.800 ; 
                RECT 90.240 306.480 99.400 306.800 ; 
                RECT 286.080 306.480 292.840 306.800 ; 
                RECT 0.160 307.840 76.280 308.160 ; 
                RECT 90.240 307.840 99.400 308.160 ; 
                RECT 286.080 307.840 292.840 308.160 ; 
                RECT 0.160 309.200 76.280 309.520 ; 
                RECT 90.240 309.200 99.400 309.520 ; 
                RECT 286.080 309.200 292.840 309.520 ; 
                RECT 0.160 310.560 99.400 310.880 ; 
                RECT 286.080 310.560 292.840 310.880 ; 
                RECT 0.160 311.920 76.280 312.240 ; 
                RECT 90.240 311.920 99.400 312.240 ; 
                RECT 286.080 311.920 292.840 312.240 ; 
                RECT 0.160 313.280 76.280 313.600 ; 
                RECT 90.240 313.280 99.400 313.600 ; 
                RECT 286.080 313.280 292.840 313.600 ; 
                RECT 0.160 314.640 76.280 314.960 ; 
                RECT 90.240 314.640 99.400 314.960 ; 
                RECT 286.080 314.640 292.840 314.960 ; 
                RECT 0.160 316.000 76.280 316.320 ; 
                RECT 90.240 316.000 99.400 316.320 ; 
                RECT 286.080 316.000 292.840 316.320 ; 
                RECT 0.160 317.360 76.280 317.680 ; 
                RECT 82.080 317.360 99.400 317.680 ; 
                RECT 286.080 317.360 292.840 317.680 ; 
                RECT 0.160 318.720 99.400 319.040 ; 
                RECT 286.080 318.720 292.840 319.040 ; 
                RECT 0.160 320.080 78.320 320.400 ; 
                RECT 90.240 320.080 99.400 320.400 ; 
                RECT 286.080 320.080 292.840 320.400 ; 
                RECT 0.160 321.440 78.320 321.760 ; 
                RECT 90.240 321.440 99.400 321.760 ; 
                RECT 286.080 321.440 292.840 321.760 ; 
                RECT 0.160 322.800 78.320 323.120 ; 
                RECT 90.240 322.800 99.400 323.120 ; 
                RECT 286.080 322.800 292.840 323.120 ; 
                RECT 0.160 324.160 78.320 324.480 ; 
                RECT 90.240 324.160 99.400 324.480 ; 
                RECT 286.080 324.160 292.840 324.480 ; 
                RECT 0.160 325.520 99.400 325.840 ; 
                RECT 286.080 325.520 292.840 325.840 ; 
                RECT 0.160 326.880 84.440 327.200 ; 
                RECT 90.240 326.880 99.400 327.200 ; 
                RECT 286.080 326.880 292.840 327.200 ; 
                RECT 0.160 328.240 78.320 328.560 ; 
                RECT 90.240 328.240 99.400 328.560 ; 
                RECT 286.080 328.240 292.840 328.560 ; 
                RECT 0.160 329.600 78.320 329.920 ; 
                RECT 90.240 329.600 99.400 329.920 ; 
                RECT 286.080 329.600 292.840 329.920 ; 
                RECT 0.160 330.960 78.320 331.280 ; 
                RECT 90.240 330.960 99.400 331.280 ; 
                RECT 286.080 330.960 292.840 331.280 ; 
                RECT 0.160 332.320 78.320 332.640 ; 
                RECT 90.240 332.320 99.400 332.640 ; 
                RECT 286.080 332.320 292.840 332.640 ; 
                RECT 0.160 333.680 99.400 334.000 ; 
                RECT 286.080 333.680 292.840 334.000 ; 
                RECT 0.160 335.040 78.320 335.360 ; 
                RECT 90.240 335.040 99.400 335.360 ; 
                RECT 286.080 335.040 292.840 335.360 ; 
                RECT 0.160 336.400 86.480 336.720 ; 
                RECT 90.240 336.400 99.400 336.720 ; 
                RECT 286.080 336.400 292.840 336.720 ; 
                RECT 0.160 337.760 78.320 338.080 ; 
                RECT 90.240 337.760 99.400 338.080 ; 
                RECT 286.080 337.760 292.840 338.080 ; 
                RECT 0.160 339.120 78.320 339.440 ; 
                RECT 90.240 339.120 99.400 339.440 ; 
                RECT 286.080 339.120 292.840 339.440 ; 
                RECT 0.160 340.480 78.320 340.800 ; 
                RECT 90.240 340.480 99.400 340.800 ; 
                RECT 286.080 340.480 292.840 340.800 ; 
                RECT 0.160 341.840 99.400 342.160 ; 
                RECT 286.080 341.840 292.840 342.160 ; 
                RECT 0.160 343.200 79.000 343.520 ; 
                RECT 90.240 343.200 99.400 343.520 ; 
                RECT 286.080 343.200 292.840 343.520 ; 
                RECT 0.160 344.560 79.000 344.880 ; 
                RECT 90.240 344.560 99.400 344.880 ; 
                RECT 286.080 344.560 292.840 344.880 ; 
                RECT 0.160 345.920 81.720 346.240 ; 
                RECT 90.240 345.920 99.400 346.240 ; 
                RECT 286.080 345.920 292.840 346.240 ; 
                RECT 0.160 347.280 79.000 347.600 ; 
                RECT 90.240 347.280 99.400 347.600 ; 
                RECT 286.080 347.280 292.840 347.600 ; 
                RECT 0.160 348.640 79.000 348.960 ; 
                RECT 90.240 348.640 99.400 348.960 ; 
                RECT 286.080 348.640 292.840 348.960 ; 
                RECT 0.160 350.000 99.400 350.320 ; 
                RECT 286.080 350.000 292.840 350.320 ; 
                RECT 0.160 351.360 79.000 351.680 ; 
                RECT 90.240 351.360 99.400 351.680 ; 
                RECT 286.080 351.360 292.840 351.680 ; 
                RECT 0.160 352.720 79.000 353.040 ; 
                RECT 90.240 352.720 99.400 353.040 ; 
                RECT 286.080 352.720 292.840 353.040 ; 
                RECT 0.160 354.080 79.000 354.400 ; 
                RECT 90.240 354.080 99.400 354.400 ; 
                RECT 286.080 354.080 292.840 354.400 ; 
                RECT 0.160 355.440 83.760 355.760 ; 
                RECT 90.240 355.440 99.400 355.760 ; 
                RECT 286.080 355.440 292.840 355.760 ; 
                RECT 0.160 356.800 79.000 357.120 ; 
                RECT 90.240 356.800 99.400 357.120 ; 
                RECT 286.080 356.800 292.840 357.120 ; 
                RECT 0.160 358.160 99.400 358.480 ; 
                RECT 286.080 358.160 292.840 358.480 ; 
                RECT 0.160 359.520 79.000 359.840 ; 
                RECT 90.240 359.520 99.400 359.840 ; 
                RECT 286.080 359.520 292.840 359.840 ; 
                RECT 0.160 360.880 79.000 361.200 ; 
                RECT 90.240 360.880 99.400 361.200 ; 
                RECT 286.080 360.880 292.840 361.200 ; 
                RECT 0.160 362.240 79.000 362.560 ; 
                RECT 90.240 362.240 99.400 362.560 ; 
                RECT 286.080 362.240 292.840 362.560 ; 
                RECT 0.160 363.600 79.000 363.920 ; 
                RECT 90.240 363.600 99.400 363.920 ; 
                RECT 286.080 363.600 292.840 363.920 ; 
                RECT 0.160 364.960 99.400 365.280 ; 
                RECT 286.080 364.960 292.840 365.280 ; 
                RECT 0.160 366.320 86.480 366.640 ; 
                RECT 90.240 366.320 99.400 366.640 ; 
                RECT 286.080 366.320 292.840 366.640 ; 
                RECT 0.160 367.680 79.000 368.000 ; 
                RECT 90.240 367.680 99.400 368.000 ; 
                RECT 286.080 367.680 292.840 368.000 ; 
                RECT 0.160 369.040 79.000 369.360 ; 
                RECT 90.240 369.040 99.400 369.360 ; 
                RECT 286.080 369.040 292.840 369.360 ; 
                RECT 0.160 370.400 79.000 370.720 ; 
                RECT 90.240 370.400 99.400 370.720 ; 
                RECT 286.080 370.400 292.840 370.720 ; 
                RECT 0.160 371.760 79.000 372.080 ; 
                RECT 90.240 371.760 99.400 372.080 ; 
                RECT 286.080 371.760 292.840 372.080 ; 
                RECT 0.160 373.120 99.400 373.440 ; 
                RECT 286.080 373.120 292.840 373.440 ; 
                RECT 0.160 374.480 80.360 374.800 ; 
                RECT 90.240 374.480 99.400 374.800 ; 
                RECT 286.080 374.480 292.840 374.800 ; 
                RECT 0.160 375.840 81.040 376.160 ; 
                RECT 90.240 375.840 99.400 376.160 ; 
                RECT 286.080 375.840 292.840 376.160 ; 
                RECT 0.160 377.200 79.680 377.520 ; 
                RECT 90.240 377.200 99.400 377.520 ; 
                RECT 286.080 377.200 292.840 377.520 ; 
                RECT 0.160 378.560 79.680 378.880 ; 
                RECT 90.240 378.560 99.400 378.880 ; 
                RECT 286.080 378.560 292.840 378.880 ; 
                RECT 0.160 379.920 79.680 380.240 ; 
                RECT 90.240 379.920 99.400 380.240 ; 
                RECT 286.080 379.920 292.840 380.240 ; 
                RECT 0.160 381.280 99.400 381.600 ; 
                RECT 286.080 381.280 292.840 381.600 ; 
                RECT 0.160 382.640 79.680 382.960 ; 
                RECT 90.240 382.640 99.400 382.960 ; 
                RECT 286.080 382.640 292.840 382.960 ; 
                RECT 0.160 384.000 79.680 384.320 ; 
                RECT 90.240 384.000 99.400 384.320 ; 
                RECT 286.080 384.000 292.840 384.320 ; 
                RECT 0.160 385.360 83.080 385.680 ; 
                RECT 90.240 385.360 99.400 385.680 ; 
                RECT 286.080 385.360 292.840 385.680 ; 
                RECT 0.160 386.720 79.680 387.040 ; 
                RECT 90.240 386.720 99.400 387.040 ; 
                RECT 286.080 386.720 292.840 387.040 ; 
                RECT 0.160 388.080 79.680 388.400 ; 
                RECT 90.240 388.080 99.400 388.400 ; 
                RECT 286.080 388.080 292.840 388.400 ; 
                RECT 0.160 389.440 99.400 389.760 ; 
                RECT 286.080 389.440 292.840 389.760 ; 
                RECT 0.160 390.800 79.680 391.120 ; 
                RECT 90.240 390.800 99.400 391.120 ; 
                RECT 286.080 390.800 292.840 391.120 ; 
                RECT 0.160 392.160 79.680 392.480 ; 
                RECT 90.240 392.160 99.400 392.480 ; 
                RECT 286.080 392.160 292.840 392.480 ; 
                RECT 0.160 393.520 79.680 393.840 ; 
                RECT 90.240 393.520 99.400 393.840 ; 
                RECT 286.080 393.520 292.840 393.840 ; 
                RECT 0.160 394.880 85.800 395.200 ; 
                RECT 90.240 394.880 99.400 395.200 ; 
                RECT 286.080 394.880 292.840 395.200 ; 
                RECT 0.160 396.240 79.680 396.560 ; 
                RECT 90.240 396.240 99.400 396.560 ; 
                RECT 286.080 396.240 292.840 396.560 ; 
                RECT 0.160 397.600 99.400 397.920 ; 
                RECT 286.080 397.600 292.840 397.920 ; 
                RECT 0.160 398.960 79.680 399.280 ; 
                RECT 90.240 398.960 99.400 399.280 ; 
                RECT 286.080 398.960 292.840 399.280 ; 
                RECT 0.160 400.320 79.680 400.640 ; 
                RECT 90.240 400.320 99.400 400.640 ; 
                RECT 286.080 400.320 292.840 400.640 ; 
                RECT 0.160 401.680 79.680 402.000 ; 
                RECT 90.240 401.680 99.400 402.000 ; 
                RECT 286.080 401.680 292.840 402.000 ; 
                RECT 0.160 403.040 79.680 403.360 ; 
                RECT 90.240 403.040 99.400 403.360 ; 
                RECT 286.080 403.040 292.840 403.360 ; 
                RECT 0.160 404.400 99.400 404.720 ; 
                RECT 286.080 404.400 292.840 404.720 ; 
                RECT 0.160 405.760 80.360 406.080 ; 
                RECT 90.240 405.760 99.400 406.080 ; 
                RECT 286.080 405.760 292.840 406.080 ; 
                RECT 0.160 407.120 80.360 407.440 ; 
                RECT 90.240 407.120 99.400 407.440 ; 
                RECT 286.080 407.120 292.840 407.440 ; 
                RECT 0.160 408.480 80.360 408.800 ; 
                RECT 90.240 408.480 99.400 408.800 ; 
                RECT 286.080 408.480 292.840 408.800 ; 
                RECT 0.160 409.840 80.360 410.160 ; 
                RECT 90.240 409.840 99.400 410.160 ; 
                RECT 286.080 409.840 292.840 410.160 ; 
                RECT 0.160 411.200 80.360 411.520 ; 
                RECT 90.240 411.200 99.400 411.520 ; 
                RECT 286.080 411.200 292.840 411.520 ; 
                RECT 0.160 412.560 99.400 412.880 ; 
                RECT 286.080 412.560 292.840 412.880 ; 
                RECT 0.160 413.920 82.400 414.240 ; 
                RECT 90.240 413.920 99.400 414.240 ; 
                RECT 286.080 413.920 292.840 414.240 ; 
                RECT 0.160 415.280 80.360 415.600 ; 
                RECT 90.240 415.280 99.400 415.600 ; 
                RECT 286.080 415.280 292.840 415.600 ; 
                RECT 0.160 416.640 80.360 416.960 ; 
                RECT 90.240 416.640 99.400 416.960 ; 
                RECT 286.080 416.640 292.840 416.960 ; 
                RECT 0.160 418.000 80.360 418.320 ; 
                RECT 90.240 418.000 99.400 418.320 ; 
                RECT 286.080 418.000 292.840 418.320 ; 
                RECT 0.160 419.360 80.360 419.680 ; 
                RECT 90.240 419.360 99.400 419.680 ; 
                RECT 286.080 419.360 292.840 419.680 ; 
                RECT 0.160 420.720 99.400 421.040 ; 
                RECT 286.080 420.720 292.840 421.040 ; 
                RECT 0.160 422.080 80.360 422.400 ; 
                RECT 90.240 422.080 99.400 422.400 ; 
                RECT 286.080 422.080 292.840 422.400 ; 
                RECT 0.160 423.440 85.120 423.760 ; 
                RECT 90.240 423.440 99.400 423.760 ; 
                RECT 286.080 423.440 292.840 423.760 ; 
                RECT 0.160 424.800 85.120 425.120 ; 
                RECT 90.240 424.800 99.400 425.120 ; 
                RECT 286.080 424.800 292.840 425.120 ; 
                RECT 0.160 426.160 80.360 426.480 ; 
                RECT 90.240 426.160 99.400 426.480 ; 
                RECT 286.080 426.160 292.840 426.480 ; 
                RECT 0.160 427.520 80.360 427.840 ; 
                RECT 90.240 427.520 99.400 427.840 ; 
                RECT 286.080 427.520 292.840 427.840 ; 
                RECT 0.160 428.880 99.400 429.200 ; 
                RECT 286.080 428.880 292.840 429.200 ; 
                RECT 0.160 430.240 80.360 430.560 ; 
                RECT 90.240 430.240 99.400 430.560 ; 
                RECT 286.080 430.240 292.840 430.560 ; 
                RECT 0.160 431.600 80.360 431.920 ; 
                RECT 90.240 431.600 99.400 431.920 ; 
                RECT 286.080 431.600 292.840 431.920 ; 
                RECT 0.160 432.960 87.160 433.280 ; 
                RECT 90.240 432.960 99.400 433.280 ; 
                RECT 286.080 432.960 292.840 433.280 ; 
                RECT 0.160 434.320 87.840 434.640 ; 
                RECT 90.240 434.320 99.400 434.640 ; 
                RECT 286.080 434.320 292.840 434.640 ; 
                RECT 0.160 435.680 80.360 436.000 ; 
                RECT 90.240 435.680 99.400 436.000 ; 
                RECT 286.080 435.680 292.840 436.000 ; 
                RECT 0.160 437.040 99.400 437.360 ; 
                RECT 286.080 437.040 292.840 437.360 ; 
                RECT 0.160 438.400 178.960 438.720 ; 
                RECT 286.080 438.400 292.840 438.720 ; 
                RECT 0.160 439.760 178.960 440.080 ; 
                RECT 286.080 439.760 292.840 440.080 ; 
                RECT 0.160 441.120 178.960 441.440 ; 
                RECT 286.080 441.120 292.840 441.440 ; 
                RECT 0.160 442.480 292.840 442.800 ; 
                RECT 0.160 443.840 292.840 444.160 ; 
                RECT 0.160 445.200 292.840 445.520 ; 
                RECT 0.160 446.560 292.840 446.880 ; 
                RECT 0.160 0.160 292.840 1.520 ; 
                RECT 0.160 451.280 292.840 452.640 ; 
                RECT 183.100 35.005 188.900 36.375 ; 
                RECT 275.800 35.005 281.600 36.375 ; 
                RECT 183.100 39.720 188.900 40.840 ; 
                RECT 275.800 39.720 281.600 40.840 ; 
                RECT 183.100 44.945 188.900 46.745 ; 
                RECT 275.800 44.945 281.600 46.745 ; 
                RECT 183.100 51.185 188.900 52.985 ; 
                RECT 275.800 51.185 281.600 52.985 ; 
                RECT 183.100 79.260 281.600 80.060 ; 
                RECT 183.100 166.545 281.600 170.145 ; 
                RECT 183.100 129.205 281.600 131.005 ; 
                RECT 183.100 97.165 281.600 97.455 ; 
                RECT 183.100 74.370 281.600 75.170 ; 
                RECT 183.100 59.890 281.600 61.690 ; 
                RECT 183.100 89.785 281.600 93.385 ; 
                RECT 183.100 71.360 281.600 72.160 ; 
                RECT 183.100 19.250 281.600 21.050 ; 
                RECT 103.750 183.115 105.670 437.495 ; 
                RECT 113.320 183.115 115.240 437.495 ; 
                RECT 117.160 183.115 119.080 437.495 ; 
                RECT 129.985 183.115 131.905 437.495 ; 
                RECT 133.825 183.115 135.745 437.495 ; 
                RECT 137.665 183.115 139.585 437.495 ; 
                RECT 155.280 183.115 157.200 437.495 ; 
                RECT 159.120 183.115 161.040 437.495 ; 
                RECT 162.960 183.115 164.880 437.495 ; 
                RECT 166.800 183.115 168.720 437.495 ; 
                RECT 170.640 183.115 172.560 437.495 ; 
                RECT 174.480 183.115 176.400 437.495 ; 
                RECT 130.600 55.565 132.520 108.165 ; 
                RECT 137.575 55.565 139.495 108.165 ; 
                RECT 146.930 55.565 148.850 108.165 ; 
                RECT 150.770 55.565 152.690 108.165 ; 
                RECT 135.715 150.940 137.255 176.480 ; 
                RECT 141.725 150.940 143.475 176.480 ; 
                RECT 150.120 150.940 152.040 176.480 ; 
                RECT 151.195 139.780 153.115 144.940 ; 
                RECT 151.495 44.405 153.245 49.565 ; 
                RECT 26.500 185.385 35.660 186.135 ; 
                RECT 26.500 190.785 35.660 192.705 ; 
                RECT 67.340 173.095 83.380 173.945 ; 
                RECT 45.740 172.795 65.380 175.505 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 194.600 5.560 ; 
                RECT 196.320 5.240 205.480 5.560 ; 
                RECT 207.200 5.240 216.360 5.560 ; 
                RECT 218.080 5.240 227.240 5.560 ; 
                RECT 228.960 5.240 238.120 5.560 ; 
                RECT 239.840 5.240 249.000 5.560 ; 
                RECT 250.720 5.240 259.880 5.560 ; 
                RECT 261.600 5.240 270.760 5.560 ; 
                RECT 272.480 5.240 290.120 5.560 ; 
                RECT 2.880 6.600 290.120 6.920 ; 
                RECT 2.880 7.960 290.120 8.280 ; 
                RECT 2.880 9.320 155.160 9.640 ; 
                RECT 187.480 9.320 290.120 9.640 ; 
                RECT 2.880 10.680 290.120 11.000 ; 
                RECT 2.880 12.040 290.120 12.360 ; 
                RECT 2.880 13.400 80.360 13.720 ; 
                RECT 156.200 13.400 181.680 13.720 ; 
                RECT 283.360 13.400 290.120 13.720 ; 
                RECT 2.880 14.760 181.680 15.080 ; 
                RECT 283.360 14.760 290.120 15.080 ; 
                RECT 2.880 16.120 181.680 16.440 ; 
                RECT 283.360 16.120 290.120 16.440 ; 
                RECT 2.880 17.480 80.360 17.800 ; 
                RECT 155.520 17.480 181.680 17.800 ; 
                RECT 283.360 17.480 290.120 17.800 ; 
                RECT 2.880 18.840 181.680 19.160 ; 
                RECT 283.360 18.840 290.120 19.160 ; 
                RECT 2.880 20.200 181.680 20.520 ; 
                RECT 283.360 20.200 290.120 20.520 ; 
                RECT 2.880 21.560 181.680 21.880 ; 
                RECT 283.360 21.560 290.120 21.880 ; 
                RECT 2.880 22.920 181.680 23.240 ; 
                RECT 283.360 22.920 290.120 23.240 ; 
                RECT 2.880 24.280 181.680 24.600 ; 
                RECT 283.360 24.280 290.120 24.600 ; 
                RECT 2.880 25.640 181.680 25.960 ; 
                RECT 283.360 25.640 290.120 25.960 ; 
                RECT 2.880 27.000 181.680 27.320 ; 
                RECT 283.360 27.000 290.120 27.320 ; 
                RECT 2.880 28.360 181.680 28.680 ; 
                RECT 283.360 28.360 290.120 28.680 ; 
                RECT 2.880 29.720 181.680 30.040 ; 
                RECT 283.360 29.720 290.120 30.040 ; 
                RECT 2.880 31.080 181.000 31.400 ; 
                RECT 283.360 31.080 290.120 31.400 ; 
                RECT 2.880 32.440 181.680 32.760 ; 
                RECT 283.360 32.440 290.120 32.760 ; 
                RECT 2.880 33.800 181.680 34.120 ; 
                RECT 283.360 33.800 290.120 34.120 ; 
                RECT 2.880 35.160 114.360 35.480 ; 
                RECT 126.960 35.160 181.680 35.480 ; 
                RECT 283.360 35.160 290.120 35.480 ; 
                RECT 2.880 36.520 113.000 36.840 ; 
                RECT 133.080 36.520 181.680 36.840 ; 
                RECT 283.360 36.520 290.120 36.840 ; 
                RECT 2.880 37.880 111.640 38.200 ; 
                RECT 139.200 37.880 181.680 38.200 ; 
                RECT 283.360 37.880 290.120 38.200 ; 
                RECT 2.880 39.240 92.600 39.560 ; 
                RECT 156.200 39.240 181.680 39.560 ; 
                RECT 283.360 39.240 290.120 39.560 ; 
                RECT 2.880 40.600 91.240 40.920 ; 
                RECT 152.120 40.600 181.680 40.920 ; 
                RECT 283.360 40.600 290.120 40.920 ; 
                RECT 2.880 41.960 181.680 42.280 ; 
                RECT 283.360 41.960 290.120 42.280 ; 
                RECT 2.880 43.320 181.680 43.640 ; 
                RECT 283.360 43.320 290.120 43.640 ; 
                RECT 2.880 44.680 148.360 45.000 ; 
                RECT 154.160 44.680 181.680 45.000 ; 
                RECT 283.360 44.680 290.120 45.000 ; 
                RECT 2.880 46.040 148.360 46.360 ; 
                RECT 283.360 46.040 290.120 46.360 ; 
                RECT 2.880 47.400 148.360 47.720 ; 
                RECT 283.360 47.400 290.120 47.720 ; 
                RECT 2.880 48.760 110.280 49.080 ; 
                RECT 145.320 48.760 148.360 49.080 ; 
                RECT 154.160 48.760 181.680 49.080 ; 
                RECT 283.360 48.760 290.120 49.080 ; 
                RECT 2.880 50.120 181.680 50.440 ; 
                RECT 283.360 50.120 290.120 50.440 ; 
                RECT 2.880 51.480 181.680 51.800 ; 
                RECT 283.360 51.480 290.120 51.800 ; 
                RECT 2.880 52.840 181.680 53.160 ; 
                RECT 283.360 52.840 290.120 53.160 ; 
                RECT 2.880 54.200 181.680 54.520 ; 
                RECT 283.360 54.200 290.120 54.520 ; 
                RECT 2.880 55.560 126.600 55.880 ; 
                RECT 153.480 55.560 181.680 55.880 ; 
                RECT 283.360 55.560 290.120 55.880 ; 
                RECT 2.880 56.920 112.320 57.240 ; 
                RECT 119.480 56.920 126.600 57.240 ; 
                RECT 163.000 56.920 181.680 57.240 ; 
                RECT 283.360 56.920 290.120 57.240 ; 
                RECT 2.880 58.280 113.680 58.600 ; 
                RECT 118.800 58.280 126.600 58.600 ; 
                RECT 161.640 58.280 181.680 58.600 ; 
                RECT 283.360 58.280 290.120 58.600 ; 
                RECT 2.880 59.640 115.040 59.960 ; 
                RECT 118.120 59.640 126.600 59.960 ; 
                RECT 163.000 59.640 181.680 59.960 ; 
                RECT 283.360 59.640 290.120 59.960 ; 
                RECT 2.880 61.000 126.600 61.320 ; 
                RECT 163.000 61.000 181.680 61.320 ; 
                RECT 283.360 61.000 290.120 61.320 ; 
                RECT 2.880 62.360 126.600 62.680 ; 
                RECT 161.640 62.360 181.680 62.680 ; 
                RECT 283.360 62.360 290.120 62.680 ; 
                RECT 2.880 63.720 126.600 64.040 ; 
                RECT 165.720 63.720 181.680 64.040 ; 
                RECT 283.360 63.720 290.120 64.040 ; 
                RECT 2.880 65.080 126.600 65.400 ; 
                RECT 153.480 65.080 181.680 65.400 ; 
                RECT 283.360 65.080 290.120 65.400 ; 
                RECT 2.880 66.440 126.600 66.760 ; 
                RECT 165.720 66.440 181.680 66.760 ; 
                RECT 283.360 66.440 290.120 66.760 ; 
                RECT 2.880 67.800 126.600 68.120 ; 
                RECT 165.720 67.800 181.680 68.120 ; 
                RECT 283.360 67.800 290.120 68.120 ; 
                RECT 2.880 69.160 126.600 69.480 ; 
                RECT 168.440 69.160 181.680 69.480 ; 
                RECT 283.360 69.160 290.120 69.480 ; 
                RECT 2.880 70.520 126.600 70.840 ; 
                RECT 167.080 70.520 181.680 70.840 ; 
                RECT 283.360 70.520 290.120 70.840 ; 
                RECT 2.880 71.880 126.600 72.200 ; 
                RECT 168.440 71.880 181.680 72.200 ; 
                RECT 283.360 71.880 290.120 72.200 ; 
                RECT 2.880 73.240 126.600 73.560 ; 
                RECT 153.480 73.240 181.680 73.560 ; 
                RECT 283.360 73.240 290.120 73.560 ; 
                RECT 2.880 74.600 126.600 74.920 ; 
                RECT 168.440 74.600 181.680 74.920 ; 
                RECT 283.360 74.600 290.120 74.920 ; 
                RECT 2.880 75.960 126.600 76.280 ; 
                RECT 171.160 75.960 181.680 76.280 ; 
                RECT 283.360 75.960 290.120 76.280 ; 
                RECT 2.880 77.320 126.600 77.640 ; 
                RECT 169.800 77.320 181.680 77.640 ; 
                RECT 283.360 77.320 290.120 77.640 ; 
                RECT 2.880 78.680 126.600 79.000 ; 
                RECT 171.160 78.680 181.680 79.000 ; 
                RECT 283.360 78.680 290.120 79.000 ; 
                RECT 2.880 80.040 126.600 80.360 ; 
                RECT 171.160 80.040 181.680 80.360 ; 
                RECT 283.360 80.040 290.120 80.360 ; 
                RECT 2.880 81.400 126.600 81.720 ; 
                RECT 169.800 81.400 181.680 81.720 ; 
                RECT 283.360 81.400 290.120 81.720 ; 
                RECT 2.880 82.760 87.840 83.080 ; 
                RECT 99.080 82.760 126.600 83.080 ; 
                RECT 173.880 82.760 181.680 83.080 ; 
                RECT 283.360 82.760 290.120 83.080 ; 
                RECT 2.880 84.120 89.200 84.440 ; 
                RECT 95.000 84.120 102.800 84.440 ; 
                RECT 105.200 84.120 126.600 84.440 ; 
                RECT 172.520 84.120 181.680 84.440 ; 
                RECT 283.360 84.120 290.120 84.440 ; 
                RECT 2.880 85.480 90.560 85.800 ; 
                RECT 94.320 85.480 126.600 85.800 ; 
                RECT 173.880 85.480 181.680 85.800 ; 
                RECT 283.360 85.480 290.120 85.800 ; 
                RECT 2.880 86.840 126.600 87.160 ; 
                RECT 173.880 86.840 181.680 87.160 ; 
                RECT 283.360 86.840 290.120 87.160 ; 
                RECT 2.880 88.200 97.360 88.520 ; 
                RECT 105.880 88.200 126.600 88.520 ; 
                RECT 153.480 88.200 181.680 88.520 ; 
                RECT 283.360 88.200 290.120 88.520 ; 
                RECT 2.880 89.560 89.880 89.880 ; 
                RECT 99.080 89.560 126.600 89.880 ; 
                RECT 175.240 89.560 181.680 89.880 ; 
                RECT 283.360 89.560 290.120 89.880 ; 
                RECT 2.880 90.920 93.280 91.240 ; 
                RECT 98.400 90.920 126.600 91.240 ; 
                RECT 153.480 90.920 181.680 91.240 ; 
                RECT 283.360 90.920 290.120 91.240 ; 
                RECT 2.880 92.280 126.600 92.600 ; 
                RECT 176.600 92.280 181.680 92.600 ; 
                RECT 283.360 92.280 290.120 92.600 ; 
                RECT 2.880 93.640 87.160 93.960 ; 
                RECT 99.080 93.640 126.600 93.960 ; 
                RECT 176.600 93.640 181.680 93.960 ; 
                RECT 283.360 93.640 290.120 93.960 ; 
                RECT 2.880 95.000 96.000 95.320 ; 
                RECT 104.520 95.000 126.600 95.320 ; 
                RECT 179.320 95.000 181.680 95.320 ; 
                RECT 283.360 95.000 290.120 95.320 ; 
                RECT 2.880 96.360 126.600 96.680 ; 
                RECT 177.960 96.360 181.680 96.680 ; 
                RECT 283.360 96.360 290.120 96.680 ; 
                RECT 2.880 97.720 97.360 98.040 ; 
                RECT 103.160 97.720 126.600 98.040 ; 
                RECT 179.320 97.720 181.680 98.040 ; 
                RECT 283.360 97.720 290.120 98.040 ; 
                RECT 2.880 99.080 100.080 99.400 ; 
                RECT 105.200 99.080 126.600 99.400 ; 
                RECT 153.480 99.080 181.680 99.400 ; 
                RECT 283.360 99.080 290.120 99.400 ; 
                RECT 2.880 100.440 93.960 100.760 ; 
                RECT 99.080 100.440 126.600 100.760 ; 
                RECT 179.320 100.440 181.680 100.760 ; 
                RECT 283.360 100.440 290.120 100.760 ; 
                RECT 2.880 101.800 126.600 102.120 ; 
                RECT 283.360 101.800 290.120 102.120 ; 
                RECT 2.880 103.160 87.160 103.480 ; 
                RECT 99.080 103.160 100.080 103.480 ; 
                RECT 109.960 103.160 126.600 103.480 ; 
                RECT 283.360 103.160 290.120 103.480 ; 
                RECT 2.880 104.520 97.360 104.840 ; 
                RECT 105.200 104.520 126.600 104.840 ; 
                RECT 283.360 104.520 290.120 104.840 ; 
                RECT 2.880 105.880 96.000 106.200 ; 
                RECT 99.080 105.880 104.160 106.200 ; 
                RECT 112.000 105.880 126.600 106.200 ; 
                RECT 283.360 105.880 290.120 106.200 ; 
                RECT 2.880 107.240 87.840 107.560 ; 
                RECT 101.800 107.240 126.600 107.560 ; 
                RECT 283.360 107.240 290.120 107.560 ; 
                RECT 2.880 108.600 96.680 108.920 ; 
                RECT 105.200 108.600 181.680 108.920 ; 
                RECT 283.360 108.600 290.120 108.920 ; 
                RECT 2.880 109.960 93.960 110.280 ; 
                RECT 98.400 109.960 181.680 110.280 ; 
                RECT 283.360 109.960 290.120 110.280 ; 
                RECT 2.880 111.320 97.360 111.640 ; 
                RECT 105.880 111.320 157.200 111.640 ; 
                RECT 283.360 111.320 290.120 111.640 ; 
                RECT 2.880 112.680 178.960 113.000 ; 
                RECT 283.360 112.680 290.120 113.000 ; 
                RECT 2.880 114.040 89.880 114.360 ; 
                RECT 92.960 114.040 176.240 114.360 ; 
                RECT 283.360 114.040 290.120 114.360 ; 
                RECT 2.880 115.400 89.880 115.720 ; 
                RECT 99.080 115.400 173.520 115.720 ; 
                RECT 283.360 115.400 290.120 115.720 ; 
                RECT 2.880 116.760 170.800 117.080 ; 
                RECT 283.360 116.760 290.120 117.080 ; 
                RECT 2.880 118.120 168.080 118.440 ; 
                RECT 283.360 118.120 290.120 118.440 ; 
                RECT 2.880 119.480 96.000 119.800 ; 
                RECT 98.400 119.480 162.640 119.800 ; 
                RECT 283.360 119.480 290.120 119.800 ; 
                RECT 2.880 120.840 89.200 121.160 ; 
                RECT 104.520 120.840 159.920 121.160 ; 
                RECT 283.360 120.840 290.120 121.160 ; 
                RECT 2.880 122.200 96.000 122.520 ; 
                RECT 98.400 122.200 159.920 122.520 ; 
                RECT 283.360 122.200 290.120 122.520 ; 
                RECT 2.880 123.560 181.680 123.880 ; 
                RECT 283.360 123.560 290.120 123.880 ; 
                RECT 2.880 124.920 66.080 125.240 ; 
                RECT 84.800 124.920 91.240 125.240 ; 
                RECT 99.080 124.920 181.680 125.240 ; 
                RECT 283.360 124.920 290.120 125.240 ; 
                RECT 2.880 126.280 66.080 126.600 ; 
                RECT 84.800 126.280 87.840 126.600 ; 
                RECT 99.080 126.280 181.680 126.600 ; 
                RECT 283.360 126.280 290.120 126.600 ; 
                RECT 2.880 127.640 66.080 127.960 ; 
                RECT 84.800 127.640 93.280 127.960 ; 
                RECT 105.200 127.640 181.680 127.960 ; 
                RECT 283.360 127.640 290.120 127.960 ; 
                RECT 2.880 129.000 66.080 129.320 ; 
                RECT 84.800 129.000 87.160 129.320 ; 
                RECT 95.000 129.000 181.680 129.320 ; 
                RECT 283.360 129.000 290.120 129.320 ; 
                RECT 2.880 130.360 66.080 130.680 ; 
                RECT 101.800 130.360 181.680 130.680 ; 
                RECT 283.360 130.360 290.120 130.680 ; 
                RECT 2.880 131.720 66.080 132.040 ; 
                RECT 84.800 131.720 181.680 132.040 ; 
                RECT 283.360 131.720 290.120 132.040 ; 
                RECT 2.880 133.080 66.080 133.400 ; 
                RECT 84.800 133.080 181.680 133.400 ; 
                RECT 283.360 133.080 290.120 133.400 ; 
                RECT 2.880 134.440 66.080 134.760 ; 
                RECT 84.800 134.440 181.680 134.760 ; 
                RECT 283.360 134.440 290.120 134.760 ; 
                RECT 2.880 135.800 66.080 136.120 ; 
                RECT 84.800 135.800 100.080 136.120 ; 
                RECT 105.880 135.800 181.680 136.120 ; 
                RECT 283.360 135.800 290.120 136.120 ; 
                RECT 2.880 137.160 66.080 137.480 ; 
                RECT 84.800 137.160 181.680 137.480 ; 
                RECT 283.360 137.160 290.120 137.480 ; 
                RECT 2.880 138.520 66.080 138.840 ; 
                RECT 84.800 138.520 181.680 138.840 ; 
                RECT 283.360 138.520 290.120 138.840 ; 
                RECT 2.880 139.880 66.080 140.200 ; 
                RECT 84.800 139.880 87.160 140.200 ; 
                RECT 92.960 139.880 110.960 140.200 ; 
                RECT 153.480 139.880 181.680 140.200 ; 
                RECT 283.360 139.880 290.120 140.200 ; 
                RECT 2.880 141.240 66.080 141.560 ; 
                RECT 84.800 141.240 147.680 141.560 ; 
                RECT 153.480 141.240 181.680 141.560 ; 
                RECT 283.360 141.240 290.120 141.560 ; 
                RECT 2.880 142.600 66.080 142.920 ; 
                RECT 84.800 142.600 147.680 142.920 ; 
                RECT 153.480 142.600 181.680 142.920 ; 
                RECT 283.360 142.600 290.120 142.920 ; 
                RECT 2.880 143.960 66.080 144.280 ; 
                RECT 84.800 143.960 147.680 144.280 ; 
                RECT 153.480 143.960 181.680 144.280 ; 
                RECT 283.360 143.960 290.120 144.280 ; 
                RECT 2.880 145.320 66.080 145.640 ; 
                RECT 84.800 145.320 181.680 145.640 ; 
                RECT 283.360 145.320 290.120 145.640 ; 
                RECT 2.880 146.680 66.080 147.000 ; 
                RECT 84.800 146.680 92.600 147.000 ; 
                RECT 105.200 146.680 181.680 147.000 ; 
                RECT 283.360 146.680 290.120 147.000 ; 
                RECT 2.880 148.040 66.080 148.360 ; 
                RECT 84.800 148.040 161.280 148.360 ; 
                RECT 283.360 148.040 290.120 148.360 ; 
                RECT 2.880 149.400 66.080 149.720 ; 
                RECT 84.800 149.400 89.880 149.720 ; 
                RECT 94.320 149.400 161.280 149.720 ; 
                RECT 283.360 149.400 290.120 149.720 ; 
                RECT 2.880 150.760 66.080 151.080 ; 
                RECT 84.800 150.760 132.720 151.080 ; 
                RECT 152.800 150.760 164.000 151.080 ; 
                RECT 283.360 150.760 290.120 151.080 ; 
                RECT 2.880 152.120 66.080 152.440 ; 
                RECT 84.800 152.120 132.720 152.440 ; 
                RECT 152.800 152.120 169.440 152.440 ; 
                RECT 283.360 152.120 290.120 152.440 ; 
                RECT 2.880 153.480 66.080 153.800 ; 
                RECT 84.800 153.480 132.720 153.800 ; 
                RECT 152.800 153.480 172.160 153.800 ; 
                RECT 283.360 153.480 290.120 153.800 ; 
                RECT 2.880 154.840 66.080 155.160 ; 
                RECT 84.800 154.840 92.600 155.160 ; 
                RECT 95.000 154.840 132.720 155.160 ; 
                RECT 152.800 154.840 174.880 155.160 ; 
                RECT 283.360 154.840 290.120 155.160 ; 
                RECT 2.880 156.200 66.080 156.520 ; 
                RECT 84.800 156.200 89.200 156.520 ; 
                RECT 92.280 156.200 102.800 156.520 ; 
                RECT 105.880 156.200 132.720 156.520 ; 
                RECT 152.800 156.200 177.600 156.520 ; 
                RECT 283.360 156.200 290.120 156.520 ; 
                RECT 2.880 157.560 66.080 157.880 ; 
                RECT 84.800 157.560 132.720 157.880 ; 
                RECT 152.800 157.560 180.320 157.880 ; 
                RECT 283.360 157.560 290.120 157.880 ; 
                RECT 2.880 158.920 66.080 159.240 ; 
                RECT 84.800 158.920 132.720 159.240 ; 
                RECT 283.360 158.920 290.120 159.240 ; 
                RECT 2.880 160.280 66.080 160.600 ; 
                RECT 84.800 160.280 132.720 160.600 ; 
                RECT 152.800 160.280 181.680 160.600 ; 
                RECT 283.360 160.280 290.120 160.600 ; 
                RECT 2.880 161.640 66.080 161.960 ; 
                RECT 84.800 161.640 132.720 161.960 ; 
                RECT 152.800 161.640 181.680 161.960 ; 
                RECT 283.360 161.640 290.120 161.960 ; 
                RECT 2.880 163.000 66.080 163.320 ; 
                RECT 84.800 163.000 132.720 163.320 ; 
                RECT 152.800 163.000 181.680 163.320 ; 
                RECT 283.360 163.000 290.120 163.320 ; 
                RECT 2.880 164.360 66.080 164.680 ; 
                RECT 84.800 164.360 96.000 164.680 ; 
                RECT 104.520 164.360 132.720 164.680 ; 
                RECT 152.800 164.360 181.680 164.680 ; 
                RECT 283.360 164.360 290.120 164.680 ; 
                RECT 2.880 165.720 91.240 166.040 ; 
                RECT 95.000 165.720 132.720 166.040 ; 
                RECT 152.800 165.720 181.680 166.040 ; 
                RECT 283.360 165.720 290.120 166.040 ; 
                RECT 2.880 167.080 132.720 167.400 ; 
                RECT 152.800 167.080 181.680 167.400 ; 
                RECT 283.360 167.080 290.120 167.400 ; 
                RECT 2.880 168.440 45.000 168.760 ; 
                RECT 65.760 168.440 132.720 168.760 ; 
                RECT 152.800 168.440 181.680 168.760 ; 
                RECT 283.360 168.440 290.120 168.760 ; 
                RECT 2.880 169.800 45.000 170.120 ; 
                RECT 65.760 169.800 93.280 170.120 ; 
                RECT 99.080 169.800 132.720 170.120 ; 
                RECT 152.800 169.800 181.680 170.120 ; 
                RECT 283.360 169.800 290.120 170.120 ; 
                RECT 2.880 171.160 45.000 171.480 ; 
                RECT 65.760 171.160 72.200 171.480 ; 
                RECT 79.360 171.160 132.720 171.480 ; 
                RECT 152.800 171.160 181.680 171.480 ; 
                RECT 283.360 171.160 290.120 171.480 ; 
                RECT 2.880 172.520 45.000 172.840 ; 
                RECT 65.760 172.520 66.760 172.840 ; 
                RECT 84.120 172.520 132.720 172.840 ; 
                RECT 152.800 172.520 181.680 172.840 ; 
                RECT 283.360 172.520 290.120 172.840 ; 
                RECT 2.880 173.880 45.000 174.200 ; 
                RECT 65.760 173.880 66.760 174.200 ; 
                RECT 84.120 173.880 132.720 174.200 ; 
                RECT 283.360 173.880 290.120 174.200 ; 
                RECT 2.880 175.240 45.000 175.560 ; 
                RECT 65.760 175.240 72.200 175.560 ; 
                RECT 79.360 175.240 87.840 175.560 ; 
                RECT 97.720 175.240 132.720 175.560 ; 
                RECT 283.360 175.240 290.120 175.560 ; 
                RECT 2.880 176.600 32.760 176.920 ; 
                RECT 78.680 176.600 132.720 176.920 ; 
                RECT 152.800 176.600 290.120 176.920 ; 
                RECT 2.880 177.960 78.320 178.280 ; 
                RECT 129.680 177.960 290.120 178.280 ; 
                RECT 2.880 179.320 178.960 179.640 ; 
                RECT 286.080 179.320 290.120 179.640 ; 
                RECT 2.880 180.680 178.960 181.000 ; 
                RECT 286.080 180.680 290.120 181.000 ; 
                RECT 2.880 182.040 178.960 182.360 ; 
                RECT 286.080 182.040 290.120 182.360 ; 
                RECT 2.880 183.400 28.000 183.720 ; 
                RECT 34.480 183.400 36.160 183.720 ; 
                RECT 49.440 183.400 99.400 183.720 ; 
                RECT 286.080 183.400 290.120 183.720 ; 
                RECT 2.880 184.760 25.960 185.080 ; 
                RECT 48.080 184.760 59.960 185.080 ; 
                RECT 61.680 184.760 76.280 185.080 ; 
                RECT 90.240 184.760 99.400 185.080 ; 
                RECT 286.080 184.760 290.120 185.080 ; 
                RECT 2.880 186.120 25.960 186.440 ; 
                RECT 36.520 186.120 59.960 186.440 ; 
                RECT 63.720 186.120 76.280 186.440 ; 
                RECT 90.240 186.120 99.400 186.440 ; 
                RECT 286.080 186.120 290.120 186.440 ; 
                RECT 2.880 187.480 25.960 187.800 ; 
                RECT 36.520 187.480 59.960 187.800 ; 
                RECT 64.400 187.480 76.280 187.800 ; 
                RECT 90.240 187.480 99.400 187.800 ; 
                RECT 286.080 187.480 290.120 187.800 ; 
                RECT 2.880 188.840 25.960 189.160 ; 
                RECT 36.520 188.840 59.960 189.160 ; 
                RECT 65.080 188.840 76.280 189.160 ; 
                RECT 90.240 188.840 99.400 189.160 ; 
                RECT 286.080 188.840 290.120 189.160 ; 
                RECT 2.880 190.200 25.960 190.520 ; 
                RECT 36.520 190.200 59.960 190.520 ; 
                RECT 61.680 190.200 76.280 190.520 ; 
                RECT 90.240 190.200 99.400 190.520 ; 
                RECT 286.080 190.200 290.120 190.520 ; 
                RECT 2.880 191.560 25.960 191.880 ; 
                RECT 36.520 191.560 99.400 191.880 ; 
                RECT 286.080 191.560 290.120 191.880 ; 
                RECT 2.880 192.920 25.960 193.240 ; 
                RECT 36.520 192.920 76.280 193.240 ; 
                RECT 90.240 192.920 99.400 193.240 ; 
                RECT 286.080 192.920 290.120 193.240 ; 
                RECT 2.880 194.280 76.280 194.600 ; 
                RECT 90.240 194.280 99.400 194.600 ; 
                RECT 286.080 194.280 290.120 194.600 ; 
                RECT 2.880 195.640 76.280 195.960 ; 
                RECT 90.240 195.640 99.400 195.960 ; 
                RECT 286.080 195.640 290.120 195.960 ; 
                RECT 2.880 197.000 19.160 197.320 ; 
                RECT 21.560 197.000 76.280 197.320 ; 
                RECT 90.240 197.000 99.400 197.320 ; 
                RECT 286.080 197.000 290.120 197.320 ; 
                RECT 2.880 198.360 76.280 198.680 ; 
                RECT 90.240 198.360 99.400 198.680 ; 
                RECT 286.080 198.360 290.120 198.680 ; 
                RECT 2.880 199.720 18.480 200.040 ; 
                RECT 21.560 199.720 34.800 200.040 ; 
                RECT 48.760 199.720 99.400 200.040 ; 
                RECT 286.080 199.720 290.120 200.040 ; 
                RECT 2.880 201.080 17.800 201.400 ; 
                RECT 21.560 201.080 34.800 201.400 ; 
                RECT 48.080 201.080 59.960 201.400 ; 
                RECT 61.680 201.080 76.280 201.400 ; 
                RECT 90.240 201.080 99.400 201.400 ; 
                RECT 286.080 201.080 290.120 201.400 ; 
                RECT 2.880 202.440 17.120 202.760 ; 
                RECT 21.560 202.440 34.800 202.760 ; 
                RECT 39.240 202.440 59.960 202.760 ; 
                RECT 61.680 202.440 76.280 202.760 ; 
                RECT 90.240 202.440 99.400 202.760 ; 
                RECT 286.080 202.440 290.120 202.760 ; 
                RECT 2.880 203.800 59.960 204.120 ; 
                RECT 62.360 203.800 76.280 204.120 ; 
                RECT 90.240 203.800 99.400 204.120 ; 
                RECT 286.080 203.800 290.120 204.120 ; 
                RECT 2.880 205.160 16.440 205.480 ; 
                RECT 21.560 205.160 34.800 205.480 ; 
                RECT 39.920 205.160 59.960 205.480 ; 
                RECT 63.040 205.160 76.280 205.480 ; 
                RECT 90.240 205.160 99.400 205.480 ; 
                RECT 286.080 205.160 290.120 205.480 ; 
                RECT 2.880 206.520 15.760 206.840 ; 
                RECT 21.560 206.520 34.800 206.840 ; 
                RECT 40.600 206.520 59.960 206.840 ; 
                RECT 63.040 206.520 76.280 206.840 ; 
                RECT 90.240 206.520 99.400 206.840 ; 
                RECT 286.080 206.520 290.120 206.840 ; 
                RECT 2.880 207.880 15.080 208.200 ; 
                RECT 21.560 207.880 99.400 208.200 ; 
                RECT 286.080 207.880 290.120 208.200 ; 
                RECT 2.880 209.240 14.400 209.560 ; 
                RECT 21.560 209.240 76.280 209.560 ; 
                RECT 90.240 209.240 99.400 209.560 ; 
                RECT 286.080 209.240 290.120 209.560 ; 
                RECT 2.880 210.600 76.280 210.920 ; 
                RECT 90.240 210.600 99.400 210.920 ; 
                RECT 286.080 210.600 290.120 210.920 ; 
                RECT 2.880 211.960 13.720 212.280 ; 
                RECT 21.560 211.960 76.280 212.280 ; 
                RECT 90.240 211.960 99.400 212.280 ; 
                RECT 286.080 211.960 290.120 212.280 ; 
                RECT 2.880 213.320 13.040 213.640 ; 
                RECT 21.560 213.320 76.280 213.640 ; 
                RECT 90.240 213.320 99.400 213.640 ; 
                RECT 286.080 213.320 290.120 213.640 ; 
                RECT 2.880 214.680 76.280 215.000 ; 
                RECT 85.480 214.680 99.400 215.000 ; 
                RECT 286.080 214.680 290.120 215.000 ; 
                RECT 2.880 216.040 12.360 216.360 ; 
                RECT 21.560 216.040 34.800 216.360 ; 
                RECT 39.240 216.040 80.360 216.360 ; 
                RECT 90.240 216.040 99.400 216.360 ; 
                RECT 286.080 216.040 290.120 216.360 ; 
                RECT 2.880 217.400 11.680 217.720 ; 
                RECT 21.560 217.400 34.800 217.720 ; 
                RECT 38.560 217.400 76.280 217.720 ; 
                RECT 90.240 217.400 99.400 217.720 ; 
                RECT 286.080 217.400 290.120 217.720 ; 
                RECT 2.880 218.760 76.280 219.080 ; 
                RECT 90.240 218.760 99.400 219.080 ; 
                RECT 286.080 218.760 290.120 219.080 ; 
                RECT 2.880 220.120 11.000 220.440 ; 
                RECT 21.560 220.120 34.800 220.440 ; 
                RECT 37.880 220.120 76.280 220.440 ; 
                RECT 90.240 220.120 99.400 220.440 ; 
                RECT 286.080 220.120 290.120 220.440 ; 
                RECT 2.880 221.480 10.320 221.800 ; 
                RECT 21.560 221.480 34.800 221.800 ; 
                RECT 37.200 221.480 76.280 221.800 ; 
                RECT 90.240 221.480 99.400 221.800 ; 
                RECT 286.080 221.480 290.120 221.800 ; 
                RECT 2.880 222.840 76.280 223.160 ; 
                RECT 86.840 222.840 99.400 223.160 ; 
                RECT 286.080 222.840 290.120 223.160 ; 
                RECT 2.880 224.200 76.280 224.520 ; 
                RECT 90.240 224.200 99.400 224.520 ; 
                RECT 286.080 224.200 290.120 224.520 ; 
                RECT 2.880 225.560 76.280 225.880 ; 
                RECT 90.240 225.560 99.400 225.880 ; 
                RECT 286.080 225.560 290.120 225.880 ; 
                RECT 2.880 226.920 76.280 227.240 ; 
                RECT 90.240 226.920 99.400 227.240 ; 
                RECT 286.080 226.920 290.120 227.240 ; 
                RECT 2.880 228.280 76.280 228.600 ; 
                RECT 90.240 228.280 99.400 228.600 ; 
                RECT 286.080 228.280 290.120 228.600 ; 
                RECT 2.880 229.640 76.280 229.960 ; 
                RECT 90.240 229.640 99.400 229.960 ; 
                RECT 286.080 229.640 290.120 229.960 ; 
                RECT 2.880 231.000 76.280 231.320 ; 
                RECT 87.520 231.000 99.400 231.320 ; 
                RECT 286.080 231.000 290.120 231.320 ; 
                RECT 2.880 232.360 76.280 232.680 ; 
                RECT 90.240 232.360 99.400 232.680 ; 
                RECT 286.080 232.360 290.120 232.680 ; 
                RECT 2.880 233.720 76.280 234.040 ; 
                RECT 90.240 233.720 99.400 234.040 ; 
                RECT 286.080 233.720 290.120 234.040 ; 
                RECT 2.880 235.080 76.280 235.400 ; 
                RECT 90.240 235.080 99.400 235.400 ; 
                RECT 286.080 235.080 290.120 235.400 ; 
                RECT 2.880 236.440 76.280 236.760 ; 
                RECT 90.240 236.440 99.400 236.760 ; 
                RECT 286.080 236.440 290.120 236.760 ; 
                RECT 2.880 237.800 76.280 238.120 ; 
                RECT 90.240 237.800 99.400 238.120 ; 
                RECT 286.080 237.800 290.120 238.120 ; 
                RECT 2.880 239.160 99.400 239.480 ; 
                RECT 286.080 239.160 290.120 239.480 ; 
                RECT 2.880 240.520 76.280 240.840 ; 
                RECT 90.240 240.520 99.400 240.840 ; 
                RECT 286.080 240.520 290.120 240.840 ; 
                RECT 2.880 241.880 76.280 242.200 ; 
                RECT 90.240 241.880 99.400 242.200 ; 
                RECT 286.080 241.880 290.120 242.200 ; 
                RECT 2.880 243.240 76.280 243.560 ; 
                RECT 90.240 243.240 99.400 243.560 ; 
                RECT 286.080 243.240 290.120 243.560 ; 
                RECT 2.880 244.600 76.280 244.920 ; 
                RECT 90.240 244.600 99.400 244.920 ; 
                RECT 286.080 244.600 290.120 244.920 ; 
                RECT 2.880 245.960 76.280 246.280 ; 
                RECT 90.240 245.960 99.400 246.280 ; 
                RECT 286.080 245.960 290.120 246.280 ; 
                RECT 2.880 247.320 99.400 247.640 ; 
                RECT 286.080 247.320 290.120 247.640 ; 
                RECT 2.880 248.680 77.640 249.000 ; 
                RECT 90.240 248.680 99.400 249.000 ; 
                RECT 286.080 248.680 290.120 249.000 ; 
                RECT 2.880 250.040 77.640 250.360 ; 
                RECT 90.240 250.040 99.400 250.360 ; 
                RECT 286.080 250.040 290.120 250.360 ; 
                RECT 2.880 251.400 77.640 251.720 ; 
                RECT 90.240 251.400 99.400 251.720 ; 
                RECT 286.080 251.400 290.120 251.720 ; 
                RECT 2.880 252.760 81.720 253.080 ; 
                RECT 90.240 252.760 99.400 253.080 ; 
                RECT 286.080 252.760 290.120 253.080 ; 
                RECT 2.880 254.120 77.640 254.440 ; 
                RECT 90.240 254.120 99.400 254.440 ; 
                RECT 286.080 254.120 290.120 254.440 ; 
                RECT 2.880 255.480 38.880 255.800 ; 
                RECT 65.080 255.480 99.400 255.800 ; 
                RECT 286.080 255.480 290.120 255.800 ; 
                RECT 2.880 256.840 37.520 257.160 ; 
                RECT 64.400 256.840 76.280 257.160 ; 
                RECT 90.240 256.840 99.400 257.160 ; 
                RECT 286.080 256.840 290.120 257.160 ; 
                RECT 2.880 258.200 36.160 258.520 ; 
                RECT 63.040 258.200 76.280 258.520 ; 
                RECT 90.240 258.200 99.400 258.520 ; 
                RECT 286.080 258.200 290.120 258.520 ; 
                RECT 2.880 259.560 77.640 259.880 ; 
                RECT 90.240 259.560 99.400 259.880 ; 
                RECT 286.080 259.560 290.120 259.880 ; 
                RECT 2.880 260.920 76.280 261.240 ; 
                RECT 90.240 260.920 99.400 261.240 ; 
                RECT 286.080 260.920 290.120 261.240 ; 
                RECT 2.880 262.280 76.280 262.600 ; 
                RECT 78.680 262.280 99.400 262.600 ; 
                RECT 286.080 262.280 290.120 262.600 ; 
                RECT 2.880 263.640 84.440 263.960 ; 
                RECT 90.240 263.640 99.400 263.960 ; 
                RECT 286.080 263.640 290.120 263.960 ; 
                RECT 2.880 265.000 76.280 265.320 ; 
                RECT 90.240 265.000 99.400 265.320 ; 
                RECT 286.080 265.000 290.120 265.320 ; 
                RECT 2.880 266.360 76.280 266.680 ; 
                RECT 90.240 266.360 99.400 266.680 ; 
                RECT 286.080 266.360 290.120 266.680 ; 
                RECT 2.880 267.720 76.280 268.040 ; 
                RECT 90.240 267.720 99.400 268.040 ; 
                RECT 286.080 267.720 290.120 268.040 ; 
                RECT 2.880 269.080 76.280 269.400 ; 
                RECT 90.240 269.080 99.400 269.400 ; 
                RECT 286.080 269.080 290.120 269.400 ; 
                RECT 2.880 270.440 76.280 270.760 ; 
                RECT 78.680 270.440 99.400 270.760 ; 
                RECT 286.080 270.440 290.120 270.760 ; 
                RECT 2.880 271.800 86.480 272.120 ; 
                RECT 90.240 271.800 99.400 272.120 ; 
                RECT 286.080 271.800 290.120 272.120 ; 
                RECT 2.880 273.160 76.280 273.480 ; 
                RECT 90.240 273.160 99.400 273.480 ; 
                RECT 286.080 273.160 290.120 273.480 ; 
                RECT 2.880 274.520 76.280 274.840 ; 
                RECT 90.240 274.520 99.400 274.840 ; 
                RECT 286.080 274.520 290.120 274.840 ; 
                RECT 2.880 275.880 76.280 276.200 ; 
                RECT 90.240 275.880 99.400 276.200 ; 
                RECT 286.080 275.880 290.120 276.200 ; 
                RECT 2.880 277.240 76.280 277.560 ; 
                RECT 90.240 277.240 99.400 277.560 ; 
                RECT 286.080 277.240 290.120 277.560 ; 
                RECT 2.880 278.600 99.400 278.920 ; 
                RECT 286.080 278.600 290.120 278.920 ; 
                RECT 2.880 279.960 78.320 280.280 ; 
                RECT 90.240 279.960 99.400 280.280 ; 
                RECT 286.080 279.960 290.120 280.280 ; 
                RECT 2.880 281.320 76.280 281.640 ; 
                RECT 90.240 281.320 99.400 281.640 ; 
                RECT 286.080 281.320 290.120 281.640 ; 
                RECT 2.880 282.680 76.280 283.000 ; 
                RECT 90.240 282.680 99.400 283.000 ; 
                RECT 286.080 282.680 290.120 283.000 ; 
                RECT 2.880 284.040 76.280 284.360 ; 
                RECT 90.240 284.040 99.400 284.360 ; 
                RECT 286.080 284.040 290.120 284.360 ; 
                RECT 2.880 285.400 76.280 285.720 ; 
                RECT 90.240 285.400 99.400 285.720 ; 
                RECT 286.080 285.400 290.120 285.720 ; 
                RECT 2.880 286.760 99.400 287.080 ; 
                RECT 286.080 286.760 290.120 287.080 ; 
                RECT 2.880 288.120 78.320 288.440 ; 
                RECT 90.240 288.120 99.400 288.440 ; 
                RECT 286.080 288.120 290.120 288.440 ; 
                RECT 2.880 289.480 76.280 289.800 ; 
                RECT 90.240 289.480 99.400 289.800 ; 
                RECT 286.080 289.480 290.120 289.800 ; 
                RECT 2.880 290.840 76.280 291.160 ; 
                RECT 90.240 290.840 99.400 291.160 ; 
                RECT 286.080 290.840 290.120 291.160 ; 
                RECT 2.880 292.200 76.280 292.520 ; 
                RECT 90.240 292.200 99.400 292.520 ; 
                RECT 286.080 292.200 290.120 292.520 ; 
                RECT 2.880 293.560 76.280 293.880 ; 
                RECT 90.240 293.560 99.400 293.880 ; 
                RECT 286.080 293.560 290.120 293.880 ; 
                RECT 2.880 294.920 99.400 295.240 ; 
                RECT 286.080 294.920 290.120 295.240 ; 
                RECT 2.880 296.280 76.280 296.600 ; 
                RECT 90.240 296.280 99.400 296.600 ; 
                RECT 286.080 296.280 290.120 296.600 ; 
                RECT 2.880 297.640 76.280 297.960 ; 
                RECT 90.240 297.640 99.400 297.960 ; 
                RECT 286.080 297.640 290.120 297.960 ; 
                RECT 2.880 299.000 78.320 299.320 ; 
                RECT 90.240 299.000 99.400 299.320 ; 
                RECT 286.080 299.000 290.120 299.320 ; 
                RECT 2.880 300.360 76.280 300.680 ; 
                RECT 90.240 300.360 99.400 300.680 ; 
                RECT 286.080 300.360 290.120 300.680 ; 
                RECT 2.880 301.720 76.280 302.040 ; 
                RECT 80.720 301.720 99.400 302.040 ; 
                RECT 286.080 301.720 290.120 302.040 ; 
                RECT 2.880 303.080 86.480 303.400 ; 
                RECT 90.240 303.080 99.400 303.400 ; 
                RECT 286.080 303.080 290.120 303.400 ; 
                RECT 2.880 304.440 76.280 304.760 ; 
                RECT 90.240 304.440 99.400 304.760 ; 
                RECT 286.080 304.440 290.120 304.760 ; 
                RECT 2.880 305.800 76.280 306.120 ; 
                RECT 90.240 305.800 99.400 306.120 ; 
                RECT 286.080 305.800 290.120 306.120 ; 
                RECT 2.880 307.160 76.280 307.480 ; 
                RECT 90.240 307.160 99.400 307.480 ; 
                RECT 286.080 307.160 290.120 307.480 ; 
                RECT 2.880 308.520 76.280 308.840 ; 
                RECT 90.240 308.520 99.400 308.840 ; 
                RECT 286.080 308.520 290.120 308.840 ; 
                RECT 2.880 309.880 76.280 310.200 ; 
                RECT 81.400 309.880 99.400 310.200 ; 
                RECT 286.080 309.880 290.120 310.200 ; 
                RECT 2.880 311.240 80.360 311.560 ; 
                RECT 90.240 311.240 99.400 311.560 ; 
                RECT 286.080 311.240 290.120 311.560 ; 
                RECT 2.880 312.600 76.280 312.920 ; 
                RECT 90.240 312.600 99.400 312.920 ; 
                RECT 286.080 312.600 290.120 312.920 ; 
                RECT 2.880 313.960 76.280 314.280 ; 
                RECT 90.240 313.960 99.400 314.280 ; 
                RECT 286.080 313.960 290.120 314.280 ; 
                RECT 2.880 315.320 76.280 315.640 ; 
                RECT 90.240 315.320 99.400 315.640 ; 
                RECT 286.080 315.320 290.120 315.640 ; 
                RECT 2.880 316.680 76.280 317.000 ; 
                RECT 90.240 316.680 99.400 317.000 ; 
                RECT 286.080 316.680 290.120 317.000 ; 
                RECT 2.880 318.040 99.400 318.360 ; 
                RECT 286.080 318.040 290.120 318.360 ; 
                RECT 2.880 319.400 78.320 319.720 ; 
                RECT 90.240 319.400 99.400 319.720 ; 
                RECT 286.080 319.400 290.120 319.720 ; 
                RECT 2.880 320.760 83.080 321.080 ; 
                RECT 90.240 320.760 99.400 321.080 ; 
                RECT 286.080 320.760 290.120 321.080 ; 
                RECT 2.880 322.120 83.080 322.440 ; 
                RECT 90.240 322.120 99.400 322.440 ; 
                RECT 286.080 322.120 290.120 322.440 ; 
                RECT 2.880 323.480 78.320 323.800 ; 
                RECT 90.240 323.480 99.400 323.800 ; 
                RECT 286.080 323.480 290.120 323.800 ; 
                RECT 2.880 324.840 78.320 325.160 ; 
                RECT 90.240 324.840 99.400 325.160 ; 
                RECT 286.080 324.840 290.120 325.160 ; 
                RECT 2.880 326.200 99.400 326.520 ; 
                RECT 286.080 326.200 290.120 326.520 ; 
                RECT 2.880 327.560 78.320 327.880 ; 
                RECT 90.240 327.560 99.400 327.880 ; 
                RECT 286.080 327.560 290.120 327.880 ; 
                RECT 2.880 328.920 78.320 329.240 ; 
                RECT 90.240 328.920 99.400 329.240 ; 
                RECT 286.080 328.920 290.120 329.240 ; 
                RECT 2.880 330.280 78.320 330.600 ; 
                RECT 90.240 330.280 99.400 330.600 ; 
                RECT 286.080 330.280 290.120 330.600 ; 
                RECT 2.880 331.640 85.800 331.960 ; 
                RECT 90.240 331.640 99.400 331.960 ; 
                RECT 286.080 331.640 290.120 331.960 ; 
                RECT 2.880 333.000 78.320 333.320 ; 
                RECT 90.240 333.000 99.400 333.320 ; 
                RECT 286.080 333.000 290.120 333.320 ; 
                RECT 2.880 334.360 99.400 334.680 ; 
                RECT 286.080 334.360 290.120 334.680 ; 
                RECT 2.880 335.720 78.320 336.040 ; 
                RECT 90.240 335.720 99.400 336.040 ; 
                RECT 286.080 335.720 290.120 336.040 ; 
                RECT 2.880 337.080 78.320 337.400 ; 
                RECT 90.240 337.080 99.400 337.400 ; 
                RECT 286.080 337.080 290.120 337.400 ; 
                RECT 2.880 338.440 78.320 338.760 ; 
                RECT 90.240 338.440 99.400 338.760 ; 
                RECT 286.080 338.440 290.120 338.760 ; 
                RECT 2.880 339.800 78.320 340.120 ; 
                RECT 90.240 339.800 99.400 340.120 ; 
                RECT 286.080 339.800 290.120 340.120 ; 
                RECT 2.880 341.160 99.400 341.480 ; 
                RECT 286.080 341.160 290.120 341.480 ; 
                RECT 2.880 342.520 80.360 342.840 ; 
                RECT 90.240 342.520 99.400 342.840 ; 
                RECT 286.080 342.520 290.120 342.840 ; 
                RECT 2.880 343.880 79.000 344.200 ; 
                RECT 90.240 343.880 99.400 344.200 ; 
                RECT 286.080 343.880 290.120 344.200 ; 
                RECT 2.880 345.240 79.000 345.560 ; 
                RECT 90.240 345.240 99.400 345.560 ; 
                RECT 286.080 345.240 290.120 345.560 ; 
                RECT 2.880 346.600 79.000 346.920 ; 
                RECT 90.240 346.600 99.400 346.920 ; 
                RECT 286.080 346.600 290.120 346.920 ; 
                RECT 2.880 347.960 79.000 348.280 ; 
                RECT 90.240 347.960 99.400 348.280 ; 
                RECT 286.080 347.960 290.120 348.280 ; 
                RECT 2.880 349.320 99.400 349.640 ; 
                RECT 286.080 349.320 290.120 349.640 ; 
                RECT 2.880 350.680 82.400 351.000 ; 
                RECT 90.240 350.680 99.400 351.000 ; 
                RECT 286.080 350.680 290.120 351.000 ; 
                RECT 2.880 352.040 79.000 352.360 ; 
                RECT 90.240 352.040 99.400 352.360 ; 
                RECT 286.080 352.040 290.120 352.360 ; 
                RECT 2.880 353.400 79.000 353.720 ; 
                RECT 90.240 353.400 99.400 353.720 ; 
                RECT 286.080 353.400 290.120 353.720 ; 
                RECT 2.880 354.760 79.000 355.080 ; 
                RECT 90.240 354.760 99.400 355.080 ; 
                RECT 286.080 354.760 290.120 355.080 ; 
                RECT 2.880 356.120 79.000 356.440 ; 
                RECT 90.240 356.120 99.400 356.440 ; 
                RECT 286.080 356.120 290.120 356.440 ; 
                RECT 2.880 357.480 99.400 357.800 ; 
                RECT 286.080 357.480 290.120 357.800 ; 
                RECT 2.880 358.840 79.000 359.160 ; 
                RECT 90.240 358.840 99.400 359.160 ; 
                RECT 286.080 358.840 290.120 359.160 ; 
                RECT 2.880 360.200 85.120 360.520 ; 
                RECT 90.240 360.200 99.400 360.520 ; 
                RECT 286.080 360.200 290.120 360.520 ; 
                RECT 2.880 361.560 79.000 361.880 ; 
                RECT 90.240 361.560 99.400 361.880 ; 
                RECT 286.080 361.560 290.120 361.880 ; 
                RECT 2.880 362.920 79.000 363.240 ; 
                RECT 90.240 362.920 99.400 363.240 ; 
                RECT 286.080 362.920 290.120 363.240 ; 
                RECT 2.880 364.280 79.000 364.600 ; 
                RECT 90.240 364.280 99.400 364.600 ; 
                RECT 286.080 364.280 290.120 364.600 ; 
                RECT 2.880 365.640 99.400 365.960 ; 
                RECT 286.080 365.640 290.120 365.960 ; 
                RECT 2.880 367.000 79.000 367.320 ; 
                RECT 90.240 367.000 99.400 367.320 ; 
                RECT 286.080 367.000 290.120 367.320 ; 
                RECT 2.880 368.360 79.000 368.680 ; 
                RECT 90.240 368.360 99.400 368.680 ; 
                RECT 286.080 368.360 290.120 368.680 ; 
                RECT 2.880 369.720 87.160 370.040 ; 
                RECT 90.240 369.720 99.400 370.040 ; 
                RECT 286.080 369.720 290.120 370.040 ; 
                RECT 2.880 371.080 87.840 371.400 ; 
                RECT 90.240 371.080 99.400 371.400 ; 
                RECT 286.080 371.080 290.120 371.400 ; 
                RECT 2.880 372.440 79.000 372.760 ; 
                RECT 90.240 372.440 99.400 372.760 ; 
                RECT 286.080 372.440 290.120 372.760 ; 
                RECT 2.880 373.800 99.400 374.120 ; 
                RECT 286.080 373.800 290.120 374.120 ; 
                RECT 2.880 375.160 79.680 375.480 ; 
                RECT 90.240 375.160 99.400 375.480 ; 
                RECT 286.080 375.160 290.120 375.480 ; 
                RECT 2.880 376.520 79.680 376.840 ; 
                RECT 90.240 376.520 99.400 376.840 ; 
                RECT 286.080 376.520 290.120 376.840 ; 
                RECT 2.880 377.880 79.680 378.200 ; 
                RECT 90.240 377.880 99.400 378.200 ; 
                RECT 286.080 377.880 290.120 378.200 ; 
                RECT 2.880 379.240 81.720 379.560 ; 
                RECT 90.240 379.240 99.400 379.560 ; 
                RECT 286.080 379.240 290.120 379.560 ; 
                RECT 2.880 380.600 99.400 380.920 ; 
                RECT 286.080 380.600 290.120 380.920 ; 
                RECT 2.880 381.960 82.400 382.280 ; 
                RECT 90.240 381.960 99.400 382.280 ; 
                RECT 286.080 381.960 290.120 382.280 ; 
                RECT 2.880 383.320 79.680 383.640 ; 
                RECT 90.240 383.320 99.400 383.640 ; 
                RECT 286.080 383.320 290.120 383.640 ; 
                RECT 2.880 384.680 79.680 385.000 ; 
                RECT 90.240 384.680 99.400 385.000 ; 
                RECT 286.080 384.680 290.120 385.000 ; 
                RECT 2.880 386.040 79.680 386.360 ; 
                RECT 90.240 386.040 99.400 386.360 ; 
                RECT 286.080 386.040 290.120 386.360 ; 
                RECT 2.880 387.400 79.680 387.720 ; 
                RECT 90.240 387.400 99.400 387.720 ; 
                RECT 286.080 387.400 290.120 387.720 ; 
                RECT 2.880 388.760 99.400 389.080 ; 
                RECT 286.080 388.760 290.120 389.080 ; 
                RECT 2.880 390.120 84.440 390.440 ; 
                RECT 90.240 390.120 99.400 390.440 ; 
                RECT 286.080 390.120 290.120 390.440 ; 
                RECT 2.880 391.480 79.680 391.800 ; 
                RECT 90.240 391.480 99.400 391.800 ; 
                RECT 286.080 391.480 290.120 391.800 ; 
                RECT 2.880 392.840 79.680 393.160 ; 
                RECT 90.240 392.840 99.400 393.160 ; 
                RECT 286.080 392.840 290.120 393.160 ; 
                RECT 2.880 394.200 79.680 394.520 ; 
                RECT 90.240 394.200 99.400 394.520 ; 
                RECT 286.080 394.200 290.120 394.520 ; 
                RECT 2.880 395.560 79.680 395.880 ; 
                RECT 90.240 395.560 99.400 395.880 ; 
                RECT 286.080 395.560 290.120 395.880 ; 
                RECT 2.880 396.920 99.400 397.240 ; 
                RECT 286.080 396.920 290.120 397.240 ; 
                RECT 2.880 398.280 79.680 398.600 ; 
                RECT 90.240 398.280 99.400 398.600 ; 
                RECT 286.080 398.280 290.120 398.600 ; 
                RECT 2.880 399.640 86.480 399.960 ; 
                RECT 90.240 399.640 99.400 399.960 ; 
                RECT 286.080 399.640 290.120 399.960 ; 
                RECT 2.880 401.000 79.680 401.320 ; 
                RECT 90.240 401.000 99.400 401.320 ; 
                RECT 286.080 401.000 290.120 401.320 ; 
                RECT 2.880 402.360 79.680 402.680 ; 
                RECT 90.240 402.360 99.400 402.680 ; 
                RECT 286.080 402.360 290.120 402.680 ; 
                RECT 2.880 403.720 79.680 404.040 ; 
                RECT 90.240 403.720 99.400 404.040 ; 
                RECT 286.080 403.720 290.120 404.040 ; 
                RECT 2.880 405.080 99.400 405.400 ; 
                RECT 286.080 405.080 290.120 405.400 ; 
                RECT 2.880 406.440 80.360 406.760 ; 
                RECT 90.240 406.440 99.400 406.760 ; 
                RECT 286.080 406.440 290.120 406.760 ; 
                RECT 2.880 407.800 80.360 408.120 ; 
                RECT 90.240 407.800 99.400 408.120 ; 
                RECT 286.080 407.800 290.120 408.120 ; 
                RECT 2.880 409.160 81.720 409.480 ; 
                RECT 90.240 409.160 99.400 409.480 ; 
                RECT 286.080 409.160 290.120 409.480 ; 
                RECT 2.880 410.520 80.360 410.840 ; 
                RECT 90.240 410.520 99.400 410.840 ; 
                RECT 286.080 410.520 290.120 410.840 ; 
                RECT 2.880 411.880 80.360 412.200 ; 
                RECT 90.240 411.880 99.400 412.200 ; 
                RECT 286.080 411.880 290.120 412.200 ; 
                RECT 2.880 413.240 99.400 413.560 ; 
                RECT 286.080 413.240 290.120 413.560 ; 
                RECT 2.880 414.600 80.360 414.920 ; 
                RECT 90.240 414.600 99.400 414.920 ; 
                RECT 286.080 414.600 290.120 414.920 ; 
                RECT 2.880 415.960 80.360 416.280 ; 
                RECT 90.240 415.960 99.400 416.280 ; 
                RECT 286.080 415.960 290.120 416.280 ; 
                RECT 2.880 417.320 80.360 417.640 ; 
                RECT 90.240 417.320 99.400 417.640 ; 
                RECT 286.080 417.320 290.120 417.640 ; 
                RECT 2.880 418.680 83.760 419.000 ; 
                RECT 90.240 418.680 99.400 419.000 ; 
                RECT 286.080 418.680 290.120 419.000 ; 
                RECT 2.880 420.040 80.360 420.360 ; 
                RECT 90.240 420.040 99.400 420.360 ; 
                RECT 286.080 420.040 290.120 420.360 ; 
                RECT 2.880 421.400 99.400 421.720 ; 
                RECT 286.080 421.400 290.120 421.720 ; 
                RECT 2.880 422.760 80.360 423.080 ; 
                RECT 90.240 422.760 99.400 423.080 ; 
                RECT 286.080 422.760 290.120 423.080 ; 
                RECT 2.880 424.120 80.360 424.440 ; 
                RECT 90.240 424.120 99.400 424.440 ; 
                RECT 286.080 424.120 290.120 424.440 ; 
                RECT 2.880 425.480 80.360 425.800 ; 
                RECT 90.240 425.480 99.400 425.800 ; 
                RECT 286.080 425.480 290.120 425.800 ; 
                RECT 2.880 426.840 80.360 427.160 ; 
                RECT 90.240 426.840 99.400 427.160 ; 
                RECT 286.080 426.840 290.120 427.160 ; 
                RECT 2.880 428.200 99.400 428.520 ; 
                RECT 286.080 428.200 290.120 428.520 ; 
                RECT 2.880 429.560 86.480 429.880 ; 
                RECT 90.240 429.560 99.400 429.880 ; 
                RECT 286.080 429.560 290.120 429.880 ; 
                RECT 2.880 430.920 80.360 431.240 ; 
                RECT 90.240 430.920 99.400 431.240 ; 
                RECT 286.080 430.920 290.120 431.240 ; 
                RECT 2.880 432.280 80.360 432.600 ; 
                RECT 90.240 432.280 99.400 432.600 ; 
                RECT 286.080 432.280 290.120 432.600 ; 
                RECT 2.880 433.640 80.360 433.960 ; 
                RECT 90.240 433.640 99.400 433.960 ; 
                RECT 286.080 433.640 290.120 433.960 ; 
                RECT 2.880 435.000 80.360 435.320 ; 
                RECT 90.240 435.000 99.400 435.320 ; 
                RECT 286.080 435.000 290.120 435.320 ; 
                RECT 2.880 436.360 99.400 436.680 ; 
                RECT 286.080 436.360 290.120 436.680 ; 
                RECT 2.880 437.720 99.400 438.040 ; 
                RECT 286.080 437.720 290.120 438.040 ; 
                RECT 2.880 439.080 178.960 439.400 ; 
                RECT 286.080 439.080 290.120 439.400 ; 
                RECT 2.880 440.440 178.960 440.760 ; 
                RECT 286.080 440.440 290.120 440.760 ; 
                RECT 2.880 441.800 290.120 442.120 ; 
                RECT 2.880 443.160 290.120 443.480 ; 
                RECT 2.880 444.520 290.120 444.840 ; 
                RECT 2.880 445.880 290.120 446.200 ; 
                RECT 2.880 447.240 290.120 447.560 ; 
                RECT 2.880 2.880 290.120 4.240 ; 
                RECT 2.880 448.560 290.120 449.920 ; 
                RECT 183.100 32.360 188.900 33.480 ; 
                RECT 275.800 32.360 281.600 33.480 ; 
                RECT 183.100 38.100 188.900 38.620 ; 
                RECT 275.800 38.100 281.600 38.620 ; 
                RECT 183.100 42.575 188.900 43.375 ; 
                RECT 275.800 42.575 281.600 43.375 ; 
                RECT 183.100 48.815 188.900 49.615 ; 
                RECT 275.800 48.815 281.600 49.615 ; 
                RECT 183.100 77.370 281.600 78.170 ; 
                RECT 183.100 109.725 281.600 110.015 ; 
                RECT 183.100 80.580 281.600 81.380 ; 
                RECT 183.100 72.680 281.600 73.480 ; 
                RECT 183.100 84.265 281.600 87.865 ; 
                RECT 183.100 75.690 281.600 76.490 ; 
                RECT 183.100 63.630 281.600 65.430 ; 
                RECT 183.100 141.935 281.600 143.735 ; 
                RECT 183.100 22.990 281.600 24.790 ; 
                RECT 100.155 183.115 101.265 437.495 ; 
                RECT 108.960 183.115 110.710 437.495 ; 
                RECT 123.375 183.115 125.295 437.495 ; 
                RECT 144.985 183.115 146.905 437.495 ; 
                RECT 148.825 183.115 150.745 437.495 ; 
                RECT 127.435 55.565 128.545 108.165 ; 
                RECT 134.950 55.565 135.840 108.165 ; 
                RECT 142.270 55.565 144.190 108.165 ; 
                RECT 133.330 150.940 134.220 176.480 ; 
                RECT 139.230 150.940 140.120 176.480 ; 
                RECT 145.775 150.940 147.095 176.480 ; 
                RECT 148.570 139.780 149.460 144.940 ; 
                RECT 149.000 44.405 149.890 49.565 ; 
                RECT 26.500 184.180 35.660 184.550 ; 
                RECT 26.500 187.620 35.660 188.730 ; 
                RECT 45.740 168.640 65.380 169.310 ; 
                RECT 45.740 169.975 65.380 171.665 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 293.000 452.800 ; 
        LAYER met2 ;
            RECT 0.000 0.000 293.000 452.800 ; 
    END 
END sram22_1024x8m8w1 
END LIBRARY 

