VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_1024x32m8w8
    CLASS BLOCK  ;
    FOREIGN sram22_1024x32m8w8   ;
    SIZE 764.240 BY 460.280 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 404.710 0.000 404.850 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 415.610 0.000 415.750 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 426.510 0.000 426.650 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 437.410 0.000 437.550 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 448.310 0.000 448.450 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 459.210 0.000 459.350 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 470.110 0.000 470.250 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 481.010 0.000 481.150 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 491.910 0.000 492.050 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 502.810 0.000 502.950 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 513.710 0.000 513.850 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 524.610 0.000 524.750 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 535.510 0.000 535.650 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 546.410 0.000 546.550 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 557.310 0.000 557.450 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 568.210 0.000 568.350 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 579.110 0.000 579.250 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 590.010 0.000 590.150 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 600.910 0.000 601.050 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 611.810 0.000 611.950 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 622.710 0.000 622.850 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 633.610 0.000 633.750 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 644.510 0.000 644.650 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 655.410 0.000 655.550 0.140 ; 
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 666.310 0.000 666.450 0.140 ; 
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 677.210 0.000 677.350 0.140 ; 
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 688.110 0.000 688.250 0.140 ; 
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 699.010 0.000 699.150 0.140 ; 
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 709.910 0.000 710.050 0.140 ; 
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 720.810 0.000 720.950 0.140 ; 
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 731.710 0.000 731.850 0.140 ; 
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 742.610 0.000 742.750 0.140 ; 
        END 
    END dout[31] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 404.290 0.000 404.430 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 415.190 0.000 415.330 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 426.090 0.000 426.230 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 436.990 0.000 437.130 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 447.890 0.000 448.030 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 458.790 0.000 458.930 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 469.690 0.000 469.830 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 480.590 0.000 480.730 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 491.490 0.000 491.630 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 502.390 0.000 502.530 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 513.290 0.000 513.430 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 524.190 0.000 524.330 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 535.090 0.000 535.230 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 545.990 0.000 546.130 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 556.890 0.000 557.030 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 567.790 0.000 567.930 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 578.690 0.000 578.830 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 589.590 0.000 589.730 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 600.490 0.000 600.630 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 611.390 0.000 611.530 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 622.290 0.000 622.430 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 633.190 0.000 633.330 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 644.090 0.000 644.230 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 654.990 0.000 655.130 0.140 ; 
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 665.890 0.000 666.030 0.140 ; 
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 676.790 0.000 676.930 0.140 ; 
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 687.690 0.000 687.830 0.140 ; 
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 698.590 0.000 698.730 0.140 ; 
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 709.490 0.000 709.630 0.140 ; 
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 720.390 0.000 720.530 0.140 ; 
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 731.290 0.000 731.430 0.140 ; 
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.858800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 742.190 0.000 742.330 0.140 ; 
        END 
    END din[31] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.669200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 403.940 0.000 404.080 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.669200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 491.140 0.000 491.280 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.669200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 578.340 0.000 578.480 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.669200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 665.540 0.000 665.680 0.140 ; 
        END 
    END wmask[3] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 347.960 0.000 348.280 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 341.840 0.000 342.160 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 335.720 0.000 336.040 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 329.600 0.000 329.920 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 323.480 0.000 323.800 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 318.040 0.000 318.360 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 311.920 0.000 312.240 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 305.800 0.000 306.120 0.320 ; 
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 299.680 0.000 300.000 0.320 ; 
        END 
    END addr[8] 
    PIN addr[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 293.560 0.000 293.880 0.320 ; 
        END 
    END addr[9] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 360.200 0.000 360.520 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.184700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 354.080 0.000 354.400 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 22.878000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 363.600 0.000 363.920 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 26.784000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 364.280 0.000 364.600 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 404.040 6.240 ; 
                RECT 743.720 5.920 764.080 6.240 ; 
                RECT 0.160 7.280 764.080 7.600 ; 
                RECT 0.160 8.640 764.080 8.960 ; 
                RECT 0.160 10.000 363.920 10.320 ; 
                RECT 666.200 10.000 764.080 10.320 ; 
                RECT 0.160 11.360 391.120 11.680 ; 
                RECT 754.600 11.360 764.080 11.680 ; 
                RECT 0.160 12.720 391.120 13.040 ; 
                RECT 754.600 12.720 764.080 13.040 ; 
                RECT 0.160 14.080 391.120 14.400 ; 
                RECT 754.600 14.080 764.080 14.400 ; 
                RECT 0.160 15.440 391.120 15.760 ; 
                RECT 754.600 15.440 764.080 15.760 ; 
                RECT 0.160 16.800 391.120 17.120 ; 
                RECT 754.600 16.800 764.080 17.120 ; 
                RECT 0.160 18.160 391.120 18.480 ; 
                RECT 754.600 18.160 764.080 18.480 ; 
                RECT 0.160 19.520 391.120 19.840 ; 
                RECT 754.600 19.520 764.080 19.840 ; 
                RECT 0.160 20.880 289.120 21.200 ; 
                RECT 364.960 20.880 391.120 21.200 ; 
                RECT 754.600 20.880 764.080 21.200 ; 
                RECT 0.160 22.240 391.120 22.560 ; 
                RECT 754.600 22.240 764.080 22.560 ; 
                RECT 0.160 23.600 391.120 23.920 ; 
                RECT 754.600 23.600 764.080 23.920 ; 
                RECT 0.160 24.960 289.120 25.280 ; 
                RECT 364.280 24.960 391.120 25.280 ; 
                RECT 754.600 24.960 764.080 25.280 ; 
                RECT 0.160 26.320 391.120 26.640 ; 
                RECT 754.600 26.320 764.080 26.640 ; 
                RECT 0.160 27.680 390.440 28.000 ; 
                RECT 754.600 27.680 764.080 28.000 ; 
                RECT 0.160 29.040 391.120 29.360 ; 
                RECT 754.600 29.040 764.080 29.360 ; 
                RECT 0.160 30.400 391.120 30.720 ; 
                RECT 754.600 30.400 764.080 30.720 ; 
                RECT 0.160 31.760 391.120 32.080 ; 
                RECT 754.600 31.760 764.080 32.080 ; 
                RECT 0.160 33.120 391.120 33.440 ; 
                RECT 754.600 33.120 764.080 33.440 ; 
                RECT 0.160 34.480 391.120 34.800 ; 
                RECT 754.600 34.480 764.080 34.800 ; 
                RECT 0.160 35.840 391.120 36.160 ; 
                RECT 754.600 35.840 764.080 36.160 ; 
                RECT 0.160 37.200 391.120 37.520 ; 
                RECT 754.600 37.200 764.080 37.520 ; 
                RECT 0.160 38.560 391.120 38.880 ; 
                RECT 754.600 38.560 764.080 38.880 ; 
                RECT 0.160 39.920 391.120 40.240 ; 
                RECT 754.600 39.920 764.080 40.240 ; 
                RECT 0.160 41.280 391.120 41.600 ; 
                RECT 754.600 41.280 764.080 41.600 ; 
                RECT 0.160 42.640 251.720 42.960 ; 
                RECT 337.080 42.640 391.120 42.960 ; 
                RECT 754.600 42.640 764.080 42.960 ; 
                RECT 0.160 44.000 250.360 44.320 ; 
                RECT 343.200 44.000 391.120 44.320 ; 
                RECT 754.600 44.000 764.080 44.320 ; 
                RECT 0.160 45.360 249.000 45.680 ; 
                RECT 349.320 45.360 391.120 45.680 ; 
                RECT 754.600 45.360 764.080 45.680 ; 
                RECT 0.160 46.720 225.880 47.040 ; 
                RECT 364.280 46.720 391.120 47.040 ; 
                RECT 754.600 46.720 764.080 47.040 ; 
                RECT 0.160 48.080 227.240 48.400 ; 
                RECT 354.760 48.080 391.120 48.400 ; 
                RECT 754.600 48.080 764.080 48.400 ; 
                RECT 0.160 49.440 391.120 49.760 ; 
                RECT 754.600 49.440 764.080 49.760 ; 
                RECT 0.160 50.800 391.120 51.120 ; 
                RECT 754.600 50.800 764.080 51.120 ; 
                RECT 0.160 52.160 355.760 52.480 ; 
                RECT 362.240 52.160 391.120 52.480 ; 
                RECT 754.600 52.160 764.080 52.480 ; 
                RECT 0.160 53.520 355.760 53.840 ; 
                RECT 754.600 53.520 764.080 53.840 ; 
                RECT 0.160 54.880 246.960 55.200 ; 
                RECT 352.720 54.880 355.760 55.200 ; 
                RECT 362.240 54.880 391.120 55.200 ; 
                RECT 754.600 54.880 764.080 55.200 ; 
                RECT 0.160 56.240 391.120 56.560 ; 
                RECT 754.600 56.240 764.080 56.560 ; 
                RECT 0.160 57.600 391.120 57.920 ; 
                RECT 754.600 57.600 764.080 57.920 ; 
                RECT 0.160 58.960 391.120 59.280 ; 
                RECT 754.600 58.960 764.080 59.280 ; 
                RECT 0.160 60.320 391.120 60.640 ; 
                RECT 754.600 60.320 764.080 60.640 ; 
                RECT 0.160 61.680 248.320 62.000 ; 
                RECT 256.840 61.680 263.280 62.000 ; 
                RECT 361.560 61.680 391.120 62.000 ; 
                RECT 754.600 61.680 764.080 62.000 ; 
                RECT 0.160 63.040 249.680 63.360 ; 
                RECT 255.480 63.040 263.280 63.360 ; 
                RECT 372.440 63.040 391.120 63.360 ; 
                RECT 754.600 63.040 764.080 63.360 ; 
                RECT 0.160 64.400 251.040 64.720 ; 
                RECT 254.800 64.400 263.280 64.720 ; 
                RECT 371.080 64.400 391.120 64.720 ; 
                RECT 754.600 64.400 764.080 64.720 ; 
                RECT 0.160 65.760 263.280 66.080 ; 
                RECT 372.440 65.760 391.120 66.080 ; 
                RECT 754.600 65.760 764.080 66.080 ; 
                RECT 0.160 67.120 263.280 67.440 ; 
                RECT 372.440 67.120 391.120 67.440 ; 
                RECT 754.600 67.120 764.080 67.440 ; 
                RECT 0.160 68.480 263.280 68.800 ; 
                RECT 375.160 68.480 391.120 68.800 ; 
                RECT 754.600 68.480 764.080 68.800 ; 
                RECT 0.160 69.840 263.280 70.160 ; 
                RECT 373.800 69.840 391.120 70.160 ; 
                RECT 754.600 69.840 764.080 70.160 ; 
                RECT 0.160 71.200 263.280 71.520 ; 
                RECT 361.560 71.200 391.120 71.520 ; 
                RECT 754.600 71.200 764.080 71.520 ; 
                RECT 0.160 72.560 263.280 72.880 ; 
                RECT 375.160 72.560 391.120 72.880 ; 
                RECT 754.600 72.560 764.080 72.880 ; 
                RECT 0.160 73.920 263.280 74.240 ; 
                RECT 375.160 73.920 391.120 74.240 ; 
                RECT 754.600 73.920 764.080 74.240 ; 
                RECT 0.160 75.280 263.280 75.600 ; 
                RECT 377.880 75.280 391.120 75.600 ; 
                RECT 754.600 75.280 764.080 75.600 ; 
                RECT 0.160 76.640 263.280 76.960 ; 
                RECT 376.520 76.640 391.120 76.960 ; 
                RECT 754.600 76.640 764.080 76.960 ; 
                RECT 0.160 78.000 263.280 78.320 ; 
                RECT 377.880 78.000 391.120 78.320 ; 
                RECT 754.600 78.000 764.080 78.320 ; 
                RECT 0.160 79.360 263.280 79.680 ; 
                RECT 361.560 79.360 391.120 79.680 ; 
                RECT 754.600 79.360 764.080 79.680 ; 
                RECT 0.160 80.720 263.280 81.040 ; 
                RECT 377.880 80.720 391.120 81.040 ; 
                RECT 754.600 80.720 764.080 81.040 ; 
                RECT 0.160 82.080 263.280 82.400 ; 
                RECT 380.600 82.080 391.120 82.400 ; 
                RECT 754.600 82.080 764.080 82.400 ; 
                RECT 0.160 83.440 263.280 83.760 ; 
                RECT 379.240 83.440 391.120 83.760 ; 
                RECT 754.600 83.440 764.080 83.760 ; 
                RECT 0.160 84.800 263.280 85.120 ; 
                RECT 380.600 84.800 391.120 85.120 ; 
                RECT 754.600 84.800 764.080 85.120 ; 
                RECT 0.160 86.160 223.840 86.480 ; 
                RECT 235.080 86.160 263.280 86.480 ; 
                RECT 380.600 86.160 391.120 86.480 ; 
                RECT 754.600 86.160 764.080 86.480 ; 
                RECT 0.160 87.520 225.200 87.840 ; 
                RECT 228.960 87.520 263.280 87.840 ; 
                RECT 361.560 87.520 391.120 87.840 ; 
                RECT 754.600 87.520 764.080 87.840 ; 
                RECT 0.160 88.880 227.240 89.200 ; 
                RECT 231.680 88.880 238.800 89.200 ; 
                RECT 241.200 88.880 263.280 89.200 ; 
                RECT 383.320 88.880 391.120 89.200 ; 
                RECT 754.600 88.880 764.080 89.200 ; 
                RECT 0.160 90.240 263.280 90.560 ; 
                RECT 381.960 90.240 391.120 90.560 ; 
                RECT 754.600 90.240 764.080 90.560 ; 
                RECT 0.160 91.600 233.360 91.920 ; 
                RECT 241.880 91.600 263.280 91.920 ; 
                RECT 383.320 91.600 391.120 91.920 ; 
                RECT 754.600 91.600 764.080 91.920 ; 
                RECT 0.160 92.960 228.600 93.280 ; 
                RECT 235.080 92.960 263.280 93.280 ; 
                RECT 383.320 92.960 391.120 93.280 ; 
                RECT 754.600 92.960 764.080 93.280 ; 
                RECT 0.160 94.320 225.880 94.640 ; 
                RECT 235.080 94.320 263.280 94.640 ; 
                RECT 386.040 94.320 391.120 94.640 ; 
                RECT 754.600 94.320 764.080 94.640 ; 
                RECT 0.160 95.680 263.280 96.000 ; 
                RECT 384.680 95.680 391.120 96.000 ; 
                RECT 754.600 95.680 764.080 96.000 ; 
                RECT 0.160 97.040 223.160 97.360 ; 
                RECT 235.080 97.040 263.280 97.360 ; 
                RECT 361.560 97.040 391.120 97.360 ; 
                RECT 754.600 97.040 764.080 97.360 ; 
                RECT 0.160 98.400 233.360 98.720 ; 
                RECT 241.200 98.400 263.280 98.720 ; 
                RECT 384.680 98.400 391.120 98.720 ; 
                RECT 754.600 98.400 764.080 98.720 ; 
                RECT 0.160 99.760 232.680 100.080 ; 
                RECT 235.080 99.760 263.280 100.080 ; 
                RECT 386.040 99.760 391.120 100.080 ; 
                RECT 754.600 99.760 764.080 100.080 ; 
                RECT 0.160 101.120 263.280 101.440 ; 
                RECT 388.760 101.120 391.120 101.440 ; 
                RECT 754.600 101.120 764.080 101.440 ; 
                RECT 0.160 102.480 233.360 102.800 ; 
                RECT 241.200 102.480 263.280 102.800 ; 
                RECT 387.400 102.480 391.120 102.800 ; 
                RECT 754.600 102.480 764.080 102.800 ; 
                RECT 0.160 103.840 229.960 104.160 ; 
                RECT 235.080 103.840 263.280 104.160 ; 
                RECT 388.760 103.840 391.120 104.160 ; 
                RECT 754.600 103.840 764.080 104.160 ; 
                RECT 0.160 105.200 232.680 105.520 ; 
                RECT 235.080 105.200 263.280 105.520 ; 
                RECT 361.560 105.200 391.120 105.520 ; 
                RECT 754.600 105.200 764.080 105.520 ; 
                RECT 0.160 106.560 236.080 106.880 ; 
                RECT 246.640 106.560 263.280 106.880 ; 
                RECT 388.760 106.560 391.120 106.880 ; 
                RECT 754.600 106.560 764.080 106.880 ; 
                RECT 0.160 107.920 223.840 108.240 ; 
                RECT 241.200 107.920 263.280 108.240 ; 
                RECT 754.600 107.920 764.080 108.240 ; 
                RECT 0.160 109.280 232.680 109.600 ; 
                RECT 235.080 109.280 240.840 109.600 ; 
                RECT 248.000 109.280 263.280 109.600 ; 
                RECT 754.600 109.280 764.080 109.600 ; 
                RECT 0.160 110.640 244.920 110.960 ; 
                RECT 248.680 110.640 263.280 110.960 ; 
                RECT 754.600 110.640 764.080 110.960 ; 
                RECT 0.160 112.000 223.840 112.320 ; 
                RECT 237.800 112.000 263.280 112.320 ; 
                RECT 754.600 112.000 764.080 112.320 ; 
                RECT 0.160 113.360 232.680 113.680 ; 
                RECT 241.200 113.360 263.280 113.680 ; 
                RECT 361.560 113.360 391.120 113.680 ; 
                RECT 754.600 113.360 764.080 113.680 ; 
                RECT 0.160 114.720 230.640 115.040 ; 
                RECT 241.880 114.720 391.120 115.040 ; 
                RECT 754.600 114.720 764.080 115.040 ; 
                RECT 0.160 116.080 391.120 116.400 ; 
                RECT 754.600 116.080 764.080 116.400 ; 
                RECT 0.160 117.440 226.560 117.760 ; 
                RECT 228.960 117.440 366.640 117.760 ; 
                RECT 754.600 117.440 764.080 117.760 ; 
                RECT 0.160 118.800 225.880 119.120 ; 
                RECT 235.080 118.800 388.400 119.120 ; 
                RECT 754.600 118.800 764.080 119.120 ; 
                RECT 0.160 120.160 228.600 120.480 ; 
                RECT 232.360 120.160 385.680 120.480 ; 
                RECT 754.600 120.160 764.080 120.480 ; 
                RECT 0.160 121.520 382.960 121.840 ; 
                RECT 754.600 121.520 764.080 121.840 ; 
                RECT 0.160 122.880 232.680 123.200 ; 
                RECT 234.400 122.880 380.240 123.200 ; 
                RECT 754.600 122.880 764.080 123.200 ; 
                RECT 0.160 124.240 225.200 124.560 ; 
                RECT 240.520 124.240 374.800 124.560 ; 
                RECT 754.600 124.240 764.080 124.560 ; 
                RECT 0.160 125.600 372.080 125.920 ; 
                RECT 754.600 125.600 764.080 125.920 ; 
                RECT 0.160 126.960 232.680 127.280 ; 
                RECT 234.400 126.960 369.360 127.280 ; 
                RECT 754.600 126.960 764.080 127.280 ; 
                RECT 0.160 128.320 227.240 128.640 ; 
                RECT 235.080 128.320 369.360 128.640 ; 
                RECT 754.600 128.320 764.080 128.640 ; 
                RECT 0.160 129.680 223.840 130.000 ; 
                RECT 231.680 129.680 232.680 130.000 ; 
                RECT 235.760 129.680 391.120 130.000 ; 
                RECT 754.600 129.680 764.080 130.000 ; 
                RECT 0.160 131.040 391.120 131.360 ; 
                RECT 754.600 131.040 764.080 131.360 ; 
                RECT 0.160 132.400 202.760 132.720 ; 
                RECT 220.800 132.400 223.160 132.720 ; 
                RECT 241.200 132.400 391.120 132.720 ; 
                RECT 754.600 132.400 764.080 132.720 ; 
                RECT 0.160 133.760 202.760 134.080 ; 
                RECT 234.400 133.760 391.120 134.080 ; 
                RECT 754.600 133.760 764.080 134.080 ; 
                RECT 0.160 135.120 202.760 135.440 ; 
                RECT 220.800 135.120 223.840 135.440 ; 
                RECT 237.800 135.120 391.120 135.440 ; 
                RECT 754.600 135.120 764.080 135.440 ; 
                RECT 0.160 136.480 202.760 136.800 ; 
                RECT 220.800 136.480 391.120 136.800 ; 
                RECT 754.600 136.480 764.080 136.800 ; 
                RECT 0.160 137.840 202.760 138.160 ; 
                RECT 220.800 137.840 391.120 138.160 ; 
                RECT 754.600 137.840 764.080 138.160 ; 
                RECT 0.160 139.200 202.760 139.520 ; 
                RECT 220.800 139.200 236.080 139.520 ; 
                RECT 242.560 139.200 391.120 139.520 ; 
                RECT 754.600 139.200 764.080 139.520 ; 
                RECT 0.160 140.560 202.760 140.880 ; 
                RECT 220.800 140.560 239.480 140.880 ; 
                RECT 241.200 140.560 391.120 140.880 ; 
                RECT 754.600 140.560 764.080 140.880 ; 
                RECT 0.160 141.920 202.760 142.240 ; 
                RECT 220.800 141.920 310.200 142.240 ; 
                RECT 360.880 141.920 391.120 142.240 ; 
                RECT 754.600 141.920 764.080 142.240 ; 
                RECT 0.160 143.280 202.760 143.600 ; 
                RECT 220.800 143.280 225.880 143.600 ; 
                RECT 228.960 143.280 310.200 143.600 ; 
                RECT 360.880 143.280 391.120 143.600 ; 
                RECT 754.600 143.280 764.080 143.600 ; 
                RECT 0.160 144.640 202.760 144.960 ; 
                RECT 220.800 144.640 223.840 144.960 ; 
                RECT 227.600 144.640 310.200 144.960 ; 
                RECT 360.880 144.640 391.120 144.960 ; 
                RECT 754.600 144.640 764.080 144.960 ; 
                RECT 0.160 146.000 202.760 146.320 ; 
                RECT 220.800 146.000 310.200 146.320 ; 
                RECT 360.880 146.000 391.120 146.320 ; 
                RECT 754.600 146.000 764.080 146.320 ; 
                RECT 0.160 147.360 202.760 147.680 ; 
                RECT 220.800 147.360 310.200 147.680 ; 
                RECT 360.880 147.360 391.120 147.680 ; 
                RECT 754.600 147.360 764.080 147.680 ; 
                RECT 0.160 148.720 202.760 149.040 ; 
                RECT 220.800 148.720 391.120 149.040 ; 
                RECT 754.600 148.720 764.080 149.040 ; 
                RECT 0.160 150.080 202.760 150.400 ; 
                RECT 220.800 150.080 391.120 150.400 ; 
                RECT 754.600 150.080 764.080 150.400 ; 
                RECT 0.160 151.440 202.760 151.760 ; 
                RECT 220.800 151.440 229.280 151.760 ; 
                RECT 241.200 151.440 391.120 151.760 ; 
                RECT 754.600 151.440 764.080 151.760 ; 
                RECT 0.160 152.800 202.760 153.120 ; 
                RECT 220.800 152.800 225.880 153.120 ; 
                RECT 231.000 152.800 391.120 153.120 ; 
                RECT 754.600 152.800 764.080 153.120 ; 
                RECT 0.160 154.160 202.760 154.480 ; 
                RECT 220.800 154.160 297.280 154.480 ; 
                RECT 360.880 154.160 370.720 154.480 ; 
                RECT 754.600 154.160 764.080 154.480 ; 
                RECT 0.160 155.520 202.760 155.840 ; 
                RECT 220.800 155.520 297.280 155.840 ; 
                RECT 360.880 155.520 370.720 155.840 ; 
                RECT 754.600 155.520 764.080 155.840 ; 
                RECT 0.160 156.880 202.760 157.200 ; 
                RECT 220.800 156.880 297.280 157.200 ; 
                RECT 360.880 156.880 376.160 157.200 ; 
                RECT 754.600 156.880 764.080 157.200 ; 
                RECT 0.160 158.240 202.760 158.560 ; 
                RECT 220.800 158.240 297.280 158.560 ; 
                RECT 360.880 158.240 378.880 158.560 ; 
                RECT 754.600 158.240 764.080 158.560 ; 
                RECT 0.160 159.600 202.760 159.920 ; 
                RECT 220.800 159.600 225.200 159.920 ; 
                RECT 228.960 159.600 239.480 159.920 ; 
                RECT 241.880 159.600 297.280 159.920 ; 
                RECT 360.880 159.600 381.600 159.920 ; 
                RECT 754.600 159.600 764.080 159.920 ; 
                RECT 0.160 160.960 202.760 161.280 ; 
                RECT 220.800 160.960 297.280 161.280 ; 
                RECT 360.880 160.960 384.320 161.280 ; 
                RECT 754.600 160.960 764.080 161.280 ; 
                RECT 0.160 162.320 202.760 162.640 ; 
                RECT 220.800 162.320 228.600 162.640 ; 
                RECT 231.680 162.320 297.280 162.640 ; 
                RECT 360.880 162.320 387.040 162.640 ; 
                RECT 754.600 162.320 764.080 162.640 ; 
                RECT 0.160 163.680 202.760 164.000 ; 
                RECT 220.800 163.680 297.280 164.000 ; 
                RECT 360.880 163.680 389.760 164.000 ; 
                RECT 754.600 163.680 764.080 164.000 ; 
                RECT 0.160 165.040 202.760 165.360 ; 
                RECT 220.800 165.040 297.280 165.360 ; 
                RECT 754.600 165.040 764.080 165.360 ; 
                RECT 0.160 166.400 202.760 166.720 ; 
                RECT 220.800 166.400 297.280 166.720 ; 
                RECT 754.600 166.400 764.080 166.720 ; 
                RECT 0.160 167.760 202.760 168.080 ; 
                RECT 220.800 167.760 297.280 168.080 ; 
                RECT 360.880 167.760 391.120 168.080 ; 
                RECT 754.600 167.760 764.080 168.080 ; 
                RECT 0.160 169.120 202.760 169.440 ; 
                RECT 220.800 169.120 232.680 169.440 ; 
                RECT 241.200 169.120 297.280 169.440 ; 
                RECT 360.880 169.120 391.120 169.440 ; 
                RECT 754.600 169.120 764.080 169.440 ; 
                RECT 0.160 170.480 202.760 170.800 ; 
                RECT 220.800 170.480 297.280 170.800 ; 
                RECT 360.880 170.480 391.120 170.800 ; 
                RECT 754.600 170.480 764.080 170.800 ; 
                RECT 0.160 171.840 202.760 172.160 ; 
                RECT 220.800 171.840 297.280 172.160 ; 
                RECT 360.880 171.840 391.120 172.160 ; 
                RECT 754.600 171.840 764.080 172.160 ; 
                RECT 0.160 173.200 227.240 173.520 ; 
                RECT 231.680 173.200 297.280 173.520 ; 
                RECT 360.880 173.200 391.120 173.520 ; 
                RECT 754.600 173.200 764.080 173.520 ; 
                RECT 0.160 174.560 297.280 174.880 ; 
                RECT 360.880 174.560 391.120 174.880 ; 
                RECT 754.600 174.560 764.080 174.880 ; 
                RECT 0.160 175.920 181.680 176.240 ; 
                RECT 202.440 175.920 297.280 176.240 ; 
                RECT 360.880 175.920 391.120 176.240 ; 
                RECT 754.600 175.920 764.080 176.240 ; 
                RECT 0.160 177.280 181.680 177.600 ; 
                RECT 202.440 177.280 229.960 177.600 ; 
                RECT 235.760 177.280 297.280 177.600 ; 
                RECT 360.880 177.280 391.120 177.600 ; 
                RECT 754.600 177.280 764.080 177.600 ; 
                RECT 0.160 178.640 181.680 178.960 ; 
                RECT 202.440 178.640 208.200 178.960 ; 
                RECT 216.040 178.640 297.280 178.960 ; 
                RECT 360.880 178.640 391.120 178.960 ; 
                RECT 754.600 178.640 764.080 178.960 ; 
                RECT 0.160 180.000 181.680 180.320 ; 
                RECT 220.120 180.000 297.280 180.320 ; 
                RECT 360.880 180.000 391.120 180.320 ; 
                RECT 754.600 180.000 764.080 180.320 ; 
                RECT 0.160 181.360 181.680 181.680 ; 
                RECT 220.120 181.360 297.280 181.680 ; 
                RECT 754.600 181.360 764.080 181.680 ; 
                RECT 0.160 182.720 181.680 183.040 ; 
                RECT 202.440 182.720 208.200 183.040 ; 
                RECT 216.040 182.720 223.840 183.040 ; 
                RECT 234.400 182.720 297.280 183.040 ; 
                RECT 754.600 182.720 764.080 183.040 ; 
                RECT 0.160 184.080 168.760 184.400 ; 
                RECT 215.360 184.080 297.280 184.400 ; 
                RECT 360.880 184.080 764.080 184.400 ; 
                RECT 0.160 185.440 215.000 185.760 ; 
                RECT 294.920 185.440 764.080 185.760 ; 
                RECT 0.160 186.800 388.400 187.120 ; 
                RECT 756.640 186.800 764.080 187.120 ; 
                RECT 0.160 188.160 388.400 188.480 ; 
                RECT 756.640 188.160 764.080 188.480 ; 
                RECT 0.160 189.520 388.400 189.840 ; 
                RECT 756.640 189.520 764.080 189.840 ; 
                RECT 0.160 190.880 27.320 191.200 ; 
                RECT 33.800 190.880 36.160 191.200 ; 
                RECT 48.760 190.880 99.400 191.200 ; 
                RECT 756.640 190.880 764.080 191.200 ; 
                RECT 0.160 192.240 25.280 192.560 ; 
                RECT 35.840 192.240 37.520 192.560 ; 
                RECT 48.080 192.240 59.280 192.560 ; 
                RECT 61.000 192.240 75.600 192.560 ; 
                RECT 89.560 192.240 99.400 192.560 ; 
                RECT 756.640 192.240 764.080 192.560 ; 
                RECT 0.160 193.600 25.280 193.920 ; 
                RECT 35.840 193.600 59.280 193.920 ; 
                RECT 63.720 193.600 75.600 193.920 ; 
                RECT 89.560 193.600 99.400 193.920 ; 
                RECT 756.640 193.600 764.080 193.920 ; 
                RECT 0.160 194.960 25.280 195.280 ; 
                RECT 35.840 194.960 59.280 195.280 ; 
                RECT 63.720 194.960 75.600 195.280 ; 
                RECT 89.560 194.960 99.400 195.280 ; 
                RECT 756.640 194.960 764.080 195.280 ; 
                RECT 0.160 196.320 25.280 196.640 ; 
                RECT 35.840 196.320 59.280 196.640 ; 
                RECT 64.400 196.320 75.600 196.640 ; 
                RECT 89.560 196.320 99.400 196.640 ; 
                RECT 756.640 196.320 764.080 196.640 ; 
                RECT 0.160 197.680 25.280 198.000 ; 
                RECT 35.840 197.680 59.280 198.000 ; 
                RECT 61.000 197.680 75.600 198.000 ; 
                RECT 89.560 197.680 99.400 198.000 ; 
                RECT 756.640 197.680 764.080 198.000 ; 
                RECT 0.160 199.040 25.280 199.360 ; 
                RECT 35.840 199.040 99.400 199.360 ; 
                RECT 756.640 199.040 764.080 199.360 ; 
                RECT 0.160 200.400 25.280 200.720 ; 
                RECT 35.840 200.400 75.600 200.720 ; 
                RECT 89.560 200.400 99.400 200.720 ; 
                RECT 756.640 200.400 764.080 200.720 ; 
                RECT 0.160 201.760 75.600 202.080 ; 
                RECT 89.560 201.760 99.400 202.080 ; 
                RECT 756.640 201.760 764.080 202.080 ; 
                RECT 0.160 203.120 75.600 203.440 ; 
                RECT 89.560 203.120 99.400 203.440 ; 
                RECT 756.640 203.120 764.080 203.440 ; 
                RECT 0.160 204.480 18.480 204.800 ; 
                RECT 20.880 204.480 75.600 204.800 ; 
                RECT 89.560 204.480 99.400 204.800 ; 
                RECT 756.640 204.480 764.080 204.800 ; 
                RECT 0.160 205.840 75.600 206.160 ; 
                RECT 89.560 205.840 99.400 206.160 ; 
                RECT 756.640 205.840 764.080 206.160 ; 
                RECT 0.160 207.200 17.800 207.520 ; 
                RECT 20.880 207.200 34.120 207.520 ; 
                RECT 48.760 207.200 99.400 207.520 ; 
                RECT 756.640 207.200 764.080 207.520 ; 
                RECT 0.160 208.560 17.120 208.880 ; 
                RECT 20.880 208.560 34.120 208.880 ; 
                RECT 47.400 208.560 59.280 208.880 ; 
                RECT 61.000 208.560 75.600 208.880 ; 
                RECT 89.560 208.560 99.400 208.880 ; 
                RECT 756.640 208.560 764.080 208.880 ; 
                RECT 0.160 209.920 16.440 210.240 ; 
                RECT 20.880 209.920 34.120 210.240 ; 
                RECT 39.240 209.920 59.280 210.240 ; 
                RECT 61.680 209.920 75.600 210.240 ; 
                RECT 89.560 209.920 99.400 210.240 ; 
                RECT 756.640 209.920 764.080 210.240 ; 
                RECT 0.160 211.280 59.280 211.600 ; 
                RECT 62.360 211.280 75.600 211.600 ; 
                RECT 89.560 211.280 99.400 211.600 ; 
                RECT 756.640 211.280 764.080 211.600 ; 
                RECT 0.160 212.640 15.760 212.960 ; 
                RECT 20.880 212.640 34.120 212.960 ; 
                RECT 39.920 212.640 59.280 212.960 ; 
                RECT 62.360 212.640 75.600 212.960 ; 
                RECT 89.560 212.640 99.400 212.960 ; 
                RECT 756.640 212.640 764.080 212.960 ; 
                RECT 0.160 214.000 15.080 214.320 ; 
                RECT 20.880 214.000 34.120 214.320 ; 
                RECT 40.600 214.000 59.280 214.320 ; 
                RECT 63.040 214.000 75.600 214.320 ; 
                RECT 89.560 214.000 99.400 214.320 ; 
                RECT 756.640 214.000 764.080 214.320 ; 
                RECT 0.160 215.360 14.400 215.680 ; 
                RECT 20.880 215.360 99.400 215.680 ; 
                RECT 756.640 215.360 764.080 215.680 ; 
                RECT 0.160 216.720 13.720 217.040 ; 
                RECT 20.880 216.720 75.600 217.040 ; 
                RECT 89.560 216.720 99.400 217.040 ; 
                RECT 756.640 216.720 764.080 217.040 ; 
                RECT 0.160 218.080 75.600 218.400 ; 
                RECT 89.560 218.080 99.400 218.400 ; 
                RECT 756.640 218.080 764.080 218.400 ; 
                RECT 0.160 219.440 13.040 219.760 ; 
                RECT 20.880 219.440 75.600 219.760 ; 
                RECT 89.560 219.440 99.400 219.760 ; 
                RECT 756.640 219.440 764.080 219.760 ; 
                RECT 0.160 220.800 12.360 221.120 ; 
                RECT 20.880 220.800 75.600 221.120 ; 
                RECT 89.560 220.800 99.400 221.120 ; 
                RECT 756.640 220.800 764.080 221.120 ; 
                RECT 0.160 222.160 75.600 222.480 ; 
                RECT 85.480 222.160 99.400 222.480 ; 
                RECT 756.640 222.160 764.080 222.480 ; 
                RECT 0.160 223.520 11.680 223.840 ; 
                RECT 20.880 223.520 34.120 223.840 ; 
                RECT 39.240 223.520 80.360 223.840 ; 
                RECT 89.560 223.520 99.400 223.840 ; 
                RECT 756.640 223.520 764.080 223.840 ; 
                RECT 0.160 224.880 11.000 225.200 ; 
                RECT 20.880 224.880 34.120 225.200 ; 
                RECT 38.560 224.880 75.600 225.200 ; 
                RECT 89.560 224.880 99.400 225.200 ; 
                RECT 756.640 224.880 764.080 225.200 ; 
                RECT 0.160 226.240 75.600 226.560 ; 
                RECT 89.560 226.240 99.400 226.560 ; 
                RECT 756.640 226.240 764.080 226.560 ; 
                RECT 0.160 227.600 10.320 227.920 ; 
                RECT 20.880 227.600 34.120 227.920 ; 
                RECT 37.880 227.600 75.600 227.920 ; 
                RECT 89.560 227.600 99.400 227.920 ; 
                RECT 756.640 227.600 764.080 227.920 ; 
                RECT 0.160 228.960 9.640 229.280 ; 
                RECT 20.880 228.960 34.120 229.280 ; 
                RECT 37.200 228.960 75.600 229.280 ; 
                RECT 89.560 228.960 99.400 229.280 ; 
                RECT 756.640 228.960 764.080 229.280 ; 
                RECT 0.160 230.320 75.600 230.640 ; 
                RECT 86.160 230.320 99.400 230.640 ; 
                RECT 756.640 230.320 764.080 230.640 ; 
                RECT 0.160 231.680 75.600 232.000 ; 
                RECT 89.560 231.680 99.400 232.000 ; 
                RECT 756.640 231.680 764.080 232.000 ; 
                RECT 0.160 233.040 75.600 233.360 ; 
                RECT 89.560 233.040 99.400 233.360 ; 
                RECT 756.640 233.040 764.080 233.360 ; 
                RECT 0.160 234.400 75.600 234.720 ; 
                RECT 89.560 234.400 99.400 234.720 ; 
                RECT 756.640 234.400 764.080 234.720 ; 
                RECT 0.160 235.760 75.600 236.080 ; 
                RECT 89.560 235.760 99.400 236.080 ; 
                RECT 756.640 235.760 764.080 236.080 ; 
                RECT 0.160 237.120 75.600 237.440 ; 
                RECT 89.560 237.120 99.400 237.440 ; 
                RECT 756.640 237.120 764.080 237.440 ; 
                RECT 0.160 238.480 75.600 238.800 ; 
                RECT 87.520 238.480 99.400 238.800 ; 
                RECT 756.640 238.480 764.080 238.800 ; 
                RECT 0.160 239.840 75.600 240.160 ; 
                RECT 89.560 239.840 99.400 240.160 ; 
                RECT 756.640 239.840 764.080 240.160 ; 
                RECT 0.160 241.200 75.600 241.520 ; 
                RECT 89.560 241.200 99.400 241.520 ; 
                RECT 756.640 241.200 764.080 241.520 ; 
                RECT 0.160 242.560 75.600 242.880 ; 
                RECT 89.560 242.560 99.400 242.880 ; 
                RECT 756.640 242.560 764.080 242.880 ; 
                RECT 0.160 243.920 75.600 244.240 ; 
                RECT 89.560 243.920 99.400 244.240 ; 
                RECT 756.640 243.920 764.080 244.240 ; 
                RECT 0.160 245.280 75.600 245.600 ; 
                RECT 89.560 245.280 99.400 245.600 ; 
                RECT 756.640 245.280 764.080 245.600 ; 
                RECT 0.160 246.640 99.400 246.960 ; 
                RECT 756.640 246.640 764.080 246.960 ; 
                RECT 0.160 248.000 75.600 248.320 ; 
                RECT 89.560 248.000 99.400 248.320 ; 
                RECT 756.640 248.000 764.080 248.320 ; 
                RECT 0.160 249.360 75.600 249.680 ; 
                RECT 89.560 249.360 99.400 249.680 ; 
                RECT 756.640 249.360 764.080 249.680 ; 
                RECT 0.160 250.720 75.600 251.040 ; 
                RECT 89.560 250.720 99.400 251.040 ; 
                RECT 756.640 250.720 764.080 251.040 ; 
                RECT 0.160 252.080 75.600 252.400 ; 
                RECT 89.560 252.080 99.400 252.400 ; 
                RECT 756.640 252.080 764.080 252.400 ; 
                RECT 0.160 253.440 75.600 253.760 ; 
                RECT 89.560 253.440 99.400 253.760 ; 
                RECT 756.640 253.440 764.080 253.760 ; 
                RECT 0.160 254.800 99.400 255.120 ; 
                RECT 756.640 254.800 764.080 255.120 ; 
                RECT 0.160 256.160 77.640 256.480 ; 
                RECT 89.560 256.160 99.400 256.480 ; 
                RECT 756.640 256.160 764.080 256.480 ; 
                RECT 0.160 257.520 77.640 257.840 ; 
                RECT 89.560 257.520 99.400 257.840 ; 
                RECT 756.640 257.520 764.080 257.840 ; 
                RECT 0.160 258.880 77.640 259.200 ; 
                RECT 89.560 258.880 99.400 259.200 ; 
                RECT 756.640 258.880 764.080 259.200 ; 
                RECT 0.160 260.240 81.720 260.560 ; 
                RECT 89.560 260.240 99.400 260.560 ; 
                RECT 756.640 260.240 764.080 260.560 ; 
                RECT 0.160 261.600 77.640 261.920 ; 
                RECT 89.560 261.600 99.400 261.920 ; 
                RECT 756.640 261.600 764.080 261.920 ; 
                RECT 0.160 262.960 38.880 263.280 ; 
                RECT 65.080 262.960 99.400 263.280 ; 
                RECT 756.640 262.960 764.080 263.280 ; 
                RECT 0.160 264.320 37.520 264.640 ; 
                RECT 63.720 264.320 75.600 264.640 ; 
                RECT 89.560 264.320 99.400 264.640 ; 
                RECT 756.640 264.320 764.080 264.640 ; 
                RECT 0.160 265.680 36.160 266.000 ; 
                RECT 63.040 265.680 75.600 266.000 ; 
                RECT 89.560 265.680 99.400 266.000 ; 
                RECT 756.640 265.680 764.080 266.000 ; 
                RECT 0.160 267.040 77.640 267.360 ; 
                RECT 89.560 267.040 99.400 267.360 ; 
                RECT 756.640 267.040 764.080 267.360 ; 
                RECT 0.160 268.400 75.600 268.720 ; 
                RECT 89.560 268.400 99.400 268.720 ; 
                RECT 756.640 268.400 764.080 268.720 ; 
                RECT 0.160 269.760 75.600 270.080 ; 
                RECT 78.000 269.760 99.400 270.080 ; 
                RECT 756.640 269.760 764.080 270.080 ; 
                RECT 0.160 271.120 83.760 271.440 ; 
                RECT 89.560 271.120 99.400 271.440 ; 
                RECT 756.640 271.120 764.080 271.440 ; 
                RECT 0.160 272.480 75.600 272.800 ; 
                RECT 89.560 272.480 99.400 272.800 ; 
                RECT 756.640 272.480 764.080 272.800 ; 
                RECT 0.160 273.840 75.600 274.160 ; 
                RECT 89.560 273.840 99.400 274.160 ; 
                RECT 756.640 273.840 764.080 274.160 ; 
                RECT 0.160 275.200 75.600 275.520 ; 
                RECT 89.560 275.200 99.400 275.520 ; 
                RECT 756.640 275.200 764.080 275.520 ; 
                RECT 0.160 276.560 75.600 276.880 ; 
                RECT 89.560 276.560 99.400 276.880 ; 
                RECT 756.640 276.560 764.080 276.880 ; 
                RECT 0.160 277.920 75.600 278.240 ; 
                RECT 78.680 277.920 99.400 278.240 ; 
                RECT 756.640 277.920 764.080 278.240 ; 
                RECT 0.160 279.280 85.800 279.600 ; 
                RECT 89.560 279.280 99.400 279.600 ; 
                RECT 756.640 279.280 764.080 279.600 ; 
                RECT 0.160 280.640 75.600 280.960 ; 
                RECT 89.560 280.640 99.400 280.960 ; 
                RECT 756.640 280.640 764.080 280.960 ; 
                RECT 0.160 282.000 75.600 282.320 ; 
                RECT 89.560 282.000 99.400 282.320 ; 
                RECT 756.640 282.000 764.080 282.320 ; 
                RECT 0.160 283.360 75.600 283.680 ; 
                RECT 89.560 283.360 99.400 283.680 ; 
                RECT 756.640 283.360 764.080 283.680 ; 
                RECT 0.160 284.720 75.600 285.040 ; 
                RECT 89.560 284.720 99.400 285.040 ; 
                RECT 756.640 284.720 764.080 285.040 ; 
                RECT 0.160 286.080 99.400 286.400 ; 
                RECT 756.640 286.080 764.080 286.400 ; 
                RECT 0.160 287.440 77.640 287.760 ; 
                RECT 89.560 287.440 99.400 287.760 ; 
                RECT 756.640 287.440 764.080 287.760 ; 
                RECT 0.160 288.800 75.600 289.120 ; 
                RECT 89.560 288.800 99.400 289.120 ; 
                RECT 756.640 288.800 764.080 289.120 ; 
                RECT 0.160 290.160 75.600 290.480 ; 
                RECT 89.560 290.160 99.400 290.480 ; 
                RECT 756.640 290.160 764.080 290.480 ; 
                RECT 0.160 291.520 75.600 291.840 ; 
                RECT 89.560 291.520 99.400 291.840 ; 
                RECT 756.640 291.520 764.080 291.840 ; 
                RECT 0.160 292.880 75.600 293.200 ; 
                RECT 89.560 292.880 99.400 293.200 ; 
                RECT 756.640 292.880 764.080 293.200 ; 
                RECT 0.160 294.240 99.400 294.560 ; 
                RECT 756.640 294.240 764.080 294.560 ; 
                RECT 0.160 295.600 77.640 295.920 ; 
                RECT 89.560 295.600 99.400 295.920 ; 
                RECT 756.640 295.600 764.080 295.920 ; 
                RECT 0.160 296.960 75.600 297.280 ; 
                RECT 89.560 296.960 99.400 297.280 ; 
                RECT 756.640 296.960 764.080 297.280 ; 
                RECT 0.160 298.320 75.600 298.640 ; 
                RECT 89.560 298.320 99.400 298.640 ; 
                RECT 756.640 298.320 764.080 298.640 ; 
                RECT 0.160 299.680 75.600 300.000 ; 
                RECT 89.560 299.680 99.400 300.000 ; 
                RECT 756.640 299.680 764.080 300.000 ; 
                RECT 0.160 301.040 75.600 301.360 ; 
                RECT 89.560 301.040 99.400 301.360 ; 
                RECT 756.640 301.040 764.080 301.360 ; 
                RECT 0.160 302.400 99.400 302.720 ; 
                RECT 756.640 302.400 764.080 302.720 ; 
                RECT 0.160 303.760 75.600 304.080 ; 
                RECT 89.560 303.760 99.400 304.080 ; 
                RECT 756.640 303.760 764.080 304.080 ; 
                RECT 0.160 305.120 75.600 305.440 ; 
                RECT 89.560 305.120 99.400 305.440 ; 
                RECT 756.640 305.120 764.080 305.440 ; 
                RECT 0.160 306.480 77.640 306.800 ; 
                RECT 89.560 306.480 99.400 306.800 ; 
                RECT 756.640 306.480 764.080 306.800 ; 
                RECT 0.160 307.840 75.600 308.160 ; 
                RECT 89.560 307.840 99.400 308.160 ; 
                RECT 756.640 307.840 764.080 308.160 ; 
                RECT 0.160 309.200 75.600 309.520 ; 
                RECT 80.720 309.200 99.400 309.520 ; 
                RECT 756.640 309.200 764.080 309.520 ; 
                RECT 0.160 310.560 85.800 310.880 ; 
                RECT 89.560 310.560 99.400 310.880 ; 
                RECT 756.640 310.560 764.080 310.880 ; 
                RECT 0.160 311.920 75.600 312.240 ; 
                RECT 89.560 311.920 99.400 312.240 ; 
                RECT 756.640 311.920 764.080 312.240 ; 
                RECT 0.160 313.280 75.600 313.600 ; 
                RECT 89.560 313.280 99.400 313.600 ; 
                RECT 756.640 313.280 764.080 313.600 ; 
                RECT 0.160 314.640 75.600 314.960 ; 
                RECT 89.560 314.640 99.400 314.960 ; 
                RECT 756.640 314.640 764.080 314.960 ; 
                RECT 0.160 316.000 75.600 316.320 ; 
                RECT 89.560 316.000 99.400 316.320 ; 
                RECT 756.640 316.000 764.080 316.320 ; 
                RECT 0.160 317.360 75.600 317.680 ; 
                RECT 80.720 317.360 99.400 317.680 ; 
                RECT 756.640 317.360 764.080 317.680 ; 
                RECT 0.160 318.720 80.360 319.040 ; 
                RECT 89.560 318.720 99.400 319.040 ; 
                RECT 756.640 318.720 764.080 319.040 ; 
                RECT 0.160 320.080 75.600 320.400 ; 
                RECT 89.560 320.080 99.400 320.400 ; 
                RECT 756.640 320.080 764.080 320.400 ; 
                RECT 0.160 321.440 75.600 321.760 ; 
                RECT 89.560 321.440 99.400 321.760 ; 
                RECT 756.640 321.440 764.080 321.760 ; 
                RECT 0.160 322.800 75.600 323.120 ; 
                RECT 89.560 322.800 99.400 323.120 ; 
                RECT 756.640 322.800 764.080 323.120 ; 
                RECT 0.160 324.160 75.600 324.480 ; 
                RECT 89.560 324.160 99.400 324.480 ; 
                RECT 756.640 324.160 764.080 324.480 ; 
                RECT 0.160 325.520 99.400 325.840 ; 
                RECT 756.640 325.520 764.080 325.840 ; 
                RECT 0.160 326.880 78.320 327.200 ; 
                RECT 89.560 326.880 99.400 327.200 ; 
                RECT 756.640 326.880 764.080 327.200 ; 
                RECT 0.160 328.240 82.400 328.560 ; 
                RECT 89.560 328.240 99.400 328.560 ; 
                RECT 756.640 328.240 764.080 328.560 ; 
                RECT 0.160 329.600 83.080 329.920 ; 
                RECT 89.560 329.600 99.400 329.920 ; 
                RECT 756.640 329.600 764.080 329.920 ; 
                RECT 0.160 330.960 78.320 331.280 ; 
                RECT 89.560 330.960 99.400 331.280 ; 
                RECT 756.640 330.960 764.080 331.280 ; 
                RECT 0.160 332.320 78.320 332.640 ; 
                RECT 89.560 332.320 99.400 332.640 ; 
                RECT 756.640 332.320 764.080 332.640 ; 
                RECT 0.160 333.680 99.400 334.000 ; 
                RECT 756.640 333.680 764.080 334.000 ; 
                RECT 0.160 335.040 78.320 335.360 ; 
                RECT 89.560 335.040 99.400 335.360 ; 
                RECT 756.640 335.040 764.080 335.360 ; 
                RECT 0.160 336.400 78.320 336.720 ; 
                RECT 89.560 336.400 99.400 336.720 ; 
                RECT 756.640 336.400 764.080 336.720 ; 
                RECT 0.160 337.760 78.320 338.080 ; 
                RECT 89.560 337.760 99.400 338.080 ; 
                RECT 756.640 337.760 764.080 338.080 ; 
                RECT 0.160 339.120 85.800 339.440 ; 
                RECT 89.560 339.120 99.400 339.440 ; 
                RECT 756.640 339.120 764.080 339.440 ; 
                RECT 0.160 340.480 78.320 340.800 ; 
                RECT 89.560 340.480 99.400 340.800 ; 
                RECT 756.640 340.480 764.080 340.800 ; 
                RECT 0.160 341.840 99.400 342.160 ; 
                RECT 756.640 341.840 764.080 342.160 ; 
                RECT 0.160 343.200 78.320 343.520 ; 
                RECT 89.560 343.200 99.400 343.520 ; 
                RECT 756.640 343.200 764.080 343.520 ; 
                RECT 0.160 344.560 78.320 344.880 ; 
                RECT 89.560 344.560 99.400 344.880 ; 
                RECT 756.640 344.560 764.080 344.880 ; 
                RECT 0.160 345.920 78.320 346.240 ; 
                RECT 89.560 345.920 99.400 346.240 ; 
                RECT 756.640 345.920 764.080 346.240 ; 
                RECT 0.160 347.280 78.320 347.600 ; 
                RECT 89.560 347.280 99.400 347.600 ; 
                RECT 756.640 347.280 764.080 347.600 ; 
                RECT 0.160 348.640 99.400 348.960 ; 
                RECT 756.640 348.640 764.080 348.960 ; 
                RECT 0.160 350.000 80.360 350.320 ; 
                RECT 89.560 350.000 99.400 350.320 ; 
                RECT 756.640 350.000 764.080 350.320 ; 
                RECT 0.160 351.360 79.000 351.680 ; 
                RECT 89.560 351.360 99.400 351.680 ; 
                RECT 756.640 351.360 764.080 351.680 ; 
                RECT 0.160 352.720 79.000 353.040 ; 
                RECT 89.560 352.720 99.400 353.040 ; 
                RECT 756.640 352.720 764.080 353.040 ; 
                RECT 0.160 354.080 79.000 354.400 ; 
                RECT 89.560 354.080 99.400 354.400 ; 
                RECT 756.640 354.080 764.080 354.400 ; 
                RECT 0.160 355.440 79.000 355.760 ; 
                RECT 89.560 355.440 99.400 355.760 ; 
                RECT 756.640 355.440 764.080 355.760 ; 
                RECT 0.160 356.800 99.400 357.120 ; 
                RECT 756.640 356.800 764.080 357.120 ; 
                RECT 0.160 358.160 82.400 358.480 ; 
                RECT 89.560 358.160 99.400 358.480 ; 
                RECT 756.640 358.160 764.080 358.480 ; 
                RECT 0.160 359.520 79.000 359.840 ; 
                RECT 89.560 359.520 99.400 359.840 ; 
                RECT 756.640 359.520 764.080 359.840 ; 
                RECT 0.160 360.880 79.000 361.200 ; 
                RECT 89.560 360.880 99.400 361.200 ; 
                RECT 756.640 360.880 764.080 361.200 ; 
                RECT 0.160 362.240 79.000 362.560 ; 
                RECT 89.560 362.240 99.400 362.560 ; 
                RECT 756.640 362.240 764.080 362.560 ; 
                RECT 0.160 363.600 79.000 363.920 ; 
                RECT 89.560 363.600 99.400 363.920 ; 
                RECT 756.640 363.600 764.080 363.920 ; 
                RECT 0.160 364.960 99.400 365.280 ; 
                RECT 756.640 364.960 764.080 365.280 ; 
                RECT 0.160 366.320 79.000 366.640 ; 
                RECT 89.560 366.320 99.400 366.640 ; 
                RECT 756.640 366.320 764.080 366.640 ; 
                RECT 0.160 367.680 84.440 368.000 ; 
                RECT 89.560 367.680 99.400 368.000 ; 
                RECT 756.640 367.680 764.080 368.000 ; 
                RECT 0.160 369.040 79.000 369.360 ; 
                RECT 89.560 369.040 99.400 369.360 ; 
                RECT 756.640 369.040 764.080 369.360 ; 
                RECT 0.160 370.400 79.000 370.720 ; 
                RECT 89.560 370.400 99.400 370.720 ; 
                RECT 756.640 370.400 764.080 370.720 ; 
                RECT 0.160 371.760 79.000 372.080 ; 
                RECT 89.560 371.760 99.400 372.080 ; 
                RECT 756.640 371.760 764.080 372.080 ; 
                RECT 0.160 373.120 99.400 373.440 ; 
                RECT 756.640 373.120 764.080 373.440 ; 
                RECT 0.160 374.480 79.000 374.800 ; 
                RECT 89.560 374.480 99.400 374.800 ; 
                RECT 756.640 374.480 764.080 374.800 ; 
                RECT 0.160 375.840 79.000 376.160 ; 
                RECT 89.560 375.840 99.400 376.160 ; 
                RECT 756.640 375.840 764.080 376.160 ; 
                RECT 0.160 377.200 87.160 377.520 ; 
                RECT 89.560 377.200 99.400 377.520 ; 
                RECT 756.640 377.200 764.080 377.520 ; 
                RECT 0.160 378.560 87.160 378.880 ; 
                RECT 89.560 378.560 99.400 378.880 ; 
                RECT 756.640 378.560 764.080 378.880 ; 
                RECT 0.160 379.920 79.000 380.240 ; 
                RECT 89.560 379.920 99.400 380.240 ; 
                RECT 756.640 379.920 764.080 380.240 ; 
                RECT 0.160 381.280 99.400 381.600 ; 
                RECT 756.640 381.280 764.080 381.600 ; 
                RECT 0.160 382.640 79.000 382.960 ; 
                RECT 89.560 382.640 99.400 382.960 ; 
                RECT 756.640 382.640 764.080 382.960 ; 
                RECT 0.160 384.000 79.000 384.320 ; 
                RECT 89.560 384.000 99.400 384.320 ; 
                RECT 756.640 384.000 764.080 384.320 ; 
                RECT 0.160 385.360 79.000 385.680 ; 
                RECT 89.560 385.360 99.400 385.680 ; 
                RECT 756.640 385.360 764.080 385.680 ; 
                RECT 0.160 386.720 81.720 387.040 ; 
                RECT 89.560 386.720 99.400 387.040 ; 
                RECT 756.640 386.720 764.080 387.040 ; 
                RECT 0.160 388.080 99.400 388.400 ; 
                RECT 756.640 388.080 764.080 388.400 ; 
                RECT 0.160 389.440 82.400 389.760 ; 
                RECT 89.560 389.440 99.400 389.760 ; 
                RECT 756.640 389.440 764.080 389.760 ; 
                RECT 0.160 390.800 79.000 391.120 ; 
                RECT 89.560 390.800 99.400 391.120 ; 
                RECT 756.640 390.800 764.080 391.120 ; 
                RECT 0.160 392.160 79.000 392.480 ; 
                RECT 89.560 392.160 99.400 392.480 ; 
                RECT 756.640 392.160 764.080 392.480 ; 
                RECT 0.160 393.520 79.000 393.840 ; 
                RECT 89.560 393.520 99.400 393.840 ; 
                RECT 756.640 393.520 764.080 393.840 ; 
                RECT 0.160 394.880 79.000 395.200 ; 
                RECT 89.560 394.880 99.400 395.200 ; 
                RECT 756.640 394.880 764.080 395.200 ; 
                RECT 0.160 396.240 99.400 396.560 ; 
                RECT 756.640 396.240 764.080 396.560 ; 
                RECT 0.160 397.600 83.760 397.920 ; 
                RECT 89.560 397.600 99.400 397.920 ; 
                RECT 756.640 397.600 764.080 397.920 ; 
                RECT 0.160 398.960 79.000 399.280 ; 
                RECT 89.560 398.960 99.400 399.280 ; 
                RECT 756.640 398.960 764.080 399.280 ; 
                RECT 0.160 400.320 79.000 400.640 ; 
                RECT 89.560 400.320 99.400 400.640 ; 
                RECT 756.640 400.320 764.080 400.640 ; 
                RECT 0.160 401.680 79.000 402.000 ; 
                RECT 89.560 401.680 99.400 402.000 ; 
                RECT 756.640 401.680 764.080 402.000 ; 
                RECT 0.160 403.040 79.000 403.360 ; 
                RECT 89.560 403.040 99.400 403.360 ; 
                RECT 756.640 403.040 764.080 403.360 ; 
                RECT 0.160 404.400 99.400 404.720 ; 
                RECT 756.640 404.400 764.080 404.720 ; 
                RECT 0.160 405.760 79.000 406.080 ; 
                RECT 89.560 405.760 99.400 406.080 ; 
                RECT 756.640 405.760 764.080 406.080 ; 
                RECT 0.160 407.120 86.480 407.440 ; 
                RECT 89.560 407.120 99.400 407.440 ; 
                RECT 756.640 407.120 764.080 407.440 ; 
                RECT 0.160 408.480 79.000 408.800 ; 
                RECT 89.560 408.480 99.400 408.800 ; 
                RECT 756.640 408.480 764.080 408.800 ; 
                RECT 0.160 409.840 79.000 410.160 ; 
                RECT 89.560 409.840 99.400 410.160 ; 
                RECT 756.640 409.840 764.080 410.160 ; 
                RECT 0.160 411.200 79.000 411.520 ; 
                RECT 89.560 411.200 99.400 411.520 ; 
                RECT 756.640 411.200 764.080 411.520 ; 
                RECT 0.160 412.560 99.400 412.880 ; 
                RECT 756.640 412.560 764.080 412.880 ; 
                RECT 0.160 413.920 79.680 414.240 ; 
                RECT 89.560 413.920 99.400 414.240 ; 
                RECT 756.640 413.920 764.080 414.240 ; 
                RECT 0.160 415.280 79.680 415.600 ; 
                RECT 89.560 415.280 99.400 415.600 ; 
                RECT 756.640 415.280 764.080 415.600 ; 
                RECT 0.160 416.640 81.040 416.960 ; 
                RECT 89.560 416.640 99.400 416.960 ; 
                RECT 756.640 416.640 764.080 416.960 ; 
                RECT 0.160 418.000 79.680 418.320 ; 
                RECT 89.560 418.000 99.400 418.320 ; 
                RECT 756.640 418.000 764.080 418.320 ; 
                RECT 0.160 419.360 79.680 419.680 ; 
                RECT 89.560 419.360 99.400 419.680 ; 
                RECT 756.640 419.360 764.080 419.680 ; 
                RECT 0.160 420.720 99.400 421.040 ; 
                RECT 756.640 420.720 764.080 421.040 ; 
                RECT 0.160 422.080 79.680 422.400 ; 
                RECT 89.560 422.080 99.400 422.400 ; 
                RECT 756.640 422.080 764.080 422.400 ; 
                RECT 0.160 423.440 79.680 423.760 ; 
                RECT 89.560 423.440 99.400 423.760 ; 
                RECT 756.640 423.440 764.080 423.760 ; 
                RECT 0.160 424.800 79.680 425.120 ; 
                RECT 89.560 424.800 99.400 425.120 ; 
                RECT 756.640 424.800 764.080 425.120 ; 
                RECT 0.160 426.160 83.760 426.480 ; 
                RECT 89.560 426.160 99.400 426.480 ; 
                RECT 756.640 426.160 764.080 426.480 ; 
                RECT 0.160 427.520 79.680 427.840 ; 
                RECT 89.560 427.520 99.400 427.840 ; 
                RECT 756.640 427.520 764.080 427.840 ; 
                RECT 0.160 428.880 99.400 429.200 ; 
                RECT 756.640 428.880 764.080 429.200 ; 
                RECT 0.160 430.240 79.680 430.560 ; 
                RECT 89.560 430.240 99.400 430.560 ; 
                RECT 756.640 430.240 764.080 430.560 ; 
                RECT 0.160 431.600 79.680 431.920 ; 
                RECT 89.560 431.600 99.400 431.920 ; 
                RECT 756.640 431.600 764.080 431.920 ; 
                RECT 0.160 432.960 79.680 433.280 ; 
                RECT 89.560 432.960 99.400 433.280 ; 
                RECT 756.640 432.960 764.080 433.280 ; 
                RECT 0.160 434.320 79.680 434.640 ; 
                RECT 89.560 434.320 99.400 434.640 ; 
                RECT 756.640 434.320 764.080 434.640 ; 
                RECT 0.160 435.680 99.400 436.000 ; 
                RECT 756.640 435.680 764.080 436.000 ; 
                RECT 0.160 437.040 85.800 437.360 ; 
                RECT 89.560 437.040 99.400 437.360 ; 
                RECT 756.640 437.040 764.080 437.360 ; 
                RECT 0.160 438.400 79.680 438.720 ; 
                RECT 89.560 438.400 99.400 438.720 ; 
                RECT 756.640 438.400 764.080 438.720 ; 
                RECT 0.160 439.760 79.680 440.080 ; 
                RECT 89.560 439.760 99.400 440.080 ; 
                RECT 756.640 439.760 764.080 440.080 ; 
                RECT 0.160 441.120 79.680 441.440 ; 
                RECT 89.560 441.120 99.400 441.440 ; 
                RECT 756.640 441.120 764.080 441.440 ; 
                RECT 0.160 442.480 79.680 442.800 ; 
                RECT 89.560 442.480 99.400 442.800 ; 
                RECT 756.640 442.480 764.080 442.800 ; 
                RECT 0.160 443.840 99.400 444.160 ; 
                RECT 756.640 443.840 764.080 444.160 ; 
                RECT 0.160 445.200 99.400 445.520 ; 
                RECT 756.640 445.200 764.080 445.520 ; 
                RECT 0.160 446.560 388.400 446.880 ; 
                RECT 756.640 446.560 764.080 446.880 ; 
                RECT 0.160 447.920 388.400 448.240 ; 
                RECT 756.640 447.920 764.080 448.240 ; 
                RECT 0.160 449.280 764.080 449.600 ; 
                RECT 0.160 450.640 764.080 450.960 ; 
                RECT 0.160 452.000 764.080 452.320 ; 
                RECT 0.160 453.360 764.080 453.680 ; 
                RECT 0.160 454.720 764.080 455.040 ; 
                RECT 0.160 0.160 764.080 1.520 ; 
                RECT 0.160 458.760 764.080 460.120 ; 
                RECT 392.540 32.420 398.340 33.790 ; 
                RECT 746.840 32.420 752.640 33.790 ; 
                RECT 392.540 37.455 398.340 38.815 ; 
                RECT 746.840 37.455 752.640 38.815 ; 
                RECT 392.540 42.520 398.340 43.920 ; 
                RECT 746.840 42.520 752.640 43.920 ; 
                RECT 392.540 47.695 398.340 49.135 ; 
                RECT 746.840 47.695 752.640 49.135 ; 
                RECT 392.540 52.790 398.340 54.120 ; 
                RECT 746.840 52.790 752.640 54.120 ; 
                RECT 392.540 57.720 398.340 59.050 ; 
                RECT 746.840 57.720 752.640 59.050 ; 
                RECT 392.540 65.860 752.640 67.660 ; 
                RECT 392.540 135.175 752.640 136.975 ; 
                RECT 392.540 103.135 752.640 103.425 ; 
                RECT 392.540 173.365 752.640 176.965 ; 
                RECT 392.540 95.755 752.640 99.355 ; 
                RECT 392.540 80.340 752.640 81.140 ; 
                RECT 392.540 85.230 752.640 86.030 ; 
                RECT 392.540 77.330 752.640 78.130 ; 
                RECT 392.540 16.665 752.640 18.465 ; 
                RECT 103.590 190.595 105.510 444.975 ; 
                RECT 113.805 190.595 115.725 444.975 ; 
                RECT 117.645 190.595 119.565 444.975 ; 
                RECT 130.055 190.595 131.975 444.975 ; 
                RECT 133.895 190.595 135.815 444.975 ; 
                RECT 137.735 190.595 139.655 444.975 ; 
                RECT 141.575 190.595 143.495 444.975 ; 
                RECT 159.220 190.595 161.140 444.975 ; 
                RECT 163.060 190.595 164.980 444.975 ; 
                RECT 166.900 190.595 168.820 444.975 ; 
                RECT 170.740 190.595 172.660 444.975 ; 
                RECT 174.580 190.595 176.500 444.975 ; 
                RECT 178.420 190.595 180.340 444.975 ; 
                RECT 182.260 190.595 184.180 444.975 ; 
                RECT 209.070 190.595 210.990 444.975 ; 
                RECT 212.910 190.595 214.830 444.975 ; 
                RECT 216.750 190.595 218.670 444.975 ; 
                RECT 220.590 190.595 222.510 444.975 ; 
                RECT 224.430 190.595 226.350 444.975 ; 
                RECT 228.270 190.595 230.190 444.975 ; 
                RECT 232.110 190.595 234.030 444.975 ; 
                RECT 235.950 190.595 237.870 444.975 ; 
                RECT 239.790 190.595 241.710 444.975 ; 
                RECT 243.630 190.595 245.550 444.975 ; 
                RECT 247.470 190.595 249.390 444.975 ; 
                RECT 251.310 190.595 253.230 444.975 ; 
                RECT 255.150 190.595 257.070 444.975 ; 
                RECT 298.970 190.595 300.890 444.975 ; 
                RECT 302.810 190.595 304.730 444.975 ; 
                RECT 306.650 190.595 308.570 444.975 ; 
                RECT 310.490 190.595 312.410 444.975 ; 
                RECT 314.330 190.595 316.250 444.975 ; 
                RECT 318.170 190.595 320.090 444.975 ; 
                RECT 322.010 190.595 323.930 444.975 ; 
                RECT 325.850 190.595 327.770 444.975 ; 
                RECT 329.690 190.595 331.610 444.975 ; 
                RECT 333.530 190.595 335.450 444.975 ; 
                RECT 337.370 190.595 339.290 444.975 ; 
                RECT 341.210 190.595 343.130 444.975 ; 
                RECT 345.050 190.595 346.970 444.975 ; 
                RECT 348.890 190.595 350.810 444.975 ; 
                RECT 352.730 190.595 354.650 444.975 ; 
                RECT 356.570 190.595 358.490 444.975 ; 
                RECT 360.410 190.595 362.330 444.975 ; 
                RECT 364.250 190.595 366.170 444.975 ; 
                RECT 368.090 190.595 370.010 444.975 ; 
                RECT 371.930 190.595 373.850 444.975 ; 
                RECT 375.770 190.595 377.690 444.975 ; 
                RECT 379.610 190.595 381.530 444.975 ; 
                RECT 383.450 190.595 385.370 444.975 ; 
                RECT 266.265 61.535 268.185 114.135 ; 
                RECT 272.785 61.535 274.325 114.135 ; 
                RECT 281.720 61.535 283.640 114.135 ; 
                RECT 294.975 61.535 296.895 114.135 ; 
                RECT 298.815 61.535 300.735 114.135 ; 
                RECT 302.655 61.535 304.575 114.135 ; 
                RECT 306.495 61.535 308.415 114.135 ; 
                RECT 328.040 61.535 329.960 114.135 ; 
                RECT 331.880 61.535 333.800 114.135 ; 
                RECT 335.720 61.535 337.640 114.135 ; 
                RECT 339.560 61.535 341.480 114.135 ; 
                RECT 343.400 61.535 345.320 114.135 ; 
                RECT 347.240 61.535 349.160 114.135 ; 
                RECT 351.080 61.535 353.000 114.135 ; 
                RECT 354.920 61.535 356.840 114.135 ; 
                RECT 358.760 61.535 360.680 114.135 ; 
                RECT 301.720 153.680 303.640 183.960 ; 
                RECT 309.125 153.680 311.045 183.960 ; 
                RECT 315.755 153.680 317.505 183.960 ; 
                RECT 323.950 153.680 325.870 183.960 ; 
                RECT 327.790 153.680 329.710 183.960 ; 
                RECT 343.225 153.680 345.145 183.960 ; 
                RECT 347.065 153.680 348.985 183.960 ; 
                RECT 350.905 153.680 352.825 183.960 ; 
                RECT 354.745 153.680 356.665 183.960 ; 
                RECT 358.585 153.680 360.505 183.960 ; 
                RECT 314.380 142.520 316.300 147.680 ; 
                RECT 323.520 142.520 325.440 147.680 ; 
                RECT 327.360 142.520 329.280 147.680 ; 
                RECT 343.010 142.520 344.930 147.680 ; 
                RECT 346.850 142.520 348.770 147.680 ; 
                RECT 350.690 142.520 352.610 147.680 ; 
                RECT 354.530 142.520 356.450 147.680 ; 
                RECT 358.370 142.520 360.290 147.680 ; 
                RECT 359.525 51.955 361.445 55.535 ; 
                RECT 26.230 192.865 35.390 193.615 ; 
                RECT 26.230 198.265 35.390 200.185 ; 
                RECT 203.650 180.575 219.690 181.425 ; 
                RECT 182.050 180.275 201.690 182.985 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 404.040 5.560 ; 
                RECT 743.720 5.240 761.360 5.560 ; 
                RECT 2.880 6.600 761.360 6.920 ; 
                RECT 2.880 7.960 761.360 8.280 ; 
                RECT 2.880 9.320 761.360 9.640 ; 
                RECT 2.880 10.680 363.240 11.000 ; 
                RECT 754.600 10.680 761.360 11.000 ; 
                RECT 2.880 12.040 391.120 12.360 ; 
                RECT 754.600 12.040 761.360 12.360 ; 
                RECT 2.880 13.400 391.120 13.720 ; 
                RECT 754.600 13.400 761.360 13.720 ; 
                RECT 2.880 14.760 391.120 15.080 ; 
                RECT 754.600 14.760 761.360 15.080 ; 
                RECT 2.880 16.120 391.120 16.440 ; 
                RECT 754.600 16.120 761.360 16.440 ; 
                RECT 2.880 17.480 391.120 17.800 ; 
                RECT 754.600 17.480 761.360 17.800 ; 
                RECT 2.880 18.840 391.120 19.160 ; 
                RECT 754.600 18.840 761.360 19.160 ; 
                RECT 2.880 20.200 289.120 20.520 ; 
                RECT 364.960 20.200 391.120 20.520 ; 
                RECT 754.600 20.200 761.360 20.520 ; 
                RECT 2.880 21.560 391.120 21.880 ; 
                RECT 754.600 21.560 761.360 21.880 ; 
                RECT 2.880 22.920 391.120 23.240 ; 
                RECT 754.600 22.920 761.360 23.240 ; 
                RECT 2.880 24.280 391.120 24.600 ; 
                RECT 754.600 24.280 761.360 24.600 ; 
                RECT 2.880 25.640 289.120 25.960 ; 
                RECT 364.280 25.640 391.120 25.960 ; 
                RECT 754.600 25.640 761.360 25.960 ; 
                RECT 2.880 27.000 391.120 27.320 ; 
                RECT 754.600 27.000 761.360 27.320 ; 
                RECT 2.880 28.360 390.440 28.680 ; 
                RECT 754.600 28.360 761.360 28.680 ; 
                RECT 2.880 29.720 391.120 30.040 ; 
                RECT 754.600 29.720 761.360 30.040 ; 
                RECT 2.880 31.080 391.120 31.400 ; 
                RECT 754.600 31.080 761.360 31.400 ; 
                RECT 2.880 32.440 391.120 32.760 ; 
                RECT 754.600 32.440 761.360 32.760 ; 
                RECT 2.880 33.800 391.120 34.120 ; 
                RECT 754.600 33.800 761.360 34.120 ; 
                RECT 2.880 35.160 391.120 35.480 ; 
                RECT 754.600 35.160 761.360 35.480 ; 
                RECT 2.880 36.520 391.120 36.840 ; 
                RECT 754.600 36.520 761.360 36.840 ; 
                RECT 2.880 37.880 391.120 38.200 ; 
                RECT 754.600 37.880 761.360 38.200 ; 
                RECT 2.880 39.240 391.120 39.560 ; 
                RECT 754.600 39.240 761.360 39.560 ; 
                RECT 2.880 40.600 391.120 40.920 ; 
                RECT 754.600 40.600 761.360 40.920 ; 
                RECT 2.880 41.960 391.120 42.280 ; 
                RECT 754.600 41.960 761.360 42.280 ; 
                RECT 2.880 43.320 251.040 43.640 ; 
                RECT 335.720 43.320 391.120 43.640 ; 
                RECT 754.600 43.320 761.360 43.640 ; 
                RECT 2.880 44.680 249.680 45.000 ; 
                RECT 341.840 44.680 391.120 45.000 ; 
                RECT 754.600 44.680 761.360 45.000 ; 
                RECT 2.880 46.040 248.320 46.360 ; 
                RECT 347.960 46.040 391.120 46.360 ; 
                RECT 754.600 46.040 761.360 46.360 ; 
                RECT 2.880 47.400 228.600 47.720 ; 
                RECT 364.960 47.400 391.120 47.720 ; 
                RECT 754.600 47.400 761.360 47.720 ; 
                RECT 2.880 48.760 227.920 49.080 ; 
                RECT 360.880 48.760 391.120 49.080 ; 
                RECT 754.600 48.760 761.360 49.080 ; 
                RECT 2.880 50.120 391.120 50.440 ; 
                RECT 754.600 50.120 761.360 50.440 ; 
                RECT 2.880 51.480 355.760 51.800 ; 
                RECT 362.240 51.480 391.120 51.800 ; 
                RECT 754.600 51.480 761.360 51.800 ; 
                RECT 2.880 52.840 355.760 53.160 ; 
                RECT 362.240 52.840 391.120 53.160 ; 
                RECT 754.600 52.840 761.360 53.160 ; 
                RECT 2.880 54.200 355.760 54.520 ; 
                RECT 362.240 54.200 391.120 54.520 ; 
                RECT 754.600 54.200 761.360 54.520 ; 
                RECT 2.880 55.560 355.760 55.880 ; 
                RECT 362.240 55.560 391.120 55.880 ; 
                RECT 754.600 55.560 761.360 55.880 ; 
                RECT 2.880 56.920 391.120 57.240 ; 
                RECT 754.600 56.920 761.360 57.240 ; 
                RECT 2.880 58.280 391.120 58.600 ; 
                RECT 754.600 58.280 761.360 58.600 ; 
                RECT 2.880 59.640 391.120 59.960 ; 
                RECT 754.600 59.640 761.360 59.960 ; 
                RECT 2.880 61.000 263.280 61.320 ; 
                RECT 361.560 61.000 391.120 61.320 ; 
                RECT 754.600 61.000 761.360 61.320 ; 
                RECT 2.880 62.360 249.000 62.680 ; 
                RECT 256.160 62.360 263.280 62.680 ; 
                RECT 361.560 62.360 391.120 62.680 ; 
                RECT 754.600 62.360 761.360 62.680 ; 
                RECT 2.880 63.720 250.360 64.040 ; 
                RECT 254.800 63.720 263.280 64.040 ; 
                RECT 372.440 63.720 391.120 64.040 ; 
                RECT 754.600 63.720 761.360 64.040 ; 
                RECT 2.880 65.080 251.720 65.400 ; 
                RECT 254.120 65.080 263.280 65.400 ; 
                RECT 372.440 65.080 391.120 65.400 ; 
                RECT 754.600 65.080 761.360 65.400 ; 
                RECT 2.880 66.440 263.280 66.760 ; 
                RECT 361.560 66.440 391.120 66.760 ; 
                RECT 754.600 66.440 761.360 66.760 ; 
                RECT 2.880 67.800 263.280 68.120 ; 
                RECT 371.080 67.800 391.120 68.120 ; 
                RECT 754.600 67.800 761.360 68.120 ; 
                RECT 2.880 69.160 263.280 69.480 ; 
                RECT 375.160 69.160 391.120 69.480 ; 
                RECT 754.600 69.160 761.360 69.480 ; 
                RECT 2.880 70.520 263.280 70.840 ; 
                RECT 361.560 70.520 391.120 70.840 ; 
                RECT 754.600 70.520 761.360 70.840 ; 
                RECT 2.880 71.880 263.280 72.200 ; 
                RECT 375.160 71.880 391.120 72.200 ; 
                RECT 754.600 71.880 761.360 72.200 ; 
                RECT 2.880 73.240 263.280 73.560 ; 
                RECT 375.160 73.240 391.120 73.560 ; 
                RECT 754.600 73.240 761.360 73.560 ; 
                RECT 2.880 74.600 263.280 74.920 ; 
                RECT 373.800 74.600 391.120 74.920 ; 
                RECT 754.600 74.600 761.360 74.920 ; 
                RECT 2.880 75.960 263.280 76.280 ; 
                RECT 377.880 75.960 391.120 76.280 ; 
                RECT 754.600 75.960 761.360 76.280 ; 
                RECT 2.880 77.320 263.280 77.640 ; 
                RECT 377.880 77.320 391.120 77.640 ; 
                RECT 754.600 77.320 761.360 77.640 ; 
                RECT 2.880 78.680 263.280 79.000 ; 
                RECT 376.520 78.680 391.120 79.000 ; 
                RECT 754.600 78.680 761.360 79.000 ; 
                RECT 2.880 80.040 263.280 80.360 ; 
                RECT 377.880 80.040 391.120 80.360 ; 
                RECT 754.600 80.040 761.360 80.360 ; 
                RECT 2.880 81.400 263.280 81.720 ; 
                RECT 376.520 81.400 391.120 81.720 ; 
                RECT 754.600 81.400 761.360 81.720 ; 
                RECT 2.880 82.760 263.280 83.080 ; 
                RECT 380.600 82.760 391.120 83.080 ; 
                RECT 754.600 82.760 761.360 83.080 ; 
                RECT 2.880 84.120 263.280 84.440 ; 
                RECT 380.600 84.120 391.120 84.440 ; 
                RECT 754.600 84.120 761.360 84.440 ; 
                RECT 2.880 85.480 263.280 85.800 ; 
                RECT 379.240 85.480 391.120 85.800 ; 
                RECT 754.600 85.480 761.360 85.800 ; 
                RECT 2.880 86.840 223.840 87.160 ; 
                RECT 235.080 86.840 263.280 87.160 ; 
                RECT 380.600 86.840 391.120 87.160 ; 
                RECT 754.600 86.840 761.360 87.160 ; 
                RECT 2.880 88.200 225.200 88.520 ; 
                RECT 231.680 88.200 238.800 88.520 ; 
                RECT 241.200 88.200 263.280 88.520 ; 
                RECT 361.560 88.200 391.120 88.520 ; 
                RECT 754.600 88.200 761.360 88.520 ; 
                RECT 2.880 89.560 227.240 89.880 ; 
                RECT 230.320 89.560 263.280 89.880 ; 
                RECT 383.320 89.560 391.120 89.880 ; 
                RECT 754.600 89.560 761.360 89.880 ; 
                RECT 2.880 90.920 233.360 91.240 ; 
                RECT 240.520 90.920 263.280 91.240 ; 
                RECT 383.320 90.920 391.120 91.240 ; 
                RECT 754.600 90.920 761.360 91.240 ; 
                RECT 2.880 92.280 228.600 92.600 ; 
                RECT 235.080 92.280 236.080 92.600 ; 
                RECT 241.880 92.280 263.280 92.600 ; 
                RECT 361.560 92.280 391.120 92.600 ; 
                RECT 754.600 92.280 761.360 92.600 ; 
                RECT 2.880 93.640 225.880 93.960 ; 
                RECT 235.080 93.640 263.280 93.960 ; 
                RECT 381.960 93.640 391.120 93.960 ; 
                RECT 754.600 93.640 761.360 93.960 ; 
                RECT 2.880 95.000 263.280 95.320 ; 
                RECT 386.040 95.000 391.120 95.320 ; 
                RECT 754.600 95.000 761.360 95.320 ; 
                RECT 2.880 96.360 225.200 96.680 ; 
                RECT 228.280 96.360 263.280 96.680 ; 
                RECT 361.560 96.360 391.120 96.680 ; 
                RECT 754.600 96.360 761.360 96.680 ; 
                RECT 2.880 97.720 223.160 98.040 ; 
                RECT 241.200 97.720 263.280 98.040 ; 
                RECT 386.040 97.720 391.120 98.040 ; 
                RECT 754.600 97.720 761.360 98.040 ; 
                RECT 2.880 99.080 232.680 99.400 ; 
                RECT 235.080 99.080 263.280 99.400 ; 
                RECT 386.040 99.080 391.120 99.400 ; 
                RECT 754.600 99.080 761.360 99.400 ; 
                RECT 2.880 100.440 263.280 100.760 ; 
                RECT 384.680 100.440 391.120 100.760 ; 
                RECT 754.600 100.440 761.360 100.760 ; 
                RECT 2.880 101.800 233.360 102.120 ; 
                RECT 241.200 101.800 263.280 102.120 ; 
                RECT 388.760 101.800 391.120 102.120 ; 
                RECT 754.600 101.800 761.360 102.120 ; 
                RECT 2.880 103.160 229.960 103.480 ; 
                RECT 235.080 103.160 263.280 103.480 ; 
                RECT 388.760 103.160 391.120 103.480 ; 
                RECT 754.600 103.160 761.360 103.480 ; 
                RECT 2.880 104.520 232.680 104.840 ; 
                RECT 235.080 104.520 263.280 104.840 ; 
                RECT 387.400 104.520 391.120 104.840 ; 
                RECT 754.600 104.520 761.360 104.840 ; 
                RECT 2.880 105.880 263.280 106.200 ; 
                RECT 388.760 105.880 391.120 106.200 ; 
                RECT 754.600 105.880 761.360 106.200 ; 
                RECT 2.880 107.240 223.840 107.560 ; 
                RECT 246.640 107.240 263.280 107.560 ; 
                RECT 387.400 107.240 391.120 107.560 ; 
                RECT 754.600 107.240 761.360 107.560 ; 
                RECT 2.880 108.600 263.280 108.920 ; 
                RECT 754.600 108.600 761.360 108.920 ; 
                RECT 2.880 109.960 232.680 110.280 ; 
                RECT 235.080 109.960 240.840 110.280 ; 
                RECT 248.680 109.960 263.280 110.280 ; 
                RECT 754.600 109.960 761.360 110.280 ; 
                RECT 2.880 111.320 223.840 111.640 ; 
                RECT 237.800 111.320 263.280 111.640 ; 
                RECT 754.600 111.320 761.360 111.640 ; 
                RECT 2.880 112.680 232.680 113.000 ; 
                RECT 241.200 112.680 263.280 113.000 ; 
                RECT 754.600 112.680 761.360 113.000 ; 
                RECT 2.880 114.040 230.640 114.360 ; 
                RECT 234.400 114.040 263.280 114.360 ; 
                RECT 361.560 114.040 391.120 114.360 ; 
                RECT 754.600 114.040 761.360 114.360 ; 
                RECT 2.880 115.400 233.360 115.720 ; 
                RECT 241.880 115.400 391.120 115.720 ; 
                RECT 754.600 115.400 761.360 115.720 ; 
                RECT 2.880 116.760 366.640 117.080 ; 
                RECT 754.600 116.760 761.360 117.080 ; 
                RECT 2.880 118.120 226.560 118.440 ; 
                RECT 228.960 118.120 388.400 118.440 ; 
                RECT 754.600 118.120 761.360 118.440 ; 
                RECT 2.880 119.480 225.880 119.800 ; 
                RECT 235.080 119.480 385.680 119.800 ; 
                RECT 754.600 119.480 761.360 119.800 ; 
                RECT 2.880 120.840 382.960 121.160 ; 
                RECT 754.600 120.840 761.360 121.160 ; 
                RECT 2.880 122.200 232.680 122.520 ; 
                RECT 234.400 122.200 380.240 122.520 ; 
                RECT 754.600 122.200 761.360 122.520 ; 
                RECT 2.880 123.560 225.200 123.880 ; 
                RECT 235.760 123.560 377.520 123.880 ; 
                RECT 754.600 123.560 761.360 123.880 ; 
                RECT 2.880 124.920 229.960 125.240 ; 
                RECT 240.520 124.920 374.800 125.240 ; 
                RECT 754.600 124.920 761.360 125.240 ; 
                RECT 2.880 126.280 232.680 126.600 ; 
                RECT 234.400 126.280 372.080 126.600 ; 
                RECT 754.600 126.280 761.360 126.600 ; 
                RECT 2.880 127.640 227.240 127.960 ; 
                RECT 235.080 127.640 369.360 127.960 ; 
                RECT 754.600 127.640 761.360 127.960 ; 
                RECT 2.880 129.000 232.680 129.320 ; 
                RECT 235.760 129.000 391.120 129.320 ; 
                RECT 754.600 129.000 761.360 129.320 ; 
                RECT 2.880 130.360 223.840 130.680 ; 
                RECT 231.680 130.360 391.120 130.680 ; 
                RECT 754.600 130.360 761.360 130.680 ; 
                RECT 2.880 131.720 223.160 132.040 ; 
                RECT 241.200 131.720 391.120 132.040 ; 
                RECT 754.600 131.720 761.360 132.040 ; 
                RECT 2.880 133.080 202.760 133.400 ; 
                RECT 234.400 133.080 391.120 133.400 ; 
                RECT 754.600 133.080 761.360 133.400 ; 
                RECT 2.880 134.440 202.760 134.760 ; 
                RECT 220.800 134.440 223.840 134.760 ; 
                RECT 237.800 134.440 391.120 134.760 ; 
                RECT 754.600 134.440 761.360 134.760 ; 
                RECT 2.880 135.800 202.760 136.120 ; 
                RECT 220.800 135.800 391.120 136.120 ; 
                RECT 754.600 135.800 761.360 136.120 ; 
                RECT 2.880 137.160 202.760 137.480 ; 
                RECT 220.800 137.160 391.120 137.480 ; 
                RECT 754.600 137.160 761.360 137.480 ; 
                RECT 2.880 138.520 202.760 138.840 ; 
                RECT 220.800 138.520 236.080 138.840 ; 
                RECT 242.560 138.520 391.120 138.840 ; 
                RECT 754.600 138.520 761.360 138.840 ; 
                RECT 2.880 139.880 202.760 140.200 ; 
                RECT 220.800 139.880 239.480 140.200 ; 
                RECT 241.200 139.880 391.120 140.200 ; 
                RECT 754.600 139.880 761.360 140.200 ; 
                RECT 2.880 141.240 202.760 141.560 ; 
                RECT 220.800 141.240 391.120 141.560 ; 
                RECT 754.600 141.240 761.360 141.560 ; 
                RECT 2.880 142.600 202.760 142.920 ; 
                RECT 220.800 142.600 247.640 142.920 ; 
                RECT 307.160 142.600 310.200 142.920 ; 
                RECT 360.880 142.600 391.120 142.920 ; 
                RECT 754.600 142.600 761.360 142.920 ; 
                RECT 2.880 143.960 202.760 144.280 ; 
                RECT 220.800 143.960 223.840 144.280 ; 
                RECT 228.960 143.960 310.200 144.280 ; 
                RECT 360.880 143.960 391.120 144.280 ; 
                RECT 754.600 143.960 761.360 144.280 ; 
                RECT 2.880 145.320 202.760 145.640 ; 
                RECT 220.800 145.320 310.200 145.640 ; 
                RECT 360.880 145.320 391.120 145.640 ; 
                RECT 754.600 145.320 761.360 145.640 ; 
                RECT 2.880 146.680 202.760 147.000 ; 
                RECT 220.800 146.680 310.200 147.000 ; 
                RECT 360.880 146.680 391.120 147.000 ; 
                RECT 754.600 146.680 761.360 147.000 ; 
                RECT 2.880 148.040 202.760 148.360 ; 
                RECT 220.800 148.040 391.120 148.360 ; 
                RECT 754.600 148.040 761.360 148.360 ; 
                RECT 2.880 149.400 202.760 149.720 ; 
                RECT 220.800 149.400 391.120 149.720 ; 
                RECT 754.600 149.400 761.360 149.720 ; 
                RECT 2.880 150.760 202.760 151.080 ; 
                RECT 221.480 150.760 229.280 151.080 ; 
                RECT 241.200 150.760 391.120 151.080 ; 
                RECT 754.600 150.760 761.360 151.080 ; 
                RECT 2.880 152.120 202.760 152.440 ; 
                RECT 220.800 152.120 391.120 152.440 ; 
                RECT 754.600 152.120 761.360 152.440 ; 
                RECT 2.880 153.480 202.760 153.800 ; 
                RECT 220.800 153.480 225.880 153.800 ; 
                RECT 231.000 153.480 297.280 153.800 ; 
                RECT 360.880 153.480 391.120 153.800 ; 
                RECT 754.600 153.480 761.360 153.800 ; 
                RECT 2.880 154.840 202.760 155.160 ; 
                RECT 220.800 154.840 297.280 155.160 ; 
                RECT 360.880 154.840 370.720 155.160 ; 
                RECT 754.600 154.840 761.360 155.160 ; 
                RECT 2.880 156.200 202.760 156.520 ; 
                RECT 220.800 156.200 297.280 156.520 ; 
                RECT 360.880 156.200 373.440 156.520 ; 
                RECT 754.600 156.200 761.360 156.520 ; 
                RECT 2.880 157.560 202.760 157.880 ; 
                RECT 220.800 157.560 297.280 157.880 ; 
                RECT 360.880 157.560 376.160 157.880 ; 
                RECT 754.600 157.560 761.360 157.880 ; 
                RECT 2.880 158.920 202.760 159.240 ; 
                RECT 220.800 158.920 297.280 159.240 ; 
                RECT 360.880 158.920 378.880 159.240 ; 
                RECT 754.600 158.920 761.360 159.240 ; 
                RECT 2.880 160.280 202.760 160.600 ; 
                RECT 220.800 160.280 225.200 160.600 ; 
                RECT 228.960 160.280 239.480 160.600 ; 
                RECT 241.880 160.280 297.280 160.600 ; 
                RECT 360.880 160.280 381.600 160.600 ; 
                RECT 754.600 160.280 761.360 160.600 ; 
                RECT 2.880 161.640 202.760 161.960 ; 
                RECT 220.800 161.640 228.600 161.960 ; 
                RECT 231.680 161.640 297.280 161.960 ; 
                RECT 360.880 161.640 384.320 161.960 ; 
                RECT 754.600 161.640 761.360 161.960 ; 
                RECT 2.880 163.000 202.760 163.320 ; 
                RECT 220.800 163.000 297.280 163.320 ; 
                RECT 360.880 163.000 387.040 163.320 ; 
                RECT 754.600 163.000 761.360 163.320 ; 
                RECT 2.880 164.360 202.760 164.680 ; 
                RECT 220.800 164.360 297.280 164.680 ; 
                RECT 754.600 164.360 761.360 164.680 ; 
                RECT 2.880 165.720 202.760 166.040 ; 
                RECT 220.800 165.720 297.280 166.040 ; 
                RECT 754.600 165.720 761.360 166.040 ; 
                RECT 2.880 167.080 202.760 167.400 ; 
                RECT 220.800 167.080 297.280 167.400 ; 
                RECT 360.880 167.080 391.120 167.400 ; 
                RECT 754.600 167.080 761.360 167.400 ; 
                RECT 2.880 168.440 202.760 168.760 ; 
                RECT 220.800 168.440 232.680 168.760 ; 
                RECT 241.200 168.440 297.280 168.760 ; 
                RECT 360.880 168.440 391.120 168.760 ; 
                RECT 754.600 168.440 761.360 168.760 ; 
                RECT 2.880 169.800 202.760 170.120 ; 
                RECT 220.800 169.800 297.280 170.120 ; 
                RECT 360.880 169.800 391.120 170.120 ; 
                RECT 754.600 169.800 761.360 170.120 ; 
                RECT 2.880 171.160 202.760 171.480 ; 
                RECT 220.800 171.160 297.280 171.480 ; 
                RECT 360.880 171.160 391.120 171.480 ; 
                RECT 754.600 171.160 761.360 171.480 ; 
                RECT 2.880 172.520 227.240 172.840 ; 
                RECT 231.680 172.520 297.280 172.840 ; 
                RECT 360.880 172.520 391.120 172.840 ; 
                RECT 754.600 172.520 761.360 172.840 ; 
                RECT 2.880 173.880 297.280 174.200 ; 
                RECT 360.880 173.880 391.120 174.200 ; 
                RECT 754.600 173.880 761.360 174.200 ; 
                RECT 2.880 175.240 297.280 175.560 ; 
                RECT 360.880 175.240 391.120 175.560 ; 
                RECT 754.600 175.240 761.360 175.560 ; 
                RECT 2.880 176.600 181.680 176.920 ; 
                RECT 202.440 176.600 297.280 176.920 ; 
                RECT 360.880 176.600 391.120 176.920 ; 
                RECT 754.600 176.600 761.360 176.920 ; 
                RECT 2.880 177.960 181.680 178.280 ; 
                RECT 202.440 177.960 229.960 178.280 ; 
                RECT 235.760 177.960 297.280 178.280 ; 
                RECT 360.880 177.960 391.120 178.280 ; 
                RECT 754.600 177.960 761.360 178.280 ; 
                RECT 2.880 179.320 181.680 179.640 ; 
                RECT 202.440 179.320 208.200 179.640 ; 
                RECT 216.040 179.320 297.280 179.640 ; 
                RECT 360.880 179.320 391.120 179.640 ; 
                RECT 754.600 179.320 761.360 179.640 ; 
                RECT 2.880 180.680 181.680 181.000 ; 
                RECT 220.120 180.680 297.280 181.000 ; 
                RECT 754.600 180.680 761.360 181.000 ; 
                RECT 2.880 182.040 181.680 182.360 ; 
                RECT 202.440 182.040 297.280 182.360 ; 
                RECT 754.600 182.040 761.360 182.360 ; 
                RECT 2.880 183.400 168.760 183.720 ; 
                RECT 216.040 183.400 223.840 183.720 ; 
                RECT 234.400 183.400 297.280 183.720 ; 
                RECT 360.880 183.400 391.120 183.720 ; 
                RECT 754.600 183.400 761.360 183.720 ; 
                RECT 2.880 184.760 208.200 185.080 ; 
                RECT 228.960 184.760 761.360 185.080 ; 
                RECT 2.880 186.120 32.080 186.440 ; 
                RECT 227.600 186.120 761.360 186.440 ; 
                RECT 2.880 187.480 388.400 187.800 ; 
                RECT 756.640 187.480 761.360 187.800 ; 
                RECT 2.880 188.840 388.400 189.160 ; 
                RECT 756.640 188.840 761.360 189.160 ; 
                RECT 2.880 190.200 27.320 190.520 ; 
                RECT 33.800 190.200 99.400 190.520 ; 
                RECT 756.640 190.200 761.360 190.520 ; 
                RECT 2.880 191.560 25.280 191.880 ; 
                RECT 48.760 191.560 99.400 191.880 ; 
                RECT 756.640 191.560 761.360 191.880 ; 
                RECT 2.880 192.920 25.280 193.240 ; 
                RECT 47.400 192.920 59.280 193.240 ; 
                RECT 61.000 192.920 75.600 193.240 ; 
                RECT 89.560 192.920 99.400 193.240 ; 
                RECT 756.640 192.920 761.360 193.240 ; 
                RECT 2.880 194.280 59.280 194.600 ; 
                RECT 61.000 194.280 75.600 194.600 ; 
                RECT 89.560 194.280 99.400 194.600 ; 
                RECT 756.640 194.280 761.360 194.600 ; 
                RECT 2.880 195.640 25.280 195.960 ; 
                RECT 35.840 195.640 59.280 195.960 ; 
                RECT 63.720 195.640 75.600 195.960 ; 
                RECT 89.560 195.640 99.400 195.960 ; 
                RECT 756.640 195.640 761.360 195.960 ; 
                RECT 2.880 197.000 59.280 197.320 ; 
                RECT 64.400 197.000 75.600 197.320 ; 
                RECT 89.560 197.000 99.400 197.320 ; 
                RECT 756.640 197.000 761.360 197.320 ; 
                RECT 2.880 198.360 25.280 198.680 ; 
                RECT 35.840 198.360 59.280 198.680 ; 
                RECT 65.080 198.360 75.600 198.680 ; 
                RECT 89.560 198.360 99.400 198.680 ; 
                RECT 756.640 198.360 761.360 198.680 ; 
                RECT 2.880 199.720 25.280 200.040 ; 
                RECT 35.840 199.720 99.400 200.040 ; 
                RECT 756.640 199.720 761.360 200.040 ; 
                RECT 2.880 201.080 75.600 201.400 ; 
                RECT 89.560 201.080 99.400 201.400 ; 
                RECT 756.640 201.080 761.360 201.400 ; 
                RECT 2.880 202.440 75.600 202.760 ; 
                RECT 89.560 202.440 99.400 202.760 ; 
                RECT 756.640 202.440 761.360 202.760 ; 
                RECT 2.880 203.800 75.600 204.120 ; 
                RECT 89.560 203.800 99.400 204.120 ; 
                RECT 756.640 203.800 761.360 204.120 ; 
                RECT 2.880 205.160 18.480 205.480 ; 
                RECT 20.880 205.160 34.120 205.480 ; 
                RECT 37.200 205.160 75.600 205.480 ; 
                RECT 89.560 205.160 99.400 205.480 ; 
                RECT 756.640 205.160 761.360 205.480 ; 
                RECT 2.880 206.520 17.800 206.840 ; 
                RECT 20.880 206.520 38.880 206.840 ; 
                RECT 48.760 206.520 75.600 206.840 ; 
                RECT 83.440 206.520 99.400 206.840 ; 
                RECT 756.640 206.520 761.360 206.840 ; 
                RECT 2.880 207.880 17.120 208.200 ; 
                RECT 20.880 207.880 40.240 208.200 ; 
                RECT 48.080 207.880 83.760 208.200 ; 
                RECT 89.560 207.880 99.400 208.200 ; 
                RECT 756.640 207.880 761.360 208.200 ; 
                RECT 2.880 209.240 16.440 209.560 ; 
                RECT 20.880 209.240 59.280 209.560 ; 
                RECT 61.680 209.240 75.600 209.560 ; 
                RECT 89.560 209.240 99.400 209.560 ; 
                RECT 756.640 209.240 761.360 209.560 ; 
                RECT 2.880 210.600 59.280 210.920 ; 
                RECT 62.360 210.600 75.600 210.920 ; 
                RECT 89.560 210.600 99.400 210.920 ; 
                RECT 756.640 210.600 761.360 210.920 ; 
                RECT 2.880 211.960 15.760 212.280 ; 
                RECT 20.880 211.960 59.280 212.280 ; 
                RECT 62.360 211.960 75.600 212.280 ; 
                RECT 89.560 211.960 99.400 212.280 ; 
                RECT 756.640 211.960 761.360 212.280 ; 
                RECT 2.880 213.320 15.080 213.640 ; 
                RECT 20.880 213.320 59.280 213.640 ; 
                RECT 61.000 213.320 75.600 213.640 ; 
                RECT 89.560 213.320 99.400 213.640 ; 
                RECT 756.640 213.320 761.360 213.640 ; 
                RECT 2.880 214.680 59.280 215.000 ; 
                RECT 63.040 214.680 75.600 215.000 ; 
                RECT 84.120 214.680 99.400 215.000 ; 
                RECT 756.640 214.680 761.360 215.000 ; 
                RECT 2.880 216.040 14.400 216.360 ; 
                RECT 20.880 216.040 34.120 216.360 ; 
                RECT 41.280 216.040 75.600 216.360 ; 
                RECT 89.560 216.040 99.400 216.360 ; 
                RECT 756.640 216.040 761.360 216.360 ; 
                RECT 2.880 217.400 13.720 217.720 ; 
                RECT 20.880 217.400 34.120 217.720 ; 
                RECT 41.960 217.400 75.600 217.720 ; 
                RECT 89.560 217.400 99.400 217.720 ; 
                RECT 756.640 217.400 761.360 217.720 ; 
                RECT 2.880 218.760 75.600 219.080 ; 
                RECT 89.560 218.760 99.400 219.080 ; 
                RECT 756.640 218.760 761.360 219.080 ; 
                RECT 2.880 220.120 13.040 220.440 ; 
                RECT 20.880 220.120 34.120 220.440 ; 
                RECT 40.600 220.120 75.600 220.440 ; 
                RECT 89.560 220.120 99.400 220.440 ; 
                RECT 756.640 220.120 761.360 220.440 ; 
                RECT 2.880 221.480 12.360 221.800 ; 
                RECT 20.880 221.480 34.120 221.800 ; 
                RECT 39.920 221.480 75.600 221.800 ; 
                RECT 89.560 221.480 99.400 221.800 ; 
                RECT 756.640 221.480 761.360 221.800 ; 
                RECT 2.880 222.840 11.680 223.160 ; 
                RECT 20.880 222.840 99.400 223.160 ; 
                RECT 756.640 222.840 761.360 223.160 ; 
                RECT 2.880 224.200 11.000 224.520 ; 
                RECT 20.880 224.200 75.600 224.520 ; 
                RECT 89.560 224.200 99.400 224.520 ; 
                RECT 756.640 224.200 761.360 224.520 ; 
                RECT 2.880 225.560 75.600 225.880 ; 
                RECT 89.560 225.560 99.400 225.880 ; 
                RECT 756.640 225.560 761.360 225.880 ; 
                RECT 2.880 226.920 10.320 227.240 ; 
                RECT 20.880 226.920 75.600 227.240 ; 
                RECT 89.560 226.920 99.400 227.240 ; 
                RECT 756.640 226.920 761.360 227.240 ; 
                RECT 2.880 228.280 9.640 228.600 ; 
                RECT 20.880 228.280 75.600 228.600 ; 
                RECT 89.560 228.280 99.400 228.600 ; 
                RECT 756.640 228.280 761.360 228.600 ; 
                RECT 2.880 229.640 75.600 229.960 ; 
                RECT 89.560 229.640 99.400 229.960 ; 
                RECT 756.640 229.640 761.360 229.960 ; 
                RECT 2.880 231.000 99.400 231.320 ; 
                RECT 756.640 231.000 761.360 231.320 ; 
                RECT 2.880 232.360 75.600 232.680 ; 
                RECT 89.560 232.360 99.400 232.680 ; 
                RECT 756.640 232.360 761.360 232.680 ; 
                RECT 2.880 233.720 75.600 234.040 ; 
                RECT 89.560 233.720 99.400 234.040 ; 
                RECT 756.640 233.720 761.360 234.040 ; 
                RECT 2.880 235.080 75.600 235.400 ; 
                RECT 89.560 235.080 99.400 235.400 ; 
                RECT 756.640 235.080 761.360 235.400 ; 
                RECT 2.880 236.440 75.600 236.760 ; 
                RECT 89.560 236.440 99.400 236.760 ; 
                RECT 756.640 236.440 761.360 236.760 ; 
                RECT 2.880 237.800 75.600 238.120 ; 
                RECT 89.560 237.800 99.400 238.120 ; 
                RECT 756.640 237.800 761.360 238.120 ; 
                RECT 2.880 239.160 99.400 239.480 ; 
                RECT 756.640 239.160 761.360 239.480 ; 
                RECT 2.880 240.520 75.600 240.840 ; 
                RECT 89.560 240.520 99.400 240.840 ; 
                RECT 756.640 240.520 761.360 240.840 ; 
                RECT 2.880 241.880 75.600 242.200 ; 
                RECT 89.560 241.880 99.400 242.200 ; 
                RECT 756.640 241.880 761.360 242.200 ; 
                RECT 2.880 243.240 75.600 243.560 ; 
                RECT 89.560 243.240 99.400 243.560 ; 
                RECT 756.640 243.240 761.360 243.560 ; 
                RECT 2.880 244.600 75.600 244.920 ; 
                RECT 89.560 244.600 99.400 244.920 ; 
                RECT 756.640 244.600 761.360 244.920 ; 
                RECT 2.880 245.960 75.600 246.280 ; 
                RECT 88.200 245.960 99.400 246.280 ; 
                RECT 756.640 245.960 761.360 246.280 ; 
                RECT 2.880 247.320 85.800 247.640 ; 
                RECT 89.560 247.320 99.400 247.640 ; 
                RECT 756.640 247.320 761.360 247.640 ; 
                RECT 2.880 248.680 75.600 249.000 ; 
                RECT 89.560 248.680 99.400 249.000 ; 
                RECT 756.640 248.680 761.360 249.000 ; 
                RECT 2.880 250.040 75.600 250.360 ; 
                RECT 89.560 250.040 99.400 250.360 ; 
                RECT 756.640 250.040 761.360 250.360 ; 
                RECT 2.880 251.400 75.600 251.720 ; 
                RECT 89.560 251.400 99.400 251.720 ; 
                RECT 756.640 251.400 761.360 251.720 ; 
                RECT 2.880 252.760 75.600 253.080 ; 
                RECT 89.560 252.760 99.400 253.080 ; 
                RECT 756.640 252.760 761.360 253.080 ; 
                RECT 2.880 254.120 75.600 254.440 ; 
                RECT 88.880 254.120 99.400 254.440 ; 
                RECT 756.640 254.120 761.360 254.440 ; 
                RECT 2.880 255.480 80.360 255.800 ; 
                RECT 89.560 255.480 99.400 255.800 ; 
                RECT 756.640 255.480 761.360 255.800 ; 
                RECT 2.880 256.840 77.640 257.160 ; 
                RECT 89.560 256.840 99.400 257.160 ; 
                RECT 756.640 256.840 761.360 257.160 ; 
                RECT 2.880 258.200 77.640 258.520 ; 
                RECT 89.560 258.200 99.400 258.520 ; 
                RECT 756.640 258.200 761.360 258.520 ; 
                RECT 2.880 259.560 77.640 259.880 ; 
                RECT 89.560 259.560 99.400 259.880 ; 
                RECT 756.640 259.560 761.360 259.880 ; 
                RECT 2.880 260.920 77.640 261.240 ; 
                RECT 89.560 260.920 99.400 261.240 ; 
                RECT 756.640 260.920 761.360 261.240 ; 
                RECT 2.880 262.280 39.560 262.600 ; 
                RECT 65.080 262.280 99.400 262.600 ; 
                RECT 756.640 262.280 761.360 262.600 ; 
                RECT 2.880 263.640 38.200 263.960 ; 
                RECT 64.400 263.640 77.640 263.960 ; 
                RECT 89.560 263.640 99.400 263.960 ; 
                RECT 756.640 263.640 761.360 263.960 ; 
                RECT 2.880 265.000 36.840 265.320 ; 
                RECT 63.040 265.000 75.600 265.320 ; 
                RECT 89.560 265.000 99.400 265.320 ; 
                RECT 756.640 265.000 761.360 265.320 ; 
                RECT 2.880 266.360 75.600 266.680 ; 
                RECT 89.560 266.360 99.400 266.680 ; 
                RECT 756.640 266.360 761.360 266.680 ; 
                RECT 2.880 267.720 75.600 268.040 ; 
                RECT 89.560 267.720 99.400 268.040 ; 
                RECT 756.640 267.720 761.360 268.040 ; 
                RECT 2.880 269.080 75.600 269.400 ; 
                RECT 89.560 269.080 99.400 269.400 ; 
                RECT 756.640 269.080 761.360 269.400 ; 
                RECT 2.880 270.440 99.400 270.760 ; 
                RECT 756.640 270.440 761.360 270.760 ; 
                RECT 2.880 271.800 77.640 272.120 ; 
                RECT 89.560 271.800 99.400 272.120 ; 
                RECT 756.640 271.800 761.360 272.120 ; 
                RECT 2.880 273.160 75.600 273.480 ; 
                RECT 89.560 273.160 99.400 273.480 ; 
                RECT 756.640 273.160 761.360 273.480 ; 
                RECT 2.880 274.520 75.600 274.840 ; 
                RECT 89.560 274.520 99.400 274.840 ; 
                RECT 756.640 274.520 761.360 274.840 ; 
                RECT 2.880 275.880 75.600 276.200 ; 
                RECT 89.560 275.880 99.400 276.200 ; 
                RECT 756.640 275.880 761.360 276.200 ; 
                RECT 2.880 277.240 75.600 277.560 ; 
                RECT 89.560 277.240 99.400 277.560 ; 
                RECT 756.640 277.240 761.360 277.560 ; 
                RECT 2.880 278.600 99.400 278.920 ; 
                RECT 756.640 278.600 761.360 278.920 ; 
                RECT 2.880 279.960 75.600 280.280 ; 
                RECT 89.560 279.960 99.400 280.280 ; 
                RECT 756.640 279.960 761.360 280.280 ; 
                RECT 2.880 281.320 75.600 281.640 ; 
                RECT 89.560 281.320 99.400 281.640 ; 
                RECT 756.640 281.320 761.360 281.640 ; 
                RECT 2.880 282.680 75.600 283.000 ; 
                RECT 89.560 282.680 99.400 283.000 ; 
                RECT 756.640 282.680 761.360 283.000 ; 
                RECT 2.880 284.040 75.600 284.360 ; 
                RECT 89.560 284.040 99.400 284.360 ; 
                RECT 756.640 284.040 761.360 284.360 ; 
                RECT 2.880 285.400 75.600 285.720 ; 
                RECT 79.360 285.400 99.400 285.720 ; 
                RECT 756.640 285.400 761.360 285.720 ; 
                RECT 2.880 286.760 80.360 287.080 ; 
                RECT 89.560 286.760 99.400 287.080 ; 
                RECT 756.640 286.760 761.360 287.080 ; 
                RECT 2.880 288.120 75.600 288.440 ; 
                RECT 89.560 288.120 99.400 288.440 ; 
                RECT 756.640 288.120 761.360 288.440 ; 
                RECT 2.880 289.480 75.600 289.800 ; 
                RECT 89.560 289.480 99.400 289.800 ; 
                RECT 756.640 289.480 761.360 289.800 ; 
                RECT 2.880 290.840 77.640 291.160 ; 
                RECT 89.560 290.840 99.400 291.160 ; 
                RECT 756.640 290.840 761.360 291.160 ; 
                RECT 2.880 292.200 75.600 292.520 ; 
                RECT 89.560 292.200 99.400 292.520 ; 
                RECT 756.640 292.200 761.360 292.520 ; 
                RECT 2.880 293.560 75.600 293.880 ; 
                RECT 79.360 293.560 99.400 293.880 ; 
                RECT 756.640 293.560 761.360 293.880 ; 
                RECT 2.880 294.920 82.400 295.240 ; 
                RECT 89.560 294.920 99.400 295.240 ; 
                RECT 756.640 294.920 761.360 295.240 ; 
                RECT 2.880 296.280 75.600 296.600 ; 
                RECT 89.560 296.280 99.400 296.600 ; 
                RECT 756.640 296.280 761.360 296.600 ; 
                RECT 2.880 297.640 75.600 297.960 ; 
                RECT 89.560 297.640 99.400 297.960 ; 
                RECT 756.640 297.640 761.360 297.960 ; 
                RECT 2.880 299.000 75.600 299.320 ; 
                RECT 89.560 299.000 99.400 299.320 ; 
                RECT 756.640 299.000 761.360 299.320 ; 
                RECT 2.880 300.360 75.600 300.680 ; 
                RECT 89.560 300.360 99.400 300.680 ; 
                RECT 756.640 300.360 761.360 300.680 ; 
                RECT 2.880 301.720 99.400 302.040 ; 
                RECT 756.640 301.720 761.360 302.040 ; 
                RECT 2.880 303.080 77.640 303.400 ; 
                RECT 89.560 303.080 99.400 303.400 ; 
                RECT 756.640 303.080 761.360 303.400 ; 
                RECT 2.880 304.440 75.600 304.760 ; 
                RECT 89.560 304.440 99.400 304.760 ; 
                RECT 756.640 304.440 761.360 304.760 ; 
                RECT 2.880 305.800 75.600 306.120 ; 
                RECT 89.560 305.800 99.400 306.120 ; 
                RECT 756.640 305.800 761.360 306.120 ; 
                RECT 2.880 307.160 75.600 307.480 ; 
                RECT 89.560 307.160 99.400 307.480 ; 
                RECT 756.640 307.160 761.360 307.480 ; 
                RECT 2.880 308.520 75.600 308.840 ; 
                RECT 89.560 308.520 99.400 308.840 ; 
                RECT 756.640 308.520 761.360 308.840 ; 
                RECT 2.880 309.880 99.400 310.200 ; 
                RECT 756.640 309.880 761.360 310.200 ; 
                RECT 2.880 311.240 77.640 311.560 ; 
                RECT 89.560 311.240 99.400 311.560 ; 
                RECT 756.640 311.240 761.360 311.560 ; 
                RECT 2.880 312.600 75.600 312.920 ; 
                RECT 89.560 312.600 99.400 312.920 ; 
                RECT 756.640 312.600 761.360 312.920 ; 
                RECT 2.880 313.960 75.600 314.280 ; 
                RECT 89.560 313.960 99.400 314.280 ; 
                RECT 756.640 313.960 761.360 314.280 ; 
                RECT 2.880 315.320 75.600 315.640 ; 
                RECT 89.560 315.320 99.400 315.640 ; 
                RECT 756.640 315.320 761.360 315.640 ; 
                RECT 2.880 316.680 75.600 317.000 ; 
                RECT 89.560 316.680 99.400 317.000 ; 
                RECT 756.640 316.680 761.360 317.000 ; 
                RECT 2.880 318.040 99.400 318.360 ; 
                RECT 756.640 318.040 761.360 318.360 ; 
                RECT 2.880 319.400 75.600 319.720 ; 
                RECT 89.560 319.400 99.400 319.720 ; 
                RECT 756.640 319.400 761.360 319.720 ; 
                RECT 2.880 320.760 75.600 321.080 ; 
                RECT 89.560 320.760 99.400 321.080 ; 
                RECT 756.640 320.760 761.360 321.080 ; 
                RECT 2.880 322.120 75.600 322.440 ; 
                RECT 89.560 322.120 99.400 322.440 ; 
                RECT 756.640 322.120 761.360 322.440 ; 
                RECT 2.880 323.480 75.600 323.800 ; 
                RECT 89.560 323.480 99.400 323.800 ; 
                RECT 756.640 323.480 761.360 323.800 ; 
                RECT 2.880 324.840 75.600 325.160 ; 
                RECT 81.400 324.840 99.400 325.160 ; 
                RECT 756.640 324.840 761.360 325.160 ; 
                RECT 2.880 326.200 99.400 326.520 ; 
                RECT 756.640 326.200 761.360 326.520 ; 
                RECT 2.880 327.560 78.320 327.880 ; 
                RECT 89.560 327.560 99.400 327.880 ; 
                RECT 756.640 327.560 761.360 327.880 ; 
                RECT 2.880 328.920 78.320 329.240 ; 
                RECT 89.560 328.920 99.400 329.240 ; 
                RECT 756.640 328.920 761.360 329.240 ; 
                RECT 2.880 330.280 78.320 330.600 ; 
                RECT 89.560 330.280 99.400 330.600 ; 
                RECT 756.640 330.280 761.360 330.600 ; 
                RECT 2.880 331.640 78.320 331.960 ; 
                RECT 89.560 331.640 99.400 331.960 ; 
                RECT 756.640 331.640 761.360 331.960 ; 
                RECT 2.880 333.000 99.400 333.320 ; 
                RECT 756.640 333.000 761.360 333.320 ; 
                RECT 2.880 334.360 83.760 334.680 ; 
                RECT 89.560 334.360 99.400 334.680 ; 
                RECT 756.640 334.360 761.360 334.680 ; 
                RECT 2.880 335.720 78.320 336.040 ; 
                RECT 89.560 335.720 99.400 336.040 ; 
                RECT 756.640 335.720 761.360 336.040 ; 
                RECT 2.880 337.080 78.320 337.400 ; 
                RECT 89.560 337.080 99.400 337.400 ; 
                RECT 756.640 337.080 761.360 337.400 ; 
                RECT 2.880 338.440 78.320 338.760 ; 
                RECT 89.560 338.440 99.400 338.760 ; 
                RECT 756.640 338.440 761.360 338.760 ; 
                RECT 2.880 339.800 78.320 340.120 ; 
                RECT 89.560 339.800 99.400 340.120 ; 
                RECT 756.640 339.800 761.360 340.120 ; 
                RECT 2.880 341.160 99.400 341.480 ; 
                RECT 756.640 341.160 761.360 341.480 ; 
                RECT 2.880 342.520 78.320 342.840 ; 
                RECT 89.560 342.520 99.400 342.840 ; 
                RECT 756.640 342.520 761.360 342.840 ; 
                RECT 2.880 343.880 86.480 344.200 ; 
                RECT 89.560 343.880 99.400 344.200 ; 
                RECT 756.640 343.880 761.360 344.200 ; 
                RECT 2.880 345.240 78.320 345.560 ; 
                RECT 89.560 345.240 99.400 345.560 ; 
                RECT 756.640 345.240 761.360 345.560 ; 
                RECT 2.880 346.600 78.320 346.920 ; 
                RECT 89.560 346.600 99.400 346.920 ; 
                RECT 756.640 346.600 761.360 346.920 ; 
                RECT 2.880 347.960 78.320 348.280 ; 
                RECT 89.560 347.960 99.400 348.280 ; 
                RECT 756.640 347.960 761.360 348.280 ; 
                RECT 2.880 349.320 99.400 349.640 ; 
                RECT 756.640 349.320 761.360 349.640 ; 
                RECT 2.880 350.680 79.000 351.000 ; 
                RECT 89.560 350.680 99.400 351.000 ; 
                RECT 756.640 350.680 761.360 351.000 ; 
                RECT 2.880 352.040 79.000 352.360 ; 
                RECT 89.560 352.040 99.400 352.360 ; 
                RECT 756.640 352.040 761.360 352.360 ; 
                RECT 2.880 353.400 81.040 353.720 ; 
                RECT 89.560 353.400 99.400 353.720 ; 
                RECT 756.640 353.400 761.360 353.720 ; 
                RECT 2.880 354.760 79.000 355.080 ; 
                RECT 89.560 354.760 99.400 355.080 ; 
                RECT 756.640 354.760 761.360 355.080 ; 
                RECT 2.880 356.120 79.000 356.440 ; 
                RECT 89.560 356.120 99.400 356.440 ; 
                RECT 756.640 356.120 761.360 356.440 ; 
                RECT 2.880 357.480 99.400 357.800 ; 
                RECT 756.640 357.480 761.360 357.800 ; 
                RECT 2.880 358.840 79.000 359.160 ; 
                RECT 89.560 358.840 99.400 359.160 ; 
                RECT 756.640 358.840 761.360 359.160 ; 
                RECT 2.880 360.200 79.000 360.520 ; 
                RECT 89.560 360.200 99.400 360.520 ; 
                RECT 756.640 360.200 761.360 360.520 ; 
                RECT 2.880 361.560 79.000 361.880 ; 
                RECT 89.560 361.560 99.400 361.880 ; 
                RECT 756.640 361.560 761.360 361.880 ; 
                RECT 2.880 362.920 83.760 363.240 ; 
                RECT 89.560 362.920 99.400 363.240 ; 
                RECT 756.640 362.920 761.360 363.240 ; 
                RECT 2.880 364.280 79.000 364.600 ; 
                RECT 89.560 364.280 99.400 364.600 ; 
                RECT 756.640 364.280 761.360 364.600 ; 
                RECT 2.880 365.640 99.400 365.960 ; 
                RECT 756.640 365.640 761.360 365.960 ; 
                RECT 2.880 367.000 79.000 367.320 ; 
                RECT 89.560 367.000 99.400 367.320 ; 
                RECT 756.640 367.000 761.360 367.320 ; 
                RECT 2.880 368.360 79.000 368.680 ; 
                RECT 89.560 368.360 99.400 368.680 ; 
                RECT 756.640 368.360 761.360 368.680 ; 
                RECT 2.880 369.720 79.000 370.040 ; 
                RECT 89.560 369.720 99.400 370.040 ; 
                RECT 756.640 369.720 761.360 370.040 ; 
                RECT 2.880 371.080 79.000 371.400 ; 
                RECT 89.560 371.080 99.400 371.400 ; 
                RECT 756.640 371.080 761.360 371.400 ; 
                RECT 2.880 372.440 99.400 372.760 ; 
                RECT 756.640 372.440 761.360 372.760 ; 
                RECT 2.880 373.800 85.800 374.120 ; 
                RECT 89.560 373.800 99.400 374.120 ; 
                RECT 756.640 373.800 761.360 374.120 ; 
                RECT 2.880 375.160 79.000 375.480 ; 
                RECT 89.560 375.160 99.400 375.480 ; 
                RECT 756.640 375.160 761.360 375.480 ; 
                RECT 2.880 376.520 79.000 376.840 ; 
                RECT 89.560 376.520 99.400 376.840 ; 
                RECT 756.640 376.520 761.360 376.840 ; 
                RECT 2.880 377.880 79.000 378.200 ; 
                RECT 89.560 377.880 99.400 378.200 ; 
                RECT 756.640 377.880 761.360 378.200 ; 
                RECT 2.880 379.240 79.000 379.560 ; 
                RECT 89.560 379.240 99.400 379.560 ; 
                RECT 756.640 379.240 761.360 379.560 ; 
                RECT 2.880 380.600 99.400 380.920 ; 
                RECT 756.640 380.600 761.360 380.920 ; 
                RECT 2.880 381.960 80.360 382.280 ; 
                RECT 89.560 381.960 99.400 382.280 ; 
                RECT 756.640 381.960 761.360 382.280 ; 
                RECT 2.880 383.320 81.040 383.640 ; 
                RECT 89.560 383.320 99.400 383.640 ; 
                RECT 756.640 383.320 761.360 383.640 ; 
                RECT 2.880 384.680 79.000 385.000 ; 
                RECT 89.560 384.680 99.400 385.000 ; 
                RECT 756.640 384.680 761.360 385.000 ; 
                RECT 2.880 386.040 79.000 386.360 ; 
                RECT 89.560 386.040 99.400 386.360 ; 
                RECT 756.640 386.040 761.360 386.360 ; 
                RECT 2.880 387.400 79.000 387.720 ; 
                RECT 89.560 387.400 99.400 387.720 ; 
                RECT 756.640 387.400 761.360 387.720 ; 
                RECT 2.880 388.760 99.400 389.080 ; 
                RECT 756.640 388.760 761.360 389.080 ; 
                RECT 2.880 390.120 79.000 390.440 ; 
                RECT 89.560 390.120 99.400 390.440 ; 
                RECT 756.640 390.120 761.360 390.440 ; 
                RECT 2.880 391.480 79.000 391.800 ; 
                RECT 89.560 391.480 99.400 391.800 ; 
                RECT 756.640 391.480 761.360 391.800 ; 
                RECT 2.880 392.840 83.080 393.160 ; 
                RECT 89.560 392.840 99.400 393.160 ; 
                RECT 756.640 392.840 761.360 393.160 ; 
                RECT 2.880 394.200 79.000 394.520 ; 
                RECT 89.560 394.200 99.400 394.520 ; 
                RECT 756.640 394.200 761.360 394.520 ; 
                RECT 2.880 395.560 79.000 395.880 ; 
                RECT 89.560 395.560 99.400 395.880 ; 
                RECT 756.640 395.560 761.360 395.880 ; 
                RECT 2.880 396.920 99.400 397.240 ; 
                RECT 756.640 396.920 761.360 397.240 ; 
                RECT 2.880 398.280 79.000 398.600 ; 
                RECT 89.560 398.280 99.400 398.600 ; 
                RECT 756.640 398.280 761.360 398.600 ; 
                RECT 2.880 399.640 79.000 399.960 ; 
                RECT 89.560 399.640 99.400 399.960 ; 
                RECT 756.640 399.640 761.360 399.960 ; 
                RECT 2.880 401.000 79.000 401.320 ; 
                RECT 89.560 401.000 99.400 401.320 ; 
                RECT 756.640 401.000 761.360 401.320 ; 
                RECT 2.880 402.360 85.800 402.680 ; 
                RECT 89.560 402.360 99.400 402.680 ; 
                RECT 756.640 402.360 761.360 402.680 ; 
                RECT 2.880 403.720 79.000 404.040 ; 
                RECT 89.560 403.720 99.400 404.040 ; 
                RECT 756.640 403.720 761.360 404.040 ; 
                RECT 2.880 405.080 99.400 405.400 ; 
                RECT 756.640 405.080 761.360 405.400 ; 
                RECT 2.880 406.440 79.000 406.760 ; 
                RECT 89.560 406.440 99.400 406.760 ; 
                RECT 756.640 406.440 761.360 406.760 ; 
                RECT 2.880 407.800 79.000 408.120 ; 
                RECT 89.560 407.800 99.400 408.120 ; 
                RECT 756.640 407.800 761.360 408.120 ; 
                RECT 2.880 409.160 79.000 409.480 ; 
                RECT 89.560 409.160 99.400 409.480 ; 
                RECT 756.640 409.160 761.360 409.480 ; 
                RECT 2.880 410.520 79.000 410.840 ; 
                RECT 89.560 410.520 99.400 410.840 ; 
                RECT 756.640 410.520 761.360 410.840 ; 
                RECT 2.880 411.880 99.400 412.200 ; 
                RECT 756.640 411.880 761.360 412.200 ; 
                RECT 2.880 413.240 80.360 413.560 ; 
                RECT 89.560 413.240 99.400 413.560 ; 
                RECT 756.640 413.240 761.360 413.560 ; 
                RECT 2.880 414.600 79.680 414.920 ; 
                RECT 89.560 414.600 99.400 414.920 ; 
                RECT 756.640 414.600 761.360 414.920 ; 
                RECT 2.880 415.960 79.680 416.280 ; 
                RECT 89.560 415.960 99.400 416.280 ; 
                RECT 756.640 415.960 761.360 416.280 ; 
                RECT 2.880 417.320 79.680 417.640 ; 
                RECT 89.560 417.320 99.400 417.640 ; 
                RECT 756.640 417.320 761.360 417.640 ; 
                RECT 2.880 418.680 79.680 419.000 ; 
                RECT 89.560 418.680 99.400 419.000 ; 
                RECT 756.640 418.680 761.360 419.000 ; 
                RECT 2.880 420.040 99.400 420.360 ; 
                RECT 756.640 420.040 761.360 420.360 ; 
                RECT 2.880 421.400 82.400 421.720 ; 
                RECT 89.560 421.400 99.400 421.720 ; 
                RECT 756.640 421.400 761.360 421.720 ; 
                RECT 2.880 422.760 79.680 423.080 ; 
                RECT 89.560 422.760 99.400 423.080 ; 
                RECT 756.640 422.760 761.360 423.080 ; 
                RECT 2.880 424.120 79.680 424.440 ; 
                RECT 89.560 424.120 99.400 424.440 ; 
                RECT 756.640 424.120 761.360 424.440 ; 
                RECT 2.880 425.480 79.680 425.800 ; 
                RECT 89.560 425.480 99.400 425.800 ; 
                RECT 756.640 425.480 761.360 425.800 ; 
                RECT 2.880 426.840 79.680 427.160 ; 
                RECT 89.560 426.840 99.400 427.160 ; 
                RECT 756.640 426.840 761.360 427.160 ; 
                RECT 2.880 428.200 99.400 428.520 ; 
                RECT 756.640 428.200 761.360 428.520 ; 
                RECT 2.880 429.560 79.680 429.880 ; 
                RECT 89.560 429.560 99.400 429.880 ; 
                RECT 756.640 429.560 761.360 429.880 ; 
                RECT 2.880 430.920 84.440 431.240 ; 
                RECT 89.560 430.920 99.400 431.240 ; 
                RECT 756.640 430.920 761.360 431.240 ; 
                RECT 2.880 432.280 85.120 432.600 ; 
                RECT 89.560 432.280 99.400 432.600 ; 
                RECT 756.640 432.280 761.360 432.600 ; 
                RECT 2.880 433.640 79.680 433.960 ; 
                RECT 89.560 433.640 99.400 433.960 ; 
                RECT 756.640 433.640 761.360 433.960 ; 
                RECT 2.880 435.000 79.680 435.320 ; 
                RECT 89.560 435.000 99.400 435.320 ; 
                RECT 756.640 435.000 761.360 435.320 ; 
                RECT 2.880 436.360 99.400 436.680 ; 
                RECT 756.640 436.360 761.360 436.680 ; 
                RECT 2.880 437.720 79.680 438.040 ; 
                RECT 89.560 437.720 99.400 438.040 ; 
                RECT 756.640 437.720 761.360 438.040 ; 
                RECT 2.880 439.080 79.680 439.400 ; 
                RECT 89.560 439.080 99.400 439.400 ; 
                RECT 756.640 439.080 761.360 439.400 ; 
                RECT 2.880 440.440 87.160 440.760 ; 
                RECT 89.560 440.440 99.400 440.760 ; 
                RECT 756.640 440.440 761.360 440.760 ; 
                RECT 2.880 441.800 87.160 442.120 ; 
                RECT 89.560 441.800 99.400 442.120 ; 
                RECT 756.640 441.800 761.360 442.120 ; 
                RECT 2.880 443.160 79.680 443.480 ; 
                RECT 89.560 443.160 99.400 443.480 ; 
                RECT 756.640 443.160 761.360 443.480 ; 
                RECT 2.880 444.520 99.400 444.840 ; 
                RECT 756.640 444.520 761.360 444.840 ; 
                RECT 2.880 445.880 388.400 446.200 ; 
                RECT 756.640 445.880 761.360 446.200 ; 
                RECT 2.880 447.240 388.400 447.560 ; 
                RECT 756.640 447.240 761.360 447.560 ; 
                RECT 2.880 448.600 388.400 448.920 ; 
                RECT 756.640 448.600 761.360 448.920 ; 
                RECT 2.880 449.960 761.360 450.280 ; 
                RECT 2.880 451.320 761.360 451.640 ; 
                RECT 2.880 452.680 761.360 453.000 ; 
                RECT 2.880 454.040 761.360 454.360 ; 
                RECT 2.880 2.880 761.360 4.240 ; 
                RECT 2.880 456.040 761.360 457.400 ; 
                RECT 392.540 29.775 398.340 30.895 ; 
                RECT 746.840 29.775 752.640 30.895 ; 
                RECT 392.540 35.565 398.340 36.185 ; 
                RECT 746.840 35.565 752.640 36.185 ; 
                RECT 392.540 40.590 398.340 41.230 ; 
                RECT 746.840 40.590 752.640 41.230 ; 
                RECT 392.540 45.720 398.340 46.370 ; 
                RECT 746.840 45.720 752.640 46.370 ; 
                RECT 392.540 50.935 398.340 51.545 ; 
                RECT 746.840 50.935 752.640 51.545 ; 
                RECT 392.540 55.865 398.340 56.475 ; 
                RECT 746.840 55.865 752.640 56.475 ; 
                RECT 392.540 81.660 752.640 82.460 ; 
                RECT 392.540 90.235 752.640 93.835 ; 
                RECT 392.540 86.550 752.640 87.350 ; 
                RECT 392.540 147.905 752.640 149.705 ; 
                RECT 392.540 115.695 752.640 115.985 ; 
                RECT 392.540 78.650 752.640 79.450 ; 
                RECT 392.540 69.600 752.640 71.400 ; 
                RECT 392.540 83.340 752.640 84.140 ; 
                RECT 392.540 20.405 752.640 22.205 ; 
                RECT 99.995 190.595 101.105 444.975 ; 
                RECT 108.930 190.595 110.850 444.975 ; 
                RECT 124.290 190.595 126.210 444.975 ; 
                RECT 146.560 190.595 148.480 444.975 ; 
                RECT 150.400 190.595 152.320 444.975 ; 
                RECT 154.240 190.595 156.160 444.975 ; 
                RECT 188.395 190.595 190.315 444.975 ; 
                RECT 192.235 190.595 194.155 444.975 ; 
                RECT 196.075 190.595 197.995 444.975 ; 
                RECT 199.915 190.595 201.835 444.975 ; 
                RECT 203.755 190.595 205.675 444.975 ; 
                RECT 261.435 190.595 263.355 444.975 ; 
                RECT 265.275 190.595 267.195 444.975 ; 
                RECT 269.115 190.595 271.035 444.975 ; 
                RECT 272.955 190.595 274.875 444.975 ; 
                RECT 276.795 190.595 278.715 444.975 ; 
                RECT 280.635 190.595 282.555 444.975 ; 
                RECT 284.475 190.595 286.395 444.975 ; 
                RECT 288.315 190.595 290.235 444.975 ; 
                RECT 292.155 190.595 294.075 444.975 ; 
                RECT 263.640 61.535 264.530 114.135 ; 
                RECT 270.400 61.535 271.290 114.135 ; 
                RECT 276.620 61.535 278.160 114.135 ; 
                RECT 289.210 61.535 291.130 114.135 ; 
                RECT 313.200 61.535 315.120 114.135 ; 
                RECT 317.040 61.535 318.960 114.135 ; 
                RECT 320.880 61.535 322.800 114.135 ; 
                RECT 298.125 153.680 299.235 183.960 ; 
                RECT 306.500 153.680 307.390 183.960 ; 
                RECT 313.260 153.680 314.150 183.960 ; 
                RECT 320.020 153.680 321.770 183.960 ; 
                RECT 333.160 153.680 335.080 183.960 ; 
                RECT 337.000 153.680 338.920 183.960 ; 
                RECT 310.785 142.520 311.895 147.680 ; 
                RECT 319.590 142.520 321.340 147.680 ; 
                RECT 332.730 142.520 334.650 147.680 ; 
                RECT 336.570 142.520 338.490 147.680 ; 
                RECT 356.145 51.955 357.255 55.535 ; 
                RECT 26.230 191.660 35.390 192.030 ; 
                RECT 26.230 195.100 35.390 196.210 ; 
                RECT 182.050 176.120 201.690 176.790 ; 
                RECT 182.050 177.455 201.690 179.145 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 764.240 460.280 ; 
        LAYER met2 ;
            RECT 0.000 0.000 764.240 460.280 ; 
    END 
END sram22_1024x32m8w8 
END LIBRARY 

