VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sramgen_sram_1024x32m8w8_replica_v1
  CLASS BLOCK ;
  ORIGIN 84.035 353.63 ;
  FOREIGN sramgen_sram_1024x32m8w8_replica_v1 -84.035 -353.63 ;
  SIZE 746.495 BY 365.345 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -78.6 -353.23 -78.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -77 -353.23 -76.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -75.4 -353.23 -75 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.8 -353.23 -73.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.2 -353.23 -71.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.6 -323.62 -70.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -69 -340.58 -68.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -339.52 -67 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -353.23 -67 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.8 -353.23 -65.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -335.28 -63.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -353.23 -63.8 -342.06 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.6 -339.52 -62.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -61 -353.23 -60.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -334.22 -59 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -353.23 -59 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.8 -340.58 -57.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -339.52 -55.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -353.23 -55.8 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.6 -353.23 -54.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -333.16 -52.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -353.23 -52.6 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.4 -340.58 -51 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -339.52 -49.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -353.23 -49.4 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.2 -353.23 -47.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -333.16 -46.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -353.23 -46.2 -342.06 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -339.52 -44.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -353.23 -44.6 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.4 -353.23 -43 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -331.04 -41.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -353.23 -41.4 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.2 -340.58 -39.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -339.52 -38.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -353.23 -38.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -37 -353.23 -36.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -329.98 -35 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -353.23 -35 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.8 -340.58 -33.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.2 -353.23 -31.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -328.92 -30.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -353.23 -30.2 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -329.98 -28.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -353.23 -28.6 -342.06 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -339.52 -27 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -353.23 -27 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.8 -353.23 -25.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -327.86 -23.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -353.23 -23.8 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.6 -340.58 -22.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -339.52 -20.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -353.23 -20.6 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.4 -353.23 -19 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -326.8 -17.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -353.23 -17.4 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.2 -340.58 -15.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.6 -353.23 -14.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -325.74 -12.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -353.23 -12.6 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -326.8 -11 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -353.23 -11 -342.06 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -212.32 -9.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -339.52 -9.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -353.23 -9.4 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.2 -353.23 -7.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -321.5 -6.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -353.23 -6.2 -342.06 ;
    END
    PORT
      LAYER met3 ;
        RECT -5 -353.23 -4.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.4 -353.23 -3 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 2.86 -1.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 -353.23 -1.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 2.86 0.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 -353.23 0.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 2.86 1.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 -353.23 1.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 2.86 3.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 -353.23 3.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 2.86 5 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 -353.23 5 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 2.86 6.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -353.23 6.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 2.86 8.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -353.23 8.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 2.86 9.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -353.23 9.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 2.86 11.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -258.96 11.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -353.23 11.4 -303.9 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 2.86 13 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -221.86 13 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -295 13 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 2.86 14.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -232.46 14.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -353.23 14.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 2.86 16.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 -353.23 16.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 2.86 17.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 -353.23 17.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 2.86 19.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -353.23 19.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 2.86 21 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -353.23 21 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 2.86 22.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 -301.36 22.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 2.86 24.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 -300.3 24.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 2.86 25.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 -353.23 25.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 2.86 27.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 -353.23 27.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 2.86 29 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -353.23 29 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 2.86 30.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -353.23 30.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 2.86 32.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 -353.23 32.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 2.86 33.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -221.86 33.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -295 33.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 2.86 35.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -221.86 35.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -353.23 35.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 2.86 37 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -237.76 37 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -353.23 37 -318.74 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 2.86 38.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -353.23 38.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 2.86 40.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -353.23 40.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 2.86 41.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 -353.23 41.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 2.86 43.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 -353.23 43.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 2.86 45 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 -353.23 45 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 2.86 46.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 -353.23 46.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 2.86 48.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -353.23 48.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 2.86 49.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -353.23 49.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 2.86 51.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 -353.23 51.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 2.86 53 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -221.86 53 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -295 53 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 2.86 54.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -232.46 54.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -353.23 54.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 2.86 56.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 -353.23 56.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 2.86 57.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 -353.23 57.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 2.86 59.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -353.23 59.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 2.86 61 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -353.23 61 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 2.86 62.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 -301.36 62.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 2.86 64.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -300.3 64.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -353.23 64.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 2.86 65.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 -353.23 65.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 2.86 67.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 -353.23 67.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 2.86 69 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -353.23 69 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 2.86 70.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -353.23 70.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 2.86 72.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 -353.23 72.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 2.86 73.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -221.86 73.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -295 73.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 2.86 75.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -221.86 75.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -353.23 75.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 2.86 77 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 -353.23 77 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 2.86 78.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -353.23 78.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 2.86 80.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -353.23 80.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 2.86 81.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 -353.23 81.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 2.86 83.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 -353.23 83.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 2.86 85 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 -353.23 85 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 2.86 86.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 -353.23 86.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 2.86 88.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -353.23 88.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 2.86 89.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -353.23 89.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 2.86 91.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 -353.23 91.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 2.86 93 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -221.86 93 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -295 93 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 2.86 94.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -232.46 94.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -353.23 94.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 2.86 96.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 -353.23 96.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 2.86 97.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 -353.23 97.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 2.86 99.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -353.23 99.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 2.86 101 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -353.23 101 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 2.86 102.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 -301.36 102.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 2.86 104.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -300.3 104.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -353.23 104.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 2.86 105.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 -353.23 105.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 2.86 107.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 -353.23 107.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 2.86 109 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -353.23 109 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 2.86 110.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -353.23 110.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 2.86 112.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 -353.23 112.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 2.86 113.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -221.86 113.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -295 113.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 2.86 115.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -221.86 115.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -353.23 115.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 2.86 117 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 -353.23 117 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 2.86 118.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -353.23 118.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 2.86 120.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -353.23 120.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 2.86 121.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 -353.23 121.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 2.86 123.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 -353.23 123.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 2.86 125 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 -353.23 125 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 2.86 126.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 -353.23 126.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 2.86 128.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -353.23 128.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 2.86 129.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -353.23 129.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 2.86 131.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 -353.23 131.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 2.86 133 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -221.86 133 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -295 133 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 2.86 134.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -232.46 134.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -353.23 134.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 2.86 136.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 -353.23 136.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 2.86 137.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 -353.23 137.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 2.86 139.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -353.23 139.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 2.86 141 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -353.23 141 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 2.86 142.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 -301.36 142.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 2.86 144.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -300.3 144.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -353.23 144.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 2.86 145.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 -353.23 145.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 2.86 147.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 -353.23 147.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 2.86 149 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -353.23 149 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 2.86 150.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -353.23 150.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 2.86 152.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 -353.23 152.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 2.86 153.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -221.86 153.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -295 153.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 2.86 155.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -221.86 155.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -353.23 155.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 2.86 157 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 -353.23 157 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 2.86 158.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -353.23 158.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 2.86 160.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -353.23 160.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 2.86 161.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 -353.23 161.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 2.86 163.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 -353.23 163.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 2.86 165 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 -353.23 165 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 2.86 166.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 -353.23 166.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 2.86 168.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -353.23 168.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 2.86 169.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -353.23 169.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 2.86 171.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 -353.23 171.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 2.86 173 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -221.86 173 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -295 173 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 2.86 174.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -232.46 174.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -353.23 174.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 2.86 176.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 -353.23 176.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 2.86 177.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 -353.23 177.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 2.86 179.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 -353.23 179.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 2.86 181 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 -353.23 181 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 2.86 182.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 -301.36 182.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 2.86 184.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 -300.3 184.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 2.86 185.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 -353.23 185.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 2.86 187.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 -353.23 187.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 2.86 189 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 -353.23 189 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 2.86 190.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 -353.23 190.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 2.86 192.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 -353.23 192.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 2.86 193.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -221.86 193.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -295 193.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 2.86 195.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -221.86 195.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -353.23 195.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 2.86 197 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 -237.76 197 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 -353.23 197 -318.74 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 2.86 198.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 -353.23 198.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 2.86 200.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 -353.23 200.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 2.86 201.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 -353.23 201.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 2.86 203.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 -353.23 203.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 2.86 205 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 -353.23 205 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 2.86 206.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 -353.23 206.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 2.86 208.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 -353.23 208.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 2.86 209.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 -353.23 209.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 2.86 211.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 -353.23 211.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 2.86 213 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 -221.86 213 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 -295 213 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 2.86 214.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 -232.46 214.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 -353.23 214.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 2.86 216.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 -353.23 216.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 2.86 217.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 -353.23 217.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 2.86 219.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 -353.23 219.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 2.86 221 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 -353.23 221 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 2.86 222.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 -301.36 222.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 2.86 224.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 -300.3 224.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 -353.23 224.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 2.86 225.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 -353.23 225.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 2.86 227.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 -353.23 227.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 2.86 229 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 -353.23 229 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 2.86 230.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 -353.23 230.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 2.86 232.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 -353.23 232.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 2.86 233.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -221.86 233.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -295 233.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 2.86 235.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 -221.86 235.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 -353.23 235.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 2.86 237 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 -353.23 237 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 2.86 238.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 -353.23 238.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 2.86 240.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 -353.23 240.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 2.86 241.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 -353.23 241.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 2.86 243.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 -353.23 243.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 2.86 245 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 -353.23 245 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 2.86 246.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 -353.23 246.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 2.86 248.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 -353.23 248.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 2.86 249.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -353.23 249.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 2.86 251.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 -353.23 251.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 2.86 253 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 -221.86 253 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 -295 253 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 2.86 254.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 -232.46 254.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 -353.23 254.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 2.86 256.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 -353.23 256.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 2.86 257.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 -353.23 257.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 2.86 259.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 -353.23 259.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 2.86 261 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 -353.23 261 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 2.86 262.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 -301.36 262.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 2.86 264.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 -300.3 264.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 -353.23 264.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 2.86 265.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 -353.23 265.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 2.86 267.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 -353.23 267.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 2.86 269 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 -353.23 269 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 2.86 270.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 -353.23 270.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 2.86 272.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 -353.23 272.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 2.86 273.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -221.86 273.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -295 273.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 2.86 275.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 -221.86 275.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 -353.23 275.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 2.86 277 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 -353.23 277 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 2.86 278.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 -353.23 278.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 2.86 280.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 -353.23 280.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 2.86 281.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 -353.23 281.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 2.86 283.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 -353.23 283.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 2.86 285 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 -353.23 285 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 2.86 286.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 -353.23 286.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 2.86 288.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 -353.23 288.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 2.86 289.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 -353.23 289.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 2.86 291.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 -353.23 291.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 2.86 293 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 -221.86 293 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 -295 293 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 2.86 294.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 -232.46 294.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 -353.23 294.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 2.86 296.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 -353.23 296.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 2.86 297.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 -353.23 297.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 2.86 299.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 -353.23 299.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 2.86 301 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 -353.23 301 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 2.86 302.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 -301.36 302.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 2.86 304.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 -300.3 304.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 -353.23 304.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 2.86 305.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 -353.23 305.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 2.86 307.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 -353.23 307.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 2.86 309 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 -353.23 309 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 2.86 310.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 -353.23 310.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 2.86 312.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 -353.23 312.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 2.86 313.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -221.86 313.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -295 313.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 2.86 315.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 -221.86 315.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 -353.23 315.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 2.86 317 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 -353.23 317 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 2.86 318.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 -353.23 318.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 2.86 320.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 -353.23 320.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 2.86 321.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 -353.23 321.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 2.86 323.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 -353.23 323.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 2.86 325 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 -353.23 325 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 2.86 326.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 -353.23 326.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 2.86 328.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 -353.23 328.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 2.86 329.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 -353.23 329.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 331 2.86 331.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 331 -353.23 331.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 2.86 333 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 -221.86 333 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 -295 333 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 2.86 334.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 -232.46 334.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 -353.23 334.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.8 2.86 336.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.8 -353.23 336.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.4 2.86 337.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.4 -353.23 337.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 339 2.86 339.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 339 -353.23 339.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.6 2.86 341 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.6 -353.23 341 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.2 2.86 342.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.2 -301.36 342.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.8 2.86 344.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.8 -300.3 344.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.4 2.86 345.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.4 -353.23 345.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 347 2.86 347.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 347 -353.23 347.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.6 2.86 349 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.6 -353.23 349 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.2 2.86 350.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.2 -353.23 350.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.8 2.86 352.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.8 -353.23 352.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 2.86 353.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 -221.86 353.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.4 -295 353.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 2.86 355.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 -221.86 355.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 355 -353.23 355.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 2.86 357 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 -237.76 357 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.6 -353.23 357 -318.74 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.2 2.86 358.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.2 -353.23 358.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.8 2.86 360.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.8 -353.23 360.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.4 2.86 361.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.4 -353.23 361.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 363 2.86 363.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 363 -353.23 363.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.6 2.86 365 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.6 -353.23 365 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.2 2.86 366.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.2 -353.23 366.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.8 2.86 368.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.8 -353.23 368.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.4 2.86 369.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.4 -353.23 369.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 371 2.86 371.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 371 -353.23 371.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 2.86 373 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 -221.86 373 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.6 -295 373 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 2.86 374.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 -232.46 374.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.2 -353.23 374.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.8 2.86 376.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.8 -353.23 376.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.4 2.86 377.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.4 -353.23 377.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 379 2.86 379.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 379 -353.23 379.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.6 2.86 381 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.6 -353.23 381 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.2 2.86 382.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.2 -301.36 382.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 2.86 384.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 -300.3 384.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.8 -353.23 384.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.4 2.86 385.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.4 -353.23 385.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 387 2.86 387.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 387 -353.23 387.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.6 2.86 389 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.6 -353.23 389 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.2 2.86 390.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.2 -353.23 390.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.8 2.86 392.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.8 -353.23 392.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 2.86 393.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 -221.86 393.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.4 -295 393.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 2.86 395.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 -221.86 395.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 395 -353.23 395.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.6 2.86 397 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.6 -353.23 397 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.2 2.86 398.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.2 -353.23 398.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.8 2.86 400.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.8 -353.23 400.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.4 2.86 401.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.4 -353.23 401.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 403 2.86 403.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 403 -353.23 403.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.6 2.86 405 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 404.6 -353.23 405 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.2 2.86 406.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.2 -353.23 406.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.8 2.86 408.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 407.8 -353.23 408.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.4 2.86 409.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.4 -353.23 409.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 411 2.86 411.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 411 -353.23 411.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 2.86 413 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 -221.86 413 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.6 -295 413 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 2.86 414.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 -232.46 414.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 414.2 -353.23 414.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.8 2.86 416.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 415.8 -353.23 416.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.4 2.86 417.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 417.4 -353.23 417.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 419 2.86 419.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 419 -353.23 419.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.6 2.86 421 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.6 -353.23 421 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.2 2.86 422.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 422.2 -301.36 422.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 2.86 424.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 -300.3 424.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 423.8 -353.23 424.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.4 2.86 425.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 425.4 -353.23 425.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 427 2.86 427.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 427 -353.23 427.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.6 2.86 429 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.6 -353.23 429 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.2 2.86 430.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.2 -353.23 430.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.8 2.86 432.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 431.8 -353.23 432.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 2.86 433.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 -221.86 433.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 433.4 -295 433.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 2.86 435.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 -221.86 435.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 435 -353.23 435.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.6 2.86 437 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.6 -353.23 437 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.2 2.86 438.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.2 -353.23 438.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.8 2.86 440.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.8 -353.23 440.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.4 2.86 441.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 441.4 -353.23 441.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 443 2.86 443.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 443 -353.23 443.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.6 2.86 445 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 444.6 -353.23 445 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.2 2.86 446.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 446.2 -353.23 446.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.8 2.86 448.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 447.8 -353.23 448.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.4 2.86 449.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.4 -353.23 449.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 451 2.86 451.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 451 -353.23 451.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 2.86 453 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 -221.86 453 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 452.6 -295 453 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 2.86 454.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 -232.46 454.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.2 -353.23 454.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.8 2.86 456.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 455.8 -353.23 456.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.4 2.86 457.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 457.4 -353.23 457.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 459 2.86 459.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 459 -353.23 459.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.6 2.86 461 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.6 -353.23 461 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.2 2.86 462.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 462.2 -301.36 462.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 2.86 464.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 -300.3 464.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 463.8 -353.23 464.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.4 2.86 465.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 465.4 -353.23 465.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 467 2.86 467.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 467 -353.23 467.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.6 2.86 469 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.6 -353.23 469 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.2 2.86 470.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 470.2 -353.23 470.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.8 2.86 472.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 471.8 -353.23 472.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 2.86 473.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 -221.86 473.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.4 -295 473.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 2.86 475.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 -221.86 475.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 475 -353.23 475.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.6 2.86 477 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 476.6 -353.23 477 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.2 2.86 478.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.2 -353.23 478.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.8 2.86 480.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.8 -353.23 480.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.4 2.86 481.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 481.4 -353.23 481.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 483 2.86 483.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 483 -353.23 483.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.6 2.86 485 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.6 -353.23 485 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.2 2.86 486.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 486.2 -353.23 486.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.8 2.86 488.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 487.8 -353.23 488.2 -211.68 ;
        RECT 487.75 -298.355 488.2 -298.025 ;
        RECT 487.75 -312.495 488.2 -312.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.4 2.86 489.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 489.4 -353.23 489.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 491 2.86 491.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 491 -353.23 491.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 2.86 493 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 -221.86 493 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 492.6 -295 493 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 2.86 494.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 -232.46 494.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.2 -353.23 494.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.8 2.86 496.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 495.8 -353.23 496.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.4 2.86 497.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 497.4 -353.23 497.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 499 2.86 499.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 499 -353.23 499.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.6 2.86 501 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 500.6 -353.23 501 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.2 2.86 502.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.2 -301.36 502.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.8 2.86 504.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.8 -300.3 504.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.4 2.86 505.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 505.4 -353.23 505.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 507 2.86 507.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 507 -353.23 507.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.6 2.86 509 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.6 -353.23 509 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.2 2.86 510.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 510.2 -353.23 510.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.8 2.86 512.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 511.8 -353.23 512.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 2.86 513.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 -221.86 513.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.4 -295 513.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 2.86 515.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 -221.86 515.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 515 -353.23 515.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 2.86 517 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 -237.76 517 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 516.6 -353.23 517 -318.74 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.2 2.86 518.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 518.2 -353.23 518.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.8 2.86 520.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 519.8 -353.23 520.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.4 2.86 521.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 521.4 -353.23 521.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 523 2.86 523.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 523 -353.23 523.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.6 2.86 525 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.6 -353.23 525 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.2 2.86 526.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.2 -353.23 526.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.8 2.86 528.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 527.8 -353.23 528.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.4 2.86 529.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 529.4 -353.23 529.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 531 2.86 531.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 531 -353.23 531.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 2.86 533 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 -221.86 533 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.6 -295 533 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 2.86 534.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 -232.46 534.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 534.2 -353.23 534.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.8 2.86 536.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 535.8 -353.23 536.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.4 2.86 537.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 537.4 -353.23 537.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 539 2.86 539.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 539 -353.23 539.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.6 2.86 541 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 540.6 -353.23 541 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.2 2.86 542.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 542.2 -301.36 542.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 2.86 544.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 -300.3 544.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.8 -353.23 544.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.4 2.86 545.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 545.4 -353.23 545.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 547 2.86 547.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 547 -353.23 547.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.6 2.86 549 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 548.6 -353.23 549 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.2 2.86 550.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 550.2 -353.23 550.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.8 2.86 552.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 551.8 -353.23 552.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 2.86 553.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 -221.86 553.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 553.4 -295 553.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 2.86 555.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 -221.86 555.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 555 -353.23 555.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.6 2.86 557 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 556.6 -353.23 557 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.2 2.86 558.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.2 -353.23 558.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.8 2.86 560.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 559.8 -353.23 560.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.4 2.86 561.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 561.4 -353.23 561.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 563 2.86 563.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 563 -353.23 563.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.6 2.86 565 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 564.6 -353.23 565 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.2 2.86 566.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 566.2 -353.23 566.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.8 2.86 568.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 567.8 -353.23 568.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.4 2.86 569.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 569.4 -353.23 569.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 571 2.86 571.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 571 -353.23 571.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 2.86 573 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 -221.86 573 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 572.6 -295 573 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 2.86 574.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 -232.46 574.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 574.2 -353.23 574.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.8 2.86 576.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 575.8 -353.23 576.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.4 2.86 577.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.4 -353.23 577.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 579 2.86 579.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 579 -353.23 579.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.6 2.86 581 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 580.6 -353.23 581 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.2 2.86 582.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 582.2 -301.36 582.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 2.86 584.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 -300.3 584.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.8 -353.23 584.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.4 2.86 585.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 585.4 -353.23 585.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 587 2.86 587.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 587 -353.23 587.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.6 2.86 589 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.6 -353.23 589 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.2 2.86 590.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 590.2 -353.23 590.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.8 2.86 592.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 591.8 -353.23 592.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 2.86 593.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 -221.86 593.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 593.4 -295 593.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 2.86 595.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 -221.86 595.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 595 -353.23 595.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.6 2.86 597 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 596.6 -353.23 597 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.2 2.86 598.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.2 -353.23 598.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.8 2.86 600.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 599.8 -353.23 600.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.4 2.86 601.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 601.4 -353.23 601.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 603 2.86 603.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 603 -353.23 603.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.6 2.86 605 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 604.6 -353.23 605 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.2 2.86 606.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 606.2 -353.23 606.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.8 2.86 608.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.8 -353.23 608.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.4 2.86 609.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 609.4 -353.23 609.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 611 2.86 611.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 611 -353.23 611.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 2.86 613 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 -221.86 613 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 612.6 -295 613 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 2.86 614.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 -232.46 614.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 614.2 -353.23 614.6 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.8 2.86 616.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 615.8 -353.23 616.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.4 2.86 617.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.4 -353.23 617.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 619 2.86 619.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 619 -353.23 619.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.6 2.86 621 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 620.6 -353.23 621 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.2 2.86 622.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.2 -301.36 622.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 2.86 624.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 -300.3 624.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 623.8 -353.23 624.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.4 2.86 625.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 625.4 -353.23 625.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 627 2.86 627.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 627 -353.23 627.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.6 2.86 629 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.6 -353.23 629 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.2 2.86 630.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 630.2 -353.23 630.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.8 2.86 632.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 631.8 -353.23 632.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 2.86 633.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 -221.86 633.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 633.4 -295 633.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 2.86 635.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 -221.86 635.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 635 -353.23 635.4 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.6 2.86 637 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 636.6 -353.23 637 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.2 2.86 638.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 638.2 -353.23 638.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.8 2.86 640.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 639.8 -353.23 640.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.4 2.86 641.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 641.4 -353.23 641.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 643 2.86 643.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 643 -353.23 643.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.6 2.86 645 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 644.6 -353.23 645 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.2 2.86 646.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.2 -353.23 646.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.8 2.86 648.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.8 -353.23 648.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.4 2.86 649.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 649.4 -353.23 649.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 651 -353.23 651.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 652.6 -353.23 653 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 654.2 -353.23 654.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 655.8 -353.23 656.2 11.315 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -77.8 -351.69 -77.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -76.2 -351.69 -75.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.6 -351.69 -74.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -73 -351.69 -72.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.4 -351.69 -71 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.8 -323.62 -69.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -339.52 -67.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -351.69 -67.8 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.6 -351.69 -66.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -335.28 -64.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -351.69 -64.6 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.4 -340.58 -63 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -339.52 -61.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -351.69 -61.4 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.2 -351.69 -59.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -334.22 -58.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -351.69 -58.2 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -57 -340.58 -56.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.4 -351.69 -55 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -333.16 -53.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -351.69 -53.4 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.2 -333.16 -51.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -339.52 -50.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -351.69 -50.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -49 -351.69 -48.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -332.1 -47 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -351.69 -47 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.8 -340.58 -45.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -339.52 -43.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -351.69 -43.8 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.6 -351.69 -42.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -331.04 -40.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -351.69 -40.6 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.4 -339.52 -39 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.8 -351.69 -37.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -329.98 -35.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -351.69 -35.8 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.6 -331.04 -34.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -339.52 -32.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -351.69 -32.6 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.4 -351.69 -31 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -328.92 -29.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -351.69 -29.4 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.2 -340.58 -27.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -339.52 -26.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -351.69 -26.2 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -25 -351.69 -24.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -328.92 -23 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -351.69 -23 -342.06 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.8 -339.52 -21.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.2 -351.69 -19.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -326.8 -18.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -351.69 -18.2 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -17 -327.86 -16.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -339.52 -15 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -351.69 -15 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.8 -351.69 -13.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -325.74 -11.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -351.69 -11.8 -343.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -212.32 -10.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -340.58 -10.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -339.52 -8.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -351.69 -8.6 -346.3 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.4 -351.69 -7 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -321.5 -5.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -351.69 -5.4 -342.06 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.2 -351.69 -3.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.6 -351.69 -2.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 2.86 -0.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 -351.69 -0.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 2.86 1 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 -351.69 1 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 2.86 2.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 -351.69 2.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 2.86 4.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 -351.69 4.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 2.86 5.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -351.69 5.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 2.86 7.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 -351.69 7.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 2.86 9 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -351.69 9 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 2.86 10.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -351.69 10.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 2.86 12.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 -351.69 12.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 2.86 13.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -221.86 13.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -295 13.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 2.86 15.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -221.86 15.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -351.69 15.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 2.86 17 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 -351.69 17 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 2.86 18.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -351.69 18.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 2.86 20.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -351.69 20.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 2.86 21.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -301.36 21.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 2.86 23.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 -300.3 23.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 2.86 25 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 -317.26 25 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 2.86 26.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 -351.69 26.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 2.86 28.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -351.69 28.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 2.86 29.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -351.69 29.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 2.86 31.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 -351.69 31.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 2.86 33 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -221.86 33 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -295 33 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 2.86 34.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -232.46 34.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -351.69 34.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 2.86 36.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -237.76 36.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -351.69 36.2 -318.74 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 2.86 37.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 -351.69 37.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 2.86 39.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -351.69 39.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 2.86 41 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -351.69 41 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 2.86 42.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 -351.69 42.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 2.86 44.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 -351.69 44.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 2.86 45.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 -351.69 45.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 2.86 47.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 -351.69 47.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 2.86 49 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -351.69 49 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 2.86 50.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -351.69 50.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 2.86 52.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 -351.69 52.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 2.86 53.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -221.86 53.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -295 53.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 2.86 55.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -221.86 55.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -351.69 55.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 2.86 57 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 -351.69 57 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 2.86 58.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -351.69 58.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 2.86 60.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -351.69 60.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 2.86 61.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 -301.36 61.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 2.86 63.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 -300.3 63.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 2.86 65 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 -351.69 65 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 2.86 66.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 -351.69 66.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 2.86 68.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -351.69 68.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 2.86 69.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -351.69 69.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 2.86 71.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 -351.69 71.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 2.86 73 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -221.86 73 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -295 73 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 2.86 74.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -232.46 74.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -351.69 74.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 2.86 76.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 -351.69 76.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 2.86 77.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 -351.69 77.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 2.86 79.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -351.69 79.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 2.86 81 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -351.69 81 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 2.86 82.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 -351.69 82.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 2.86 84.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 -351.69 84.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 2.86 85.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 -351.69 85.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 2.86 87.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 -351.69 87.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 2.86 89 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -351.69 89 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 2.86 90.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -351.69 90.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 2.86 92.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 -351.69 92.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 2.86 93.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -221.86 93.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -295 93.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 2.86 95.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -221.86 95.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -351.69 95.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 2.86 97 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 -351.69 97 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 2.86 98.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -351.69 98.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 2.86 100.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -351.69 100.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 2.86 101.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -301.36 101.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 2.86 103.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 -300.3 103.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 2.86 105 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 -351.69 105 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 2.86 106.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 -351.69 106.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 2.86 108.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -351.69 108.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 2.86 109.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -351.69 109.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 2.86 111.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 -351.69 111.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 2.86 113 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -221.86 113 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -295 113 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 2.86 114.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -232.46 114.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -351.69 114.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 2.86 116.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 -351.69 116.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 2.86 117.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 -351.69 117.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 2.86 119.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -351.69 119.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 2.86 121 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -351.69 121 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 2.86 122.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 -351.69 122.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 2.86 124.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 -351.69 124.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 2.86 125.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 -351.69 125.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 2.86 127.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 -351.69 127.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 2.86 129 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -351.69 129 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 2.86 130.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -351.69 130.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 2.86 132.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 -351.69 132.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 2.86 133.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -221.86 133.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -295 133.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 2.86 135.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -221.86 135.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -351.69 135.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 2.86 137 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 -351.69 137 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 2.86 138.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -351.69 138.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 2.86 140.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -351.69 140.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 2.86 141.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 -301.36 141.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 2.86 143.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 -300.3 143.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 2.86 145 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 -351.69 145 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 2.86 146.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 -351.69 146.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 2.86 148.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -351.69 148.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 2.86 149.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -351.69 149.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 2.86 151.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 -351.69 151.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 2.86 153 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -221.86 153 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -295 153 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 2.86 154.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -232.46 154.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -351.69 154.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 2.86 156.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 -351.69 156.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 2.86 157.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 -351.69 157.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 2.86 159.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -351.69 159.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 2.86 161 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -351.69 161 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 2.86 162.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 -351.69 162.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 2.86 164.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 -351.69 164.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 2.86 165.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 -351.69 165.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 2.86 167.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 -351.69 167.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 2.86 169 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -351.69 169 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 2.86 170.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -351.69 170.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 2.86 172.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 -351.69 172.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 2.86 173.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -221.86 173.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -295 173.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 2.86 175.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -221.86 175.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -351.69 175.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 2.86 177 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 -351.69 177 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 2.86 178.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 -351.69 178.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 2.86 180.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 -351.69 180.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 2.86 181.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 -301.36 181.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 2.86 183.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 -300.3 183.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 2.86 185 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 -317.26 185 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 2.86 186.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 -351.69 186.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 2.86 188.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 -351.69 188.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 2.86 189.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 -351.69 189.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 2.86 191.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 -351.69 191.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 2.86 193 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 -221.86 193 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 -295 193 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 2.86 194.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 -232.46 194.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 -351.69 194.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 2.86 196.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 -237.76 196.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 -351.69 196.2 -318.74 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 2.86 197.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 -351.69 197.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 2.86 199.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 -351.69 199.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 2.86 201 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 -351.69 201 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 2.86 202.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 -351.69 202.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 2.86 204.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 -351.69 204.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 2.86 205.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 -351.69 205.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 2.86 207.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 -351.69 207.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 2.86 209 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 -351.69 209 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 2.86 210.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 -351.69 210.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 2.86 212.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 -351.69 212.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 2.86 213.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -221.86 213.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -295 213.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 2.86 215.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 -221.86 215.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 -351.69 215.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 2.86 217 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 -351.69 217 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 2.86 218.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 -351.69 218.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 2.86 220.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 -351.69 220.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 2.86 221.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 -301.36 221.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 2.86 223.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 -300.3 223.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 2.86 225 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 -351.69 225 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 2.86 226.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 -351.69 226.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 2.86 228.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 -351.69 228.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 2.86 229.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 -351.69 229.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 2.86 231.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 -351.69 231.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 2.86 233 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 -221.86 233 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 -295 233 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 2.86 234.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 -232.46 234.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 -351.69 234.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 2.86 236.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 -351.69 236.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 2.86 237.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 -351.69 237.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 2.86 239.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 -351.69 239.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 2.86 241 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 -351.69 241 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 2.86 242.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 -351.69 242.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 2.86 244.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 -351.69 244.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 2.86 245.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 -351.69 245.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 2.86 247.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 -351.69 247.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 2.86 249 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 -351.69 249 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 2.86 250.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 -351.69 250.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 2.86 252.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 -351.69 252.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 2.86 253.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -221.86 253.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -295 253.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 2.86 255.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 -221.86 255.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 -351.69 255.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 2.86 257 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 -351.69 257 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 2.86 258.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 -351.69 258.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 2.86 260.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 -351.69 260.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 2.86 261.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 -301.36 261.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 2.86 263.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 -300.3 263.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 2.86 265 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 -351.69 265 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 2.86 266.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 -351.69 266.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 2.86 268.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 -351.69 268.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 2.86 269.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 -351.69 269.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 2.86 271.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 -351.69 271.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 2.86 273 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 -221.86 273 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 -295 273 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 2.86 274.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 -232.46 274.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 -351.69 274.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 2.86 276.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 -351.69 276.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 2.86 277.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 -351.69 277.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 2.86 279.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 -351.69 279.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 2.86 281 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 -351.69 281 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 2.86 282.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 -351.69 282.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 2.86 284.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 -351.69 284.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 2.86 285.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 -351.69 285.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 2.86 287.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 -351.69 287.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 2.86 289 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 -351.69 289 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 2.86 290.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -351.69 290.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 2.86 292.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 -351.69 292.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 2.86 293.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -221.86 293.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -295 293.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 2.86 295.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 -221.86 295.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 -351.69 295.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 2.86 297 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 -351.69 297 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 2.86 298.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 -351.69 298.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 2.86 300.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 -351.69 300.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 2.86 301.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 -301.36 301.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 2.86 303.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 -300.3 303.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 2.86 305 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 -351.69 305 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 2.86 306.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 -351.69 306.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 2.86 308.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 -351.69 308.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 2.86 309.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 -351.69 309.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 2.86 311.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 -351.69 311.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 2.86 313 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 -221.86 313 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 -295 313 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 2.86 314.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 -232.46 314.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 -351.69 314.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 2.86 316.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 -351.69 316.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 2.86 317.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 -351.69 317.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 2.86 319.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 -351.69 319.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 2.86 321 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 -351.69 321 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 2.86 322.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 -351.69 322.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 2.86 324.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 -351.69 324.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 2.86 325.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 -351.69 325.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 2.86 327.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 -351.69 327.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 2.86 329 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 -351.69 329 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 2.86 330.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 -351.69 330.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.8 2.86 332.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.8 -351.69 332.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 2.86 333.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 -221.86 333.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 -295 333.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 2.86 335.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 -221.86 335.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 -351.69 335.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.6 2.86 337 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.6 -351.69 337 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.2 2.86 338.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.2 -351.69 338.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.8 2.86 340.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.8 -351.69 340.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.4 2.86 341.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.4 -301.36 341.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 343 2.86 343.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 343 -300.3 343.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.6 2.86 345 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.6 -317.26 345 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.2 2.86 346.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.2 -351.69 346.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.8 2.86 348.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.8 -351.69 348.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.4 2.86 349.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.4 -351.69 349.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 351 2.86 351.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 351 -351.69 351.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 2.86 353 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 -221.86 353 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.6 -295 353 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 2.86 354.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 -232.46 354.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.2 -351.69 354.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 2.86 356.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 -237.76 356.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.8 -351.69 356.2 -318.74 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.4 2.86 357.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.4 -351.69 357.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 359 2.86 359.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 359 -351.69 359.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.6 2.86 361 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.6 -351.69 361 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.2 2.86 362.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.2 -351.69 362.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.8 2.86 364.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.8 -351.69 364.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.4 2.86 365.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.4 -351.69 365.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 367 2.86 367.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 367 -351.69 367.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.6 2.86 369 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.6 -351.69 369 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.2 2.86 370.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.2 -351.69 370.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.8 2.86 372.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.8 -351.69 372.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 2.86 373.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 -221.86 373.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.4 -295 373.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 2.86 375.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 -221.86 375.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 375 -351.69 375.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.6 2.86 377 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.6 -351.69 377 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.2 2.86 378.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.2 -351.69 378.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.8 2.86 380.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.8 -351.69 380.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.4 2.86 381.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.4 -301.36 381.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 383 2.86 383.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 383 -300.3 383.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.6 2.86 385 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.6 -351.69 385 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.2 2.86 386.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.2 -351.69 386.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.8 2.86 388.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.8 -351.69 388.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.4 2.86 389.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.4 -351.69 389.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 391 2.86 391.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 391 -351.69 391.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 2.86 393 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 -221.86 393 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.6 -295 393 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 2.86 394.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 -232.46 394.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.2 -351.69 394.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.8 2.86 396.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.8 -351.69 396.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.4 2.86 397.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.4 -351.69 397.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 399 2.86 399.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 399 -351.69 399.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.6 2.86 401 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.6 -351.69 401 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.2 2.86 402.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.2 -351.69 402.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.8 2.86 404.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 403.8 -351.69 404.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.4 2.86 405.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.4 -351.69 405.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 407 2.86 407.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 407 -351.69 407.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.6 2.86 409 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 408.6 -351.69 409 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.2 2.86 410.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 410.2 -351.69 410.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.8 2.86 412.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 411.8 -351.69 412.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 2.86 413.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 -221.86 413.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.4 -295 413.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 2.86 415.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 -221.86 415.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 415 -351.69 415.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.6 2.86 417 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 416.6 -351.69 417 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.2 2.86 418.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.2 -351.69 418.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.8 2.86 420.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 419.8 -351.69 420.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.4 2.86 421.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 421.4 -301.36 421.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 423 2.86 423.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 423 -300.3 423.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.6 2.86 425 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.6 -351.69 425 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.2 2.86 426.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 426.2 -351.69 426.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.8 2.86 428.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 427.8 -351.69 428.2 -211.68 ;
        RECT 427.75 -321.365 428.2 -321.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.4 2.86 429.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 429.4 -351.69 429.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 431 2.86 431.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 431 -351.69 431.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 2.86 433 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 -221.86 433 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 432.6 -295 433 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 2.86 434.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 -232.46 434.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 434.2 -351.69 434.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.8 2.86 436.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.8 -351.69 436.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.4 2.86 437.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 437.4 -351.69 437.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 439 2.86 439.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 439 -351.69 439.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.6 2.86 441 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 440.6 -351.69 441 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.2 2.86 442.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.2 -351.69 442.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.8 2.86 444.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.8 -351.69 444.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.4 2.86 445.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 445.4 -351.69 445.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 447 2.86 447.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 447 -351.69 447.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.6 2.86 449 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.6 -351.69 449 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.2 2.86 450.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 450.2 -351.69 450.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.8 2.86 452.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 451.8 -351.69 452.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 2.86 453.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 -221.86 453.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 -295 453.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 2.86 455.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 -221.86 455.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 455 -351.69 455.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.6 2.86 457 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 456.6 -351.69 457 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.2 2.86 458.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.2 -351.69 458.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.8 2.86 460.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 459.8 -351.69 460.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.4 2.86 461.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 461.4 -301.36 461.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 463 2.86 463.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 463 -300.3 463.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.6 2.86 465 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.6 -351.69 465 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.2 2.86 466.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.2 -351.69 466.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.8 2.86 468.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.8 -351.69 468.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.4 2.86 469.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.4 -351.69 469.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 471 2.86 471.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 471 -351.69 471.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 2.86 473 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 -221.86 473 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.6 -295 473 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 2.86 474.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 -232.46 474.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 474.2 -351.69 474.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.8 2.86 476.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 475.8 -351.69 476.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.4 2.86 477.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 477.4 -351.69 477.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 479 2.86 479.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 479 -351.69 479.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.6 2.86 481 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 480.6 -351.69 481 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.2 2.86 482.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 482.2 -351.69 482.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.8 2.86 484.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.8 -351.69 484.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.4 2.86 485.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 485.4 -351.69 485.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 487 2.86 487.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 487 -351.69 487.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.6 2.86 489 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.6 -351.69 489 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.2 2.86 490.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.2 -351.69 490.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.8 2.86 492.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 491.8 -351.69 492.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 2.86 493.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 -221.86 493.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 493.4 -295 493.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 2.86 495.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 -221.86 495.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 495 -351.69 495.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.6 2.86 497 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.6 -351.69 497 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.2 2.86 498.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.2 -351.69 498.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.8 2.86 500.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 499.8 -351.69 500.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.4 2.86 501.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 501.4 -301.36 501.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 503 2.86 503.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 503 -300.3 503.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.6 2.86 505 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 504.6 -317.26 505 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.2 2.86 506.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 506.2 -351.69 506.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.8 2.86 508.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 507.8 -351.69 508.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.4 2.86 509.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.4 -351.69 509.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 511 2.86 511.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 511 -351.69 511.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 2.86 513 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 -221.86 513 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 512.6 -295 513 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 2.86 514.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 -232.46 514.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.2 -351.69 514.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 2.86 516.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 -237.76 516.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 515.8 -351.69 516.2 -318.74 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.4 2.86 517.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.4 -351.69 517.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 519 2.86 519.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 519 -351.69 519.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.6 2.86 521 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.6 -351.69 521 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.2 2.86 522.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 522.2 -351.69 522.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.8 2.86 524.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 523.8 -351.69 524.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.4 2.86 525.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 525.4 -351.69 525.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 527 2.86 527.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 527 -351.69 527.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.6 2.86 529 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.6 -351.69 529 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.2 2.86 530.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 530.2 -351.69 530.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.8 2.86 532.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 531.8 -351.69 532.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 2.86 533.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 -221.86 533.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 533.4 -295 533.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 2.86 535.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 -221.86 535.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 535 -351.69 535.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.6 2.86 537 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 536.6 -351.69 537 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.2 2.86 538.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.2 -351.69 538.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.8 2.86 540.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.8 -351.69 540.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.4 2.86 541.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 541.4 -301.36 541.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 543 2.86 543.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 543 -300.3 543.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.6 2.86 545 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.6 -351.69 545 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.2 2.86 546.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 546.2 -351.69 546.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.8 2.86 548.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.8 -351.69 548.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.4 2.86 549.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 549.4 -351.69 549.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 551 2.86 551.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 551 -351.69 551.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 2.86 553 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 -221.86 553 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 552.6 -295 553 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 2.86 554.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 -232.46 554.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.2 -351.69 554.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.8 2.86 556.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 555.8 -351.69 556.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 557.4 2.86 557.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 557.4 -351.69 557.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 559 2.86 559.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 559 -351.69 559.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.6 2.86 561 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 560.6 -351.69 561 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 2.86 562.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 -351.69 562.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.8 2.86 564.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 563.8 -351.69 564.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.4 2.86 565.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 565.4 -351.69 565.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 567 2.86 567.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 567 -351.69 567.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.6 2.86 569 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.6 -351.69 569 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.2 2.86 570.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 570.2 -351.69 570.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.8 2.86 572.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 571.8 -351.69 572.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 2.86 573.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 -221.86 573.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.4 -295 573.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 2.86 575.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 -221.86 575.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 575 -351.69 575.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.6 2.86 577 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 576.6 -351.69 577 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.2 2.86 578.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 578.2 -351.69 578.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.8 2.86 580.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 579.8 -351.69 580.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.4 2.86 581.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 581.4 -301.36 581.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 583 2.86 583.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 583 -300.3 583.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.6 2.86 585 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 584.6 -351.69 585 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.2 2.86 586.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 586.2 -351.69 586.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.8 2.86 588.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 587.8 -351.69 588.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.4 2.86 589.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 589.4 -351.69 589.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 591 2.86 591.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 591 -351.69 591.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 2.86 593 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 -221.86 593 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.6 -295 593 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 2.86 594.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 -232.46 594.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 594.2 -351.69 594.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.8 2.86 596.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 595.8 -351.69 596.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.4 2.86 597.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 597.4 -351.69 597.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 599 2.86 599.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 599 -351.69 599.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.6 2.86 601 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 600.6 -351.69 601 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.2 2.86 602.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.2 -351.69 602.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.8 2.86 604.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 603.8 -351.69 604.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.4 2.86 605.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 605.4 -351.69 605.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 607 2.86 607.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 607 -351.69 607.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.6 2.86 609 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 608.6 -351.69 609 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.2 2.86 610.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 610.2 -351.69 610.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.8 2.86 612.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 611.8 -351.69 612.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 2.86 613.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 -221.86 613.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.4 -295 613.8 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 2.86 615.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 -221.86 615.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 615 -351.69 615.4 -301.78 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.6 2.86 617 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 616.6 -351.69 617 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.2 2.86 618.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 618.2 -351.69 618.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.8 2.86 620.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 619.8 -351.69 620.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.4 2.86 621.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 621.4 -301.36 621.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 623 2.86 623.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 623 -300.3 623.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.6 2.86 625 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 624.6 -351.69 625 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.2 2.86 626.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 626.2 -351.69 626.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.8 2.86 628.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 627.8 -351.69 628.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.4 2.86 629.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 629.4 -351.69 629.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 631 2.86 631.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 631 -351.69 631.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 2.86 633 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 -221.86 633 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.6 -295 633 -285.88 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 2.86 634.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 -232.46 634.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 634.2 -351.69 634.6 -310.26 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.8 2.86 636.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 635.8 -351.69 636.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.4 2.86 637.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 637.4 -351.69 637.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 639 2.86 639.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 639 -351.69 639.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.6 2.86 641 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 640.6 -351.69 641 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.2 2.86 642.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.2 -351.69 642.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.8 2.86 644.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.8 -351.69 644.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.4 2.86 645.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.4 -351.69 645.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 647 2.86 647.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 647 -351.69 647.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.6 2.86 649 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.6 -351.69 649 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.2 2.86 650.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 650.2 -351.69 650.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.8 -351.69 652.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.4 -351.69 653.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 655 -351.69 655.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.6 -351.69 657 9.775 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -16.46 -353.63 -16.16 -353.33 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -22.3 -353.63 -22 -353.33 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.14 -353.63 -27.84 -353.33 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -33.98 -353.63 -33.68 -353.33 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -39.82 -353.63 -39.52 -353.33 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -45.66 -353.63 -45.36 -353.33 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -51.5 -353.63 -51.2 -353.33 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -57.34 -353.63 -57.04 -353.33 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -63.18 -353.63 -62.88 -353.33 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -69.02 -353.63 -68.72 -353.33 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -70.04 -353.63 -69.62 -353.21 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.015 -353.63 22.315 -353.33 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.015 -353.63 222.315 -353.33 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.63 -353.63 222.93 -353.33 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.015 -353.63 262.315 -353.33 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 262.63 -353.63 262.93 -353.33 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 302.015 -353.63 302.315 -353.33 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 302.63 -353.63 302.93 -353.33 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 342.015 -353.63 342.315 -353.33 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 342.63 -353.63 342.93 -353.33 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 382.015 -353.63 382.315 -353.33 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 382.63 -353.63 382.93 -353.33 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.63 -353.63 22.93 -353.33 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 422.015 -353.63 422.315 -353.33 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 422.63 -353.63 422.93 -353.33 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 462.015 -353.63 462.315 -353.33 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 462.63 -353.63 462.93 -353.33 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 502.015 -353.63 502.315 -353.33 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 502.63 -353.63 502.93 -353.33 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 542.015 -353.63 542.315 -353.33 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 542.63 -353.63 542.93 -353.33 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.015 -353.63 582.315 -353.33 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.63 -353.63 582.93 -353.33 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.015 -353.63 62.315 -353.33 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 622.015 -353.63 622.315 -353.33 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 622.63 -353.63 622.93 -353.33 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.63 -353.63 62.93 -353.33 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.015 -353.63 102.315 -353.33 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.63 -353.63 102.93 -353.33 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.015 -353.63 142.315 -353.33 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.63 -353.63 142.93 -353.33 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.015 -353.63 182.315 -353.33 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.63 -353.63 182.93 -353.33 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 13.285 -353.63 13.585 -353.33 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.285 -353.63 213.585 -353.33 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.285 -353.63 233.585 -353.33 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 253.285 -353.63 253.585 -353.33 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 273.285 -353.63 273.585 -353.33 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 293.285 -353.63 293.585 -353.33 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.285 -353.63 313.585 -353.33 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 333.285 -353.63 333.585 -353.33 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 353.285 -353.63 353.585 -353.33 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 373.285 -353.63 373.585 -353.33 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.285 -353.63 393.585 -353.33 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 33.285 -353.63 33.585 -353.33 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 413.285 -353.63 413.585 -353.33 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 433.285 -353.63 433.585 -353.33 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 453.285 -353.63 453.585 -353.33 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.285 -353.63 473.585 -353.33 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.285 -353.63 493.585 -353.33 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 513.285 -353.63 513.585 -353.33 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 533.285 -353.63 533.585 -353.33 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 553.285 -353.63 553.585 -353.33 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 573.285 -353.63 573.585 -353.33 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 593.285 -353.63 593.585 -353.33 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.285 -353.63 53.585 -353.33 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.285 -353.63 613.585 -353.33 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 633.285 -353.63 633.585 -353.33 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 73.285 -353.63 73.585 -353.33 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 93.285 -353.63 93.585 -353.33 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.285 -353.63 113.585 -353.33 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.285 -353.63 133.585 -353.33 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 153.285 -353.63 153.585 -353.33 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 173.285 -353.63 173.585 -353.33 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.285 -353.63 193.585 -353.33 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -10.62 -353.63 -10.32 -353.33 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.125 -353.63 24.425 -353.33 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 184.125 -353.63 184.425 -353.33 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 344.125 -353.63 344.425 -353.33 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 504.125 -353.63 504.425 -353.33 ;
    END
  END wmask[3]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -84.035 -353.63 662.46 11.715 ;
    LAYER met2 SPACING 0.14 ;
      RECT -84.035 -353.63 662.46 11.715 ;
    LAYER met3 SPACING 0.3 ;
      RECT 635.115 -270.01 635.445 -269.68 ;
      RECT 635.13 -285.44 635.43 -269.68 ;
      RECT 635.115 -285.44 635.445 -285.11 ;
      RECT 635.13 -266.225 635.43 -222.48 ;
      RECT 635.115 -224.455 635.445 -224.125 ;
      RECT 635.115 -265.815 635.445 -265.485 ;
      RECT 634.515 -309.33 634.815 -233.74 ;
      RECT 634.5 -234.115 634.83 -233.785 ;
      RECT 634.5 -253.595 634.83 -253.265 ;
      RECT 634.5 -309.33 634.83 -309 ;
      RECT 633.9 -248.935 634.2 -234.37 ;
      RECT 633.885 -234.745 634.215 -234.415 ;
      RECT 633.885 -248.935 634.215 -248.605 ;
      RECT 633.27 -296.415 633.6 -296.085 ;
      RECT 633.285 -352.84 633.585 -296.085 ;
      RECT 633.27 -270.47 633.6 -270.14 ;
      RECT 633.285 -285.44 633.585 -270.14 ;
      RECT 633.27 -285.44 633.6 -285.11 ;
      RECT 633.285 -266.245 633.585 -222.48 ;
      RECT 633.27 -222.855 633.6 -222.525 ;
      RECT 633.27 -266.245 633.6 -265.915 ;
      RECT 623.245 -301.805 623.575 -301.475 ;
      RECT 623.26 -345.57 623.56 -301.475 ;
      RECT 623.245 -309.045 623.575 -308.715 ;
      RECT 623.245 -345.525 623.575 -345.195 ;
      RECT 622.615 -308.245 622.945 -307.915 ;
      RECT 622.63 -352.84 622.93 -307.915 ;
      RECT 622 -302.605 622.33 -302.275 ;
      RECT 622.015 -352.84 622.315 -302.275 ;
      RECT 615.115 -270.01 615.445 -269.68 ;
      RECT 615.13 -285.44 615.43 -269.68 ;
      RECT 615.115 -285.44 615.445 -285.11 ;
      RECT 615.13 -266.225 615.43 -222.48 ;
      RECT 615.115 -224.455 615.445 -224.125 ;
      RECT 615.115 -265.815 615.445 -265.485 ;
      RECT 614.515 -301.32 614.815 -233.74 ;
      RECT 614.5 -234.115 614.83 -233.785 ;
      RECT 614.5 -253.595 614.83 -253.265 ;
      RECT 614.5 -301.32 614.83 -300.99 ;
      RECT 613.9 -248.935 614.2 -234.37 ;
      RECT 613.885 -234.745 614.215 -234.415 ;
      RECT 613.885 -248.935 614.215 -248.605 ;
      RECT 613.27 -296.415 613.6 -296.085 ;
      RECT 613.285 -352.84 613.585 -296.085 ;
      RECT 613.27 -270.47 613.6 -270.14 ;
      RECT 613.285 -285.44 613.585 -270.14 ;
      RECT 613.27 -285.44 613.6 -285.11 ;
      RECT 613.285 -266.245 613.585 -222.48 ;
      RECT 613.27 -222.855 613.6 -222.525 ;
      RECT 613.27 -266.245 613.6 -265.915 ;
      RECT 595.115 -270.01 595.445 -269.68 ;
      RECT 595.13 -285.44 595.43 -269.68 ;
      RECT 595.115 -285.44 595.445 -285.11 ;
      RECT 595.13 -266.225 595.43 -222.48 ;
      RECT 595.115 -224.455 595.445 -224.125 ;
      RECT 595.115 -265.815 595.445 -265.485 ;
      RECT 594.515 -309.33 594.815 -233.74 ;
      RECT 594.5 -234.115 594.83 -233.785 ;
      RECT 594.5 -253.595 594.83 -253.265 ;
      RECT 594.5 -309.33 594.83 -309 ;
      RECT 593.9 -248.935 594.2 -234.37 ;
      RECT 593.885 -234.745 594.215 -234.415 ;
      RECT 593.885 -248.935 594.215 -248.605 ;
      RECT 593.27 -296.415 593.6 -296.085 ;
      RECT 593.285 -352.84 593.585 -296.085 ;
      RECT 593.27 -270.47 593.6 -270.14 ;
      RECT 593.285 -285.44 593.585 -270.14 ;
      RECT 593.27 -285.44 593.6 -285.11 ;
      RECT 593.285 -266.245 593.585 -222.48 ;
      RECT 593.27 -222.855 593.6 -222.525 ;
      RECT 593.27 -266.245 593.6 -265.915 ;
      RECT 583.245 -301.805 583.575 -301.475 ;
      RECT 583.26 -345.57 583.56 -301.475 ;
      RECT 583.245 -309.045 583.575 -308.715 ;
      RECT 583.245 -345.525 583.575 -345.195 ;
      RECT 582.615 -308.245 582.945 -307.915 ;
      RECT 582.63 -352.84 582.93 -307.915 ;
      RECT 582 -302.605 582.33 -302.275 ;
      RECT 582.015 -352.84 582.315 -302.275 ;
      RECT 575.115 -270.01 575.445 -269.68 ;
      RECT 575.13 -285.44 575.43 -269.68 ;
      RECT 575.115 -285.44 575.445 -285.11 ;
      RECT 575.13 -266.225 575.43 -222.48 ;
      RECT 575.115 -224.455 575.445 -224.125 ;
      RECT 575.115 -265.815 575.445 -265.485 ;
      RECT 574.515 -301.32 574.815 -233.74 ;
      RECT 574.5 -234.115 574.83 -233.785 ;
      RECT 574.5 -253.595 574.83 -253.265 ;
      RECT 574.5 -301.32 574.83 -300.99 ;
      RECT 573.9 -248.935 574.2 -234.37 ;
      RECT 573.885 -234.745 574.215 -234.415 ;
      RECT 573.885 -248.935 574.215 -248.605 ;
      RECT 573.27 -296.415 573.6 -296.085 ;
      RECT 573.285 -352.84 573.585 -296.085 ;
      RECT 573.27 -270.47 573.6 -270.14 ;
      RECT 573.285 -285.44 573.585 -270.14 ;
      RECT 573.27 -285.44 573.6 -285.11 ;
      RECT 573.285 -266.245 573.585 -222.48 ;
      RECT 573.27 -222.855 573.6 -222.525 ;
      RECT 573.27 -266.245 573.6 -265.915 ;
      RECT 555.115 -270.01 555.445 -269.68 ;
      RECT 555.13 -285.44 555.43 -269.68 ;
      RECT 555.115 -285.44 555.445 -285.11 ;
      RECT 555.13 -266.225 555.43 -222.48 ;
      RECT 555.115 -224.455 555.445 -224.125 ;
      RECT 555.115 -265.815 555.445 -265.485 ;
      RECT 554.515 -309.33 554.815 -233.74 ;
      RECT 554.5 -234.115 554.83 -233.785 ;
      RECT 554.5 -253.595 554.83 -253.265 ;
      RECT 554.5 -309.33 554.83 -309 ;
      RECT 553.9 -248.935 554.2 -234.37 ;
      RECT 553.885 -234.745 554.215 -234.415 ;
      RECT 553.885 -248.935 554.215 -248.605 ;
      RECT 553.27 -296.415 553.6 -296.085 ;
      RECT 553.285 -352.84 553.585 -296.085 ;
      RECT 553.27 -270.47 553.6 -270.14 ;
      RECT 553.285 -285.44 553.585 -270.14 ;
      RECT 553.27 -285.44 553.6 -285.11 ;
      RECT 553.285 -266.245 553.585 -222.48 ;
      RECT 553.27 -222.855 553.6 -222.525 ;
      RECT 553.27 -266.245 553.6 -265.915 ;
      RECT 543.245 -301.805 543.575 -301.475 ;
      RECT 543.26 -345.57 543.56 -301.475 ;
      RECT 543.245 -309.045 543.575 -308.715 ;
      RECT 543.245 -345.525 543.575 -345.195 ;
      RECT 542.615 -308.245 542.945 -307.915 ;
      RECT 542.63 -352.84 542.93 -307.915 ;
      RECT 542 -302.605 542.33 -302.275 ;
      RECT 542.015 -352.84 542.315 -302.275 ;
      RECT 535.115 -270.01 535.445 -269.68 ;
      RECT 535.13 -285.44 535.43 -269.68 ;
      RECT 535.115 -285.44 535.445 -285.11 ;
      RECT 535.13 -266.225 535.43 -222.48 ;
      RECT 535.115 -224.455 535.445 -224.125 ;
      RECT 535.115 -265.815 535.445 -265.485 ;
      RECT 534.515 -301.32 534.815 -233.74 ;
      RECT 534.5 -234.115 534.83 -233.785 ;
      RECT 534.5 -253.595 534.83 -253.265 ;
      RECT 534.5 -301.32 534.83 -300.99 ;
      RECT 533.9 -248.935 534.2 -234.37 ;
      RECT 533.885 -234.745 534.215 -234.415 ;
      RECT 533.885 -248.935 534.215 -248.605 ;
      RECT 533.27 -296.415 533.6 -296.085 ;
      RECT 533.285 -352.84 533.585 -296.085 ;
      RECT 533.27 -270.47 533.6 -270.14 ;
      RECT 533.285 -285.44 533.585 -270.14 ;
      RECT 533.27 -285.44 533.6 -285.11 ;
      RECT 533.285 -266.245 533.585 -222.48 ;
      RECT 533.27 -222.855 533.6 -222.525 ;
      RECT 533.27 -266.245 533.6 -265.915 ;
      RECT 516.3 -318.17 516.6 -238.465 ;
      RECT 516.285 -238.84 516.615 -238.51 ;
      RECT 516.285 -318.17 516.615 -317.84 ;
      RECT 515.115 -270.01 515.445 -269.68 ;
      RECT 515.13 -285.44 515.43 -269.68 ;
      RECT 515.115 -285.44 515.445 -285.11 ;
      RECT 515.13 -266.225 515.43 -222.48 ;
      RECT 515.115 -224.455 515.445 -224.125 ;
      RECT 515.115 -265.815 515.445 -265.485 ;
      RECT 514.515 -309.33 514.815 -233.74 ;
      RECT 514.5 -234.115 514.83 -233.785 ;
      RECT 514.5 -253.595 514.83 -253.265 ;
      RECT 514.5 -309.33 514.83 -309 ;
      RECT 513.9 -248.935 514.2 -234.37 ;
      RECT 513.885 -234.745 514.215 -234.415 ;
      RECT 513.885 -248.935 514.215 -248.605 ;
      RECT 513.27 -296.415 513.6 -296.085 ;
      RECT 513.285 -352.84 513.585 -296.085 ;
      RECT 513.27 -270.47 513.6 -270.14 ;
      RECT 513.285 -285.44 513.585 -270.14 ;
      RECT 513.27 -285.44 513.6 -285.11 ;
      RECT 513.285 -266.245 513.585 -222.48 ;
      RECT 513.27 -222.855 513.6 -222.525 ;
      RECT 513.27 -266.245 513.6 -265.915 ;
      RECT 504.11 -318.545 504.44 -318.215 ;
      RECT 504.125 -352.84 504.425 -318.215 ;
      RECT 503.245 -301.805 503.575 -301.475 ;
      RECT 503.26 -345.57 503.56 -301.475 ;
      RECT 503.245 -309.045 503.575 -308.715 ;
      RECT 503.245 -317.745 503.575 -317.415 ;
      RECT 503.245 -345.525 503.575 -345.195 ;
      RECT 502.615 -308.245 502.945 -307.915 ;
      RECT 502.63 -352.84 502.93 -307.915 ;
      RECT 502 -302.605 502.33 -302.275 ;
      RECT 502.015 -352.84 502.315 -302.275 ;
      RECT 495.115 -270.01 495.445 -269.68 ;
      RECT 495.13 -285.44 495.43 -269.68 ;
      RECT 495.115 -285.44 495.445 -285.11 ;
      RECT 495.13 -266.225 495.43 -222.48 ;
      RECT 495.115 -224.455 495.445 -224.125 ;
      RECT 495.115 -265.815 495.445 -265.485 ;
      RECT 494.515 -301.32 494.815 -233.74 ;
      RECT 494.5 -234.115 494.83 -233.785 ;
      RECT 494.5 -253.595 494.83 -253.265 ;
      RECT 494.5 -301.32 494.83 -300.99 ;
      RECT 493.9 -248.935 494.2 -234.37 ;
      RECT 493.885 -234.745 494.215 -234.415 ;
      RECT 493.885 -248.935 494.215 -248.605 ;
      RECT 493.27 -296.415 493.6 -296.085 ;
      RECT 493.285 -352.84 493.585 -296.085 ;
      RECT 493.27 -270.47 493.6 -270.14 ;
      RECT 493.285 -285.44 493.585 -270.14 ;
      RECT 493.27 -285.44 493.6 -285.11 ;
      RECT 493.285 -266.245 493.585 -222.48 ;
      RECT 493.27 -222.855 493.6 -222.525 ;
      RECT 493.27 -266.245 493.6 -265.915 ;
      RECT 475.115 -270.01 475.445 -269.68 ;
      RECT 475.13 -285.44 475.43 -269.68 ;
      RECT 475.115 -285.44 475.445 -285.11 ;
      RECT 475.13 -266.225 475.43 -222.48 ;
      RECT 475.115 -224.455 475.445 -224.125 ;
      RECT 475.115 -265.815 475.445 -265.485 ;
      RECT 474.515 -309.33 474.815 -233.74 ;
      RECT 474.5 -234.115 474.83 -233.785 ;
      RECT 474.5 -253.595 474.83 -253.265 ;
      RECT 474.5 -309.33 474.83 -309 ;
      RECT 473.9 -248.935 474.2 -234.37 ;
      RECT 473.885 -234.745 474.215 -234.415 ;
      RECT 473.885 -248.935 474.215 -248.605 ;
      RECT 473.27 -296.415 473.6 -296.085 ;
      RECT 473.285 -352.84 473.585 -296.085 ;
      RECT 473.27 -270.47 473.6 -270.14 ;
      RECT 473.285 -285.44 473.585 -270.14 ;
      RECT 473.27 -285.44 473.6 -285.11 ;
      RECT 473.285 -266.245 473.585 -222.48 ;
      RECT 473.27 -222.855 473.6 -222.525 ;
      RECT 473.27 -266.245 473.6 -265.915 ;
      RECT 463.245 -301.805 463.575 -301.475 ;
      RECT 463.26 -345.57 463.56 -301.475 ;
      RECT 463.245 -309.045 463.575 -308.715 ;
      RECT 463.245 -345.525 463.575 -345.195 ;
      RECT 462.615 -308.245 462.945 -307.915 ;
      RECT 462.63 -352.84 462.93 -307.915 ;
      RECT 462 -302.605 462.33 -302.275 ;
      RECT 462.015 -352.84 462.315 -302.275 ;
      RECT 455.115 -270.01 455.445 -269.68 ;
      RECT 455.13 -285.44 455.43 -269.68 ;
      RECT 455.115 -285.44 455.445 -285.11 ;
      RECT 455.13 -266.225 455.43 -222.48 ;
      RECT 455.115 -224.455 455.445 -224.125 ;
      RECT 455.115 -265.815 455.445 -265.485 ;
      RECT 454.515 -301.32 454.815 -233.74 ;
      RECT 454.5 -234.115 454.83 -233.785 ;
      RECT 454.5 -253.595 454.83 -253.265 ;
      RECT 454.5 -301.32 454.83 -300.99 ;
      RECT 453.9 -248.935 454.2 -234.37 ;
      RECT 453.885 -234.745 454.215 -234.415 ;
      RECT 453.885 -248.935 454.215 -248.605 ;
      RECT 453.27 -296.415 453.6 -296.085 ;
      RECT 453.285 -352.84 453.585 -296.085 ;
      RECT 453.27 -270.47 453.6 -270.14 ;
      RECT 453.285 -285.44 453.585 -270.14 ;
      RECT 453.27 -285.44 453.6 -285.11 ;
      RECT 453.285 -266.245 453.585 -222.48 ;
      RECT 453.27 -222.855 453.6 -222.525 ;
      RECT 453.27 -266.245 453.6 -265.915 ;
      RECT 435.115 -270.01 435.445 -269.68 ;
      RECT 435.13 -285.44 435.43 -269.68 ;
      RECT 435.115 -285.44 435.445 -285.11 ;
      RECT 435.13 -266.225 435.43 -222.48 ;
      RECT 435.115 -224.455 435.445 -224.125 ;
      RECT 435.115 -265.815 435.445 -265.485 ;
      RECT 434.515 -309.33 434.815 -233.74 ;
      RECT 434.5 -234.115 434.83 -233.785 ;
      RECT 434.5 -253.595 434.83 -253.265 ;
      RECT 434.5 -309.33 434.83 -309 ;
      RECT 433.9 -248.935 434.2 -234.37 ;
      RECT 433.885 -234.745 434.215 -234.415 ;
      RECT 433.885 -248.935 434.215 -248.605 ;
      RECT 433.27 -296.415 433.6 -296.085 ;
      RECT 433.285 -352.84 433.585 -296.085 ;
      RECT 433.27 -270.47 433.6 -270.14 ;
      RECT 433.285 -285.44 433.585 -270.14 ;
      RECT 433.27 -285.44 433.6 -285.11 ;
      RECT 433.285 -266.245 433.585 -222.48 ;
      RECT 433.27 -222.855 433.6 -222.525 ;
      RECT 433.27 -266.245 433.6 -265.915 ;
      RECT 423.245 -301.805 423.575 -301.475 ;
      RECT 423.26 -345.57 423.56 -301.475 ;
      RECT 423.245 -309.045 423.575 -308.715 ;
      RECT 423.245 -345.525 423.575 -345.195 ;
      RECT 422.615 -308.245 422.945 -307.915 ;
      RECT 422.63 -352.84 422.93 -307.915 ;
      RECT 422 -302.605 422.33 -302.275 ;
      RECT 422.015 -352.84 422.315 -302.275 ;
      RECT 415.115 -270.01 415.445 -269.68 ;
      RECT 415.13 -285.44 415.43 -269.68 ;
      RECT 415.115 -285.44 415.445 -285.11 ;
      RECT 415.13 -266.225 415.43 -222.48 ;
      RECT 415.115 -224.455 415.445 -224.125 ;
      RECT 415.115 -265.815 415.445 -265.485 ;
      RECT 414.515 -301.32 414.815 -233.74 ;
      RECT 414.5 -234.115 414.83 -233.785 ;
      RECT 414.5 -253.595 414.83 -253.265 ;
      RECT 414.5 -301.32 414.83 -300.99 ;
      RECT 413.9 -248.935 414.2 -234.37 ;
      RECT 413.885 -234.745 414.215 -234.415 ;
      RECT 413.885 -248.935 414.215 -248.605 ;
      RECT 413.27 -296.415 413.6 -296.085 ;
      RECT 413.285 -352.84 413.585 -296.085 ;
      RECT 413.27 -270.47 413.6 -270.14 ;
      RECT 413.285 -285.44 413.585 -270.14 ;
      RECT 413.27 -285.44 413.6 -285.11 ;
      RECT 413.285 -266.245 413.585 -222.48 ;
      RECT 413.27 -222.855 413.6 -222.525 ;
      RECT 413.27 -266.245 413.6 -265.915 ;
      RECT 395.115 -270.01 395.445 -269.68 ;
      RECT 395.13 -285.44 395.43 -269.68 ;
      RECT 395.115 -285.44 395.445 -285.11 ;
      RECT 395.13 -266.225 395.43 -222.48 ;
      RECT 395.115 -224.455 395.445 -224.125 ;
      RECT 395.115 -265.815 395.445 -265.485 ;
      RECT 394.515 -309.33 394.815 -233.74 ;
      RECT 394.5 -234.115 394.83 -233.785 ;
      RECT 394.5 -253.595 394.83 -253.265 ;
      RECT 394.5 -309.33 394.83 -309 ;
      RECT 393.9 -248.935 394.2 -234.37 ;
      RECT 393.885 -234.745 394.215 -234.415 ;
      RECT 393.885 -248.935 394.215 -248.605 ;
      RECT 393.27 -296.415 393.6 -296.085 ;
      RECT 393.285 -352.84 393.585 -296.085 ;
      RECT 393.27 -270.47 393.6 -270.14 ;
      RECT 393.285 -285.44 393.585 -270.14 ;
      RECT 393.27 -285.44 393.6 -285.11 ;
      RECT 393.285 -266.245 393.585 -222.48 ;
      RECT 393.27 -222.855 393.6 -222.525 ;
      RECT 393.27 -266.245 393.6 -265.915 ;
      RECT 383.245 -301.805 383.575 -301.475 ;
      RECT 383.26 -345.57 383.56 -301.475 ;
      RECT 383.245 -309.045 383.575 -308.715 ;
      RECT 383.245 -345.525 383.575 -345.195 ;
      RECT 382.615 -308.245 382.945 -307.915 ;
      RECT 382.63 -352.84 382.93 -307.915 ;
      RECT 382 -302.605 382.33 -302.275 ;
      RECT 382.015 -352.84 382.315 -302.275 ;
      RECT 375.115 -270.01 375.445 -269.68 ;
      RECT 375.13 -285.44 375.43 -269.68 ;
      RECT 375.115 -285.44 375.445 -285.11 ;
      RECT 375.13 -266.225 375.43 -222.48 ;
      RECT 375.115 -224.455 375.445 -224.125 ;
      RECT 375.115 -265.815 375.445 -265.485 ;
      RECT 374.515 -301.32 374.815 -233.74 ;
      RECT 374.5 -234.115 374.83 -233.785 ;
      RECT 374.5 -253.595 374.83 -253.265 ;
      RECT 374.5 -301.32 374.83 -300.99 ;
      RECT 373.9 -248.935 374.2 -234.37 ;
      RECT 373.885 -234.745 374.215 -234.415 ;
      RECT 373.885 -248.935 374.215 -248.605 ;
      RECT 373.27 -296.415 373.6 -296.085 ;
      RECT 373.285 -352.84 373.585 -296.085 ;
      RECT 373.27 -270.47 373.6 -270.14 ;
      RECT 373.285 -285.44 373.585 -270.14 ;
      RECT 373.27 -285.44 373.6 -285.11 ;
      RECT 373.285 -266.245 373.585 -222.48 ;
      RECT 373.27 -222.855 373.6 -222.525 ;
      RECT 373.27 -266.245 373.6 -265.915 ;
      RECT 356.3 -318.17 356.6 -238.465 ;
      RECT 356.285 -238.84 356.615 -238.51 ;
      RECT 356.285 -318.17 356.615 -317.84 ;
      RECT 355.115 -270.01 355.445 -269.68 ;
      RECT 355.13 -285.44 355.43 -269.68 ;
      RECT 355.115 -285.44 355.445 -285.11 ;
      RECT 355.13 -266.225 355.43 -222.48 ;
      RECT 355.115 -224.455 355.445 -224.125 ;
      RECT 355.115 -265.815 355.445 -265.485 ;
      RECT 354.515 -309.33 354.815 -233.74 ;
      RECT 354.5 -234.115 354.83 -233.785 ;
      RECT 354.5 -253.595 354.83 -253.265 ;
      RECT 354.5 -309.33 354.83 -309 ;
      RECT 353.9 -248.935 354.2 -234.37 ;
      RECT 353.885 -234.745 354.215 -234.415 ;
      RECT 353.885 -248.935 354.215 -248.605 ;
      RECT 353.27 -296.415 353.6 -296.085 ;
      RECT 353.285 -352.84 353.585 -296.085 ;
      RECT 353.27 -270.47 353.6 -270.14 ;
      RECT 353.285 -285.44 353.585 -270.14 ;
      RECT 353.27 -285.44 353.6 -285.11 ;
      RECT 353.285 -266.245 353.585 -222.48 ;
      RECT 353.27 -222.855 353.6 -222.525 ;
      RECT 353.27 -266.245 353.6 -265.915 ;
      RECT 344.11 -318.545 344.44 -318.215 ;
      RECT 344.125 -352.84 344.425 -318.215 ;
      RECT 343.245 -301.805 343.575 -301.475 ;
      RECT 343.26 -345.57 343.56 -301.475 ;
      RECT 343.245 -309.045 343.575 -308.715 ;
      RECT 343.245 -317.745 343.575 -317.415 ;
      RECT 343.245 -345.525 343.575 -345.195 ;
      RECT 342.615 -308.245 342.945 -307.915 ;
      RECT 342.63 -352.84 342.93 -307.915 ;
      RECT 342 -302.605 342.33 -302.275 ;
      RECT 342.015 -352.84 342.315 -302.275 ;
      RECT 335.115 -270.01 335.445 -269.68 ;
      RECT 335.13 -285.44 335.43 -269.68 ;
      RECT 335.115 -285.44 335.445 -285.11 ;
      RECT 335.13 -266.225 335.43 -222.48 ;
      RECT 335.115 -224.455 335.445 -224.125 ;
      RECT 335.115 -265.815 335.445 -265.485 ;
      RECT 334.515 -301.32 334.815 -233.74 ;
      RECT 334.5 -234.115 334.83 -233.785 ;
      RECT 334.5 -253.595 334.83 -253.265 ;
      RECT 334.5 -301.32 334.83 -300.99 ;
      RECT 333.9 -248.935 334.2 -234.37 ;
      RECT 333.885 -234.745 334.215 -234.415 ;
      RECT 333.885 -248.935 334.215 -248.605 ;
      RECT 333.27 -296.415 333.6 -296.085 ;
      RECT 333.285 -352.84 333.585 -296.085 ;
      RECT 333.27 -270.47 333.6 -270.14 ;
      RECT 333.285 -285.44 333.585 -270.14 ;
      RECT 333.27 -285.44 333.6 -285.11 ;
      RECT 333.285 -266.245 333.585 -222.48 ;
      RECT 333.27 -222.855 333.6 -222.525 ;
      RECT 333.27 -266.245 333.6 -265.915 ;
      RECT 315.115 -270.01 315.445 -269.68 ;
      RECT 315.13 -285.44 315.43 -269.68 ;
      RECT 315.115 -285.44 315.445 -285.11 ;
      RECT 315.13 -266.225 315.43 -222.48 ;
      RECT 315.115 -224.455 315.445 -224.125 ;
      RECT 315.115 -265.815 315.445 -265.485 ;
      RECT 314.515 -309.33 314.815 -233.74 ;
      RECT 314.5 -234.115 314.83 -233.785 ;
      RECT 314.5 -253.595 314.83 -253.265 ;
      RECT 314.5 -309.33 314.83 -309 ;
      RECT 313.9 -248.935 314.2 -234.37 ;
      RECT 313.885 -234.745 314.215 -234.415 ;
      RECT 313.885 -248.935 314.215 -248.605 ;
      RECT 313.27 -296.415 313.6 -296.085 ;
      RECT 313.285 -352.84 313.585 -296.085 ;
      RECT 313.27 -270.47 313.6 -270.14 ;
      RECT 313.285 -285.44 313.585 -270.14 ;
      RECT 313.27 -285.44 313.6 -285.11 ;
      RECT 313.285 -266.245 313.585 -222.48 ;
      RECT 313.27 -222.855 313.6 -222.525 ;
      RECT 313.27 -266.245 313.6 -265.915 ;
      RECT 303.245 -301.805 303.575 -301.475 ;
      RECT 303.26 -345.57 303.56 -301.475 ;
      RECT 303.245 -309.045 303.575 -308.715 ;
      RECT 303.245 -345.525 303.575 -345.195 ;
      RECT 302.615 -308.245 302.945 -307.915 ;
      RECT 302.63 -352.84 302.93 -307.915 ;
      RECT 302 -302.605 302.33 -302.275 ;
      RECT 302.015 -352.84 302.315 -302.275 ;
      RECT 295.115 -270.01 295.445 -269.68 ;
      RECT 295.13 -285.44 295.43 -269.68 ;
      RECT 295.115 -285.44 295.445 -285.11 ;
      RECT 295.13 -266.225 295.43 -222.48 ;
      RECT 295.115 -224.455 295.445 -224.125 ;
      RECT 295.115 -265.815 295.445 -265.485 ;
      RECT 294.515 -301.32 294.815 -233.74 ;
      RECT 294.5 -234.115 294.83 -233.785 ;
      RECT 294.5 -253.595 294.83 -253.265 ;
      RECT 294.5 -301.32 294.83 -300.99 ;
      RECT 293.9 -248.935 294.2 -234.37 ;
      RECT 293.885 -234.745 294.215 -234.415 ;
      RECT 293.885 -248.935 294.215 -248.605 ;
      RECT 293.27 -296.415 293.6 -296.085 ;
      RECT 293.285 -352.84 293.585 -296.085 ;
      RECT 293.27 -270.47 293.6 -270.14 ;
      RECT 293.285 -285.44 293.585 -270.14 ;
      RECT 293.27 -285.44 293.6 -285.11 ;
      RECT 293.285 -266.245 293.585 -222.48 ;
      RECT 293.27 -222.855 293.6 -222.525 ;
      RECT 293.27 -266.245 293.6 -265.915 ;
      RECT 275.115 -270.01 275.445 -269.68 ;
      RECT 275.13 -285.44 275.43 -269.68 ;
      RECT 275.115 -285.44 275.445 -285.11 ;
      RECT 275.13 -266.225 275.43 -222.48 ;
      RECT 275.115 -224.455 275.445 -224.125 ;
      RECT 275.115 -265.815 275.445 -265.485 ;
      RECT 274.515 -309.33 274.815 -233.74 ;
      RECT 274.5 -234.115 274.83 -233.785 ;
      RECT 274.5 -253.595 274.83 -253.265 ;
      RECT 274.5 -309.33 274.83 -309 ;
      RECT 273.9 -248.935 274.2 -234.37 ;
      RECT 273.885 -234.745 274.215 -234.415 ;
      RECT 273.885 -248.935 274.215 -248.605 ;
      RECT 273.27 -296.415 273.6 -296.085 ;
      RECT 273.285 -352.84 273.585 -296.085 ;
      RECT 273.27 -270.47 273.6 -270.14 ;
      RECT 273.285 -285.44 273.585 -270.14 ;
      RECT 273.27 -285.44 273.6 -285.11 ;
      RECT 273.285 -266.245 273.585 -222.48 ;
      RECT 273.27 -222.855 273.6 -222.525 ;
      RECT 273.27 -266.245 273.6 -265.915 ;
      RECT 263.245 -301.805 263.575 -301.475 ;
      RECT 263.26 -345.57 263.56 -301.475 ;
      RECT 263.245 -309.045 263.575 -308.715 ;
      RECT 263.245 -345.525 263.575 -345.195 ;
      RECT 262.615 -308.245 262.945 -307.915 ;
      RECT 262.63 -352.84 262.93 -307.915 ;
      RECT 262 -302.605 262.33 -302.275 ;
      RECT 262.015 -352.84 262.315 -302.275 ;
      RECT 255.115 -270.01 255.445 -269.68 ;
      RECT 255.13 -285.44 255.43 -269.68 ;
      RECT 255.115 -285.44 255.445 -285.11 ;
      RECT 255.13 -266.225 255.43 -222.48 ;
      RECT 255.115 -224.455 255.445 -224.125 ;
      RECT 255.115 -265.815 255.445 -265.485 ;
      RECT 254.515 -301.32 254.815 -233.74 ;
      RECT 254.5 -234.115 254.83 -233.785 ;
      RECT 254.5 -253.595 254.83 -253.265 ;
      RECT 254.5 -301.32 254.83 -300.99 ;
      RECT 253.9 -248.935 254.2 -234.37 ;
      RECT 253.885 -234.745 254.215 -234.415 ;
      RECT 253.885 -248.935 254.215 -248.605 ;
      RECT 253.27 -296.415 253.6 -296.085 ;
      RECT 253.285 -352.84 253.585 -296.085 ;
      RECT 253.27 -270.47 253.6 -270.14 ;
      RECT 253.285 -285.44 253.585 -270.14 ;
      RECT 253.27 -285.44 253.6 -285.11 ;
      RECT 253.285 -266.245 253.585 -222.48 ;
      RECT 253.27 -222.855 253.6 -222.525 ;
      RECT 253.27 -266.245 253.6 -265.915 ;
      RECT 235.115 -270.01 235.445 -269.68 ;
      RECT 235.13 -285.44 235.43 -269.68 ;
      RECT 235.115 -285.44 235.445 -285.11 ;
      RECT 235.13 -266.225 235.43 -222.48 ;
      RECT 235.115 -224.455 235.445 -224.125 ;
      RECT 235.115 -265.815 235.445 -265.485 ;
      RECT 234.515 -309.33 234.815 -233.74 ;
      RECT 234.5 -234.115 234.83 -233.785 ;
      RECT 234.5 -253.595 234.83 -253.265 ;
      RECT 234.5 -309.33 234.83 -309 ;
      RECT 233.9 -248.935 234.2 -234.37 ;
      RECT 233.885 -234.745 234.215 -234.415 ;
      RECT 233.885 -248.935 234.215 -248.605 ;
      RECT 233.27 -296.415 233.6 -296.085 ;
      RECT 233.285 -352.84 233.585 -296.085 ;
      RECT 233.27 -270.47 233.6 -270.14 ;
      RECT 233.285 -285.44 233.585 -270.14 ;
      RECT 233.27 -285.44 233.6 -285.11 ;
      RECT 233.285 -266.245 233.585 -222.48 ;
      RECT 233.27 -222.855 233.6 -222.525 ;
      RECT 233.27 -266.245 233.6 -265.915 ;
      RECT 223.245 -301.805 223.575 -301.475 ;
      RECT 223.26 -345.57 223.56 -301.475 ;
      RECT 223.245 -309.045 223.575 -308.715 ;
      RECT 223.245 -345.525 223.575 -345.195 ;
      RECT 222.615 -308.245 222.945 -307.915 ;
      RECT 222.63 -352.84 222.93 -307.915 ;
      RECT 222 -302.605 222.33 -302.275 ;
      RECT 222.015 -352.84 222.315 -302.275 ;
      RECT 215.115 -270.01 215.445 -269.68 ;
      RECT 215.13 -285.44 215.43 -269.68 ;
      RECT 215.115 -285.44 215.445 -285.11 ;
      RECT 215.13 -266.225 215.43 -222.48 ;
      RECT 215.115 -224.455 215.445 -224.125 ;
      RECT 215.115 -265.815 215.445 -265.485 ;
      RECT 214.515 -301.32 214.815 -233.74 ;
      RECT 214.5 -234.115 214.83 -233.785 ;
      RECT 214.5 -253.595 214.83 -253.265 ;
      RECT 214.5 -301.32 214.83 -300.99 ;
      RECT 213.9 -248.935 214.2 -234.37 ;
      RECT 213.885 -234.745 214.215 -234.415 ;
      RECT 213.885 -248.935 214.215 -248.605 ;
      RECT 213.27 -296.415 213.6 -296.085 ;
      RECT 213.285 -352.84 213.585 -296.085 ;
      RECT 213.27 -270.47 213.6 -270.14 ;
      RECT 213.285 -285.44 213.585 -270.14 ;
      RECT 213.27 -285.44 213.6 -285.11 ;
      RECT 213.285 -266.245 213.585 -222.48 ;
      RECT 213.27 -222.855 213.6 -222.525 ;
      RECT 213.27 -266.245 213.6 -265.915 ;
      RECT 196.3 -318.17 196.6 -238.465 ;
      RECT 196.285 -238.84 196.615 -238.51 ;
      RECT 196.285 -318.17 196.615 -317.84 ;
      RECT 195.115 -270.01 195.445 -269.68 ;
      RECT 195.13 -285.44 195.43 -269.68 ;
      RECT 195.115 -285.44 195.445 -285.11 ;
      RECT 195.13 -266.225 195.43 -222.48 ;
      RECT 195.115 -224.455 195.445 -224.125 ;
      RECT 195.115 -265.815 195.445 -265.485 ;
      RECT 194.515 -309.33 194.815 -233.74 ;
      RECT 194.5 -234.115 194.83 -233.785 ;
      RECT 194.5 -253.595 194.83 -253.265 ;
      RECT 194.5 -309.33 194.83 -309 ;
      RECT 193.9 -248.935 194.2 -234.37 ;
      RECT 193.885 -234.745 194.215 -234.415 ;
      RECT 193.885 -248.935 194.215 -248.605 ;
      RECT 193.27 -296.415 193.6 -296.085 ;
      RECT 193.285 -352.84 193.585 -296.085 ;
      RECT 193.27 -270.47 193.6 -270.14 ;
      RECT 193.285 -285.44 193.585 -270.14 ;
      RECT 193.27 -285.44 193.6 -285.11 ;
      RECT 193.285 -266.245 193.585 -222.48 ;
      RECT 193.27 -222.855 193.6 -222.525 ;
      RECT 193.27 -266.245 193.6 -265.915 ;
      RECT 184.11 -318.545 184.44 -318.215 ;
      RECT 184.125 -352.84 184.425 -318.215 ;
      RECT 183.245 -301.805 183.575 -301.475 ;
      RECT 183.26 -345.57 183.56 -301.475 ;
      RECT 183.245 -309.045 183.575 -308.715 ;
      RECT 183.245 -317.745 183.575 -317.415 ;
      RECT 183.245 -345.525 183.575 -345.195 ;
      RECT 182.615 -308.245 182.945 -307.915 ;
      RECT 182.63 -352.84 182.93 -307.915 ;
      RECT 182 -302.605 182.33 -302.275 ;
      RECT 182.015 -352.84 182.315 -302.275 ;
      RECT 175.115 -270.01 175.445 -269.68 ;
      RECT 175.13 -285.44 175.43 -269.68 ;
      RECT 175.115 -285.44 175.445 -285.11 ;
      RECT 175.13 -266.225 175.43 -222.48 ;
      RECT 175.115 -224.455 175.445 -224.125 ;
      RECT 175.115 -265.815 175.445 -265.485 ;
      RECT 174.515 -301.32 174.815 -233.74 ;
      RECT 174.5 -234.115 174.83 -233.785 ;
      RECT 174.5 -253.595 174.83 -253.265 ;
      RECT 174.5 -301.32 174.83 -300.99 ;
      RECT 173.9 -248.935 174.2 -234.37 ;
      RECT 173.885 -234.745 174.215 -234.415 ;
      RECT 173.885 -248.935 174.215 -248.605 ;
      RECT 173.27 -296.415 173.6 -296.085 ;
      RECT 173.285 -352.84 173.585 -296.085 ;
      RECT 173.27 -270.47 173.6 -270.14 ;
      RECT 173.285 -285.44 173.585 -270.14 ;
      RECT 173.27 -285.44 173.6 -285.11 ;
      RECT 173.285 -266.245 173.585 -222.48 ;
      RECT 173.27 -222.855 173.6 -222.525 ;
      RECT 173.27 -266.245 173.6 -265.915 ;
      RECT 155.115 -270.01 155.445 -269.68 ;
      RECT 155.13 -285.44 155.43 -269.68 ;
      RECT 155.115 -285.44 155.445 -285.11 ;
      RECT 155.13 -266.225 155.43 -222.48 ;
      RECT 155.115 -224.455 155.445 -224.125 ;
      RECT 155.115 -265.815 155.445 -265.485 ;
      RECT 154.515 -309.33 154.815 -233.74 ;
      RECT 154.5 -234.115 154.83 -233.785 ;
      RECT 154.5 -253.595 154.83 -253.265 ;
      RECT 154.5 -309.33 154.83 -309 ;
      RECT 153.9 -248.935 154.2 -234.37 ;
      RECT 153.885 -234.745 154.215 -234.415 ;
      RECT 153.885 -248.935 154.215 -248.605 ;
      RECT 153.27 -296.415 153.6 -296.085 ;
      RECT 153.285 -352.84 153.585 -296.085 ;
      RECT 153.27 -270.47 153.6 -270.14 ;
      RECT 153.285 -285.44 153.585 -270.14 ;
      RECT 153.27 -285.44 153.6 -285.11 ;
      RECT 153.285 -266.245 153.585 -222.48 ;
      RECT 153.27 -222.855 153.6 -222.525 ;
      RECT 153.27 -266.245 153.6 -265.915 ;
      RECT 143.245 -301.805 143.575 -301.475 ;
      RECT 143.26 -345.57 143.56 -301.475 ;
      RECT 143.245 -309.045 143.575 -308.715 ;
      RECT 143.245 -345.525 143.575 -345.195 ;
      RECT 142.615 -308.245 142.945 -307.915 ;
      RECT 142.63 -352.84 142.93 -307.915 ;
      RECT 142 -302.605 142.33 -302.275 ;
      RECT 142.015 -352.84 142.315 -302.275 ;
      RECT 135.115 -270.01 135.445 -269.68 ;
      RECT 135.13 -285.44 135.43 -269.68 ;
      RECT 135.115 -285.44 135.445 -285.11 ;
      RECT 135.13 -266.225 135.43 -222.48 ;
      RECT 135.115 -224.455 135.445 -224.125 ;
      RECT 135.115 -265.815 135.445 -265.485 ;
      RECT 134.515 -301.32 134.815 -233.74 ;
      RECT 134.5 -234.115 134.83 -233.785 ;
      RECT 134.5 -253.595 134.83 -253.265 ;
      RECT 134.5 -301.32 134.83 -300.99 ;
      RECT 133.9 -248.935 134.2 -234.37 ;
      RECT 133.885 -234.745 134.215 -234.415 ;
      RECT 133.885 -248.935 134.215 -248.605 ;
      RECT 133.27 -296.415 133.6 -296.085 ;
      RECT 133.285 -352.84 133.585 -296.085 ;
      RECT 133.27 -270.47 133.6 -270.14 ;
      RECT 133.285 -285.44 133.585 -270.14 ;
      RECT 133.27 -285.44 133.6 -285.11 ;
      RECT 133.285 -266.245 133.585 -222.48 ;
      RECT 133.27 -222.855 133.6 -222.525 ;
      RECT 133.27 -266.245 133.6 -265.915 ;
      RECT 115.115 -270.01 115.445 -269.68 ;
      RECT 115.13 -285.44 115.43 -269.68 ;
      RECT 115.115 -285.44 115.445 -285.11 ;
      RECT 115.13 -266.225 115.43 -222.48 ;
      RECT 115.115 -224.455 115.445 -224.125 ;
      RECT 115.115 -265.815 115.445 -265.485 ;
      RECT 114.515 -309.33 114.815 -233.74 ;
      RECT 114.5 -234.115 114.83 -233.785 ;
      RECT 114.5 -253.595 114.83 -253.265 ;
      RECT 114.5 -309.33 114.83 -309 ;
      RECT 113.9 -248.935 114.2 -234.37 ;
      RECT 113.885 -234.745 114.215 -234.415 ;
      RECT 113.885 -248.935 114.215 -248.605 ;
      RECT 113.27 -296.415 113.6 -296.085 ;
      RECT 113.285 -352.84 113.585 -296.085 ;
      RECT 113.27 -270.47 113.6 -270.14 ;
      RECT 113.285 -285.44 113.585 -270.14 ;
      RECT 113.27 -285.44 113.6 -285.11 ;
      RECT 113.285 -266.245 113.585 -222.48 ;
      RECT 113.27 -222.855 113.6 -222.525 ;
      RECT 113.27 -266.245 113.6 -265.915 ;
      RECT 103.245 -301.805 103.575 -301.475 ;
      RECT 103.26 -345.57 103.56 -301.475 ;
      RECT 103.245 -309.045 103.575 -308.715 ;
      RECT 103.245 -345.525 103.575 -345.195 ;
      RECT 102.615 -308.245 102.945 -307.915 ;
      RECT 102.63 -352.84 102.93 -307.915 ;
      RECT 102 -302.605 102.33 -302.275 ;
      RECT 102.015 -352.84 102.315 -302.275 ;
      RECT 95.115 -270.01 95.445 -269.68 ;
      RECT 95.13 -285.44 95.43 -269.68 ;
      RECT 95.115 -285.44 95.445 -285.11 ;
      RECT 95.13 -266.225 95.43 -222.48 ;
      RECT 95.115 -224.455 95.445 -224.125 ;
      RECT 95.115 -265.815 95.445 -265.485 ;
      RECT 94.515 -301.32 94.815 -233.74 ;
      RECT 94.5 -234.115 94.83 -233.785 ;
      RECT 94.5 -253.595 94.83 -253.265 ;
      RECT 94.5 -301.32 94.83 -300.99 ;
      RECT 93.9 -248.935 94.2 -234.37 ;
      RECT 93.885 -234.745 94.215 -234.415 ;
      RECT 93.885 -248.935 94.215 -248.605 ;
      RECT 93.27 -296.415 93.6 -296.085 ;
      RECT 93.285 -352.84 93.585 -296.085 ;
      RECT 93.27 -270.47 93.6 -270.14 ;
      RECT 93.285 -285.44 93.585 -270.14 ;
      RECT 93.27 -285.44 93.6 -285.11 ;
      RECT 93.285 -266.245 93.585 -222.48 ;
      RECT 93.27 -222.855 93.6 -222.525 ;
      RECT 93.27 -266.245 93.6 -265.915 ;
      RECT 75.115 -270.01 75.445 -269.68 ;
      RECT 75.13 -285.44 75.43 -269.68 ;
      RECT 75.115 -285.44 75.445 -285.11 ;
      RECT 75.13 -266.225 75.43 -222.48 ;
      RECT 75.115 -224.455 75.445 -224.125 ;
      RECT 75.115 -265.815 75.445 -265.485 ;
      RECT 74.515 -309.33 74.815 -233.74 ;
      RECT 74.5 -234.115 74.83 -233.785 ;
      RECT 74.5 -253.595 74.83 -253.265 ;
      RECT 74.5 -309.33 74.83 -309 ;
      RECT 73.9 -248.935 74.2 -234.37 ;
      RECT 73.885 -234.745 74.215 -234.415 ;
      RECT 73.885 -248.935 74.215 -248.605 ;
      RECT 73.27 -296.415 73.6 -296.085 ;
      RECT 73.285 -352.84 73.585 -296.085 ;
      RECT 73.27 -270.47 73.6 -270.14 ;
      RECT 73.285 -285.44 73.585 -270.14 ;
      RECT 73.27 -285.44 73.6 -285.11 ;
      RECT 73.285 -266.245 73.585 -222.48 ;
      RECT 73.27 -222.855 73.6 -222.525 ;
      RECT 73.27 -266.245 73.6 -265.915 ;
      RECT 63.245 -301.805 63.575 -301.475 ;
      RECT 63.26 -345.57 63.56 -301.475 ;
      RECT 63.245 -309.045 63.575 -308.715 ;
      RECT 63.245 -345.525 63.575 -345.195 ;
      RECT 62.615 -308.245 62.945 -307.915 ;
      RECT 62.63 -352.84 62.93 -307.915 ;
      RECT 62 -302.605 62.33 -302.275 ;
      RECT 62.015 -352.84 62.315 -302.275 ;
      RECT 55.115 -270.01 55.445 -269.68 ;
      RECT 55.13 -285.44 55.43 -269.68 ;
      RECT 55.115 -285.44 55.445 -285.11 ;
      RECT 55.13 -266.225 55.43 -222.48 ;
      RECT 55.115 -224.455 55.445 -224.125 ;
      RECT 55.115 -265.815 55.445 -265.485 ;
      RECT 54.515 -301.32 54.815 -233.74 ;
      RECT 54.5 -234.115 54.83 -233.785 ;
      RECT 54.5 -253.595 54.83 -253.265 ;
      RECT 54.5 -301.32 54.83 -300.99 ;
      RECT 53.9 -248.935 54.2 -234.37 ;
      RECT 53.885 -234.745 54.215 -234.415 ;
      RECT 53.885 -248.935 54.215 -248.605 ;
      RECT 53.27 -296.415 53.6 -296.085 ;
      RECT 53.285 -352.84 53.585 -296.085 ;
      RECT 53.27 -270.47 53.6 -270.14 ;
      RECT 53.285 -285.44 53.585 -270.14 ;
      RECT 53.27 -285.44 53.6 -285.11 ;
      RECT 53.285 -266.245 53.585 -222.48 ;
      RECT 53.27 -222.855 53.6 -222.525 ;
      RECT 53.27 -266.245 53.6 -265.915 ;
      RECT 36.3 -318.17 36.6 -238.465 ;
      RECT 36.285 -238.84 36.615 -238.51 ;
      RECT 36.285 -318.17 36.615 -317.84 ;
      RECT 35.115 -270.01 35.445 -269.68 ;
      RECT 35.13 -285.44 35.43 -269.68 ;
      RECT 35.115 -285.44 35.445 -285.11 ;
      RECT 35.13 -266.225 35.43 -222.48 ;
      RECT 35.115 -224.455 35.445 -224.125 ;
      RECT 35.115 -265.815 35.445 -265.485 ;
      RECT 34.515 -309.33 34.815 -233.74 ;
      RECT 34.5 -234.115 34.83 -233.785 ;
      RECT 34.5 -253.595 34.83 -253.265 ;
      RECT 34.5 -309.33 34.83 -309 ;
      RECT 33.9 -248.935 34.2 -234.37 ;
      RECT 33.885 -234.745 34.215 -234.415 ;
      RECT 33.885 -248.935 34.215 -248.605 ;
      RECT 33.27 -296.415 33.6 -296.085 ;
      RECT 33.285 -352.84 33.585 -296.085 ;
      RECT 33.27 -270.47 33.6 -270.14 ;
      RECT 33.285 -285.44 33.585 -270.14 ;
      RECT 33.27 -285.44 33.6 -285.11 ;
      RECT 33.285 -266.245 33.585 -222.48 ;
      RECT 33.27 -222.855 33.6 -222.525 ;
      RECT 33.27 -266.245 33.6 -265.915 ;
      RECT 24.11 -318.545 24.44 -318.215 ;
      RECT 24.125 -352.84 24.425 -318.215 ;
      RECT 23.245 -301.805 23.575 -301.475 ;
      RECT 23.26 -345.57 23.56 -301.475 ;
      RECT 23.245 -309.045 23.575 -308.715 ;
      RECT 23.245 -317.745 23.575 -317.415 ;
      RECT 23.245 -345.525 23.575 -345.195 ;
      RECT 22.615 -308.245 22.945 -307.915 ;
      RECT 22.63 -352.84 22.93 -307.915 ;
      RECT 22 -302.605 22.33 -302.275 ;
      RECT 22.015 -352.84 22.315 -302.275 ;
      RECT 15.115 -270.01 15.445 -269.68 ;
      RECT 15.13 -285.44 15.43 -269.68 ;
      RECT 15.115 -285.44 15.445 -285.11 ;
      RECT 15.13 -266.225 15.43 -222.48 ;
      RECT 15.115 -224.455 15.445 -224.125 ;
      RECT 15.115 -265.815 15.445 -265.485 ;
      RECT 14.515 -301.32 14.815 -233.74 ;
      RECT 14.5 -234.115 14.83 -233.785 ;
      RECT 14.5 -253.595 14.83 -253.265 ;
      RECT 14.5 -301.32 14.83 -300.99 ;
      RECT 13.9 -248.935 14.2 -234.37 ;
      RECT 13.885 -234.745 14.215 -234.415 ;
      RECT 13.885 -248.935 14.215 -248.605 ;
      RECT 13.27 -296.415 13.6 -296.085 ;
      RECT 13.285 -352.84 13.585 -296.085 ;
      RECT 13.27 -270.47 13.6 -270.14 ;
      RECT 13.285 -285.44 13.585 -270.14 ;
      RECT 13.27 -285.44 13.6 -285.11 ;
      RECT 13.285 -266.245 13.585 -222.48 ;
      RECT 13.27 -222.855 13.6 -222.525 ;
      RECT 13.27 -266.245 13.6 -265.915 ;
      RECT 11.005 -260.23 11.335 -259.9 ;
      RECT 11.02 -302.64 11.32 -259.9 ;
      RECT 11.005 -302.64 11.335 -302.31 ;
      RECT -5.91 -323.075 -5.58 -322.745 ;
      RECT -5.895 -341.51 -5.595 -322.745 ;
      RECT -5.91 -341.51 -5.58 -341.18 ;
      RECT -9.505 -341.065 -9.175 -340.735 ;
      RECT -9.49 -345.57 -9.19 -340.735 ;
      RECT -9.505 -345.525 -9.175 -345.195 ;
      RECT -10.34 -213.02 -10.01 -212.69 ;
      RECT -10.325 -304.43 -10.025 -212.69 ;
      RECT -10.34 -304.43 -10.01 -304.1 ;
      RECT -10.635 -341.865 -10.305 -341.535 ;
      RECT -10.62 -352.84 -10.32 -341.535 ;
      RECT -11.75 -327.84 -11.42 -327.51 ;
      RECT -11.735 -341.51 -11.435 -327.51 ;
      RECT -11.75 -341.51 -11.42 -341.18 ;
      RECT -12.385 -327.34 -12.055 -327.01 ;
      RECT -12.37 -342.265 -12.07 -327.01 ;
      RECT -12.385 -342.265 -12.055 -341.935 ;
      RECT -15.345 -341.065 -15.015 -340.735 ;
      RECT -15.33 -345.57 -15.03 -340.735 ;
      RECT -15.345 -345.525 -15.015 -345.195 ;
      RECT -16.475 -341.865 -16.145 -341.535 ;
      RECT -16.46 -352.84 -16.16 -341.535 ;
      RECT -17.59 -328.84 -17.26 -328.51 ;
      RECT -17.575 -341.51 -17.275 -328.51 ;
      RECT -17.59 -341.51 -17.26 -341.18 ;
      RECT -18.225 -328.34 -17.895 -328.01 ;
      RECT -18.21 -342.265 -17.91 -328.01 ;
      RECT -18.225 -342.265 -17.895 -341.935 ;
      RECT -21.185 -341.065 -20.855 -340.735 ;
      RECT -21.17 -345.57 -20.87 -340.735 ;
      RECT -21.185 -345.525 -20.855 -345.195 ;
      RECT -22.315 -341.865 -21.985 -341.535 ;
      RECT -22.3 -352.84 -22 -341.535 ;
      RECT -23.43 -329.84 -23.1 -329.51 ;
      RECT -23.415 -341.51 -23.115 -329.51 ;
      RECT -23.43 -341.51 -23.1 -341.18 ;
      RECT -24.065 -329.34 -23.735 -329.01 ;
      RECT -24.05 -342.265 -23.75 -329.01 ;
      RECT -24.065 -342.265 -23.735 -341.935 ;
      RECT -27.025 -341.065 -26.695 -340.735 ;
      RECT -27.01 -345.57 -26.71 -340.735 ;
      RECT -27.025 -345.525 -26.695 -345.195 ;
      RECT -28.155 -341.865 -27.825 -341.535 ;
      RECT -28.14 -352.84 -27.84 -341.535 ;
      RECT -29.27 -330.84 -28.94 -330.51 ;
      RECT -29.255 -341.51 -28.955 -330.51 ;
      RECT -29.27 -341.51 -28.94 -341.18 ;
      RECT -29.905 -330.34 -29.575 -330.01 ;
      RECT -29.89 -342.265 -29.59 -330.01 ;
      RECT -29.905 -342.265 -29.575 -341.935 ;
      RECT -32.865 -341.065 -32.535 -340.735 ;
      RECT -32.85 -345.57 -32.55 -340.735 ;
      RECT -32.865 -345.525 -32.535 -345.195 ;
      RECT -33.995 -341.865 -33.665 -341.535 ;
      RECT -33.98 -352.84 -33.68 -341.535 ;
      RECT -35.11 -331.84 -34.78 -331.51 ;
      RECT -35.095 -341.51 -34.795 -331.51 ;
      RECT -35.11 -341.51 -34.78 -341.18 ;
      RECT -35.745 -331.34 -35.415 -331.01 ;
      RECT -35.73 -342.265 -35.43 -331.01 ;
      RECT -35.745 -342.265 -35.415 -341.935 ;
      RECT -38.705 -341.065 -38.375 -340.735 ;
      RECT -38.69 -345.57 -38.39 -340.735 ;
      RECT -38.705 -345.525 -38.375 -345.195 ;
      RECT -39.835 -341.865 -39.505 -341.535 ;
      RECT -39.82 -352.84 -39.52 -341.535 ;
      RECT -40.95 -332.84 -40.62 -332.51 ;
      RECT -40.935 -341.51 -40.635 -332.51 ;
      RECT -40.95 -341.51 -40.62 -341.18 ;
      RECT -41.585 -332.34 -41.255 -332.01 ;
      RECT -41.57 -342.265 -41.27 -332.01 ;
      RECT -41.585 -342.265 -41.255 -341.935 ;
      RECT -44.545 -341.065 -44.215 -340.735 ;
      RECT -44.53 -345.57 -44.23 -340.735 ;
      RECT -44.545 -345.525 -44.215 -345.195 ;
      RECT -45.675 -341.865 -45.345 -341.535 ;
      RECT -45.66 -352.84 -45.36 -341.535 ;
      RECT -46.79 -333.84 -46.46 -333.51 ;
      RECT -46.775 -341.51 -46.475 -333.51 ;
      RECT -46.79 -341.51 -46.46 -341.18 ;
      RECT -47.425 -333.34 -47.095 -333.01 ;
      RECT -47.41 -342.265 -47.11 -333.01 ;
      RECT -47.425 -342.265 -47.095 -341.935 ;
      RECT -50.385 -341.065 -50.055 -340.735 ;
      RECT -50.37 -345.57 -50.07 -340.735 ;
      RECT -50.385 -345.525 -50.055 -345.195 ;
      RECT -51.515 -341.865 -51.185 -341.535 ;
      RECT -51.5 -352.84 -51.2 -341.535 ;
      RECT -52.63 -334.84 -52.3 -334.51 ;
      RECT -52.615 -341.51 -52.315 -334.51 ;
      RECT -52.63 -341.51 -52.3 -341.18 ;
      RECT -53.265 -334.34 -52.935 -334.01 ;
      RECT -53.25 -342.265 -52.95 -334.01 ;
      RECT -53.265 -342.265 -52.935 -341.935 ;
      RECT -56.225 -341.065 -55.895 -340.735 ;
      RECT -56.21 -345.57 -55.91 -340.735 ;
      RECT -56.225 -345.525 -55.895 -345.195 ;
      RECT -57.355 -341.865 -57.025 -341.535 ;
      RECT -57.34 -352.84 -57.04 -341.535 ;
      RECT -58.47 -335.84 -58.14 -335.51 ;
      RECT -58.455 -341.51 -58.155 -335.51 ;
      RECT -58.47 -341.51 -58.14 -341.18 ;
      RECT -59.105 -335.34 -58.775 -335.01 ;
      RECT -59.09 -342.265 -58.79 -335.01 ;
      RECT -59.105 -342.265 -58.775 -341.935 ;
      RECT -62.065 -341.065 -61.735 -340.735 ;
      RECT -62.05 -345.57 -61.75 -340.735 ;
      RECT -62.065 -345.525 -61.735 -345.195 ;
      RECT -63.195 -341.865 -62.865 -341.535 ;
      RECT -63.18 -352.84 -62.88 -341.535 ;
      RECT -64.31 -336.84 -63.98 -336.51 ;
      RECT -64.295 -341.51 -63.995 -336.51 ;
      RECT -64.31 -341.51 -63.98 -341.18 ;
      RECT -64.945 -336.34 -64.615 -336.01 ;
      RECT -64.93 -342.265 -64.63 -336.01 ;
      RECT -64.945 -342.265 -64.615 -341.935 ;
      RECT -67.905 -341.065 -67.575 -340.735 ;
      RECT -67.89 -345.57 -67.59 -340.735 ;
      RECT -67.905 -345.525 -67.575 -345.195 ;
      RECT -69.035 -341.865 -68.705 -341.535 ;
      RECT -69.02 -352.84 -68.72 -341.535 ;
      RECT -69.9 -345.57 -69.5 -324.385 ;
      RECT -70.04 -352.72 -69.62 -345.15 ;
  END
END sramgen_sram_1024x32m8w8_replica_v1

END LIBRARY
