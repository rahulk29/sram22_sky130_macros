* Substrate SPICE library
* This is a generated file. Be careful when editing manually: this file may be overwritten.


.SUBCKT mos_w2300_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.300


.ENDS mos_w2300_l150_m1_nf1_id0

.SUBCKT mos_w2900_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.900


.ENDS mos_w2900_l150_m1_nf1_id1

.SUBCKT nand2_2 vdd vss a b y

  Xn1 x a vss vss mos_w2300_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2300_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2900_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2900_l150_m1_nf1_id1

.ENDS nand2_2

.SUBCKT mos_w3380_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.380


.ENDS mos_w3380_l150_m1_nf1_id1

.SUBCKT mos_w1350_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.350


.ENDS mos_w1350_l150_m1_nf1_id0

.SUBCKT folded_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w3380_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1350_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w3380_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1350_l150_m1_nf1_id0

.ENDS folded_inv_6

.SUBCKT and2_1 vdd a b y yb vss

  X0 vdd vss a b yb nand2_2
  X0_1 vdd vss yb y folded_inv_6

.ENDS and2_1

.SUBCKT mos_w700_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id1

.SUBCKT mos_w700_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id0

.SUBCKT multi_finger_inv_8 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_8

.SUBCKT multi_finger_inv_9 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_9

.SUBCKT decoder_stage_5 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] predecode_0_0 predecode_0_1 predecode_0_2 predecode_0_3 predecode_1_0 predecode_1_1 predecode_1_2 predecode_1_3

  Xgate_0_0_0 vdd predecode_0_0 predecode_1_0 x_0[0] y_b_noconn_0_0_0 vss and2_1
  Xgate_0_1_0 vdd predecode_0_1 predecode_1_0 x_0[1] y_b_noconn_0_1_0 vss and2_1
  Xgate_0_2_0 vdd predecode_0_2 predecode_1_0 x_0[2] y_b_noconn_0_2_0 vss and2_1
  Xgate_0_3_0 vdd predecode_0_3 predecode_1_0 x_0[3] y_b_noconn_0_3_0 vss and2_1
  Xgate_0_4_0 vdd predecode_0_0 predecode_1_1 x_0[4] y_b_noconn_0_4_0 vss and2_1
  Xgate_0_5_0 vdd predecode_0_1 predecode_1_1 x_0[5] y_b_noconn_0_5_0 vss and2_1
  Xgate_0_6_0 vdd predecode_0_2 predecode_1_1 x_0[6] y_b_noconn_0_6_0 vss and2_1
  Xgate_0_7_0 vdd predecode_0_3 predecode_1_1 x_0[7] y_b_noconn_0_7_0 vss and2_1
  Xgate_0_8_0 vdd predecode_0_0 predecode_1_2 x_0[8] y_b_noconn_0_8_0 vss and2_1
  Xgate_0_9_0 vdd predecode_0_1 predecode_1_2 x_0[9] y_b_noconn_0_9_0 vss and2_1
  Xgate_0_10_0 vdd predecode_0_2 predecode_1_2 x_0[10] y_b_noconn_0_10_0 vss and2_1
  Xgate_0_11_0 vdd predecode_0_3 predecode_1_2 x_0[11] y_b_noconn_0_11_0 vss and2_1
  Xgate_0_12_0 vdd predecode_0_0 predecode_1_3 x_0[12] y_b_noconn_0_12_0 vss and2_1
  Xgate_0_13_0 vdd predecode_0_1 predecode_1_3 x_0[13] y_b_noconn_0_13_0 vss and2_1
  Xgate_0_14_0 vdd predecode_0_2 predecode_1_3 x_0[14] y_b_noconn_0_14_0 vss and2_1
  Xgate_0_15_0 vdd predecode_0_3 predecode_1_3 x_0[15] y_b_noconn_0_15_0 vss and2_1
  Xgate_1_0_0 vdd vss x_0[0] y_b[0] multi_finger_inv_8
  Xgate_1_1_0 vdd vss x_0[1] y_b[1] multi_finger_inv_8
  Xgate_1_2_0 vdd vss x_0[2] y_b[2] multi_finger_inv_8
  Xgate_1_3_0 vdd vss x_0[3] y_b[3] multi_finger_inv_8
  Xgate_1_4_0 vdd vss x_0[4] y_b[4] multi_finger_inv_8
  Xgate_1_5_0 vdd vss x_0[5] y_b[5] multi_finger_inv_8
  Xgate_1_6_0 vdd vss x_0[6] y_b[6] multi_finger_inv_8
  Xgate_1_7_0 vdd vss x_0[7] y_b[7] multi_finger_inv_8
  Xgate_1_8_0 vdd vss x_0[8] y_b[8] multi_finger_inv_8
  Xgate_1_9_0 vdd vss x_0[9] y_b[9] multi_finger_inv_8
  Xgate_1_10_0 vdd vss x_0[10] y_b[10] multi_finger_inv_8
  Xgate_1_11_0 vdd vss x_0[11] y_b[11] multi_finger_inv_8
  Xgate_1_12_0 vdd vss x_0[12] y_b[12] multi_finger_inv_8
  Xgate_1_13_0 vdd vss x_0[13] y_b[13] multi_finger_inv_8
  Xgate_1_14_0 vdd vss x_0[14] y_b[14] multi_finger_inv_8
  Xgate_1_15_0 vdd vss x_0[15] y_b[15] multi_finger_inv_8
  Xgate_2_0_0 vdd vss y_b[0] y[0] multi_finger_inv_9
  Xgate_2_1_0 vdd vss y_b[1] y[1] multi_finger_inv_9
  Xgate_2_2_0 vdd vss y_b[2] y[2] multi_finger_inv_9
  Xgate_2_3_0 vdd vss y_b[3] y[3] multi_finger_inv_9
  Xgate_2_4_0 vdd vss y_b[4] y[4] multi_finger_inv_9
  Xgate_2_5_0 vdd vss y_b[5] y[5] multi_finger_inv_9
  Xgate_2_6_0 vdd vss y_b[6] y[6] multi_finger_inv_9
  Xgate_2_7_0 vdd vss y_b[7] y[7] multi_finger_inv_9
  Xgate_2_8_0 vdd vss y_b[8] y[8] multi_finger_inv_9
  Xgate_2_9_0 vdd vss y_b[9] y[9] multi_finger_inv_9
  Xgate_2_10_0 vdd vss y_b[10] y[10] multi_finger_inv_9
  Xgate_2_11_0 vdd vss y_b[11] y[11] multi_finger_inv_9
  Xgate_2_12_0 vdd vss y_b[12] y[12] multi_finger_inv_9
  Xgate_2_13_0 vdd vss y_b[13] y[13] multi_finger_inv_9
  Xgate_2_14_0 vdd vss y_b[14] y[14] multi_finger_inv_9
  Xgate_2_15_0 vdd vss y_b[15] y[15] multi_finger_inv_9

.ENDS decoder_stage_5

.SUBCKT mos_w1000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id1

.SUBCKT mos_w600_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.600


.ENDS mos_w600_l150_m1_nf1_id0

.SUBCKT folded_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w600_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w600_l150_m1_nf1_id0

.ENDS folded_inv_7

.SUBCKT sky130_fd_sc_hs__and2_4 A B VGND VNB VPB VPWR X

  X0 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X2 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X5 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X8 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X14 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X15 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_4

.SUBCKT sky130_fd_sc_hs__and2_4_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_4

.ENDS sky130_fd_sc_hs__and2_4_wrapper

.SUBCKT mos_w2000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.000


.ENDS mos_w2000_l150_m1_nf1_id0

.SUBCKT mos_w2500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.500


.ENDS mos_w2500_l150_m1_nf1_id1

.SUBCKT nand2_1 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2_1

.SUBCKT mos_w2880_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.880


.ENDS mos_w2880_l150_m1_nf1_id1

.SUBCKT mos_w1150_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.150


.ENDS mos_w1150_l150_m1_nf1_id0

.SUBCKT folded_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w2880_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1150_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2880_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1150_l150_m1_nf1_id0

.ENDS folded_inv_5

.SUBCKT decoder_stage_9 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 y_b[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 y_b[3] nand2_1
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_5
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_5
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_5
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_5

.ENDS decoder_stage_9

.SUBCKT decoder_3 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  X0 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_stage_9

.ENDS decoder_3

.SUBCKT sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_2

.SUBCKT sky130_fd_sc_hs__inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_2

.ENDS sky130_fd_sc_hs__inv_2_wrapper

.SUBCKT sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_4

.SUBCKT sky130_fd_sc_hs__inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_4

.ENDS sky130_fd_sc_hs__inv_4_wrapper

.SUBCKT inv_chain_9 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_9

.SUBCKT sram_sp_hstrap BR VDD VSS BL VNB VPB

  X0 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140

  X1 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_hstrap

.SUBCKT sram_sp_hstrap_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_hstrap

.ENDS sram_sp_hstrap_wrapper

.SUBCKT sramgen_svt_inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_2

.SUBCKT sramgen_svt_inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_2

.ENDS sramgen_svt_inv_2_wrapper

.SUBCKT sramgen_svt_inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_4

.SUBCKT sramgen_svt_inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_4

.ENDS sramgen_svt_inv_4_wrapper

.SUBCKT svt_inv_chain_18 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sramgen_svt_inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sramgen_svt_inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sramgen_svt_inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sramgen_svt_inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sramgen_svt_inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sramgen_svt_inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sramgen_svt_inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sramgen_svt_inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sramgen_svt_inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sramgen_svt_inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sramgen_svt_inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sramgen_svt_inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sramgen_svt_inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sramgen_svt_inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sramgen_svt_inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sramgen_svt_inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sramgen_svt_inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd dout sramgen_svt_inv_4_wrapper

.ENDS svt_inv_chain_18

.SUBCKT mos_w5000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=5.000


.ENDS mos_w5000_l150_m1_nf1_id1

.SUBCKT folded_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w2000_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w2000_l150_m1_nf1_id0

.ENDS folded_inv_1

.SUBCKT sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X18 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__inv_16

.SUBCKT inv_chain_2 din dout vdd vss

  Xinv0 din vss vss vdd vdd x sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_2

.SUBCKT mos_w500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id1

.SUBCKT multi_finger_inv_11 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_11

.SUBCKT mos_w1250_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.250


.ENDS mos_w1250_l150_m1_nf1_id1

.SUBCKT mos_w500_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id0

.SUBCKT folded_inv vdd vss a y

  XMP0 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w500_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w500_l150_m1_nf1_id0

.ENDS folded_inv

.SUBCKT multi_finger_inv vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv

.SUBCKT multi_finger_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_1

.SUBCKT multi_finger_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_2

.SUBCKT decoder_stage_1 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv
  Xgate_2_0_0 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_2_0_1 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_2_0_2 vdd vss x_1 y_b multi_finger_inv_1
  Xgate_3_0_0 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_1 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_2 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_3 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_4 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_5 vdd vss y_b y multi_finger_inv_2
  Xgate_3_0_6 vdd vss y_b y multi_finger_inv_2

.ENDS decoder_stage_1

.SUBCKT sram_sp_colend BR VDD VSS BL VNB VPB

  X0 BR VNB BR VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_colend

.SUBCKT sram_sp_cell BL BR VDD VSS WL VNB VPB

  X0 QB WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q QB VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 QB WL QB VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q QB VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q QB VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q QB VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell

.SUBCKT sram_sp_cell_wrapper BL BR VDD VSS WL VNB VPB

  X0 BL BR VDD VSS WL VNB VPB sram_sp_cell

.ENDS sram_sp_cell_wrapper

.SUBCKT sramgen_sp_sense_amp clk inn inp outn outp VDD VSS

  XSWOP outp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWON outn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMP midp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMN midn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XPFBP outp outn VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XPFBN outn outp VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XTAIL tail clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=4 w=1.680

  XNFBP outp outn midp VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XNFBN outn outp midn VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINP midn inp tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINN midp inn tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680


.ENDS sramgen_sp_sense_amp

.SUBCKT sramgen_sp_sense_amp_wrapper clk inn inp outn outp VDD VSS

  X0 clk inn inp outn outp VDD VSS sramgen_sp_sense_amp

.ENDS sramgen_sp_sense_amp_wrapper

.SUBCKT sky130_fd_sc_hs__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 a_1800_291# a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X1 VGND CLK a_728_331# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Q a_2363_352# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR CLK a_728_331# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 a_1499_149# a_728_331# a_1586_149# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X5 a_536_81# a_331_392# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X6 a_156_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X7 a_298_294# a_818_418# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X8 a_70_74# a_728_331# a_298_294# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X9 a_331_392# a_728_331# a_1586_149# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 a_70_74# D a_156_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X11 a_818_418# a_728_331# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_818_418# a_728_331# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_1586_149# a_818_418# a_1755_389# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X14 Q_N a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 a_298_294# a_818_418# a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X16 VGND RESET_B a_536_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X17 a_1755_389# a_1800_291# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X18 a_1586_149# a_818_418# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Q a_2363_352# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 VGND a_1586_149# Q_N VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VGND a_1586_149# a_2363_352# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X22 VPWR a_298_294# a_331_392# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X23 a_298_294# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X24 a_1499_149# a_1800_291# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X25 VPWR a_331_392# a_683_485# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X26 VPWR D a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X27 VPWR RESET_B a_1800_291# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X28 a_1974_74# a_1586_149# a_1800_291# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X29 a_70_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X30 Q_N a_1586_149# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 VPWR a_1586_149# a_2363_352# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X32 VGND a_2363_352# Q VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X33 VPWR a_1586_149# Q_N VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND RESET_B a_1974_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X35 a_683_485# a_728_331# a_298_294# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X36 VGND a_298_294# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VPWR a_2363_352# Q VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__dfrbp_2

.SUBCKT sky130_fd_sc_hs__dfrbp_2_wrapper CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 CLK D RESET_B VGND VNB VPB VPWR Q Q_N sky130_fd_sc_hs__dfrbp_2

.ENDS sky130_fd_sc_hs__dfrbp_2_wrapper

.SUBCKT dff_array_8 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_8

.SUBCKT multi_finger_inv_10 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_10

.SUBCKT mos_w1200_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.200


.ENDS mos_w1200_l150_m1_nf1_id1

.SUBCKT folded_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w2900_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1150_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2900_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1150_l150_m1_nf1_id0

.ENDS folded_inv_4

.SUBCKT sky130_fd_sc_hs__mux2_4 A0 A1 S VGND VNB VPB VPWR X

  X0 a_27_368# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 a_722_391# A0 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X2 a_722_391# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X3 VGND a_27_368# a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_193_241# A1 a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X5 a_709_119# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 a_709_119# A1 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X7 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VPWR a_27_368# a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_193_241# A0 a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X12 a_937_119# A0 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_936_391# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X14 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VPWR S a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X17 a_936_391# A1 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X18 a_193_241# A0 a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X19 a_193_241# A1 a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X20 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X21 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X22 a_27_368# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X23 a_937_119# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X24 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND S a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640


.ENDS sky130_fd_sc_hs__mux2_4

.SUBCKT sky130_fd_sc_hs__mux2_4_wrapper A0 A1 S VGND VNB VPB VPWR X

  X0 A0 A1 S VGND VNB VPB VPWR X sky130_fd_sc_hs__mux2_4

.ENDS sky130_fd_sc_hs__mux2_4_wrapper

.SUBCKT decoder_stage_8 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 y_b[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 y_b[3] nand2_1
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_4
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_4
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_4
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_4

.ENDS decoder_stage_8

.SUBCKT nand2 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2

.SUBCKT sky130_fd_sc_hs__nand2_8 A B VGND VNB VPB VPWR Y

  X0 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nand2_8

.SUBCKT inv_chain_13 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_13

.SUBCKT multi_finger_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_3

.SUBCKT multi_finger_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_5

.SUBCKT multi_finger_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_6

.SUBCKT multi_finger_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_7

.SUBCKT decoder_stage_4 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv_5
  Xgate_2_0_0 vdd vss x_1 y_b multi_finger_inv_6
  Xgate_2_0_1 vdd vss x_1 y_b multi_finger_inv_6
  Xgate_2_0_2 vdd vss x_1 y_b multi_finger_inv_6
  Xgate_2_0_3 vdd vss x_1 y_b multi_finger_inv_6
  Xgate_3_0_0 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_1 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_2 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_3 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_4 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_5 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_6 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_7 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_8 vdd vss y_b y multi_finger_inv_7
  Xgate_3_0_9 vdd vss y_b y multi_finger_inv_7

.ENDS decoder_stage_4

.SUBCKT mos_w3500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.500


.ENDS mos_w3500_l150_m1_nf1_id1

.SUBCKT mos_w1400_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.400


.ENDS mos_w1400_l150_m1_nf1_id0

.SUBCKT folded_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w3500_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1400_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w3500_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1400_l150_m1_nf1_id0

.ENDS folded_inv_2

.SUBCKT mos_w2550_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.550


.ENDS mos_w2550_l150_m1_nf1_id1

.SUBCKT mos_w1020_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.020


.ENDS mos_w1020_l150_m1_nf1_id0

.SUBCKT folded_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w2550_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1020_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2550_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1020_l150_m1_nf1_id0

.ENDS folded_inv_3

.SUBCKT decoder_stage_7 vdd vss y y_b predecode_0_0 predecode_1_0

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 x_0 nand2_1
  Xgate_1_0_0 vdd vss x_0 x_1 folded_inv_2
  Xgate_2_0_0 vdd vss x_1 y_b folded_inv_3
  Xgate_2_0_1 vdd vss x_1 y_b folded_inv_3
  Xgate_2_0_2 vdd vss x_1 y_b folded_inv_3
  Xgate_2_0_3 vdd vss x_1 y_b folded_inv_3
  Xgate_3_0_0 vdd vss y_b y folded_inv_3
  Xgate_3_0_1 vdd vss y_b y folded_inv_3
  Xgate_3_0_2 vdd vss y_b y folded_inv_3
  Xgate_3_0_3 vdd vss y_b y folded_inv_3

.ENDS decoder_stage_7

.SUBCKT mos_w800_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.800


.ENDS mos_w800_l150_m1_nf1_id0

.SUBCKT mos_w1200_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.200


.ENDS mos_w1200_l150_m1_nf1_id0

.SUBCKT mos_w1700_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.700


.ENDS mos_w1700_l150_m1_nf1_id1

.SUBCKT column_mos vdd vss bl

  Xgate_nmos vss bl vss vss mos_w800_l150_m1_nf1_id0
  Xdrain_nmos bl vss vss vss mos_w1200_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w1700_l150_m1_nf1_id1

.ENDS column_mos

.SUBCKT multi_finger_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_4

.SUBCKT decoder_stage_3 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_4

.ENDS decoder_stage_3

.SUBCKT sram_sp_cell_replica BL BR VSS VDD VPB VNB WL

  X0 VDD WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q VDD VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 VDD WL VDD VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q VDD VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q VDD VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell_replica

.SUBCKT sky130_fd_sc_hs__nor2_4 A B VGND VNB VPB VPWR Y

  X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nor2_4

.SUBCKT sky130_fd_sc_hs__nand2_8_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_8

.ENDS sky130_fd_sc_hs__nand2_8_wrapper

.SUBCKT sr_latch sb rb q qb vdd vss

  Xnand_set q0b sb vss vss vdd vdd q0 sky130_fd_sc_hs__nand2_8_wrapper
  Xnand_reset q0 rb vss vss vdd vdd q0b sky130_fd_sc_hs__nand2_8_wrapper
  Xqb_inv q0 vss vss vdd vdd qb sky130_fd_sc_hs__inv_2_wrapper
  Xq_inv q0b vss vss vdd vdd q sky130_fd_sc_hs__inv_2_wrapper

.ENDS sr_latch

.SUBCKT sky130_fd_sc_hs__inv_16_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_16

.ENDS sky130_fd_sc_hs__inv_16_wrapper

.SUBCKT inv_chain_12 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_12

.SUBCKT sky130_fd_sc_hs__and2_2 A B VGND VNB VPB VPWR X

  X0 a_31_74# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 X a_31_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 X a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_118_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 a_31_74# A a_118_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VPWR A a_31_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X6 VPWR a_31_74# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND a_31_74# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_2

.SUBCKT sky130_fd_sc_hs__and2_2_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_2

.ENDS sky130_fd_sc_hs__and2_2_wrapper

.SUBCKT edge_detector din dout vdd vss

  Xdelay_chain din delayed vdd vss inv_chain_9
  Xand din delayed vss vss vdd vdd dout sky130_fd_sc_hs__and2_4_wrapper

.ENDS edge_detector

.SUBCKT sky130_fd_sc_hs__buf_16 A VGND VNB VPB VPWR X

  X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X9 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X19 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X24 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X27 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X32 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X33 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X35 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X36 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X38 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X39 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X40 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X41 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X42 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X43 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__buf_16

.SUBCKT sky130_fd_sc_hs__buf_16_wrapper A VGND VNB VPB VPWR X

  X0 A VGND VNB VPB VPWR X sky130_fd_sc_hs__buf_16

.ENDS sky130_fd_sc_hs__buf_16_wrapper

.SUBCKT inv_chain_3 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_3

.SUBCKT inv_chain_18 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sky130_fd_sc_hs__inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sky130_fd_sc_hs__inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sky130_fd_sc_hs__inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sky130_fd_sc_hs__inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_18

.SUBCKT sky130_fd_sc_hs__nor2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nor2_4

.ENDS sky130_fd_sc_hs__nor2_4_wrapper

.SUBCKT sky130_fd_sc_hs__nand2_4 A B VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__nand2_4

.SUBCKT sky130_fd_sc_hs__nand2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_4

.ENDS sky130_fd_sc_hs__nand2_4_wrapper

.SUBCKT control_logic_replica_v2 clk ce we rstb rbl saen pc_b rwl wlen wrdrven vdd vss

  Xreset_inv rstb vss vss vdd vdd reset sky130_fd_sc_hs__inv_16_wrapper
  Xclk_delay clk clkd vdd vss inv_chain_12
  Xclk_gate clkd ce vss vss vdd vdd clk_buf sky130_fd_sc_hs__and2_2_wrapper
  Xclk_pulse clk_buf clkp0 vdd vss edge_detector
  Xclk_pulse_buf clkp0 vss vss vdd vdd clkp sky130_fd_sc_hs__buf_16_wrapper
  Xclk_pulse_inv clkp vss vss vdd vdd clkp_b sky130_fd_sc_hs__inv_16_wrapper
  Xclkp_delay clkp_b clkpd vdd vss inv_chain_3
  Xclkpd_inv clkpd vss vss vdd vdd clkpd_b sky130_fd_sc_hs__inv_2_wrapper
  Xclkpd_delay clkpd_b clkpdd vdd vss inv_chain_13
  Xmux_wlen_rst rbl_b clkpdd we vss vss vdd vdd decrepstart sky130_fd_sc_hs__mux2_4_wrapper
  Xdecoder_replica decrepstart decrepend vdd vss svt_inv_chain_18
  Xdecoder_replica_delay decrepend wlen_rst_decoderd vdd vss inv_chain_18
  Xinv_we we vss vss vdd vdd we_b sky130_fd_sc_hs__inv_2_wrapper
  Xinv_rbl rbl vss vss vdd vdd rbl_b sky130_fd_sc_hs__inv_2_wrapper
  Xwlen_grst decrepstart reset vss vss vdd vdd wlen_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xpc_set wlen_rst_decoderd reset vss vss vdd vdd pc_set_b sky130_fd_sc_hs__nor2_4_wrapper
  Xwrdrven_grst decrepend reset vss vss vdd vdd wrdrven_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xclkp_grst clkp reset vss vss vdd vdd clkp_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xnand_sense_en we_b decrepend vss vss vdd vdd saen_set_b sky130_fd_sc_hs__nand2_4_wrapper
  Xnand_wlendb_web rbl_b we_b vss vss vdd vdd wlend sky130_fd_sc_hs__nand2_4_wrapper
  Xand_wlen wlen_q wlend vss vss vdd vdd wlen sky130_fd_sc_hs__and2_4_wrapper
  Xrwl_buf wlen_q vss vss vdd vdd rwl sky130_fd_sc_hs__buf_16_wrapper
  Xwl_ctl clkpd_b wlen_grst_b wlen_q wlen_b vdd vss sr_latch
  Xsaen_ctl saen_set_b clkp_grst_b saen saen_b vdd vss sr_latch
  Xpc_ctl pc_set_b clkp_b pc pc_b0 vdd vss sr_latch
  Xpc_b_buf pc_b0 vss vss vdd vdd pc_b sky130_fd_sc_hs__buf_16_wrapper
  Xwrdrven_set clkpd we vss vss vdd vdd wrdrven_set_b0 sky130_fd_sc_hs__nand2_4_wrapper
  Xwrdrven_set_delay wrdrven_set_b0 wrdrven_set_b vdd vss inv_chain_2
  Xwrdrven_ctl wrdrven_set_b wrdrven_grst_b wrdrven wrdrven_b vdd vss sr_latch

.ENDS control_logic_replica_v2

.SUBCKT decoder_stage_2 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_3
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_3

.ENDS decoder_stage_2

.SUBCKT sram_sp_cell_replica_wrapper BL BR VSS VDD VPB VNB WL

  X0 BL BR VSS VDD VPB VNB WL sram_sp_cell_replica

.ENDS sram_sp_cell_replica_wrapper

.SUBCKT mos_w1800_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.800


.ENDS mos_w1800_l150_m1_nf1_id1

.SUBCKT mos_w1000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id0

.SUBCKT dff_array_1 vdd vss clk rb d q qn

  Xdff_0 clk d rb vss vss vdd vdd q qn sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_1

.SUBCKT mos_w800_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.800


.ENDS mos_w800_l150_m1_nf1_id1

.SUBCKT precharge_1 vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w800_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w800_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w500_l150_m1_nf1_id1

.ENDS precharge_1

.SUBCKT tgate_mux sel_b sel bl br bl_out br_out vdd vss

  XMPBL bl_out sel_b bl vdd mos_w1800_l150_m1_nf1_id1
  XMPBR br_out sel_b br vdd mos_w1800_l150_m1_nf1_id1
  XMNBL bl_out sel bl vss mos_w1200_l150_m1_nf1_id0
  XMNBR br_out sel br vss mos_w1200_l150_m1_nf1_id0

.ENDS tgate_mux

.SUBCKT tristate_inv din en en_b din_b vdd vss

  Xmn_en din_b en nint vss mos_w1200_l150_m1_nf1_id0
  Xmn_pd nint din vss vss mos_w1200_l150_m1_nf1_id0
  Xmp_en din_b en_b pint vdd mos_w1200_l150_m1_nf1_id1
  Xmp_pu pint din vdd vdd mos_w1200_l150_m1_nf1_id1

.ENDS tristate_inv

.SUBCKT write_driver en en_b data data_b bl br vdd vss

  Xbldriver data_b en en_b bl vdd vss tristate_inv
  Xbrdriver data en en_b br vdd vss tristate_inv

.ENDS write_driver

.SUBCKT diff_latch vdd vss din1 din2 dout1 dout2

  Xinbuf_1 vdd vss din1 rst folded_inv_7
  Xinbuf_2 vdd vss din2 set folded_inv_7
  Xoutbuf_1 vdd vss q dout2 folded_inv_7
  Xoutbuf_2 vdd vss qb dout1 folded_inv_7
  Xinvq_1 vdd vss q qb folded_inv_7
  Xinvq_2 vdd vss qb q folded_inv_7
  XMN10 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN11 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN20 qb set vss vss mos_w1000_l150_m1_nf1_id0
  XMN21 qb set vss vss mos_w1000_l150_m1_nf1_id0

.ENDS diff_latch

.SUBCKT column clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] br[0] br[1] br[2] br[3] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we we_b din dout sense_en

  Xprecharge_0 vdd bl[0] br[0] pc_b precharge_1
  Xmux_0 sel_b[0] sel[0] bl[0] br[0] bl_out br_out vdd vss tgate_mux
  Xprecharge_1 vdd bl[1] br[1] pc_b precharge_1
  Xmux_1 sel_b[1] sel[1] bl[1] br[1] bl_out br_out vdd vss tgate_mux
  Xprecharge_2 vdd bl[2] br[2] pc_b precharge_1
  Xmux_2 sel_b[2] sel[2] bl[2] br[2] bl_out br_out vdd vss tgate_mux
  Xprecharge_3 vdd bl[3] br[3] pc_b precharge_1
  Xmux_3 sel_b[3] sel[3] bl[3] br[3] bl_out br_out vdd vss tgate_mux
  Xwrite_driver we we_b q q_b bl_out br_out vdd vss write_driver
  Xsense_amp sense_en br_out bl_out sa_outn sa_outp vdd vss sramgen_sp_sense_amp_wrapper
  Xlatch vdd vss sa_outp sa_outn dout diff_latch_outn diff_latch
  Xdff clk din rstb vss vss vdd vdd q q_b sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS column

.SUBCKT col_peripherals clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we wmask din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21]

  Xwmask_dffs vdd vss clk rstb wmask wmask_in wmask_in_b dff_array_1
  Xwmask_and_0 vdd vss we_i we_ib we wmask_in decoder_stage_7
  Xcol_group_0 clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] br[0] br[1] br[2] br[3] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[0] dout[0] sense_en column
  Xcol_group_1 clk rstb vdd vss bl[4] bl[5] bl[6] bl[7] br[4] br[5] br[6] br[7] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[1] dout[1] sense_en column
  Xcol_group_2 clk rstb vdd vss bl[8] bl[9] bl[10] bl[11] br[8] br[9] br[10] br[11] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[2] dout[2] sense_en column
  Xcol_group_3 clk rstb vdd vss bl[12] bl[13] bl[14] bl[15] br[12] br[13] br[14] br[15] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[3] dout[3] sense_en column
  Xcol_group_4 clk rstb vdd vss bl[16] bl[17] bl[18] bl[19] br[16] br[17] br[18] br[19] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[4] dout[4] sense_en column
  Xcol_group_5 clk rstb vdd vss bl[20] bl[21] bl[22] bl[23] br[20] br[21] br[22] br[23] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[5] dout[5] sense_en column
  Xcol_group_6 clk rstb vdd vss bl[24] bl[25] bl[26] bl[27] br[24] br[25] br[26] br[27] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[6] dout[6] sense_en column
  Xcol_group_7 clk rstb vdd vss bl[28] bl[29] bl[30] bl[31] br[28] br[29] br[30] br[31] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[7] dout[7] sense_en column
  Xcol_group_8 clk rstb vdd vss bl[32] bl[33] bl[34] bl[35] br[32] br[33] br[34] br[35] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[8] dout[8] sense_en column
  Xcol_group_9 clk rstb vdd vss bl[36] bl[37] bl[38] bl[39] br[36] br[37] br[38] br[39] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[9] dout[9] sense_en column
  Xcol_group_10 clk rstb vdd vss bl[40] bl[41] bl[42] bl[43] br[40] br[41] br[42] br[43] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[10] dout[10] sense_en column
  Xcol_group_11 clk rstb vdd vss bl[44] bl[45] bl[46] bl[47] br[44] br[45] br[46] br[47] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[11] dout[11] sense_en column
  Xcol_group_12 clk rstb vdd vss bl[48] bl[49] bl[50] bl[51] br[48] br[49] br[50] br[51] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[12] dout[12] sense_en column
  Xcol_group_13 clk rstb vdd vss bl[52] bl[53] bl[54] bl[55] br[52] br[53] br[54] br[55] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[13] dout[13] sense_en column
  Xcol_group_14 clk rstb vdd vss bl[56] bl[57] bl[58] bl[59] br[56] br[57] br[58] br[59] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[14] dout[14] sense_en column
  Xcol_group_15 clk rstb vdd vss bl[60] bl[61] bl[62] bl[63] br[60] br[61] br[62] br[63] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[15] dout[15] sense_en column
  Xcol_group_16 clk rstb vdd vss bl[64] bl[65] bl[66] bl[67] br[64] br[65] br[66] br[67] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[16] dout[16] sense_en column
  Xcol_group_17 clk rstb vdd vss bl[68] bl[69] bl[70] bl[71] br[68] br[69] br[70] br[71] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[17] dout[17] sense_en column
  Xcol_group_18 clk rstb vdd vss bl[72] bl[73] bl[74] bl[75] br[72] br[73] br[74] br[75] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[18] dout[18] sense_en column
  Xcol_group_19 clk rstb vdd vss bl[76] bl[77] bl[78] bl[79] br[76] br[77] br[78] br[79] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[19] dout[19] sense_en column
  Xcol_group_20 clk rstb vdd vss bl[80] bl[81] bl[82] bl[83] br[80] br[81] br[82] br[83] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[20] dout[20] sense_en column
  Xcol_group_21 clk rstb vdd vss bl[84] bl[85] bl[86] bl[87] br[84] br[85] br[86] br[87] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i we_ib din[21] dout[21] sense_en column

.ENDS col_peripherals

.SUBCKT and2 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_1

.ENDS and2

.SUBCKT decoder_stage vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] wl_en in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7]

  Xgate_0_0_0 vdd wl_en in[0] y[0] y_b[0] vss and2
  Xgate_0_1_0 vdd wl_en in[1] y[1] y_b[1] vss and2
  Xgate_0_2_0 vdd wl_en in[2] y[2] y_b[2] vss and2
  Xgate_0_3_0 vdd wl_en in[3] y[3] y_b[3] vss and2
  Xgate_0_4_0 vdd wl_en in[4] y[4] y_b[4] vss and2
  Xgate_0_5_0 vdd wl_en in[5] y[5] y_b[5] vss and2
  Xgate_0_6_0 vdd wl_en in[6] y[6] y_b[6] vss and2
  Xgate_0_7_0 vdd wl_en in[7] y[7] y_b[7] vss and2

.ENDS decoder_stage

.SUBCKT decoder_2 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  X0 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_stage_8

.ENDS decoder_2

.SUBCKT decoder vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1

  X0 vdd vss child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_noconn_0[0] child_noconn_0[1] child_noconn_0[2] child_noconn_0[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_2
  X0_1 vdd vss child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_noconn_1[0] child_noconn_1[1] child_noconn_1[2] child_noconn_1[3] predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 decoder_3
  X0_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] decoder_stage_5

.ENDS decoder

.SUBCKT multi_finger_inv_12 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_12

.SUBCKT decoder_stage_6 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 x_0[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 x_0[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 x_0[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 x_0[3] nand2_1
  Xgate_1_0_0 vdd vss x_0[0] x_1[0] multi_finger_inv_10
  Xgate_1_1_0 vdd vss x_0[1] x_1[1] multi_finger_inv_10
  Xgate_1_2_0 vdd vss x_0[2] x_1[2] multi_finger_inv_10
  Xgate_1_3_0 vdd vss x_0[3] x_1[3] multi_finger_inv_10
  Xgate_2_0_0 vdd vss x_1[0] y_b[0] multi_finger_inv_11
  Xgate_2_0_1 vdd vss x_1[0] y_b[0] multi_finger_inv_11
  Xgate_2_1_0 vdd vss x_1[1] y_b[1] multi_finger_inv_11
  Xgate_2_1_1 vdd vss x_1[1] y_b[1] multi_finger_inv_11
  Xgate_2_2_0 vdd vss x_1[2] y_b[2] multi_finger_inv_11
  Xgate_2_2_1 vdd vss x_1[2] y_b[2] multi_finger_inv_11
  Xgate_2_3_0 vdd vss x_1[3] y_b[3] multi_finger_inv_11
  Xgate_2_3_1 vdd vss x_1[3] y_b[3] multi_finger_inv_11
  Xgate_3_0_0 vdd vss y_b[0] y[0] multi_finger_inv_12
  Xgate_3_0_1 vdd vss y_b[0] y[0] multi_finger_inv_12
  Xgate_3_0_2 vdd vss y_b[0] y[0] multi_finger_inv_12
  Xgate_3_0_3 vdd vss y_b[0] y[0] multi_finger_inv_12
  Xgate_3_1_0 vdd vss y_b[1] y[1] multi_finger_inv_12
  Xgate_3_1_1 vdd vss y_b[1] y[1] multi_finger_inv_12
  Xgate_3_1_2 vdd vss y_b[1] y[1] multi_finger_inv_12
  Xgate_3_1_3 vdd vss y_b[1] y[1] multi_finger_inv_12
  Xgate_3_2_0 vdd vss y_b[2] y[2] multi_finger_inv_12
  Xgate_3_2_1 vdd vss y_b[2] y[2] multi_finger_inv_12
  Xgate_3_2_2 vdd vss y_b[2] y[2] multi_finger_inv_12
  Xgate_3_2_3 vdd vss y_b[2] y[2] multi_finger_inv_12
  Xgate_3_3_0 vdd vss y_b[3] y[3] multi_finger_inv_12
  Xgate_3_3_1 vdd vss y_b[3] y[3] multi_finger_inv_12
  Xgate_3_3_2 vdd vss y_b[3] y[3] multi_finger_inv_12
  Xgate_3_3_3 vdd vss y_b[3] y[3] multi_finger_inv_12

.ENDS decoder_stage_6

.SUBCKT decoder_1 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  X0 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_stage_6

.ENDS decoder_1

.SUBCKT sram_sp_colend_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_colend

.ENDS sram_sp_colend_wrapper

.SUBCKT sram_sp_horiz_wlstrap_p2 VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_horiz_wlstrap_p2

.SUBCKT sram_sp_horiz_wlstrap_p2_wrapper VSS VNB

  X0 VSS VNB sram_sp_horiz_wlstrap_p2

.ENDS sram_sp_horiz_wlstrap_p2_wrapper

.SUBCKT sp_cell_array vdd vss dummy_bl dummy_br bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15]

  Xcell_0_0 bl[0] br[0] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_1 bl[1] br[1] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_2 bl[2] br[2] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_3 bl[3] br[3] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_4 bl[4] br[4] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_5 bl[5] br[5] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_6 bl[6] br[6] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_7 bl[7] br[7] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_8 bl[8] br[8] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_9 bl[9] br[9] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_10 bl[10] br[10] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_11 bl[11] br[11] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_12 bl[12] br[12] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_13 bl[13] br[13] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_14 bl[14] br[14] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_15 bl[15] br[15] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_16 bl[16] br[16] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_17 bl[17] br[17] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_18 bl[18] br[18] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_19 bl[19] br[19] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_20 bl[20] br[20] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_21 bl[21] br[21] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_22 bl[22] br[22] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_23 bl[23] br[23] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_24 bl[24] br[24] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_25 bl[25] br[25] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_26 bl[26] br[26] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_27 bl[27] br[27] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_28 bl[28] br[28] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_29 bl[29] br[29] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_30 bl[30] br[30] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_31 bl[31] br[31] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_32 bl[32] br[32] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_33 bl[33] br[33] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_34 bl[34] br[34] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_35 bl[35] br[35] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_36 bl[36] br[36] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_37 bl[37] br[37] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_38 bl[38] br[38] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_39 bl[39] br[39] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_40 bl[40] br[40] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_41 bl[41] br[41] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_42 bl[42] br[42] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_43 bl[43] br[43] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_44 bl[44] br[44] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_45 bl[45] br[45] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_46 bl[46] br[46] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_47 bl[47] br[47] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_48 bl[48] br[48] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_49 bl[49] br[49] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_50 bl[50] br[50] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_51 bl[51] br[51] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_52 bl[52] br[52] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_53 bl[53] br[53] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_54 bl[54] br[54] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_55 bl[55] br[55] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_56 bl[56] br[56] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_57 bl[57] br[57] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_58 bl[58] br[58] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_59 bl[59] br[59] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_60 bl[60] br[60] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_61 bl[61] br[61] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_62 bl[62] br[62] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_63 bl[63] br[63] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_64 bl[64] br[64] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_65 bl[65] br[65] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_66 bl[66] br[66] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_67 bl[67] br[67] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_68 bl[68] br[68] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_69 bl[69] br[69] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_70 bl[70] br[70] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_71 bl[71] br[71] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_72 bl[72] br[72] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_73 bl[73] br[73] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_74 bl[74] br[74] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_75 bl[75] br[75] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_76 bl[76] br[76] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_77 bl[77] br[77] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_78 bl[78] br[78] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_79 bl[79] br[79] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_80 bl[80] br[80] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_81 bl[81] br[81] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_82 bl[82] br[82] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_83 bl[83] br[83] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_84 bl[84] br[84] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_85 bl[85] br[85] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_86 bl[86] br[86] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_87 bl[87] br[87] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_1_0 bl[0] br[0] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_1 bl[1] br[1] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_2 bl[2] br[2] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_3 bl[3] br[3] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_4 bl[4] br[4] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_5 bl[5] br[5] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_6 bl[6] br[6] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_7 bl[7] br[7] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_8 bl[8] br[8] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_9 bl[9] br[9] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_10 bl[10] br[10] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_11 bl[11] br[11] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_12 bl[12] br[12] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_13 bl[13] br[13] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_14 bl[14] br[14] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_15 bl[15] br[15] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_16 bl[16] br[16] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_17 bl[17] br[17] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_18 bl[18] br[18] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_19 bl[19] br[19] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_20 bl[20] br[20] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_21 bl[21] br[21] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_22 bl[22] br[22] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_23 bl[23] br[23] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_24 bl[24] br[24] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_25 bl[25] br[25] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_26 bl[26] br[26] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_27 bl[27] br[27] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_28 bl[28] br[28] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_29 bl[29] br[29] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_30 bl[30] br[30] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_31 bl[31] br[31] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_32 bl[32] br[32] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_33 bl[33] br[33] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_34 bl[34] br[34] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_35 bl[35] br[35] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_36 bl[36] br[36] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_37 bl[37] br[37] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_38 bl[38] br[38] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_39 bl[39] br[39] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_40 bl[40] br[40] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_41 bl[41] br[41] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_42 bl[42] br[42] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_43 bl[43] br[43] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_44 bl[44] br[44] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_45 bl[45] br[45] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_46 bl[46] br[46] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_47 bl[47] br[47] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_48 bl[48] br[48] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_49 bl[49] br[49] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_50 bl[50] br[50] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_51 bl[51] br[51] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_52 bl[52] br[52] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_53 bl[53] br[53] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_54 bl[54] br[54] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_55 bl[55] br[55] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_56 bl[56] br[56] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_57 bl[57] br[57] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_58 bl[58] br[58] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_59 bl[59] br[59] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_60 bl[60] br[60] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_61 bl[61] br[61] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_62 bl[62] br[62] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_63 bl[63] br[63] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_64 bl[64] br[64] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_65 bl[65] br[65] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_66 bl[66] br[66] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_67 bl[67] br[67] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_68 bl[68] br[68] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_69 bl[69] br[69] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_70 bl[70] br[70] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_71 bl[71] br[71] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_72 bl[72] br[72] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_73 bl[73] br[73] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_74 bl[74] br[74] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_75 bl[75] br[75] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_76 bl[76] br[76] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_77 bl[77] br[77] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_78 bl[78] br[78] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_79 bl[79] br[79] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_80 bl[80] br[80] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_81 bl[81] br[81] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_82 bl[82] br[82] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_83 bl[83] br[83] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_84 bl[84] br[84] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_85 bl[85] br[85] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_86 bl[86] br[86] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_87 bl[87] br[87] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_2_0 bl[0] br[0] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_1 bl[1] br[1] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_2 bl[2] br[2] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_3 bl[3] br[3] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_4 bl[4] br[4] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_5 bl[5] br[5] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_6 bl[6] br[6] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_7 bl[7] br[7] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_8 bl[8] br[8] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_9 bl[9] br[9] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_10 bl[10] br[10] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_11 bl[11] br[11] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_12 bl[12] br[12] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_13 bl[13] br[13] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_14 bl[14] br[14] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_15 bl[15] br[15] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_16 bl[16] br[16] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_17 bl[17] br[17] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_18 bl[18] br[18] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_19 bl[19] br[19] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_20 bl[20] br[20] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_21 bl[21] br[21] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_22 bl[22] br[22] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_23 bl[23] br[23] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_24 bl[24] br[24] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_25 bl[25] br[25] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_26 bl[26] br[26] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_27 bl[27] br[27] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_28 bl[28] br[28] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_29 bl[29] br[29] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_30 bl[30] br[30] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_31 bl[31] br[31] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_32 bl[32] br[32] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_33 bl[33] br[33] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_34 bl[34] br[34] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_35 bl[35] br[35] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_36 bl[36] br[36] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_37 bl[37] br[37] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_38 bl[38] br[38] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_39 bl[39] br[39] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_40 bl[40] br[40] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_41 bl[41] br[41] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_42 bl[42] br[42] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_43 bl[43] br[43] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_44 bl[44] br[44] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_45 bl[45] br[45] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_46 bl[46] br[46] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_47 bl[47] br[47] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_48 bl[48] br[48] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_49 bl[49] br[49] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_50 bl[50] br[50] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_51 bl[51] br[51] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_52 bl[52] br[52] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_53 bl[53] br[53] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_54 bl[54] br[54] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_55 bl[55] br[55] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_56 bl[56] br[56] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_57 bl[57] br[57] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_58 bl[58] br[58] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_59 bl[59] br[59] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_60 bl[60] br[60] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_61 bl[61] br[61] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_62 bl[62] br[62] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_63 bl[63] br[63] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_64 bl[64] br[64] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_65 bl[65] br[65] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_66 bl[66] br[66] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_67 bl[67] br[67] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_68 bl[68] br[68] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_69 bl[69] br[69] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_70 bl[70] br[70] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_71 bl[71] br[71] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_72 bl[72] br[72] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_73 bl[73] br[73] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_74 bl[74] br[74] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_75 bl[75] br[75] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_76 bl[76] br[76] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_77 bl[77] br[77] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_78 bl[78] br[78] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_79 bl[79] br[79] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_80 bl[80] br[80] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_81 bl[81] br[81] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_82 bl[82] br[82] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_83 bl[83] br[83] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_84 bl[84] br[84] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_85 bl[85] br[85] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_86 bl[86] br[86] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_87 bl[87] br[87] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_3_0 bl[0] br[0] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_1 bl[1] br[1] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_2 bl[2] br[2] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_3 bl[3] br[3] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_4 bl[4] br[4] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_5 bl[5] br[5] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_6 bl[6] br[6] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_7 bl[7] br[7] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_8 bl[8] br[8] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_9 bl[9] br[9] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_10 bl[10] br[10] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_11 bl[11] br[11] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_12 bl[12] br[12] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_13 bl[13] br[13] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_14 bl[14] br[14] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_15 bl[15] br[15] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_16 bl[16] br[16] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_17 bl[17] br[17] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_18 bl[18] br[18] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_19 bl[19] br[19] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_20 bl[20] br[20] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_21 bl[21] br[21] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_22 bl[22] br[22] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_23 bl[23] br[23] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_24 bl[24] br[24] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_25 bl[25] br[25] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_26 bl[26] br[26] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_27 bl[27] br[27] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_28 bl[28] br[28] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_29 bl[29] br[29] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_30 bl[30] br[30] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_31 bl[31] br[31] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_32 bl[32] br[32] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_33 bl[33] br[33] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_34 bl[34] br[34] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_35 bl[35] br[35] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_36 bl[36] br[36] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_37 bl[37] br[37] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_38 bl[38] br[38] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_39 bl[39] br[39] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_40 bl[40] br[40] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_41 bl[41] br[41] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_42 bl[42] br[42] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_43 bl[43] br[43] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_44 bl[44] br[44] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_45 bl[45] br[45] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_46 bl[46] br[46] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_47 bl[47] br[47] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_48 bl[48] br[48] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_49 bl[49] br[49] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_50 bl[50] br[50] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_51 bl[51] br[51] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_52 bl[52] br[52] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_53 bl[53] br[53] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_54 bl[54] br[54] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_55 bl[55] br[55] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_56 bl[56] br[56] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_57 bl[57] br[57] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_58 bl[58] br[58] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_59 bl[59] br[59] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_60 bl[60] br[60] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_61 bl[61] br[61] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_62 bl[62] br[62] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_63 bl[63] br[63] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_64 bl[64] br[64] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_65 bl[65] br[65] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_66 bl[66] br[66] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_67 bl[67] br[67] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_68 bl[68] br[68] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_69 bl[69] br[69] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_70 bl[70] br[70] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_71 bl[71] br[71] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_72 bl[72] br[72] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_73 bl[73] br[73] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_74 bl[74] br[74] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_75 bl[75] br[75] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_76 bl[76] br[76] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_77 bl[77] br[77] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_78 bl[78] br[78] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_79 bl[79] br[79] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_80 bl[80] br[80] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_81 bl[81] br[81] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_82 bl[82] br[82] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_83 bl[83] br[83] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_84 bl[84] br[84] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_85 bl[85] br[85] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_86 bl[86] br[86] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_87 bl[87] br[87] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_4_0 bl[0] br[0] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_1 bl[1] br[1] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_2 bl[2] br[2] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_3 bl[3] br[3] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_4 bl[4] br[4] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_5 bl[5] br[5] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_6 bl[6] br[6] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_7 bl[7] br[7] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_8 bl[8] br[8] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_9 bl[9] br[9] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_10 bl[10] br[10] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_11 bl[11] br[11] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_12 bl[12] br[12] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_13 bl[13] br[13] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_14 bl[14] br[14] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_15 bl[15] br[15] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_16 bl[16] br[16] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_17 bl[17] br[17] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_18 bl[18] br[18] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_19 bl[19] br[19] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_20 bl[20] br[20] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_21 bl[21] br[21] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_22 bl[22] br[22] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_23 bl[23] br[23] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_24 bl[24] br[24] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_25 bl[25] br[25] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_26 bl[26] br[26] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_27 bl[27] br[27] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_28 bl[28] br[28] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_29 bl[29] br[29] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_30 bl[30] br[30] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_31 bl[31] br[31] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_32 bl[32] br[32] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_33 bl[33] br[33] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_34 bl[34] br[34] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_35 bl[35] br[35] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_36 bl[36] br[36] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_37 bl[37] br[37] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_38 bl[38] br[38] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_39 bl[39] br[39] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_40 bl[40] br[40] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_41 bl[41] br[41] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_42 bl[42] br[42] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_43 bl[43] br[43] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_44 bl[44] br[44] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_45 bl[45] br[45] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_46 bl[46] br[46] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_47 bl[47] br[47] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_48 bl[48] br[48] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_49 bl[49] br[49] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_50 bl[50] br[50] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_51 bl[51] br[51] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_52 bl[52] br[52] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_53 bl[53] br[53] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_54 bl[54] br[54] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_55 bl[55] br[55] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_56 bl[56] br[56] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_57 bl[57] br[57] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_58 bl[58] br[58] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_59 bl[59] br[59] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_60 bl[60] br[60] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_61 bl[61] br[61] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_62 bl[62] br[62] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_63 bl[63] br[63] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_64 bl[64] br[64] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_65 bl[65] br[65] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_66 bl[66] br[66] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_67 bl[67] br[67] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_68 bl[68] br[68] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_69 bl[69] br[69] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_70 bl[70] br[70] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_71 bl[71] br[71] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_72 bl[72] br[72] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_73 bl[73] br[73] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_74 bl[74] br[74] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_75 bl[75] br[75] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_76 bl[76] br[76] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_77 bl[77] br[77] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_78 bl[78] br[78] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_79 bl[79] br[79] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_80 bl[80] br[80] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_81 bl[81] br[81] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_82 bl[82] br[82] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_83 bl[83] br[83] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_84 bl[84] br[84] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_85 bl[85] br[85] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_86 bl[86] br[86] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_87 bl[87] br[87] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_5_0 bl[0] br[0] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_1 bl[1] br[1] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_2 bl[2] br[2] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_3 bl[3] br[3] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_4 bl[4] br[4] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_5 bl[5] br[5] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_6 bl[6] br[6] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_7 bl[7] br[7] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_8 bl[8] br[8] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_9 bl[9] br[9] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_10 bl[10] br[10] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_11 bl[11] br[11] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_12 bl[12] br[12] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_13 bl[13] br[13] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_14 bl[14] br[14] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_15 bl[15] br[15] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_16 bl[16] br[16] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_17 bl[17] br[17] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_18 bl[18] br[18] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_19 bl[19] br[19] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_20 bl[20] br[20] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_21 bl[21] br[21] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_22 bl[22] br[22] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_23 bl[23] br[23] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_24 bl[24] br[24] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_25 bl[25] br[25] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_26 bl[26] br[26] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_27 bl[27] br[27] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_28 bl[28] br[28] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_29 bl[29] br[29] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_30 bl[30] br[30] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_31 bl[31] br[31] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_32 bl[32] br[32] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_33 bl[33] br[33] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_34 bl[34] br[34] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_35 bl[35] br[35] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_36 bl[36] br[36] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_37 bl[37] br[37] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_38 bl[38] br[38] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_39 bl[39] br[39] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_40 bl[40] br[40] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_41 bl[41] br[41] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_42 bl[42] br[42] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_43 bl[43] br[43] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_44 bl[44] br[44] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_45 bl[45] br[45] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_46 bl[46] br[46] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_47 bl[47] br[47] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_48 bl[48] br[48] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_49 bl[49] br[49] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_50 bl[50] br[50] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_51 bl[51] br[51] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_52 bl[52] br[52] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_53 bl[53] br[53] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_54 bl[54] br[54] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_55 bl[55] br[55] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_56 bl[56] br[56] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_57 bl[57] br[57] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_58 bl[58] br[58] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_59 bl[59] br[59] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_60 bl[60] br[60] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_61 bl[61] br[61] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_62 bl[62] br[62] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_63 bl[63] br[63] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_64 bl[64] br[64] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_65 bl[65] br[65] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_66 bl[66] br[66] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_67 bl[67] br[67] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_68 bl[68] br[68] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_69 bl[69] br[69] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_70 bl[70] br[70] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_71 bl[71] br[71] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_72 bl[72] br[72] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_73 bl[73] br[73] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_74 bl[74] br[74] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_75 bl[75] br[75] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_76 bl[76] br[76] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_77 bl[77] br[77] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_78 bl[78] br[78] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_79 bl[79] br[79] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_80 bl[80] br[80] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_81 bl[81] br[81] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_82 bl[82] br[82] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_83 bl[83] br[83] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_84 bl[84] br[84] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_85 bl[85] br[85] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_86 bl[86] br[86] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_87 bl[87] br[87] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_6_0 bl[0] br[0] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_1 bl[1] br[1] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_2 bl[2] br[2] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_3 bl[3] br[3] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_4 bl[4] br[4] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_5 bl[5] br[5] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_6 bl[6] br[6] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_7 bl[7] br[7] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_8 bl[8] br[8] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_9 bl[9] br[9] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_10 bl[10] br[10] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_11 bl[11] br[11] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_12 bl[12] br[12] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_13 bl[13] br[13] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_14 bl[14] br[14] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_15 bl[15] br[15] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_16 bl[16] br[16] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_17 bl[17] br[17] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_18 bl[18] br[18] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_19 bl[19] br[19] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_20 bl[20] br[20] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_21 bl[21] br[21] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_22 bl[22] br[22] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_23 bl[23] br[23] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_24 bl[24] br[24] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_25 bl[25] br[25] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_26 bl[26] br[26] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_27 bl[27] br[27] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_28 bl[28] br[28] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_29 bl[29] br[29] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_30 bl[30] br[30] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_31 bl[31] br[31] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_32 bl[32] br[32] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_33 bl[33] br[33] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_34 bl[34] br[34] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_35 bl[35] br[35] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_36 bl[36] br[36] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_37 bl[37] br[37] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_38 bl[38] br[38] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_39 bl[39] br[39] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_40 bl[40] br[40] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_41 bl[41] br[41] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_42 bl[42] br[42] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_43 bl[43] br[43] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_44 bl[44] br[44] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_45 bl[45] br[45] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_46 bl[46] br[46] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_47 bl[47] br[47] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_48 bl[48] br[48] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_49 bl[49] br[49] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_50 bl[50] br[50] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_51 bl[51] br[51] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_52 bl[52] br[52] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_53 bl[53] br[53] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_54 bl[54] br[54] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_55 bl[55] br[55] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_56 bl[56] br[56] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_57 bl[57] br[57] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_58 bl[58] br[58] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_59 bl[59] br[59] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_60 bl[60] br[60] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_61 bl[61] br[61] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_62 bl[62] br[62] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_63 bl[63] br[63] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_64 bl[64] br[64] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_65 bl[65] br[65] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_66 bl[66] br[66] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_67 bl[67] br[67] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_68 bl[68] br[68] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_69 bl[69] br[69] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_70 bl[70] br[70] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_71 bl[71] br[71] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_72 bl[72] br[72] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_73 bl[73] br[73] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_74 bl[74] br[74] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_75 bl[75] br[75] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_76 bl[76] br[76] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_77 bl[77] br[77] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_78 bl[78] br[78] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_79 bl[79] br[79] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_80 bl[80] br[80] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_81 bl[81] br[81] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_82 bl[82] br[82] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_83 bl[83] br[83] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_84 bl[84] br[84] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_85 bl[85] br[85] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_86 bl[86] br[86] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_87 bl[87] br[87] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_7_0 bl[0] br[0] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_1 bl[1] br[1] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_2 bl[2] br[2] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_3 bl[3] br[3] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_4 bl[4] br[4] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_5 bl[5] br[5] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_6 bl[6] br[6] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_7 bl[7] br[7] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_8 bl[8] br[8] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_9 bl[9] br[9] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_10 bl[10] br[10] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_11 bl[11] br[11] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_12 bl[12] br[12] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_13 bl[13] br[13] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_14 bl[14] br[14] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_15 bl[15] br[15] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_16 bl[16] br[16] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_17 bl[17] br[17] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_18 bl[18] br[18] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_19 bl[19] br[19] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_20 bl[20] br[20] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_21 bl[21] br[21] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_22 bl[22] br[22] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_23 bl[23] br[23] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_24 bl[24] br[24] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_25 bl[25] br[25] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_26 bl[26] br[26] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_27 bl[27] br[27] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_28 bl[28] br[28] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_29 bl[29] br[29] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_30 bl[30] br[30] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_31 bl[31] br[31] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_32 bl[32] br[32] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_33 bl[33] br[33] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_34 bl[34] br[34] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_35 bl[35] br[35] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_36 bl[36] br[36] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_37 bl[37] br[37] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_38 bl[38] br[38] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_39 bl[39] br[39] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_40 bl[40] br[40] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_41 bl[41] br[41] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_42 bl[42] br[42] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_43 bl[43] br[43] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_44 bl[44] br[44] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_45 bl[45] br[45] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_46 bl[46] br[46] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_47 bl[47] br[47] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_48 bl[48] br[48] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_49 bl[49] br[49] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_50 bl[50] br[50] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_51 bl[51] br[51] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_52 bl[52] br[52] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_53 bl[53] br[53] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_54 bl[54] br[54] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_55 bl[55] br[55] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_56 bl[56] br[56] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_57 bl[57] br[57] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_58 bl[58] br[58] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_59 bl[59] br[59] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_60 bl[60] br[60] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_61 bl[61] br[61] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_62 bl[62] br[62] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_63 bl[63] br[63] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_64 bl[64] br[64] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_65 bl[65] br[65] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_66 bl[66] br[66] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_67 bl[67] br[67] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_68 bl[68] br[68] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_69 bl[69] br[69] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_70 bl[70] br[70] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_71 bl[71] br[71] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_72 bl[72] br[72] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_73 bl[73] br[73] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_74 bl[74] br[74] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_75 bl[75] br[75] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_76 bl[76] br[76] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_77 bl[77] br[77] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_78 bl[78] br[78] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_79 bl[79] br[79] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_80 bl[80] br[80] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_81 bl[81] br[81] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_82 bl[82] br[82] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_83 bl[83] br[83] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_84 bl[84] br[84] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_85 bl[85] br[85] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_86 bl[86] br[86] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_87 bl[87] br[87] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_8_0 bl[0] br[0] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_1 bl[1] br[1] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_2 bl[2] br[2] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_3 bl[3] br[3] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_4 bl[4] br[4] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_5 bl[5] br[5] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_6 bl[6] br[6] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_7 bl[7] br[7] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_8 bl[8] br[8] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_9 bl[9] br[9] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_10 bl[10] br[10] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_11 bl[11] br[11] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_12 bl[12] br[12] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_13 bl[13] br[13] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_14 bl[14] br[14] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_15 bl[15] br[15] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_16 bl[16] br[16] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_17 bl[17] br[17] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_18 bl[18] br[18] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_19 bl[19] br[19] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_20 bl[20] br[20] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_21 bl[21] br[21] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_22 bl[22] br[22] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_23 bl[23] br[23] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_24 bl[24] br[24] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_25 bl[25] br[25] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_26 bl[26] br[26] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_27 bl[27] br[27] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_28 bl[28] br[28] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_29 bl[29] br[29] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_30 bl[30] br[30] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_31 bl[31] br[31] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_32 bl[32] br[32] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_33 bl[33] br[33] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_34 bl[34] br[34] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_35 bl[35] br[35] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_36 bl[36] br[36] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_37 bl[37] br[37] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_38 bl[38] br[38] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_39 bl[39] br[39] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_40 bl[40] br[40] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_41 bl[41] br[41] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_42 bl[42] br[42] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_43 bl[43] br[43] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_44 bl[44] br[44] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_45 bl[45] br[45] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_46 bl[46] br[46] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_47 bl[47] br[47] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_48 bl[48] br[48] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_49 bl[49] br[49] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_50 bl[50] br[50] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_51 bl[51] br[51] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_52 bl[52] br[52] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_53 bl[53] br[53] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_54 bl[54] br[54] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_55 bl[55] br[55] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_56 bl[56] br[56] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_57 bl[57] br[57] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_58 bl[58] br[58] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_59 bl[59] br[59] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_60 bl[60] br[60] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_61 bl[61] br[61] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_62 bl[62] br[62] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_63 bl[63] br[63] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_64 bl[64] br[64] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_65 bl[65] br[65] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_66 bl[66] br[66] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_67 bl[67] br[67] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_68 bl[68] br[68] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_69 bl[69] br[69] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_70 bl[70] br[70] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_71 bl[71] br[71] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_72 bl[72] br[72] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_73 bl[73] br[73] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_74 bl[74] br[74] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_75 bl[75] br[75] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_76 bl[76] br[76] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_77 bl[77] br[77] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_78 bl[78] br[78] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_79 bl[79] br[79] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_80 bl[80] br[80] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_81 bl[81] br[81] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_82 bl[82] br[82] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_83 bl[83] br[83] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_84 bl[84] br[84] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_85 bl[85] br[85] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_86 bl[86] br[86] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_87 bl[87] br[87] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_9_0 bl[0] br[0] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_1 bl[1] br[1] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_2 bl[2] br[2] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_3 bl[3] br[3] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_4 bl[4] br[4] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_5 bl[5] br[5] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_6 bl[6] br[6] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_7 bl[7] br[7] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_8 bl[8] br[8] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_9 bl[9] br[9] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_10 bl[10] br[10] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_11 bl[11] br[11] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_12 bl[12] br[12] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_13 bl[13] br[13] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_14 bl[14] br[14] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_15 bl[15] br[15] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_16 bl[16] br[16] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_17 bl[17] br[17] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_18 bl[18] br[18] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_19 bl[19] br[19] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_20 bl[20] br[20] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_21 bl[21] br[21] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_22 bl[22] br[22] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_23 bl[23] br[23] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_24 bl[24] br[24] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_25 bl[25] br[25] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_26 bl[26] br[26] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_27 bl[27] br[27] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_28 bl[28] br[28] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_29 bl[29] br[29] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_30 bl[30] br[30] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_31 bl[31] br[31] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_32 bl[32] br[32] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_33 bl[33] br[33] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_34 bl[34] br[34] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_35 bl[35] br[35] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_36 bl[36] br[36] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_37 bl[37] br[37] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_38 bl[38] br[38] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_39 bl[39] br[39] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_40 bl[40] br[40] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_41 bl[41] br[41] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_42 bl[42] br[42] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_43 bl[43] br[43] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_44 bl[44] br[44] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_45 bl[45] br[45] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_46 bl[46] br[46] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_47 bl[47] br[47] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_48 bl[48] br[48] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_49 bl[49] br[49] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_50 bl[50] br[50] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_51 bl[51] br[51] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_52 bl[52] br[52] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_53 bl[53] br[53] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_54 bl[54] br[54] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_55 bl[55] br[55] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_56 bl[56] br[56] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_57 bl[57] br[57] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_58 bl[58] br[58] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_59 bl[59] br[59] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_60 bl[60] br[60] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_61 bl[61] br[61] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_62 bl[62] br[62] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_63 bl[63] br[63] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_64 bl[64] br[64] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_65 bl[65] br[65] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_66 bl[66] br[66] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_67 bl[67] br[67] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_68 bl[68] br[68] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_69 bl[69] br[69] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_70 bl[70] br[70] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_71 bl[71] br[71] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_72 bl[72] br[72] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_73 bl[73] br[73] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_74 bl[74] br[74] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_75 bl[75] br[75] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_76 bl[76] br[76] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_77 bl[77] br[77] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_78 bl[78] br[78] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_79 bl[79] br[79] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_80 bl[80] br[80] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_81 bl[81] br[81] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_82 bl[82] br[82] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_83 bl[83] br[83] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_84 bl[84] br[84] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_85 bl[85] br[85] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_86 bl[86] br[86] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_87 bl[87] br[87] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_10_0 bl[0] br[0] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_1 bl[1] br[1] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_2 bl[2] br[2] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_3 bl[3] br[3] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_4 bl[4] br[4] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_5 bl[5] br[5] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_6 bl[6] br[6] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_7 bl[7] br[7] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_8 bl[8] br[8] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_9 bl[9] br[9] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_10 bl[10] br[10] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_11 bl[11] br[11] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_12 bl[12] br[12] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_13 bl[13] br[13] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_14 bl[14] br[14] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_15 bl[15] br[15] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_16 bl[16] br[16] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_17 bl[17] br[17] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_18 bl[18] br[18] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_19 bl[19] br[19] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_20 bl[20] br[20] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_21 bl[21] br[21] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_22 bl[22] br[22] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_23 bl[23] br[23] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_24 bl[24] br[24] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_25 bl[25] br[25] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_26 bl[26] br[26] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_27 bl[27] br[27] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_28 bl[28] br[28] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_29 bl[29] br[29] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_30 bl[30] br[30] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_31 bl[31] br[31] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_32 bl[32] br[32] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_33 bl[33] br[33] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_34 bl[34] br[34] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_35 bl[35] br[35] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_36 bl[36] br[36] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_37 bl[37] br[37] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_38 bl[38] br[38] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_39 bl[39] br[39] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_40 bl[40] br[40] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_41 bl[41] br[41] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_42 bl[42] br[42] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_43 bl[43] br[43] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_44 bl[44] br[44] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_45 bl[45] br[45] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_46 bl[46] br[46] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_47 bl[47] br[47] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_48 bl[48] br[48] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_49 bl[49] br[49] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_50 bl[50] br[50] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_51 bl[51] br[51] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_52 bl[52] br[52] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_53 bl[53] br[53] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_54 bl[54] br[54] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_55 bl[55] br[55] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_56 bl[56] br[56] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_57 bl[57] br[57] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_58 bl[58] br[58] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_59 bl[59] br[59] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_60 bl[60] br[60] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_61 bl[61] br[61] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_62 bl[62] br[62] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_63 bl[63] br[63] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_64 bl[64] br[64] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_65 bl[65] br[65] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_66 bl[66] br[66] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_67 bl[67] br[67] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_68 bl[68] br[68] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_69 bl[69] br[69] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_70 bl[70] br[70] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_71 bl[71] br[71] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_72 bl[72] br[72] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_73 bl[73] br[73] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_74 bl[74] br[74] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_75 bl[75] br[75] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_76 bl[76] br[76] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_77 bl[77] br[77] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_78 bl[78] br[78] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_79 bl[79] br[79] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_80 bl[80] br[80] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_81 bl[81] br[81] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_82 bl[82] br[82] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_83 bl[83] br[83] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_84 bl[84] br[84] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_85 bl[85] br[85] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_86 bl[86] br[86] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_87 bl[87] br[87] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_11_0 bl[0] br[0] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_1 bl[1] br[1] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_2 bl[2] br[2] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_3 bl[3] br[3] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_4 bl[4] br[4] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_5 bl[5] br[5] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_6 bl[6] br[6] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_7 bl[7] br[7] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_8 bl[8] br[8] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_9 bl[9] br[9] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_10 bl[10] br[10] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_11 bl[11] br[11] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_12 bl[12] br[12] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_13 bl[13] br[13] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_14 bl[14] br[14] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_15 bl[15] br[15] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_16 bl[16] br[16] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_17 bl[17] br[17] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_18 bl[18] br[18] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_19 bl[19] br[19] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_20 bl[20] br[20] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_21 bl[21] br[21] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_22 bl[22] br[22] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_23 bl[23] br[23] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_24 bl[24] br[24] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_25 bl[25] br[25] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_26 bl[26] br[26] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_27 bl[27] br[27] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_28 bl[28] br[28] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_29 bl[29] br[29] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_30 bl[30] br[30] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_31 bl[31] br[31] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_32 bl[32] br[32] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_33 bl[33] br[33] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_34 bl[34] br[34] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_35 bl[35] br[35] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_36 bl[36] br[36] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_37 bl[37] br[37] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_38 bl[38] br[38] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_39 bl[39] br[39] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_40 bl[40] br[40] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_41 bl[41] br[41] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_42 bl[42] br[42] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_43 bl[43] br[43] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_44 bl[44] br[44] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_45 bl[45] br[45] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_46 bl[46] br[46] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_47 bl[47] br[47] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_48 bl[48] br[48] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_49 bl[49] br[49] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_50 bl[50] br[50] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_51 bl[51] br[51] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_52 bl[52] br[52] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_53 bl[53] br[53] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_54 bl[54] br[54] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_55 bl[55] br[55] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_56 bl[56] br[56] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_57 bl[57] br[57] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_58 bl[58] br[58] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_59 bl[59] br[59] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_60 bl[60] br[60] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_61 bl[61] br[61] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_62 bl[62] br[62] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_63 bl[63] br[63] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_64 bl[64] br[64] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_65 bl[65] br[65] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_66 bl[66] br[66] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_67 bl[67] br[67] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_68 bl[68] br[68] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_69 bl[69] br[69] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_70 bl[70] br[70] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_71 bl[71] br[71] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_72 bl[72] br[72] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_73 bl[73] br[73] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_74 bl[74] br[74] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_75 bl[75] br[75] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_76 bl[76] br[76] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_77 bl[77] br[77] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_78 bl[78] br[78] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_79 bl[79] br[79] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_80 bl[80] br[80] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_81 bl[81] br[81] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_82 bl[82] br[82] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_83 bl[83] br[83] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_84 bl[84] br[84] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_85 bl[85] br[85] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_86 bl[86] br[86] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_87 bl[87] br[87] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_12_0 bl[0] br[0] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_1 bl[1] br[1] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_2 bl[2] br[2] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_3 bl[3] br[3] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_4 bl[4] br[4] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_5 bl[5] br[5] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_6 bl[6] br[6] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_7 bl[7] br[7] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_8 bl[8] br[8] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_9 bl[9] br[9] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_10 bl[10] br[10] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_11 bl[11] br[11] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_12 bl[12] br[12] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_13 bl[13] br[13] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_14 bl[14] br[14] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_15 bl[15] br[15] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_16 bl[16] br[16] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_17 bl[17] br[17] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_18 bl[18] br[18] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_19 bl[19] br[19] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_20 bl[20] br[20] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_21 bl[21] br[21] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_22 bl[22] br[22] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_23 bl[23] br[23] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_24 bl[24] br[24] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_25 bl[25] br[25] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_26 bl[26] br[26] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_27 bl[27] br[27] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_28 bl[28] br[28] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_29 bl[29] br[29] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_30 bl[30] br[30] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_31 bl[31] br[31] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_32 bl[32] br[32] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_33 bl[33] br[33] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_34 bl[34] br[34] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_35 bl[35] br[35] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_36 bl[36] br[36] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_37 bl[37] br[37] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_38 bl[38] br[38] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_39 bl[39] br[39] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_40 bl[40] br[40] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_41 bl[41] br[41] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_42 bl[42] br[42] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_43 bl[43] br[43] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_44 bl[44] br[44] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_45 bl[45] br[45] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_46 bl[46] br[46] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_47 bl[47] br[47] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_48 bl[48] br[48] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_49 bl[49] br[49] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_50 bl[50] br[50] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_51 bl[51] br[51] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_52 bl[52] br[52] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_53 bl[53] br[53] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_54 bl[54] br[54] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_55 bl[55] br[55] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_56 bl[56] br[56] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_57 bl[57] br[57] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_58 bl[58] br[58] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_59 bl[59] br[59] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_60 bl[60] br[60] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_61 bl[61] br[61] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_62 bl[62] br[62] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_63 bl[63] br[63] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_64 bl[64] br[64] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_65 bl[65] br[65] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_66 bl[66] br[66] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_67 bl[67] br[67] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_68 bl[68] br[68] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_69 bl[69] br[69] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_70 bl[70] br[70] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_71 bl[71] br[71] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_72 bl[72] br[72] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_73 bl[73] br[73] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_74 bl[74] br[74] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_75 bl[75] br[75] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_76 bl[76] br[76] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_77 bl[77] br[77] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_78 bl[78] br[78] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_79 bl[79] br[79] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_80 bl[80] br[80] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_81 bl[81] br[81] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_82 bl[82] br[82] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_83 bl[83] br[83] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_84 bl[84] br[84] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_85 bl[85] br[85] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_86 bl[86] br[86] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_87 bl[87] br[87] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_13_0 bl[0] br[0] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_1 bl[1] br[1] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_2 bl[2] br[2] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_3 bl[3] br[3] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_4 bl[4] br[4] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_5 bl[5] br[5] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_6 bl[6] br[6] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_7 bl[7] br[7] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_8 bl[8] br[8] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_9 bl[9] br[9] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_10 bl[10] br[10] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_11 bl[11] br[11] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_12 bl[12] br[12] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_13 bl[13] br[13] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_14 bl[14] br[14] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_15 bl[15] br[15] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_16 bl[16] br[16] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_17 bl[17] br[17] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_18 bl[18] br[18] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_19 bl[19] br[19] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_20 bl[20] br[20] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_21 bl[21] br[21] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_22 bl[22] br[22] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_23 bl[23] br[23] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_24 bl[24] br[24] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_25 bl[25] br[25] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_26 bl[26] br[26] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_27 bl[27] br[27] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_28 bl[28] br[28] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_29 bl[29] br[29] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_30 bl[30] br[30] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_31 bl[31] br[31] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_32 bl[32] br[32] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_33 bl[33] br[33] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_34 bl[34] br[34] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_35 bl[35] br[35] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_36 bl[36] br[36] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_37 bl[37] br[37] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_38 bl[38] br[38] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_39 bl[39] br[39] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_40 bl[40] br[40] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_41 bl[41] br[41] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_42 bl[42] br[42] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_43 bl[43] br[43] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_44 bl[44] br[44] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_45 bl[45] br[45] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_46 bl[46] br[46] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_47 bl[47] br[47] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_48 bl[48] br[48] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_49 bl[49] br[49] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_50 bl[50] br[50] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_51 bl[51] br[51] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_52 bl[52] br[52] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_53 bl[53] br[53] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_54 bl[54] br[54] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_55 bl[55] br[55] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_56 bl[56] br[56] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_57 bl[57] br[57] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_58 bl[58] br[58] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_59 bl[59] br[59] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_60 bl[60] br[60] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_61 bl[61] br[61] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_62 bl[62] br[62] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_63 bl[63] br[63] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_64 bl[64] br[64] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_65 bl[65] br[65] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_66 bl[66] br[66] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_67 bl[67] br[67] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_68 bl[68] br[68] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_69 bl[69] br[69] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_70 bl[70] br[70] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_71 bl[71] br[71] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_72 bl[72] br[72] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_73 bl[73] br[73] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_74 bl[74] br[74] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_75 bl[75] br[75] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_76 bl[76] br[76] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_77 bl[77] br[77] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_78 bl[78] br[78] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_79 bl[79] br[79] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_80 bl[80] br[80] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_81 bl[81] br[81] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_82 bl[82] br[82] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_83 bl[83] br[83] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_84 bl[84] br[84] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_85 bl[85] br[85] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_86 bl[86] br[86] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_87 bl[87] br[87] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_14_0 bl[0] br[0] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_1 bl[1] br[1] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_2 bl[2] br[2] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_3 bl[3] br[3] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_4 bl[4] br[4] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_5 bl[5] br[5] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_6 bl[6] br[6] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_7 bl[7] br[7] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_8 bl[8] br[8] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_9 bl[9] br[9] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_10 bl[10] br[10] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_11 bl[11] br[11] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_12 bl[12] br[12] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_13 bl[13] br[13] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_14 bl[14] br[14] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_15 bl[15] br[15] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_16 bl[16] br[16] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_17 bl[17] br[17] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_18 bl[18] br[18] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_19 bl[19] br[19] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_20 bl[20] br[20] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_21 bl[21] br[21] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_22 bl[22] br[22] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_23 bl[23] br[23] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_24 bl[24] br[24] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_25 bl[25] br[25] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_26 bl[26] br[26] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_27 bl[27] br[27] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_28 bl[28] br[28] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_29 bl[29] br[29] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_30 bl[30] br[30] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_31 bl[31] br[31] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_32 bl[32] br[32] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_33 bl[33] br[33] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_34 bl[34] br[34] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_35 bl[35] br[35] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_36 bl[36] br[36] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_37 bl[37] br[37] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_38 bl[38] br[38] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_39 bl[39] br[39] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_40 bl[40] br[40] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_41 bl[41] br[41] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_42 bl[42] br[42] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_43 bl[43] br[43] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_44 bl[44] br[44] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_45 bl[45] br[45] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_46 bl[46] br[46] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_47 bl[47] br[47] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_48 bl[48] br[48] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_49 bl[49] br[49] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_50 bl[50] br[50] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_51 bl[51] br[51] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_52 bl[52] br[52] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_53 bl[53] br[53] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_54 bl[54] br[54] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_55 bl[55] br[55] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_56 bl[56] br[56] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_57 bl[57] br[57] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_58 bl[58] br[58] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_59 bl[59] br[59] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_60 bl[60] br[60] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_61 bl[61] br[61] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_62 bl[62] br[62] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_63 bl[63] br[63] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_64 bl[64] br[64] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_65 bl[65] br[65] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_66 bl[66] br[66] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_67 bl[67] br[67] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_68 bl[68] br[68] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_69 bl[69] br[69] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_70 bl[70] br[70] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_71 bl[71] br[71] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_72 bl[72] br[72] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_73 bl[73] br[73] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_74 bl[74] br[74] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_75 bl[75] br[75] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_76 bl[76] br[76] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_77 bl[77] br[77] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_78 bl[78] br[78] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_79 bl[79] br[79] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_80 bl[80] br[80] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_81 bl[81] br[81] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_82 bl[82] br[82] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_83 bl[83] br[83] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_84 bl[84] br[84] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_85 bl[85] br[85] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_86 bl[86] br[86] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_87 bl[87] br[87] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_15_0 bl[0] br[0] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_1 bl[1] br[1] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_2 bl[2] br[2] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_3 bl[3] br[3] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_4 bl[4] br[4] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_5 bl[5] br[5] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_6 bl[6] br[6] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_7 bl[7] br[7] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_8 bl[8] br[8] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_9 bl[9] br[9] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_10 bl[10] br[10] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_11 bl[11] br[11] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_12 bl[12] br[12] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_13 bl[13] br[13] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_14 bl[14] br[14] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_15 bl[15] br[15] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_16 bl[16] br[16] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_17 bl[17] br[17] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_18 bl[18] br[18] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_19 bl[19] br[19] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_20 bl[20] br[20] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_21 bl[21] br[21] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_22 bl[22] br[22] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_23 bl[23] br[23] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_24 bl[24] br[24] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_25 bl[25] br[25] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_26 bl[26] br[26] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_27 bl[27] br[27] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_28 bl[28] br[28] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_29 bl[29] br[29] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_30 bl[30] br[30] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_31 bl[31] br[31] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_32 bl[32] br[32] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_33 bl[33] br[33] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_34 bl[34] br[34] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_35 bl[35] br[35] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_36 bl[36] br[36] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_37 bl[37] br[37] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_38 bl[38] br[38] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_39 bl[39] br[39] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_40 bl[40] br[40] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_41 bl[41] br[41] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_42 bl[42] br[42] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_43 bl[43] br[43] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_44 bl[44] br[44] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_45 bl[45] br[45] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_46 bl[46] br[46] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_47 bl[47] br[47] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_48 bl[48] br[48] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_49 bl[49] br[49] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_50 bl[50] br[50] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_51 bl[51] br[51] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_52 bl[52] br[52] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_53 bl[53] br[53] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_54 bl[54] br[54] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_55 bl[55] br[55] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_56 bl[56] br[56] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_57 bl[57] br[57] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_58 bl[58] br[58] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_59 bl[59] br[59] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_60 bl[60] br[60] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_61 bl[61] br[61] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_62 bl[62] br[62] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_63 bl[63] br[63] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_64 bl[64] br[64] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_65 bl[65] br[65] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_66 bl[66] br[66] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_67 bl[67] br[67] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_68 bl[68] br[68] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_69 bl[69] br[69] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_70 bl[70] br[70] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_71 bl[71] br[71] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_72 bl[72] br[72] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_73 bl[73] br[73] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_74 bl[74] br[74] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_75 bl[75] br[75] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_76 bl[76] br[76] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_77 bl[77] br[77] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_78 bl[78] br[78] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_79 bl[79] br[79] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_80 bl[80] br[80] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_81 bl[81] br[81] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_82 bl[82] br[82] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_83 bl[83] br[83] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_84 bl[84] br[84] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_85 bl[85] br[85] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_86 bl[86] br[86] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_87 bl[87] br[87] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_0 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_0 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_1 dummy_bl dummy_br vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_1 vdd vdd vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_2 dummy_bl dummy_br vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_2 vdd vdd vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_3 dummy_bl dummy_br vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_3 vdd vdd vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_4 dummy_bl dummy_br vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_4 vdd vdd vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_5 dummy_bl dummy_br vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_5 vdd vdd vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_6 dummy_bl dummy_br vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_6 vdd vdd vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_7 dummy_bl dummy_br vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_7 vdd vdd vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_8 dummy_bl dummy_br vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_8 vdd vdd vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_9 dummy_bl dummy_br vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_9 vdd vdd vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_10 dummy_bl dummy_br vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_10 vdd vdd vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_11 dummy_bl dummy_br vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_11 vdd vdd vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_12 dummy_bl dummy_br vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_12 vdd vdd vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_13 dummy_bl dummy_br vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_13 vdd vdd vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_14 dummy_bl dummy_br vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_14 vdd vdd vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_15 dummy_bl dummy_br vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_15 vdd vdd vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_16 dummy_bl dummy_br vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_16 vdd vdd vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_17 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_17 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_64 bl[64] br[64] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_64 bl[64] br[64] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_65 bl[65] br[65] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_65 bl[65] br[65] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_66 bl[66] br[66] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_66 bl[66] br[66] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_67 bl[67] br[67] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_67 bl[67] br[67] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_68 bl[68] br[68] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_68 bl[68] br[68] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_69 bl[69] br[69] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_69 bl[69] br[69] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_70 bl[70] br[70] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_70 bl[70] br[70] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_71 bl[71] br[71] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_71 bl[71] br[71] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_72 bl[72] br[72] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_72 bl[72] br[72] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_73 bl[73] br[73] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_73 bl[73] br[73] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_74 bl[74] br[74] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_74 bl[74] br[74] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_75 bl[75] br[75] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_75 bl[75] br[75] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_76 bl[76] br[76] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_76 bl[76] br[76] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_77 bl[77] br[77] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_77 bl[77] br[77] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_78 bl[78] br[78] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_78 bl[78] br[78] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_79 bl[79] br[79] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_79 bl[79] br[79] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_80 bl[80] br[80] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_80 bl[80] br[80] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_81 bl[81] br[81] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_81 bl[81] br[81] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_82 bl[82] br[82] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_82 bl[82] br[82] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_83 bl[83] br[83] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_83 bl[83] br[83] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_84 bl[84] br[84] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_84 bl[84] br[84] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_85 bl[85] br[85] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_85 bl[85] br[85] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_86 bl[86] br[86] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_86 bl[86] br[86] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_87 bl[87] br[87] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_87 bl[87] br[87] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xcolend_top_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xcolend_bot_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xhstrap_0_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_65 br[64] vdd vss bl[64] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_65 br[64] vdd vss bl[64] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_66 br[65] vdd vss bl[65] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_66 br[65] vdd vss bl[65] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_67 br[66] vdd vss bl[66] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_67 br[66] vdd vss bl[66] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_68 br[67] vdd vss bl[67] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_68 br[67] vdd vss bl[67] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_69 br[68] vdd vss bl[68] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_69 br[68] vdd vss bl[68] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_70 br[69] vdd vss bl[69] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_70 br[69] vdd vss bl[69] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_71 br[70] vdd vss bl[70] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_71 br[70] vdd vss bl[70] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_72 br[71] vdd vss bl[71] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_72 br[71] vdd vss bl[71] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_73 br[72] vdd vss bl[72] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_73 br[72] vdd vss bl[72] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_74 br[73] vdd vss bl[73] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_74 br[73] vdd vss bl[73] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_75 br[74] vdd vss bl[74] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_75 br[74] vdd vss bl[74] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_76 br[75] vdd vss bl[75] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_76 br[75] vdd vss bl[75] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_77 br[76] vdd vss bl[76] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_77 br[76] vdd vss bl[76] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_78 br[77] vdd vss bl[77] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_78 br[77] vdd vss bl[77] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_79 br[78] vdd vss bl[78] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_79 br[78] vdd vss bl[78] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_80 br[79] vdd vss bl[79] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_80 br[79] vdd vss bl[79] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_81 br[80] vdd vss bl[80] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_81 br[80] vdd vss bl[80] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_82 br[81] vdd vss bl[81] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_82 br[81] vdd vss bl[81] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_83 br[82] vdd vss bl[82] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_83 br[82] vdd vss bl[82] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_84 br[83] vdd vss bl[83] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_84 br[83] vdd vss bl[83] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_85 br[84] vdd vss bl[84] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_85 br[84] vdd vss bl[84] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_86 br[85] vdd vss bl[85] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_86 br[85] vdd vss bl[85] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_87 br[86] vdd vss bl[86] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_87 br[86] vdd vss bl[86] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_88 br[87] vdd vss bl[87] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_88 br[87] vdd vss bl[87] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_89 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xcolend_bot_89 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xhstrap_0_89 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_89 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_89 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_89 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_89 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhoriz_wlstrap_0_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper

.ENDS sp_cell_array

.SUBCKT sram_sp_rowtapend_replica VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_rowtapend_replica

.SUBCKT sram_sp_rowtapend_replica_wrapper VSS VNB

  X0 VSS VNB sram_sp_rowtapend_replica

.ENDS sram_sp_rowtapend_replica_wrapper

.SUBCKT replica_cell_array vdd vss rbl rbr rwl

  Xcell_0_0 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_0_1 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_1_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_1_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcolend_0_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_0_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xrowtapend_0_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_0_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_0_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_0_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_1_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_1_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_1_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper

.ENDS replica_cell_array

.SUBCKT precharge vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w800_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w800_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w500_l150_m1_nf1_id1

.ENDS precharge

.SUBCKT replica_column_mos vdd vss bl

  Xunit0 vdd vss bl column_mos

.ENDS replica_column_mos

.SUBCKT sram22_inner vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] wmask din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21]

  Xaddr_gate vdd vss addr_gated[0] addr_gated[1] addr_gated[2] addr_gated[3] addr_b_gated[0] addr_b_gated[1] addr_b_gated[2] addr_b_gated[3] addr_gate_y_b_noconn[0] addr_gate_y_b_noconn[1] addr_gate_y_b_noconn[2] addr_gate_y_b_noconn[3] addr_gate_y_b_noconn[4] addr_gate_y_b_noconn[5] addr_gate_y_b_noconn[6] addr_gate_y_b_noconn[7] wl_en addr_in[2] addr_in[3] addr_in[4] addr_in[5] addr_in_b[2] addr_in_b[3] addr_in_b[4] addr_in_b[5] decoder_stage
  Xdecoder vdd vss wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl_b[0] wl_b[1] wl_b[2] wl_b[3] wl_b[4] wl_b[5] wl_b[6] wl_b[7] wl_b[8] wl_b[9] wl_b[10] wl_b[11] wl_b[12] wl_b[13] wl_b[14] wl_b[15] addr_b_gated[0] addr_gated[0] addr_b_gated[1] addr_gated[1] addr_b_gated[2] addr_gated[2] addr_b_gated[3] addr_gated[3] decoder
  Xcolumn_decoder vdd vss col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] addr_in_b[0] addr_in[0] addr_in_b[1] addr_in[1] decoder_1
  Xcontrol_logic clk ce_in we_in rstb rbl sense_en0 pc_b0 rwl wl_en0 write_driver_en0 vdd vss control_logic_replica_v2
  Xpc_b_buffer vdd vss pc_b pc pc_b0 decoder_stage_1
  Xwlen_buffer vdd vss wl_en wl_en_b wl_en0 decoder_stage_2
  Xwrite_driver_en_buffer vdd vss write_driver_en write_driver_en_b write_driver_en0 decoder_stage_3
  Xsense_en_buffer vdd vss sense_en sense_en_b sense_en0 decoder_stage_4
  Xaddr_we_ce_dffs vdd vss clk rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] we ce addr_in[0] addr_in[1] addr_in[2] addr_in[3] addr_in[4] addr_in[5] we_in ce_in addr_in_b[0] addr_in_b[1] addr_in_b[2] addr_in_b[3] addr_in_b[4] addr_in_b[5] we_in_b ce_in_b dff_array_8
  Xbitcell_array vdd vss vdd vdd bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] sp_cell_array
  Xreplica_bitcell_array vdd vss rbl rbr rwl replica_cell_array
  Xcol_circuitry clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] pc_b col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] write_driver_en wmask din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] col_peripherals
  Xreplica_precharge_0 vdd rbl rbr pc_b0 precharge
  Xreplica_precharge_1 vdd rbl rbr pc_b0 precharge
  Xreplica_mos vdd vss rbl replica_column_mos

.ENDS sram22_inner

.SUBCKT sram22_64x22m4w22 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] wmask din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21]

  X0 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] wmask din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] sram22_inner

.ENDS sram22_64x22m4w22

