VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_2048x32m8w8
    CLASS BLOCK  ;
    FOREIGN sram22_2048x32m8w8   ;
    SIZE 674.480 BY 781.920 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 314.950 0.000 315.090 0.140 ;
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 325.850 0.000 325.990 0.140 ;
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.750 0.000 336.890 0.140 ;
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 347.650 0.000 347.790 0.140 ;
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 358.550 0.000 358.690 0.140 ;
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 369.450 0.000 369.590 0.140 ;
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 380.350 0.000 380.490 0.140 ;
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 391.250 0.000 391.390 0.140 ;
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 402.150 0.000 402.290 0.140 ;
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 413.050 0.000 413.190 0.140 ;
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 423.950 0.000 424.090 0.140 ;
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 434.850 0.000 434.990 0.140 ;
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 445.750 0.000 445.890 0.140 ;
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 456.650 0.000 456.790 0.140 ;
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 467.550 0.000 467.690 0.140 ;
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 478.450 0.000 478.590 0.140 ;
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 489.350 0.000 489.490 0.140 ;
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 500.250 0.000 500.390 0.140 ;
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 511.150 0.000 511.290 0.140 ;
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 522.050 0.000 522.190 0.140 ;
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 532.950 0.000 533.090 0.140 ;
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 543.850 0.000 543.990 0.140 ;
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 554.750 0.000 554.890 0.140 ;
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 565.650 0.000 565.790 0.140 ;
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 576.550 0.000 576.690 0.140 ;
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 587.450 0.000 587.590 0.140 ;
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 598.350 0.000 598.490 0.140 ;
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 609.250 0.000 609.390 0.140 ;
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 620.150 0.000 620.290 0.140 ;
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 631.050 0.000 631.190 0.140 ;
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 641.950 0.000 642.090 0.140 ;
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 652.850 0.000 652.990 0.140 ;
        END 
    END dout[31] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 314.530 0.000 314.670 0.140 ;
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 325.430 0.000 325.570 0.140 ;
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.330 0.000 336.470 0.140 ;
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 347.230 0.000 347.370 0.140 ;
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 358.130 0.000 358.270 0.140 ;
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 369.030 0.000 369.170 0.140 ;
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 379.930 0.000 380.070 0.140 ;
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 390.830 0.000 390.970 0.140 ;
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 401.730 0.000 401.870 0.140 ;
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 412.630 0.000 412.770 0.140 ;
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 423.530 0.000 423.670 0.140 ;
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 434.430 0.000 434.570 0.140 ;
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 445.330 0.000 445.470 0.140 ;
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 456.230 0.000 456.370 0.140 ;
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 467.130 0.000 467.270 0.140 ;
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 478.030 0.000 478.170 0.140 ;
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 488.930 0.000 489.070 0.140 ;
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 499.830 0.000 499.970 0.140 ;
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 510.730 0.000 510.870 0.140 ;
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 521.630 0.000 521.770 0.140 ;
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 532.530 0.000 532.670 0.140 ;
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 543.430 0.000 543.570 0.140 ;
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 554.330 0.000 554.470 0.140 ;
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 565.230 0.000 565.370 0.140 ;
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 576.130 0.000 576.270 0.140 ;
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 587.030 0.000 587.170 0.140 ;
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 597.930 0.000 598.070 0.140 ;
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 608.830 0.000 608.970 0.140 ;
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 619.730 0.000 619.870 0.140 ;
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 630.630 0.000 630.770 0.140 ;
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 641.530 0.000 641.670 0.140 ;
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 6.402600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 652.430 0.000 652.570 0.140 ;
        END 
    END din[31] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.213000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 314.180 0.000 314.320 0.140 ;
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.213000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 401.380 0.000 401.520 0.140 ;
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.213000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 488.580 0.000 488.720 0.140 ;
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.213000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 575.780 0.000 575.920 0.140 ;
        END 
    END wmask[3] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 256.160 0.000 256.480 0.320 ;
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 250.040 0.000 250.360 0.320 ;
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 243.920 0.000 244.240 0.320 ;
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 237.800 0.000 238.120 0.320 ;
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 231.680 0.000 232.000 0.320 ;
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 225.560 0.000 225.880 0.320 ;
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 219.440 0.000 219.760 0.320 ;
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 213.320 0.000 213.640 0.320 ;
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 207.880 0.000 208.200 0.320 ;
        END 
    END addr[8] 
    PIN addr[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 201.760 0.000 202.080 0.320 ;
        END 
    END addr[9] 
    PIN addr[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 195.640 0.000 195.960 0.320 ;
        END 
    END addr[10] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 268.400 0.000 268.720 0.320 ;
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 262.280 0.000 262.600 0.320 ;
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 23.157000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 271.800 0.000 272.120 0.320 ;
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 27.063000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 272.480 0.000 272.800 0.320 ;
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 314.280 6.240 ;
                RECT 316.000 5.920 325.160 6.240 ;
                RECT 326.880 5.920 336.040 6.240 ;
                RECT 337.760 5.920 346.920 6.240 ;
                RECT 348.640 5.920 357.800 6.240 ;
                RECT 359.520 5.920 368.680 6.240 ;
                RECT 370.400 5.920 379.560 6.240 ;
                RECT 381.280 5.920 390.440 6.240 ;
                RECT 392.160 5.920 401.320 6.240 ;
                RECT 403.040 5.920 412.200 6.240 ;
                RECT 413.920 5.920 423.080 6.240 ;
                RECT 424.800 5.920 433.960 6.240 ;
                RECT 435.680 5.920 444.840 6.240 ;
                RECT 446.560 5.920 455.720 6.240 ;
                RECT 457.440 5.920 466.600 6.240 ;
                RECT 468.320 5.920 477.480 6.240 ;
                RECT 479.200 5.920 488.360 6.240 ;
                RECT 490.080 5.920 499.240 6.240 ;
                RECT 500.960 5.920 510.120 6.240 ;
                RECT 511.840 5.920 521.680 6.240 ;
                RECT 522.720 5.920 532.560 6.240 ;
                RECT 533.600 5.920 543.440 6.240 ;
                RECT 544.480 5.920 554.320 6.240 ;
                RECT 555.360 5.920 565.200 6.240 ;
                RECT 566.240 5.920 576.080 6.240 ;
                RECT 577.120 5.920 586.960 6.240 ;
                RECT 588.000 5.920 597.840 6.240 ;
                RECT 598.880 5.920 608.720 6.240 ;
                RECT 609.760 5.920 619.600 6.240 ;
                RECT 621.320 5.920 630.480 6.240 ;
                RECT 632.200 5.920 641.360 6.240 ;
                RECT 643.080 5.920 652.240 6.240 ;
                RECT 653.960 5.920 674.320 6.240 ;
                RECT 0.160 7.280 674.320 7.600 ;
                RECT 0.160 8.640 674.320 8.960 ;
                RECT 0.160 10.000 271.440 10.320 ;
                RECT 307.840 10.000 674.320 10.320 ;
                RECT 0.160 11.360 674.320 11.680 ;
                RECT 0.160 12.720 674.320 13.040 ;
                RECT 0.160 14.080 191.200 14.400 ;
                RECT 273.160 14.080 674.320 14.400 ;
                RECT 0.160 15.440 674.320 15.760 ;
                RECT 0.160 16.800 674.320 17.120 ;
                RECT 0.160 18.160 191.200 18.480 ;
                RECT 272.480 18.160 674.320 18.480 ;
                RECT 0.160 19.520 674.320 19.840 ;
                RECT 0.160 20.880 674.320 21.200 ;
                RECT 0.160 22.240 674.320 22.560 ;
                RECT 0.160 23.600 674.320 23.920 ;
                RECT 0.160 24.960 674.320 25.280 ;
                RECT 0.160 26.320 674.320 26.640 ;
                RECT 0.160 27.680 674.320 28.000 ;
                RECT 0.160 29.040 301.360 29.360 ;
                RECT 664.840 29.040 674.320 29.360 ;
                RECT 0.160 30.400 301.360 30.720 ;
                RECT 664.840 30.400 674.320 30.720 ;
                RECT 0.160 31.760 301.360 32.080 ;
                RECT 664.840 31.760 674.320 32.080 ;
                RECT 0.160 33.120 301.360 33.440 ;
                RECT 664.840 33.120 674.320 33.440 ;
                RECT 0.160 34.480 301.360 34.800 ;
                RECT 664.840 34.480 674.320 34.800 ;
                RECT 0.160 35.840 301.360 36.160 ;
                RECT 664.840 35.840 674.320 36.160 ;
                RECT 0.160 37.200 159.240 37.520 ;
                RECT 243.920 37.200 301.360 37.520 ;
                RECT 664.840 37.200 674.320 37.520 ;
                RECT 0.160 38.560 157.880 38.880 ;
                RECT 250.040 38.560 301.360 38.880 ;
                RECT 664.840 38.560 674.320 38.880 ;
                RECT 0.160 39.920 156.520 40.240 ;
                RECT 256.160 39.920 301.360 40.240 ;
                RECT 664.840 39.920 674.320 40.240 ;
                RECT 0.160 41.280 136.800 41.600 ;
                RECT 273.160 41.280 301.360 41.600 ;
                RECT 664.840 41.280 674.320 41.600 ;
                RECT 0.160 42.640 136.120 42.960 ;
                RECT 269.080 42.640 301.360 42.960 ;
                RECT 664.840 42.640 674.320 42.960 ;
                RECT 0.160 44.000 301.360 44.320 ;
                RECT 664.840 44.000 674.320 44.320 ;
                RECT 0.160 45.360 301.360 45.680 ;
                RECT 664.840 45.360 674.320 45.680 ;
                RECT 0.160 46.720 263.280 47.040 ;
                RECT 270.440 46.720 300.680 47.040 ;
                RECT 664.840 46.720 674.320 47.040 ;
                RECT 0.160 48.080 263.280 48.400 ;
                RECT 664.840 48.080 674.320 48.400 ;
                RECT 0.160 49.440 263.280 49.760 ;
                RECT 270.440 49.440 301.360 49.760 ;
                RECT 664.840 49.440 674.320 49.760 ;
                RECT 0.160 50.800 301.360 51.120 ;
                RECT 664.840 50.800 674.320 51.120 ;
                RECT 0.160 52.160 301.360 52.480 ;
                RECT 664.840 52.160 674.320 52.480 ;
                RECT 0.160 53.520 301.360 53.840 ;
                RECT 664.840 53.520 674.320 53.840 ;
                RECT 0.160 54.880 301.360 55.200 ;
                RECT 664.840 54.880 674.320 55.200 ;
                RECT 0.160 56.240 156.520 56.560 ;
                RECT 164.360 56.240 171.480 56.560 ;
                RECT 269.080 56.240 301.360 56.560 ;
                RECT 664.840 56.240 674.320 56.560 ;
                RECT 0.160 57.600 157.880 57.920 ;
                RECT 163.680 57.600 171.480 57.920 ;
                RECT 282.680 57.600 301.360 57.920 ;
                RECT 664.840 57.600 674.320 57.920 ;
                RECT 0.160 58.960 159.240 59.280 ;
                RECT 163.000 58.960 171.480 59.280 ;
                RECT 282.680 58.960 301.360 59.280 ;
                RECT 664.840 58.960 674.320 59.280 ;
                RECT 0.160 60.320 171.480 60.640 ;
                RECT 281.320 60.320 301.360 60.640 ;
                RECT 664.840 60.320 674.320 60.640 ;
                RECT 0.160 61.680 171.480 62.000 ;
                RECT 282.680 61.680 301.360 62.000 ;
                RECT 664.840 61.680 674.320 62.000 ;
                RECT 0.160 63.040 171.480 63.360 ;
                RECT 282.680 63.040 301.360 63.360 ;
                RECT 664.840 63.040 674.320 63.360 ;
                RECT 0.160 64.400 171.480 64.720 ;
                RECT 281.320 64.400 301.360 64.720 ;
                RECT 664.840 64.400 674.320 64.720 ;
                RECT 0.160 65.760 171.480 66.080 ;
                RECT 282.680 65.760 301.360 66.080 ;
                RECT 664.840 65.760 674.320 66.080 ;
                RECT 0.160 67.120 171.480 67.440 ;
                RECT 281.320 67.120 301.360 67.440 ;
                RECT 664.840 67.120 674.320 67.440 ;
                RECT 0.160 68.480 171.480 68.800 ;
                RECT 285.400 68.480 301.360 68.800 ;
                RECT 664.840 68.480 674.320 68.800 ;
                RECT 0.160 69.840 171.480 70.160 ;
                RECT 285.400 69.840 301.360 70.160 ;
                RECT 664.840 69.840 674.320 70.160 ;
                RECT 0.160 71.200 171.480 71.520 ;
                RECT 269.080 71.200 301.360 71.520 ;
                RECT 664.840 71.200 674.320 71.520 ;
                RECT 0.160 72.560 171.480 72.880 ;
                RECT 284.040 72.560 301.360 72.880 ;
                RECT 664.840 72.560 674.320 72.880 ;
                RECT 0.160 73.920 171.480 74.240 ;
                RECT 269.080 73.920 301.360 74.240 ;
                RECT 664.840 73.920 674.320 74.240 ;
                RECT 0.160 75.280 171.480 75.600 ;
                RECT 285.400 75.280 301.360 75.600 ;
                RECT 664.840 75.280 674.320 75.600 ;
                RECT 0.160 76.640 171.480 76.960 ;
                RECT 285.400 76.640 301.360 76.960 ;
                RECT 664.840 76.640 674.320 76.960 ;
                RECT 0.160 78.000 171.480 78.320 ;
                RECT 288.120 78.000 301.360 78.320 ;
                RECT 664.840 78.000 674.320 78.320 ;
                RECT 0.160 79.360 171.480 79.680 ;
                RECT 286.760 79.360 301.360 79.680 ;
                RECT 664.840 79.360 674.320 79.680 ;
                RECT 0.160 80.720 171.480 81.040 ;
                RECT 288.120 80.720 301.360 81.040 ;
                RECT 664.840 80.720 674.320 81.040 ;
                RECT 0.160 82.080 171.480 82.400 ;
                RECT 269.080 82.080 301.360 82.400 ;
                RECT 664.840 82.080 674.320 82.400 ;
                RECT 0.160 83.440 171.480 83.760 ;
                RECT 288.120 83.440 301.360 83.760 ;
                RECT 664.840 83.440 674.320 83.760 ;
                RECT 0.160 84.800 171.480 85.120 ;
                RECT 288.120 84.800 301.360 85.120 ;
                RECT 664.840 84.800 674.320 85.120 ;
                RECT 0.160 86.160 171.480 86.480 ;
                RECT 286.760 86.160 301.360 86.480 ;
                RECT 664.840 86.160 674.320 86.480 ;
                RECT 0.160 87.520 171.480 87.840 ;
                RECT 288.120 87.520 301.360 87.840 ;
                RECT 664.840 87.520 674.320 87.840 ;
                RECT 0.160 88.880 171.480 89.200 ;
                RECT 290.840 88.880 301.360 89.200 ;
                RECT 664.840 88.880 674.320 89.200 ;
                RECT 0.160 90.240 171.480 90.560 ;
                RECT 269.080 90.240 301.360 90.560 ;
                RECT 664.840 90.240 674.320 90.560 ;
                RECT 0.160 91.600 171.480 91.920 ;
                RECT 290.840 91.600 301.360 91.920 ;
                RECT 664.840 91.600 674.320 91.920 ;
                RECT 0.160 92.960 171.480 93.280 ;
                RECT 289.480 92.960 301.360 93.280 ;
                RECT 664.840 92.960 674.320 93.280 ;
                RECT 0.160 94.320 171.480 94.640 ;
                RECT 290.840 94.320 301.360 94.640 ;
                RECT 664.840 94.320 674.320 94.640 ;
                RECT 0.160 95.680 171.480 96.000 ;
                RECT 290.840 95.680 301.360 96.000 ;
                RECT 664.840 95.680 674.320 96.000 ;
                RECT 0.160 97.040 171.480 97.360 ;
                RECT 290.840 97.040 301.360 97.360 ;
                RECT 664.840 97.040 674.320 97.360 ;
                RECT 0.160 98.400 171.480 98.720 ;
                RECT 289.480 98.400 301.360 98.720 ;
                RECT 664.840 98.400 674.320 98.720 ;
                RECT 0.160 99.760 171.480 100.080 ;
                RECT 269.080 99.760 301.360 100.080 ;
                RECT 664.840 99.760 674.320 100.080 ;
                RECT 0.160 101.120 171.480 101.440 ;
                RECT 293.560 101.120 301.360 101.440 ;
                RECT 664.840 101.120 674.320 101.440 ;
                RECT 0.160 102.480 171.480 102.800 ;
                RECT 293.560 102.480 301.360 102.800 ;
                RECT 664.840 102.480 674.320 102.800 ;
                RECT 0.160 103.840 171.480 104.160 ;
                RECT 293.560 103.840 301.360 104.160 ;
                RECT 664.840 103.840 674.320 104.160 ;
                RECT 0.160 105.200 171.480 105.520 ;
                RECT 292.200 105.200 301.360 105.520 ;
                RECT 664.840 105.200 674.320 105.520 ;
                RECT 0.160 106.560 171.480 106.880 ;
                RECT 293.560 106.560 301.360 106.880 ;
                RECT 664.840 106.560 674.320 106.880 ;
                RECT 0.160 107.920 171.480 108.240 ;
                RECT 269.080 107.920 301.360 108.240 ;
                RECT 664.840 107.920 674.320 108.240 ;
                RECT 0.160 109.280 171.480 109.600 ;
                RECT 293.560 109.280 301.360 109.600 ;
                RECT 664.840 109.280 674.320 109.600 ;
                RECT 0.160 110.640 171.480 110.960 ;
                RECT 296.280 110.640 301.360 110.960 ;
                RECT 664.840 110.640 674.320 110.960 ;
                RECT 0.160 112.000 171.480 112.320 ;
                RECT 294.920 112.000 301.360 112.320 ;
                RECT 664.840 112.000 674.320 112.320 ;
                RECT 0.160 113.360 171.480 113.680 ;
                RECT 296.280 113.360 301.360 113.680 ;
                RECT 664.840 113.360 674.320 113.680 ;
                RECT 0.160 114.720 171.480 115.040 ;
                RECT 296.280 114.720 301.360 115.040 ;
                RECT 664.840 114.720 674.320 115.040 ;
                RECT 0.160 116.080 171.480 116.400 ;
                RECT 269.080 116.080 301.360 116.400 ;
                RECT 664.840 116.080 674.320 116.400 ;
                RECT 0.160 117.440 171.480 117.760 ;
                RECT 296.280 117.440 301.360 117.760 ;
                RECT 664.840 117.440 674.320 117.760 ;
                RECT 0.160 118.800 171.480 119.120 ;
                RECT 294.920 118.800 301.360 119.120 ;
                RECT 664.840 118.800 674.320 119.120 ;
                RECT 0.160 120.160 171.480 120.480 ;
                RECT 296.280 120.160 301.360 120.480 ;
                RECT 664.840 120.160 674.320 120.480 ;
                RECT 0.160 121.520 171.480 121.840 ;
                RECT 299.000 121.520 301.360 121.840 ;
                RECT 664.840 121.520 674.320 121.840 ;
                RECT 0.160 122.880 171.480 123.200 ;
                RECT 299.000 122.880 301.360 123.200 ;
                RECT 664.840 122.880 674.320 123.200 ;
                RECT 0.160 124.240 171.480 124.560 ;
                RECT 297.640 124.240 301.360 124.560 ;
                RECT 664.840 124.240 674.320 124.560 ;
                RECT 0.160 125.600 171.480 125.920 ;
                RECT 269.080 125.600 301.360 125.920 ;
                RECT 664.840 125.600 674.320 125.920 ;
                RECT 0.160 126.960 171.480 127.280 ;
                RECT 299.000 126.960 301.360 127.280 ;
                RECT 664.840 126.960 674.320 127.280 ;
                RECT 0.160 128.320 171.480 128.640 ;
                RECT 299.000 128.320 301.360 128.640 ;
                RECT 664.840 128.320 674.320 128.640 ;
                RECT 0.160 129.680 171.480 130.000 ;
                RECT 299.000 129.680 301.360 130.000 ;
                RECT 664.840 129.680 674.320 130.000 ;
                RECT 0.160 131.040 171.480 131.360 ;
                RECT 297.640 131.040 301.360 131.360 ;
                RECT 664.840 131.040 674.320 131.360 ;
                RECT 0.160 132.400 171.480 132.720 ;
                RECT 664.840 132.400 674.320 132.720 ;
                RECT 0.160 133.760 171.480 134.080 ;
                RECT 269.080 133.760 301.360 134.080 ;
                RECT 664.840 133.760 674.320 134.080 ;
                RECT 0.160 135.120 171.480 135.440 ;
                RECT 664.840 135.120 674.320 135.440 ;
                RECT 0.160 136.480 171.480 136.800 ;
                RECT 664.840 136.480 674.320 136.800 ;
                RECT 0.160 137.840 171.480 138.160 ;
                RECT 664.840 137.840 674.320 138.160 ;
                RECT 0.160 139.200 171.480 139.520 ;
                RECT 664.840 139.200 674.320 139.520 ;
                RECT 0.160 140.560 171.480 140.880 ;
                RECT 664.840 140.560 674.320 140.880 ;
                RECT 0.160 141.920 110.280 142.240 ;
                RECT 129.000 141.920 171.480 142.240 ;
                RECT 269.080 141.920 301.360 142.240 ;
                RECT 664.840 141.920 674.320 142.240 ;
                RECT 0.160 143.280 110.280 143.600 ;
                RECT 129.000 143.280 301.360 143.600 ;
                RECT 664.840 143.280 674.320 143.600 ;
                RECT 0.160 144.640 110.280 144.960 ;
                RECT 129.000 144.640 301.360 144.960 ;
                RECT 664.840 144.640 674.320 144.960 ;
                RECT 0.160 146.000 110.280 146.320 ;
                RECT 129.000 146.000 276.880 146.320 ;
                RECT 664.840 146.000 674.320 146.320 ;
                RECT 0.160 147.360 110.280 147.680 ;
                RECT 129.000 147.360 298.640 147.680 ;
                RECT 664.840 147.360 674.320 147.680 ;
                RECT 0.160 148.720 110.280 149.040 ;
                RECT 129.000 148.720 295.920 149.040 ;
                RECT 664.840 148.720 674.320 149.040 ;
                RECT 0.160 150.080 110.280 150.400 ;
                RECT 129.000 150.080 293.200 150.400 ;
                RECT 664.840 150.080 674.320 150.400 ;
                RECT 0.160 151.440 110.280 151.760 ;
                RECT 129.000 151.440 290.480 151.760 ;
                RECT 664.840 151.440 674.320 151.760 ;
                RECT 0.160 152.800 110.280 153.120 ;
                RECT 129.000 152.800 285.040 153.120 ;
                RECT 664.840 152.800 674.320 153.120 ;
                RECT 0.160 154.160 110.280 154.480 ;
                RECT 129.000 154.160 282.320 154.480 ;
                RECT 664.840 154.160 674.320 154.480 ;
                RECT 0.160 155.520 110.280 155.840 ;
                RECT 129.000 155.520 132.040 155.840 ;
                RECT 143.280 155.520 279.600 155.840 ;
                RECT 664.840 155.520 674.320 155.840 ;
                RECT 0.160 156.880 110.280 157.200 ;
                RECT 129.000 156.880 133.400 157.200 ;
                RECT 139.200 156.880 147.000 157.200 ;
                RECT 149.400 156.880 279.600 157.200 ;
                RECT 664.840 156.880 674.320 157.200 ;
                RECT 0.160 158.240 110.280 158.560 ;
                RECT 129.000 158.240 134.760 158.560 ;
                RECT 138.520 158.240 301.360 158.560 ;
                RECT 664.840 158.240 674.320 158.560 ;
                RECT 0.160 159.600 110.280 159.920 ;
                RECT 129.000 159.600 141.560 159.920 ;
                RECT 148.720 159.600 301.360 159.920 ;
                RECT 664.840 159.600 674.320 159.920 ;
                RECT 0.160 160.960 110.280 161.280 ;
                RECT 129.000 160.960 136.800 161.280 ;
                RECT 150.080 160.960 301.360 161.280 ;
                RECT 664.840 160.960 674.320 161.280 ;
                RECT 0.160 162.320 110.280 162.640 ;
                RECT 129.000 162.320 134.080 162.640 ;
                RECT 143.280 162.320 301.360 162.640 ;
                RECT 664.840 162.320 674.320 162.640 ;
                RECT 0.160 163.680 110.280 164.000 ;
                RECT 129.000 163.680 301.360 164.000 ;
                RECT 664.840 163.680 674.320 164.000 ;
                RECT 0.160 165.040 110.280 165.360 ;
                RECT 129.000 165.040 133.400 165.360 ;
                RECT 136.480 165.040 301.360 165.360 ;
                RECT 664.840 165.040 674.320 165.360 ;
                RECT 0.160 166.400 110.280 166.720 ;
                RECT 129.000 166.400 131.360 166.720 ;
                RECT 149.400 166.400 301.360 166.720 ;
                RECT 664.840 166.400 674.320 166.720 ;
                RECT 0.160 167.760 110.280 168.080 ;
                RECT 129.000 167.760 140.880 168.080 ;
                RECT 143.280 167.760 301.360 168.080 ;
                RECT 664.840 167.760 674.320 168.080 ;
                RECT 0.160 169.120 110.280 169.440 ;
                RECT 129.000 169.120 301.360 169.440 ;
                RECT 664.840 169.120 674.320 169.440 ;
                RECT 0.160 170.480 110.280 170.800 ;
                RECT 129.000 170.480 141.560 170.800 ;
                RECT 149.400 170.480 301.360 170.800 ;
                RECT 664.840 170.480 674.320 170.800 ;
                RECT 0.160 171.840 110.280 172.160 ;
                RECT 129.000 171.840 138.160 172.160 ;
                RECT 143.280 171.840 301.360 172.160 ;
                RECT 664.840 171.840 674.320 172.160 ;
                RECT 0.160 173.200 110.280 173.520 ;
                RECT 129.000 173.200 140.880 173.520 ;
                RECT 143.280 173.200 301.360 173.520 ;
                RECT 664.840 173.200 674.320 173.520 ;
                RECT 0.160 174.560 110.280 174.880 ;
                RECT 129.000 174.560 301.360 174.880 ;
                RECT 664.840 174.560 674.320 174.880 ;
                RECT 0.160 175.920 110.280 176.240 ;
                RECT 129.000 175.920 132.040 176.240 ;
                RECT 154.840 175.920 301.360 176.240 ;
                RECT 664.840 175.920 674.320 176.240 ;
                RECT 0.160 177.280 110.280 177.600 ;
                RECT 129.000 177.280 301.360 177.600 ;
                RECT 664.840 177.280 674.320 177.600 ;
                RECT 0.160 178.640 110.280 178.960 ;
                RECT 129.000 178.640 140.880 178.960 ;
                RECT 143.280 178.640 149.040 178.960 ;
                RECT 156.880 178.640 301.360 178.960 ;
                RECT 664.840 178.640 674.320 178.960 ;
                RECT 0.160 180.000 110.280 180.320 ;
                RECT 129.000 180.000 132.040 180.320 ;
                RECT 146.000 180.000 301.360 180.320 ;
                RECT 664.840 180.000 674.320 180.320 ;
                RECT 0.160 181.360 110.280 181.680 ;
                RECT 129.000 181.360 140.880 181.680 ;
                RECT 149.400 181.360 301.360 181.680 ;
                RECT 664.840 181.360 674.320 181.680 ;
                RECT 0.160 182.720 110.280 183.040 ;
                RECT 129.000 182.720 138.840 183.040 ;
                RECT 142.600 182.720 301.360 183.040 ;
                RECT 664.840 182.720 674.320 183.040 ;
                RECT 0.160 184.080 110.280 184.400 ;
                RECT 129.000 184.080 141.560 184.400 ;
                RECT 150.080 184.080 301.360 184.400 ;
                RECT 664.840 184.080 674.320 184.400 ;
                RECT 0.160 185.440 110.280 185.760 ;
                RECT 129.000 185.440 301.360 185.760 ;
                RECT 664.840 185.440 674.320 185.760 ;
                RECT 0.160 186.800 110.280 187.120 ;
                RECT 129.000 186.800 134.760 187.120 ;
                RECT 137.160 186.800 301.360 187.120 ;
                RECT 664.840 186.800 674.320 187.120 ;
                RECT 0.160 188.160 110.280 188.480 ;
                RECT 129.680 188.160 134.080 188.480 ;
                RECT 143.280 188.160 301.360 188.480 ;
                RECT 664.840 188.160 674.320 188.480 ;
                RECT 0.160 189.520 110.280 189.840 ;
                RECT 129.000 189.520 301.360 189.840 ;
                RECT 664.840 189.520 674.320 189.840 ;
                RECT 0.160 190.880 110.280 191.200 ;
                RECT 129.000 190.880 140.880 191.200 ;
                RECT 142.600 190.880 301.360 191.200 ;
                RECT 664.840 190.880 674.320 191.200 ;
                RECT 0.160 192.240 110.280 192.560 ;
                RECT 129.000 192.240 133.400 192.560 ;
                RECT 139.200 192.240 141.560 192.560 ;
                RECT 143.960 192.240 218.400 192.560 ;
                RECT 269.080 192.240 301.360 192.560 ;
                RECT 664.840 192.240 674.320 192.560 ;
                RECT 0.160 193.600 110.280 193.920 ;
                RECT 129.000 193.600 137.480 193.920 ;
                RECT 148.720 193.600 218.400 193.920 ;
                RECT 269.080 193.600 301.360 193.920 ;
                RECT 664.840 193.600 674.320 193.920 ;
                RECT 0.160 194.960 110.280 195.280 ;
                RECT 129.000 194.960 140.880 195.280 ;
                RECT 142.600 194.960 218.400 195.280 ;
                RECT 269.080 194.960 301.360 195.280 ;
                RECT 664.840 194.960 674.320 195.280 ;
                RECT 0.160 196.320 110.280 196.640 ;
                RECT 129.000 196.320 135.440 196.640 ;
                RECT 143.280 196.320 218.400 196.640 ;
                RECT 269.080 196.320 301.360 196.640 ;
                RECT 664.840 196.320 674.320 196.640 ;
                RECT 0.160 197.680 110.280 198.000 ;
                RECT 129.000 197.680 140.880 198.000 ;
                RECT 143.960 197.680 218.400 198.000 ;
                RECT 269.080 197.680 301.360 198.000 ;
                RECT 664.840 197.680 674.320 198.000 ;
                RECT 0.160 199.040 110.280 199.360 ;
                RECT 129.000 199.040 132.040 199.360 ;
                RECT 139.200 199.040 301.360 199.360 ;
                RECT 664.840 199.040 674.320 199.360 ;
                RECT 0.160 200.400 110.280 200.720 ;
                RECT 129.000 200.400 131.360 200.720 ;
                RECT 149.400 200.400 301.360 200.720 ;
                RECT 664.840 200.400 674.320 200.720 ;
                RECT 0.160 201.760 110.280 202.080 ;
                RECT 142.600 201.760 301.360 202.080 ;
                RECT 664.840 201.760 674.320 202.080 ;
                RECT 0.160 203.120 110.280 203.440 ;
                RECT 129.000 203.120 132.040 203.440 ;
                RECT 137.160 203.120 203.440 203.440 ;
                RECT 270.440 203.120 301.360 203.440 ;
                RECT 664.840 203.120 674.320 203.440 ;
                RECT 0.160 204.480 110.280 204.800 ;
                RECT 129.000 204.480 203.440 204.800 ;
                RECT 270.440 204.480 301.360 204.800 ;
                RECT 664.840 204.480 674.320 204.800 ;
                RECT 0.160 205.840 110.280 206.160 ;
                RECT 129.000 205.840 138.840 206.160 ;
                RECT 146.000 205.840 203.440 206.160 ;
                RECT 270.440 205.840 280.960 206.160 ;
                RECT 664.840 205.840 674.320 206.160 ;
                RECT 0.160 207.200 110.280 207.520 ;
                RECT 129.000 207.200 203.440 207.520 ;
                RECT 270.440 207.200 283.680 207.520 ;
                RECT 664.840 207.200 674.320 207.520 ;
                RECT 0.160 208.560 110.280 208.880 ;
                RECT 129.000 208.560 203.440 208.880 ;
                RECT 270.440 208.560 286.400 208.880 ;
                RECT 664.840 208.560 674.320 208.880 ;
                RECT 0.160 209.920 110.280 210.240 ;
                RECT 129.000 209.920 203.440 210.240 ;
                RECT 270.440 209.920 289.120 210.240 ;
                RECT 664.840 209.920 674.320 210.240 ;
                RECT 0.160 211.280 110.280 211.600 ;
                RECT 129.000 211.280 144.280 211.600 ;
                RECT 150.760 211.280 203.440 211.600 ;
                RECT 270.440 211.280 291.840 211.600 ;
                RECT 664.840 211.280 674.320 211.600 ;
                RECT 0.160 212.640 110.280 212.960 ;
                RECT 129.000 212.640 132.040 212.960 ;
                RECT 137.160 212.640 203.440 212.960 ;
                RECT 270.440 212.640 294.560 212.960 ;
                RECT 664.840 212.640 674.320 212.960 ;
                RECT 0.160 214.000 110.280 214.320 ;
                RECT 129.000 214.000 203.440 214.320 ;
                RECT 270.440 214.000 297.280 214.320 ;
                RECT 664.840 214.000 674.320 214.320 ;
                RECT 0.160 215.360 110.280 215.680 ;
                RECT 129.000 215.360 203.440 215.680 ;
                RECT 270.440 215.360 300.000 215.680 ;
                RECT 664.840 215.360 674.320 215.680 ;
                RECT 0.160 216.720 110.280 217.040 ;
                RECT 129.000 216.720 203.440 217.040 ;
                RECT 664.840 216.720 674.320 217.040 ;
                RECT 0.160 218.080 110.280 218.400 ;
                RECT 129.000 218.080 203.440 218.400 ;
                RECT 664.840 218.080 674.320 218.400 ;
                RECT 0.160 219.440 110.280 219.760 ;
                RECT 129.000 219.440 203.440 219.760 ;
                RECT 664.840 219.440 674.320 219.760 ;
                RECT 0.160 220.800 110.280 221.120 ;
                RECT 129.000 220.800 203.440 221.120 ;
                RECT 270.440 220.800 301.360 221.120 ;
                RECT 664.840 220.800 674.320 221.120 ;
                RECT 0.160 222.160 110.280 222.480 ;
                RECT 129.000 222.160 134.080 222.480 ;
                RECT 149.400 222.160 203.440 222.480 ;
                RECT 270.440 222.160 301.360 222.480 ;
                RECT 664.840 222.160 674.320 222.480 ;
                RECT 0.160 223.520 110.280 223.840 ;
                RECT 129.000 223.520 203.440 223.840 ;
                RECT 270.440 223.520 301.360 223.840 ;
                RECT 664.840 223.520 674.320 223.840 ;
                RECT 0.160 224.880 110.280 225.200 ;
                RECT 129.000 224.880 203.440 225.200 ;
                RECT 270.440 224.880 301.360 225.200 ;
                RECT 664.840 224.880 674.320 225.200 ;
                RECT 0.160 226.240 110.280 226.560 ;
                RECT 129.000 226.240 203.440 226.560 ;
                RECT 270.440 226.240 301.360 226.560 ;
                RECT 664.840 226.240 674.320 226.560 ;
                RECT 0.160 227.600 110.280 227.920 ;
                RECT 129.000 227.600 203.440 227.920 ;
                RECT 270.440 227.600 301.360 227.920 ;
                RECT 664.840 227.600 674.320 227.920 ;
                RECT 0.160 228.960 110.280 229.280 ;
                RECT 129.000 228.960 133.400 229.280 ;
                RECT 136.480 228.960 203.440 229.280 ;
                RECT 270.440 228.960 301.360 229.280 ;
                RECT 664.840 228.960 674.320 229.280 ;
                RECT 0.160 230.320 110.280 230.640 ;
                RECT 129.000 230.320 136.800 230.640 ;
                RECT 139.200 230.320 203.440 230.640 ;
                RECT 270.440 230.320 301.360 230.640 ;
                RECT 664.840 230.320 674.320 230.640 ;
                RECT 0.160 231.680 110.280 232.000 ;
                RECT 129.000 231.680 147.680 232.000 ;
                RECT 150.080 231.680 203.440 232.000 ;
                RECT 270.440 231.680 301.360 232.000 ;
                RECT 664.840 231.680 674.320 232.000 ;
                RECT 0.160 233.040 110.280 233.360 ;
                RECT 129.000 233.040 203.440 233.360 ;
                RECT 270.440 233.040 301.360 233.360 ;
                RECT 664.840 233.040 674.320 233.360 ;
                RECT 0.160 234.400 110.280 234.720 ;
                RECT 129.000 234.400 203.440 234.720 ;
                RECT 270.440 234.400 301.360 234.720 ;
                RECT 664.840 234.400 674.320 234.720 ;
                RECT 0.160 235.760 110.280 236.080 ;
                RECT 129.000 235.760 203.440 236.080 ;
                RECT 270.440 235.760 301.360 236.080 ;
                RECT 664.840 235.760 674.320 236.080 ;
                RECT 0.160 237.120 110.280 237.440 ;
                RECT 129.000 237.120 203.440 237.440 ;
                RECT 270.440 237.120 301.360 237.440 ;
                RECT 664.840 237.120 674.320 237.440 ;
                RECT 0.160 238.480 203.440 238.800 ;
                RECT 270.440 238.480 301.360 238.800 ;
                RECT 664.840 238.480 674.320 238.800 ;
                RECT 0.160 239.840 140.880 240.160 ;
                RECT 149.400 239.840 203.440 240.160 ;
                RECT 270.440 239.840 301.360 240.160 ;
                RECT 664.840 239.840 674.320 240.160 ;
                RECT 0.160 241.200 135.440 241.520 ;
                RECT 139.200 241.200 203.440 241.520 ;
                RECT 270.440 241.200 301.360 241.520 ;
                RECT 664.840 241.200 674.320 241.520 ;
                RECT 0.160 242.560 89.200 242.880 ;
                RECT 110.640 242.560 203.440 242.880 ;
                RECT 270.440 242.560 301.360 242.880 ;
                RECT 664.840 242.560 674.320 242.880 ;
                RECT 0.160 243.920 89.200 244.240 ;
                RECT 110.640 243.920 203.440 244.240 ;
                RECT 270.440 243.920 301.360 244.240 ;
                RECT 664.840 243.920 674.320 244.240 ;
                RECT 0.160 245.280 89.200 245.600 ;
                RECT 110.640 245.280 116.400 245.600 ;
                RECT 124.240 245.280 203.440 245.600 ;
                RECT 270.440 245.280 301.360 245.600 ;
                RECT 664.840 245.280 674.320 245.600 ;
                RECT 0.160 246.640 137.480 246.960 ;
                RECT 143.960 246.640 203.440 246.960 ;
                RECT 270.440 246.640 301.360 246.960 ;
                RECT 664.840 246.640 674.320 246.960 ;
                RECT 0.160 248.000 89.200 248.320 ;
                RECT 128.320 248.000 203.440 248.320 ;
                RECT 664.840 248.000 674.320 248.320 ;
                RECT 0.160 249.360 89.200 249.680 ;
                RECT 128.320 249.360 203.440 249.680 ;
                RECT 664.840 249.360 674.320 249.680 ;
                RECT 0.160 250.720 89.200 251.040 ;
                RECT 110.640 250.720 203.440 251.040 ;
                RECT 664.840 250.720 674.320 251.040 ;
                RECT 0.160 252.080 74.920 252.400 ;
                RECT 124.240 252.080 132.040 252.400 ;
                RECT 142.600 252.080 203.440 252.400 ;
                RECT 270.440 252.080 301.360 252.400 ;
                RECT 664.840 252.080 674.320 252.400 ;
                RECT 0.160 253.440 116.400 253.760 ;
                RECT 136.480 253.440 674.320 253.760 ;
                RECT 0.160 254.800 33.440 255.120 ;
                RECT 135.800 254.800 674.320 255.120 ;
                RECT 0.160 256.160 298.640 256.480 ;
                RECT 666.880 256.160 674.320 256.480 ;
                RECT 0.160 257.520 298.640 257.840 ;
                RECT 666.880 257.520 674.320 257.840 ;
                RECT 0.160 258.880 28.680 259.200 ;
                RECT 35.160 258.880 106.200 259.200 ;
                RECT 666.880 258.880 674.320 259.200 ;
                RECT 0.160 260.240 26.640 260.560 ;
                RECT 37.200 260.240 38.200 260.560 ;
                RECT 50.800 260.240 106.200 260.560 ;
                RECT 666.880 260.240 674.320 260.560 ;
                RECT 0.160 261.600 26.640 261.920 ;
                RECT 37.200 261.600 39.560 261.920 ;
                RECT 50.120 261.600 62.680 261.920 ;
                RECT 64.400 261.600 77.640 261.920 ;
                RECT 95.680 261.600 106.200 261.920 ;
                RECT 666.880 261.600 674.320 261.920 ;
                RECT 0.160 262.960 62.680 263.280 ;
                RECT 64.400 262.960 77.640 263.280 ;
                RECT 95.680 262.960 106.200 263.280 ;
                RECT 666.880 262.960 674.320 263.280 ;
                RECT 0.160 264.320 26.640 264.640 ;
                RECT 37.200 264.320 62.680 264.640 ;
                RECT 67.120 264.320 77.640 264.640 ;
                RECT 95.680 264.320 106.200 264.640 ;
                RECT 666.880 264.320 674.320 264.640 ;
                RECT 0.160 265.680 62.680 266.000 ;
                RECT 67.800 265.680 77.640 266.000 ;
                RECT 95.680 265.680 106.200 266.000 ;
                RECT 666.880 265.680 674.320 266.000 ;
                RECT 0.160 267.040 26.640 267.360 ;
                RECT 37.200 267.040 62.680 267.360 ;
                RECT 68.480 267.040 77.640 267.360 ;
                RECT 95.680 267.040 106.200 267.360 ;
                RECT 666.880 267.040 674.320 267.360 ;
                RECT 0.160 268.400 26.640 268.720 ;
                RECT 37.200 268.400 106.200 268.720 ;
                RECT 666.880 268.400 674.320 268.720 ;
                RECT 0.160 269.760 77.640 270.080 ;
                RECT 95.680 269.760 106.200 270.080 ;
                RECT 666.880 269.760 674.320 270.080 ;
                RECT 0.160 271.120 77.640 271.440 ;
                RECT 95.680 271.120 106.200 271.440 ;
                RECT 666.880 271.120 674.320 271.440 ;
                RECT 0.160 272.480 77.640 272.800 ;
                RECT 95.680 272.480 106.200 272.800 ;
                RECT 666.880 272.480 674.320 272.800 ;
                RECT 0.160 273.840 19.840 274.160 ;
                RECT 22.240 273.840 35.480 274.160 ;
                RECT 38.560 273.840 77.640 274.160 ;
                RECT 95.680 273.840 106.200 274.160 ;
                RECT 666.880 273.840 674.320 274.160 ;
                RECT 0.160 275.200 19.160 275.520 ;
                RECT 22.240 275.200 40.240 275.520 ;
                RECT 51.480 275.200 77.640 275.520 ;
                RECT 88.880 275.200 106.200 275.520 ;
                RECT 666.880 275.200 674.320 275.520 ;
                RECT 0.160 276.560 18.480 276.880 ;
                RECT 22.240 276.560 41.600 276.880 ;
                RECT 50.800 276.560 89.880 276.880 ;
                RECT 95.680 276.560 106.200 276.880 ;
                RECT 666.880 276.560 674.320 276.880 ;
                RECT 0.160 277.920 17.800 278.240 ;
                RECT 22.240 277.920 62.680 278.240 ;
                RECT 65.080 277.920 77.640 278.240 ;
                RECT 95.680 277.920 106.200 278.240 ;
                RECT 666.880 277.920 674.320 278.240 ;
                RECT 0.160 279.280 62.680 279.600 ;
                RECT 65.760 279.280 77.640 279.600 ;
                RECT 95.680 279.280 106.200 279.600 ;
                RECT 666.880 279.280 674.320 279.600 ;
                RECT 0.160 280.640 17.120 280.960 ;
                RECT 22.240 280.640 62.680 280.960 ;
                RECT 65.760 280.640 77.640 280.960 ;
                RECT 95.680 280.640 106.200 280.960 ;
                RECT 666.880 280.640 674.320 280.960 ;
                RECT 0.160 282.000 16.440 282.320 ;
                RECT 22.240 282.000 62.680 282.320 ;
                RECT 64.400 282.000 77.640 282.320 ;
                RECT 95.680 282.000 106.200 282.320 ;
                RECT 666.880 282.000 674.320 282.320 ;
                RECT 0.160 283.360 62.680 283.680 ;
                RECT 66.440 283.360 77.640 283.680 ;
                RECT 88.880 283.360 106.200 283.680 ;
                RECT 666.880 283.360 674.320 283.680 ;
                RECT 0.160 284.720 15.760 285.040 ;
                RECT 22.240 284.720 35.480 285.040 ;
                RECT 42.640 284.720 77.640 285.040 ;
                RECT 95.680 284.720 106.200 285.040 ;
                RECT 666.880 284.720 674.320 285.040 ;
                RECT 0.160 286.080 15.080 286.400 ;
                RECT 22.240 286.080 35.480 286.400 ;
                RECT 43.320 286.080 77.640 286.400 ;
                RECT 95.680 286.080 106.200 286.400 ;
                RECT 666.880 286.080 674.320 286.400 ;
                RECT 0.160 287.440 77.640 287.760 ;
                RECT 95.680 287.440 106.200 287.760 ;
                RECT 666.880 287.440 674.320 287.760 ;
                RECT 0.160 288.800 14.400 289.120 ;
                RECT 22.240 288.800 35.480 289.120 ;
                RECT 43.320 288.800 77.640 289.120 ;
                RECT 95.680 288.800 106.200 289.120 ;
                RECT 666.880 288.800 674.320 289.120 ;
                RECT 0.160 290.160 13.720 290.480 ;
                RECT 22.240 290.160 35.480 290.480 ;
                RECT 42.640 290.160 77.640 290.480 ;
                RECT 95.680 290.160 106.200 290.480 ;
                RECT 666.880 290.160 674.320 290.480 ;
                RECT 0.160 291.520 13.040 291.840 ;
                RECT 22.240 291.520 106.200 291.840 ;
                RECT 666.880 291.520 674.320 291.840 ;
                RECT 0.160 292.880 12.360 293.200 ;
                RECT 22.240 292.880 77.640 293.200 ;
                RECT 95.680 292.880 106.200 293.200 ;
                RECT 666.880 292.880 674.320 293.200 ;
                RECT 0.160 294.240 77.640 294.560 ;
                RECT 95.680 294.240 106.200 294.560 ;
                RECT 666.880 294.240 674.320 294.560 ;
                RECT 0.160 295.600 11.680 295.920 ;
                RECT 22.240 295.600 77.640 295.920 ;
                RECT 95.680 295.600 106.200 295.920 ;
                RECT 666.880 295.600 674.320 295.920 ;
                RECT 0.160 296.960 11.000 297.280 ;
                RECT 22.240 296.960 77.640 297.280 ;
                RECT 95.680 296.960 106.200 297.280 ;
                RECT 666.880 296.960 674.320 297.280 ;
                RECT 0.160 298.320 10.320 298.640 ;
                RECT 22.240 298.320 77.640 298.640 ;
                RECT 95.680 298.320 106.200 298.640 ;
                RECT 666.880 298.320 674.320 298.640 ;
                RECT 0.160 299.680 106.200 300.000 ;
                RECT 666.880 299.680 674.320 300.000 ;
                RECT 0.160 301.040 9.640 301.360 ;
                RECT 22.240 301.040 35.480 301.360 ;
                RECT 38.560 301.040 77.640 301.360 ;
                RECT 95.680 301.040 106.200 301.360 ;
                RECT 666.880 301.040 674.320 301.360 ;
                RECT 0.160 302.400 77.640 302.720 ;
                RECT 95.680 302.400 106.200 302.720 ;
                RECT 666.880 302.400 674.320 302.720 ;
                RECT 0.160 303.760 77.640 304.080 ;
                RECT 95.680 303.760 106.200 304.080 ;
                RECT 666.880 303.760 674.320 304.080 ;
                RECT 0.160 305.120 77.640 305.440 ;
                RECT 95.680 305.120 106.200 305.440 ;
                RECT 666.880 305.120 674.320 305.440 ;
                RECT 0.160 306.480 77.640 306.800 ;
                RECT 95.680 306.480 106.200 306.800 ;
                RECT 666.880 306.480 674.320 306.800 ;
                RECT 0.160 307.840 106.200 308.160 ;
                RECT 666.880 307.840 674.320 308.160 ;
                RECT 0.160 309.200 77.640 309.520 ;
                RECT 95.680 309.200 106.200 309.520 ;
                RECT 666.880 309.200 674.320 309.520 ;
                RECT 0.160 310.560 77.640 310.880 ;
                RECT 95.680 310.560 106.200 310.880 ;
                RECT 666.880 310.560 674.320 310.880 ;
                RECT 0.160 311.920 77.640 312.240 ;
                RECT 95.680 311.920 106.200 312.240 ;
                RECT 666.880 311.920 674.320 312.240 ;
                RECT 0.160 313.280 77.640 313.600 ;
                RECT 95.680 313.280 106.200 313.600 ;
                RECT 666.880 313.280 674.320 313.600 ;
                RECT 0.160 314.640 77.640 314.960 ;
                RECT 92.280 314.640 106.200 314.960 ;
                RECT 666.880 314.640 674.320 314.960 ;
                RECT 0.160 316.000 91.920 316.320 ;
                RECT 95.680 316.000 106.200 316.320 ;
                RECT 666.880 316.000 674.320 316.320 ;
                RECT 0.160 317.360 77.640 317.680 ;
                RECT 95.680 317.360 106.200 317.680 ;
                RECT 666.880 317.360 674.320 317.680 ;
                RECT 0.160 318.720 77.640 319.040 ;
                RECT 95.680 318.720 106.200 319.040 ;
                RECT 666.880 318.720 674.320 319.040 ;
                RECT 0.160 320.080 77.640 320.400 ;
                RECT 95.680 320.080 106.200 320.400 ;
                RECT 666.880 320.080 674.320 320.400 ;
                RECT 0.160 321.440 77.640 321.760 ;
                RECT 95.680 321.440 106.200 321.760 ;
                RECT 666.880 321.440 674.320 321.760 ;
                RECT 0.160 322.800 77.640 323.120 ;
                RECT 92.280 322.800 106.200 323.120 ;
                RECT 666.880 322.800 674.320 323.120 ;
                RECT 0.160 324.160 77.640 324.480 ;
                RECT 95.680 324.160 106.200 324.480 ;
                RECT 666.880 324.160 674.320 324.480 ;
                RECT 0.160 325.520 77.640 325.840 ;
                RECT 95.680 325.520 106.200 325.840 ;
                RECT 666.880 325.520 674.320 325.840 ;
                RECT 0.160 326.880 77.640 327.200 ;
                RECT 95.680 326.880 106.200 327.200 ;
                RECT 666.880 326.880 674.320 327.200 ;
                RECT 0.160 328.240 77.640 328.560 ;
                RECT 95.680 328.240 106.200 328.560 ;
                RECT 666.880 328.240 674.320 328.560 ;
                RECT 0.160 329.600 77.640 329.920 ;
                RECT 95.680 329.600 106.200 329.920 ;
                RECT 666.880 329.600 674.320 329.920 ;
                RECT 0.160 330.960 106.200 331.280 ;
                RECT 666.880 330.960 674.320 331.280 ;
                RECT 0.160 332.320 77.640 332.640 ;
                RECT 95.680 332.320 106.200 332.640 ;
                RECT 666.880 332.320 674.320 332.640 ;
                RECT 0.160 333.680 77.640 334.000 ;
                RECT 95.680 333.680 106.200 334.000 ;
                RECT 666.880 333.680 674.320 334.000 ;
                RECT 0.160 335.040 77.640 335.360 ;
                RECT 95.680 335.040 106.200 335.360 ;
                RECT 666.880 335.040 674.320 335.360 ;
                RECT 0.160 336.400 77.640 336.720 ;
                RECT 95.680 336.400 106.200 336.720 ;
                RECT 666.880 336.400 674.320 336.720 ;
                RECT 0.160 337.760 77.640 338.080 ;
                RECT 95.680 337.760 106.200 338.080 ;
                RECT 666.880 337.760 674.320 338.080 ;
                RECT 0.160 339.120 106.200 339.440 ;
                RECT 666.880 339.120 674.320 339.440 ;
                RECT 0.160 340.480 77.640 340.800 ;
                RECT 95.680 340.480 106.200 340.800 ;
                RECT 666.880 340.480 674.320 340.800 ;
                RECT 0.160 341.840 77.640 342.160 ;
                RECT 95.680 341.840 106.200 342.160 ;
                RECT 666.880 341.840 674.320 342.160 ;
                RECT 0.160 343.200 77.640 343.520 ;
                RECT 95.680 343.200 106.200 343.520 ;
                RECT 666.880 343.200 674.320 343.520 ;
                RECT 0.160 344.560 77.640 344.880 ;
                RECT 95.680 344.560 106.200 344.880 ;
                RECT 666.880 344.560 674.320 344.880 ;
                RECT 0.160 345.920 77.640 346.240 ;
                RECT 95.680 345.920 106.200 346.240 ;
                RECT 666.880 345.920 674.320 346.240 ;
                RECT 0.160 347.280 106.200 347.600 ;
                RECT 666.880 347.280 674.320 347.600 ;
                RECT 0.160 348.640 77.640 348.960 ;
                RECT 95.680 348.640 106.200 348.960 ;
                RECT 666.880 348.640 674.320 348.960 ;
                RECT 0.160 350.000 77.640 350.320 ;
                RECT 95.680 350.000 106.200 350.320 ;
                RECT 666.880 350.000 674.320 350.320 ;
                RECT 0.160 351.360 77.640 351.680 ;
                RECT 95.680 351.360 106.200 351.680 ;
                RECT 666.880 351.360 674.320 351.680 ;
                RECT 0.160 352.720 77.640 353.040 ;
                RECT 95.680 352.720 106.200 353.040 ;
                RECT 666.880 352.720 674.320 353.040 ;
                RECT 0.160 354.080 77.640 354.400 ;
                RECT 95.000 354.080 106.200 354.400 ;
                RECT 666.880 354.080 674.320 354.400 ;
                RECT 0.160 355.440 85.800 355.760 ;
                RECT 95.680 355.440 106.200 355.760 ;
                RECT 666.880 355.440 674.320 355.760 ;
                RECT 0.160 356.800 79.680 357.120 ;
                RECT 95.680 356.800 106.200 357.120 ;
                RECT 666.880 356.800 674.320 357.120 ;
                RECT 0.160 358.160 79.680 358.480 ;
                RECT 95.680 358.160 106.200 358.480 ;
                RECT 666.880 358.160 674.320 358.480 ;
                RECT 0.160 359.520 79.680 359.840 ;
                RECT 95.680 359.520 106.200 359.840 ;
                RECT 666.880 359.520 674.320 359.840 ;
                RECT 0.160 360.880 79.680 361.200 ;
                RECT 95.680 360.880 106.200 361.200 ;
                RECT 666.880 360.880 674.320 361.200 ;
                RECT 0.160 362.240 42.280 362.560 ;
                RECT 51.480 362.240 106.200 362.560 ;
                RECT 666.880 362.240 674.320 362.560 ;
                RECT 0.160 363.600 40.920 363.920 ;
                RECT 50.800 363.600 62.680 363.920 ;
                RECT 64.400 363.600 77.640 363.920 ;
                RECT 95.680 363.600 106.200 363.920 ;
                RECT 666.880 363.600 674.320 363.920 ;
                RECT 0.160 364.960 62.680 365.280 ;
                RECT 67.120 364.960 77.640 365.280 ;
                RECT 95.680 364.960 106.200 365.280 ;
                RECT 666.880 364.960 674.320 365.280 ;
                RECT 0.160 366.320 62.680 366.640 ;
                RECT 67.120 366.320 77.640 366.640 ;
                RECT 95.680 366.320 106.200 366.640 ;
                RECT 666.880 366.320 674.320 366.640 ;
                RECT 0.160 367.680 62.680 368.000 ;
                RECT 67.800 367.680 77.640 368.000 ;
                RECT 95.680 367.680 106.200 368.000 ;
                RECT 666.880 367.680 674.320 368.000 ;
                RECT 0.160 369.040 62.680 369.360 ;
                RECT 64.400 369.040 77.640 369.360 ;
                RECT 95.680 369.040 106.200 369.360 ;
                RECT 666.880 369.040 674.320 369.360 ;
                RECT 0.160 370.400 106.200 370.720 ;
                RECT 666.880 370.400 674.320 370.720 ;
                RECT 0.160 371.760 77.640 372.080 ;
                RECT 95.680 371.760 106.200 372.080 ;
                RECT 666.880 371.760 674.320 372.080 ;
                RECT 0.160 373.120 77.640 373.440 ;
                RECT 95.680 373.120 106.200 373.440 ;
                RECT 666.880 373.120 674.320 373.440 ;
                RECT 0.160 374.480 77.640 374.800 ;
                RECT 95.680 374.480 106.200 374.800 ;
                RECT 666.880 374.480 674.320 374.800 ;
                RECT 0.160 375.840 77.640 376.160 ;
                RECT 95.680 375.840 106.200 376.160 ;
                RECT 666.880 375.840 674.320 376.160 ;
                RECT 0.160 377.200 77.640 377.520 ;
                RECT 95.680 377.200 106.200 377.520 ;
                RECT 666.880 377.200 674.320 377.520 ;
                RECT 0.160 378.560 38.880 378.880 ;
                RECT 50.800 378.560 106.200 378.880 ;
                RECT 666.880 378.560 674.320 378.880 ;
                RECT 0.160 379.920 37.520 380.240 ;
                RECT 50.120 379.920 62.680 380.240 ;
                RECT 64.400 379.920 77.640 380.240 ;
                RECT 95.680 379.920 106.200 380.240 ;
                RECT 666.880 379.920 674.320 380.240 ;
                RECT 0.160 381.280 62.680 381.600 ;
                RECT 65.080 381.280 77.640 381.600 ;
                RECT 95.680 381.280 106.200 381.600 ;
                RECT 666.880 381.280 674.320 381.600 ;
                RECT 0.160 382.640 62.680 382.960 ;
                RECT 65.760 382.640 77.640 382.960 ;
                RECT 95.680 382.640 106.200 382.960 ;
                RECT 666.880 382.640 674.320 382.960 ;
                RECT 0.160 384.000 62.680 384.320 ;
                RECT 65.760 384.000 77.640 384.320 ;
                RECT 95.680 384.000 106.200 384.320 ;
                RECT 666.880 384.000 674.320 384.320 ;
                RECT 0.160 385.360 62.680 385.680 ;
                RECT 66.440 385.360 77.640 385.680 ;
                RECT 95.680 385.360 106.200 385.680 ;
                RECT 666.880 385.360 674.320 385.680 ;
                RECT 0.160 386.720 106.200 387.040 ;
                RECT 666.880 386.720 674.320 387.040 ;
                RECT 0.160 388.080 77.640 388.400 ;
                RECT 95.680 388.080 106.200 388.400 ;
                RECT 666.880 388.080 674.320 388.400 ;
                RECT 0.160 389.440 77.640 389.760 ;
                RECT 95.680 389.440 106.200 389.760 ;
                RECT 666.880 389.440 674.320 389.760 ;
                RECT 0.160 390.800 77.640 391.120 ;
                RECT 95.680 390.800 106.200 391.120 ;
                RECT 666.880 390.800 674.320 391.120 ;
                RECT 0.160 392.160 77.640 392.480 ;
                RECT 95.680 392.160 106.200 392.480 ;
                RECT 666.880 392.160 674.320 392.480 ;
                RECT 0.160 393.520 77.640 393.840 ;
                RECT 82.080 393.520 106.200 393.840 ;
                RECT 666.880 393.520 674.320 393.840 ;
                RECT 0.160 394.880 106.200 395.200 ;
                RECT 666.880 394.880 674.320 395.200 ;
                RECT 0.160 396.240 77.640 396.560 ;
                RECT 95.680 396.240 106.200 396.560 ;
                RECT 666.880 396.240 674.320 396.560 ;
                RECT 0.160 397.600 77.640 397.920 ;
                RECT 95.680 397.600 106.200 397.920 ;
                RECT 666.880 397.600 674.320 397.920 ;
                RECT 0.160 398.960 77.640 399.280 ;
                RECT 95.680 398.960 106.200 399.280 ;
                RECT 666.880 398.960 674.320 399.280 ;
                RECT 0.160 400.320 77.640 400.640 ;
                RECT 95.680 400.320 106.200 400.640 ;
                RECT 666.880 400.320 674.320 400.640 ;
                RECT 0.160 401.680 77.640 402.000 ;
                RECT 82.760 401.680 106.200 402.000 ;
                RECT 666.880 401.680 674.320 402.000 ;
                RECT 0.160 403.040 77.640 403.360 ;
                RECT 95.680 403.040 106.200 403.360 ;
                RECT 666.880 403.040 674.320 403.360 ;
                RECT 0.160 404.400 77.640 404.720 ;
                RECT 95.680 404.400 106.200 404.720 ;
                RECT 666.880 404.400 674.320 404.720 ;
                RECT 0.160 405.760 77.640 406.080 ;
                RECT 95.680 405.760 106.200 406.080 ;
                RECT 666.880 405.760 674.320 406.080 ;
                RECT 0.160 407.120 77.640 407.440 ;
                RECT 95.680 407.120 106.200 407.440 ;
                RECT 666.880 407.120 674.320 407.440 ;
                RECT 0.160 408.480 77.640 408.800 ;
                RECT 95.680 408.480 106.200 408.800 ;
                RECT 666.880 408.480 674.320 408.800 ;
                RECT 0.160 409.840 77.640 410.160 ;
                RECT 83.440 409.840 106.200 410.160 ;
                RECT 666.880 409.840 674.320 410.160 ;
                RECT 0.160 411.200 77.640 411.520 ;
                RECT 95.680 411.200 106.200 411.520 ;
                RECT 666.880 411.200 674.320 411.520 ;
                RECT 0.160 412.560 77.640 412.880 ;
                RECT 95.680 412.560 106.200 412.880 ;
                RECT 666.880 412.560 674.320 412.880 ;
                RECT 0.160 413.920 77.640 414.240 ;
                RECT 95.680 413.920 106.200 414.240 ;
                RECT 666.880 413.920 674.320 414.240 ;
                RECT 0.160 415.280 77.640 415.600 ;
                RECT 95.680 415.280 106.200 415.600 ;
                RECT 666.880 415.280 674.320 415.600 ;
                RECT 0.160 416.640 77.640 416.960 ;
                RECT 95.680 416.640 106.200 416.960 ;
                RECT 666.880 416.640 674.320 416.960 ;
                RECT 0.160 418.000 106.200 418.320 ;
                RECT 666.880 418.000 674.320 418.320 ;
                RECT 0.160 419.360 77.640 419.680 ;
                RECT 95.680 419.360 106.200 419.680 ;
                RECT 666.880 419.360 674.320 419.680 ;
                RECT 0.160 420.720 77.640 421.040 ;
                RECT 95.680 420.720 106.200 421.040 ;
                RECT 666.880 420.720 674.320 421.040 ;
                RECT 0.160 422.080 77.640 422.400 ;
                RECT 95.680 422.080 106.200 422.400 ;
                RECT 666.880 422.080 674.320 422.400 ;
                RECT 0.160 423.440 77.640 423.760 ;
                RECT 95.680 423.440 106.200 423.760 ;
                RECT 666.880 423.440 674.320 423.760 ;
                RECT 0.160 424.800 77.640 425.120 ;
                RECT 95.680 424.800 106.200 425.120 ;
                RECT 666.880 424.800 674.320 425.120 ;
                RECT 0.160 426.160 106.200 426.480 ;
                RECT 666.880 426.160 674.320 426.480 ;
                RECT 0.160 427.520 77.640 427.840 ;
                RECT 95.680 427.520 106.200 427.840 ;
                RECT 666.880 427.520 674.320 427.840 ;
                RECT 0.160 428.880 77.640 429.200 ;
                RECT 95.680 428.880 106.200 429.200 ;
                RECT 666.880 428.880 674.320 429.200 ;
                RECT 0.160 430.240 77.640 430.560 ;
                RECT 95.680 430.240 106.200 430.560 ;
                RECT 666.880 430.240 674.320 430.560 ;
                RECT 0.160 431.600 77.640 431.920 ;
                RECT 95.680 431.600 106.200 431.920 ;
                RECT 666.880 431.600 674.320 431.920 ;
                RECT 0.160 432.960 77.640 433.280 ;
                RECT 95.680 432.960 106.200 433.280 ;
                RECT 666.880 432.960 674.320 433.280 ;
                RECT 0.160 434.320 106.200 434.640 ;
                RECT 666.880 434.320 674.320 434.640 ;
                RECT 0.160 435.680 77.640 436.000 ;
                RECT 95.680 435.680 106.200 436.000 ;
                RECT 666.880 435.680 674.320 436.000 ;
                RECT 0.160 437.040 77.640 437.360 ;
                RECT 95.680 437.040 106.200 437.360 ;
                RECT 666.880 437.040 674.320 437.360 ;
                RECT 0.160 438.400 77.640 438.720 ;
                RECT 95.680 438.400 106.200 438.720 ;
                RECT 666.880 438.400 674.320 438.720 ;
                RECT 0.160 439.760 77.640 440.080 ;
                RECT 95.680 439.760 106.200 440.080 ;
                RECT 666.880 439.760 674.320 440.080 ;
                RECT 0.160 441.120 77.640 441.440 ;
                RECT 86.160 441.120 106.200 441.440 ;
                RECT 666.880 441.120 674.320 441.440 ;
                RECT 0.160 442.480 91.920 442.800 ;
                RECT 95.680 442.480 106.200 442.800 ;
                RECT 666.880 442.480 674.320 442.800 ;
                RECT 0.160 443.840 77.640 444.160 ;
                RECT 95.680 443.840 106.200 444.160 ;
                RECT 666.880 443.840 674.320 444.160 ;
                RECT 0.160 445.200 77.640 445.520 ;
                RECT 95.680 445.200 106.200 445.520 ;
                RECT 666.880 445.200 674.320 445.520 ;
                RECT 0.160 446.560 77.640 446.880 ;
                RECT 95.680 446.560 106.200 446.880 ;
                RECT 666.880 446.560 674.320 446.880 ;
                RECT 0.160 447.920 77.640 448.240 ;
                RECT 95.680 447.920 106.200 448.240 ;
                RECT 666.880 447.920 674.320 448.240 ;
                RECT 0.160 449.280 77.640 449.600 ;
                RECT 86.840 449.280 106.200 449.600 ;
                RECT 666.880 449.280 674.320 449.600 ;
                RECT 0.160 450.640 77.640 450.960 ;
                RECT 95.680 450.640 106.200 450.960 ;
                RECT 666.880 450.640 674.320 450.960 ;
                RECT 0.160 452.000 77.640 452.320 ;
                RECT 95.680 452.000 106.200 452.320 ;
                RECT 666.880 452.000 674.320 452.320 ;
                RECT 0.160 453.360 77.640 453.680 ;
                RECT 95.680 453.360 106.200 453.680 ;
                RECT 666.880 453.360 674.320 453.680 ;
                RECT 0.160 454.720 77.640 455.040 ;
                RECT 95.680 454.720 106.200 455.040 ;
                RECT 666.880 454.720 674.320 455.040 ;
                RECT 0.160 456.080 77.640 456.400 ;
                RECT 95.680 456.080 106.200 456.400 ;
                RECT 666.880 456.080 674.320 456.400 ;
                RECT 0.160 457.440 106.200 457.760 ;
                RECT 666.880 457.440 674.320 457.760 ;
                RECT 0.160 458.800 81.040 459.120 ;
                RECT 95.680 458.800 106.200 459.120 ;
                RECT 666.880 458.800 674.320 459.120 ;
                RECT 0.160 460.160 81.040 460.480 ;
                RECT 95.680 460.160 106.200 460.480 ;
                RECT 666.880 460.160 674.320 460.480 ;
                RECT 0.160 461.520 88.520 461.840 ;
                RECT 95.680 461.520 106.200 461.840 ;
                RECT 666.880 461.520 674.320 461.840 ;
                RECT 0.160 462.880 81.040 463.200 ;
                RECT 95.680 462.880 106.200 463.200 ;
                RECT 666.880 462.880 674.320 463.200 ;
                RECT 0.160 464.240 81.040 464.560 ;
                RECT 95.680 464.240 106.200 464.560 ;
                RECT 666.880 464.240 674.320 464.560 ;
                RECT 0.160 465.600 106.200 465.920 ;
                RECT 666.880 465.600 674.320 465.920 ;
                RECT 0.160 466.960 81.040 467.280 ;
                RECT 95.680 466.960 106.200 467.280 ;
                RECT 666.880 466.960 674.320 467.280 ;
                RECT 0.160 468.320 81.040 468.640 ;
                RECT 95.680 468.320 106.200 468.640 ;
                RECT 666.880 468.320 674.320 468.640 ;
                RECT 0.160 469.680 81.040 470.000 ;
                RECT 95.680 469.680 106.200 470.000 ;
                RECT 666.880 469.680 674.320 470.000 ;
                RECT 0.160 471.040 91.240 471.360 ;
                RECT 95.680 471.040 106.200 471.360 ;
                RECT 666.880 471.040 674.320 471.360 ;
                RECT 0.160 472.400 81.040 472.720 ;
                RECT 95.680 472.400 106.200 472.720 ;
                RECT 666.880 472.400 674.320 472.720 ;
                RECT 0.160 473.760 106.200 474.080 ;
                RECT 666.880 473.760 674.320 474.080 ;
                RECT 0.160 475.120 81.040 475.440 ;
                RECT 95.680 475.120 106.200 475.440 ;
                RECT 666.880 475.120 674.320 475.440 ;
                RECT 0.160 476.480 81.040 476.800 ;
                RECT 95.680 476.480 106.200 476.800 ;
                RECT 666.880 476.480 674.320 476.800 ;
                RECT 0.160 477.840 81.040 478.160 ;
                RECT 95.680 477.840 106.200 478.160 ;
                RECT 666.880 477.840 674.320 478.160 ;
                RECT 0.160 479.200 81.040 479.520 ;
                RECT 95.680 479.200 106.200 479.520 ;
                RECT 666.880 479.200 674.320 479.520 ;
                RECT 0.160 480.560 106.200 480.880 ;
                RECT 666.880 480.560 674.320 480.880 ;
                RECT 0.160 481.920 85.800 482.240 ;
                RECT 95.680 481.920 106.200 482.240 ;
                RECT 666.880 481.920 674.320 482.240 ;
                RECT 0.160 483.280 81.720 483.600 ;
                RECT 95.680 483.280 106.200 483.600 ;
                RECT 666.880 483.280 674.320 483.600 ;
                RECT 0.160 484.640 81.720 484.960 ;
                RECT 95.680 484.640 106.200 484.960 ;
                RECT 666.880 484.640 674.320 484.960 ;
                RECT 0.160 486.000 81.720 486.320 ;
                RECT 95.680 486.000 106.200 486.320 ;
                RECT 666.880 486.000 674.320 486.320 ;
                RECT 0.160 487.360 81.720 487.680 ;
                RECT 95.680 487.360 106.200 487.680 ;
                RECT 666.880 487.360 674.320 487.680 ;
                RECT 0.160 488.720 106.200 489.040 ;
                RECT 666.880 488.720 674.320 489.040 ;
                RECT 0.160 490.080 87.840 490.400 ;
                RECT 95.680 490.080 106.200 490.400 ;
                RECT 666.880 490.080 674.320 490.400 ;
                RECT 0.160 491.440 81.720 491.760 ;
                RECT 95.680 491.440 106.200 491.760 ;
                RECT 666.880 491.440 674.320 491.760 ;
                RECT 0.160 492.800 81.720 493.120 ;
                RECT 95.680 492.800 106.200 493.120 ;
                RECT 666.880 492.800 674.320 493.120 ;
                RECT 0.160 494.160 81.720 494.480 ;
                RECT 95.680 494.160 106.200 494.480 ;
                RECT 666.880 494.160 674.320 494.480 ;
                RECT 0.160 495.520 81.720 495.840 ;
                RECT 95.680 495.520 106.200 495.840 ;
                RECT 666.880 495.520 674.320 495.840 ;
                RECT 0.160 496.880 106.200 497.200 ;
                RECT 666.880 496.880 674.320 497.200 ;
                RECT 0.160 498.240 81.720 498.560 ;
                RECT 95.680 498.240 106.200 498.560 ;
                RECT 666.880 498.240 674.320 498.560 ;
                RECT 0.160 499.600 90.560 499.920 ;
                RECT 95.680 499.600 106.200 499.920 ;
                RECT 666.880 499.600 674.320 499.920 ;
                RECT 0.160 500.960 90.560 501.280 ;
                RECT 95.680 500.960 106.200 501.280 ;
                RECT 666.880 500.960 674.320 501.280 ;
                RECT 0.160 502.320 81.720 502.640 ;
                RECT 95.680 502.320 106.200 502.640 ;
                RECT 666.880 502.320 674.320 502.640 ;
                RECT 0.160 503.680 81.720 504.000 ;
                RECT 95.680 503.680 106.200 504.000 ;
                RECT 666.880 503.680 674.320 504.000 ;
                RECT 0.160 505.040 106.200 505.360 ;
                RECT 666.880 505.040 674.320 505.360 ;
                RECT 0.160 506.400 81.720 506.720 ;
                RECT 95.680 506.400 106.200 506.720 ;
                RECT 666.880 506.400 674.320 506.720 ;
                RECT 0.160 507.760 81.720 508.080 ;
                RECT 95.680 507.760 106.200 508.080 ;
                RECT 666.880 507.760 674.320 508.080 ;
                RECT 0.160 509.120 92.600 509.440 ;
                RECT 95.680 509.120 106.200 509.440 ;
                RECT 666.880 509.120 674.320 509.440 ;
                RECT 0.160 510.480 93.280 510.800 ;
                RECT 95.680 510.480 106.200 510.800 ;
                RECT 666.880 510.480 674.320 510.800 ;
                RECT 0.160 511.840 81.720 512.160 ;
                RECT 95.680 511.840 106.200 512.160 ;
                RECT 666.880 511.840 674.320 512.160 ;
                RECT 0.160 513.200 106.200 513.520 ;
                RECT 666.880 513.200 674.320 513.520 ;
                RECT 0.160 514.560 82.400 514.880 ;
                RECT 95.680 514.560 106.200 514.880 ;
                RECT 666.880 514.560 674.320 514.880 ;
                RECT 0.160 515.920 82.400 516.240 ;
                RECT 95.680 515.920 106.200 516.240 ;
                RECT 666.880 515.920 674.320 516.240 ;
                RECT 0.160 517.280 82.400 517.600 ;
                RECT 95.680 517.280 106.200 517.600 ;
                RECT 666.880 517.280 674.320 517.600 ;
                RECT 0.160 518.640 82.400 518.960 ;
                RECT 95.680 518.640 106.200 518.960 ;
                RECT 666.880 518.640 674.320 518.960 ;
                RECT 0.160 520.000 106.200 520.320 ;
                RECT 666.880 520.000 674.320 520.320 ;
                RECT 0.160 521.360 87.840 521.680 ;
                RECT 95.680 521.360 106.200 521.680 ;
                RECT 666.880 521.360 674.320 521.680 ;
                RECT 0.160 522.720 82.400 523.040 ;
                RECT 95.680 522.720 106.200 523.040 ;
                RECT 666.880 522.720 674.320 523.040 ;
                RECT 0.160 524.080 82.400 524.400 ;
                RECT 95.680 524.080 106.200 524.400 ;
                RECT 666.880 524.080 674.320 524.400 ;
                RECT 0.160 525.440 82.400 525.760 ;
                RECT 95.680 525.440 106.200 525.760 ;
                RECT 666.880 525.440 674.320 525.760 ;
                RECT 0.160 526.800 82.400 527.120 ;
                RECT 95.680 526.800 106.200 527.120 ;
                RECT 666.880 526.800 674.320 527.120 ;
                RECT 0.160 528.160 106.200 528.480 ;
                RECT 666.880 528.160 674.320 528.480 ;
                RECT 0.160 529.520 89.880 529.840 ;
                RECT 95.680 529.520 106.200 529.840 ;
                RECT 666.880 529.520 674.320 529.840 ;
                RECT 0.160 530.880 82.400 531.200 ;
                RECT 95.680 530.880 106.200 531.200 ;
                RECT 666.880 530.880 674.320 531.200 ;
                RECT 0.160 532.240 82.400 532.560 ;
                RECT 95.680 532.240 106.200 532.560 ;
                RECT 666.880 532.240 674.320 532.560 ;
                RECT 0.160 533.600 82.400 533.920 ;
                RECT 95.680 533.600 106.200 533.920 ;
                RECT 666.880 533.600 674.320 533.920 ;
                RECT 0.160 534.960 82.400 535.280 ;
                RECT 95.680 534.960 106.200 535.280 ;
                RECT 666.880 534.960 674.320 535.280 ;
                RECT 0.160 536.320 106.200 536.640 ;
                RECT 666.880 536.320 674.320 536.640 ;
                RECT 0.160 537.680 82.400 538.000 ;
                RECT 95.680 537.680 106.200 538.000 ;
                RECT 666.880 537.680 674.320 538.000 ;
                RECT 0.160 539.040 91.920 539.360 ;
                RECT 95.680 539.040 106.200 539.360 ;
                RECT 666.880 539.040 674.320 539.360 ;
                RECT 0.160 540.400 82.400 540.720 ;
                RECT 95.680 540.400 106.200 540.720 ;
                RECT 666.880 540.400 674.320 540.720 ;
                RECT 0.160 541.760 82.400 542.080 ;
                RECT 95.680 541.760 106.200 542.080 ;
                RECT 666.880 541.760 674.320 542.080 ;
                RECT 0.160 543.120 82.400 543.440 ;
                RECT 95.680 543.120 106.200 543.440 ;
                RECT 666.880 543.120 674.320 543.440 ;
                RECT 0.160 544.480 106.200 544.800 ;
                RECT 666.880 544.480 674.320 544.800 ;
                RECT 0.160 545.840 82.400 546.160 ;
                RECT 95.680 545.840 106.200 546.160 ;
                RECT 666.880 545.840 674.320 546.160 ;
                RECT 0.160 547.200 82.400 547.520 ;
                RECT 95.680 547.200 106.200 547.520 ;
                RECT 666.880 547.200 674.320 547.520 ;
                RECT 0.160 548.560 87.160 548.880 ;
                RECT 95.680 548.560 106.200 548.880 ;
                RECT 666.880 548.560 674.320 548.880 ;
                RECT 0.160 549.920 82.400 550.240 ;
                RECT 95.680 549.920 106.200 550.240 ;
                RECT 666.880 549.920 674.320 550.240 ;
                RECT 0.160 551.280 82.400 551.600 ;
                RECT 95.680 551.280 106.200 551.600 ;
                RECT 666.880 551.280 674.320 551.600 ;
                RECT 0.160 552.640 106.200 552.960 ;
                RECT 666.880 552.640 674.320 552.960 ;
                RECT 0.160 554.000 82.400 554.320 ;
                RECT 95.680 554.000 106.200 554.320 ;
                RECT 666.880 554.000 674.320 554.320 ;
                RECT 0.160 555.360 82.400 555.680 ;
                RECT 95.680 555.360 106.200 555.680 ;
                RECT 666.880 555.360 674.320 555.680 ;
                RECT 0.160 556.720 82.400 557.040 ;
                RECT 95.680 556.720 106.200 557.040 ;
                RECT 666.880 556.720 674.320 557.040 ;
                RECT 0.160 558.080 89.200 558.400 ;
                RECT 95.680 558.080 106.200 558.400 ;
                RECT 666.880 558.080 674.320 558.400 ;
                RECT 0.160 559.440 106.200 559.760 ;
                RECT 666.880 559.440 674.320 559.760 ;
                RECT 0.160 560.800 89.880 561.120 ;
                RECT 95.680 560.800 106.200 561.120 ;
                RECT 666.880 560.800 674.320 561.120 ;
                RECT 0.160 562.160 82.400 562.480 ;
                RECT 95.680 562.160 106.200 562.480 ;
                RECT 666.880 562.160 674.320 562.480 ;
                RECT 0.160 563.520 82.400 563.840 ;
                RECT 95.680 563.520 106.200 563.840 ;
                RECT 666.880 563.520 674.320 563.840 ;
                RECT 0.160 564.880 82.400 565.200 ;
                RECT 95.680 564.880 106.200 565.200 ;
                RECT 666.880 564.880 674.320 565.200 ;
                RECT 0.160 566.240 82.400 566.560 ;
                RECT 95.680 566.240 106.200 566.560 ;
                RECT 666.880 566.240 674.320 566.560 ;
                RECT 0.160 567.600 106.200 567.920 ;
                RECT 666.880 567.600 674.320 567.920 ;
                RECT 0.160 568.960 91.920 569.280 ;
                RECT 95.680 568.960 106.200 569.280 ;
                RECT 666.880 568.960 674.320 569.280 ;
                RECT 0.160 570.320 82.400 570.640 ;
                RECT 95.680 570.320 106.200 570.640 ;
                RECT 666.880 570.320 674.320 570.640 ;
                RECT 0.160 571.680 82.400 572.000 ;
                RECT 95.680 571.680 106.200 572.000 ;
                RECT 666.880 571.680 674.320 572.000 ;
                RECT 0.160 573.040 82.400 573.360 ;
                RECT 95.680 573.040 106.200 573.360 ;
                RECT 666.880 573.040 674.320 573.360 ;
                RECT 0.160 574.400 82.400 574.720 ;
                RECT 95.680 574.400 106.200 574.720 ;
                RECT 666.880 574.400 674.320 574.720 ;
                RECT 0.160 575.760 106.200 576.080 ;
                RECT 666.880 575.760 674.320 576.080 ;
                RECT 0.160 577.120 83.080 577.440 ;
                RECT 95.680 577.120 106.200 577.440 ;
                RECT 666.880 577.120 674.320 577.440 ;
                RECT 0.160 578.480 86.480 578.800 ;
                RECT 95.680 578.480 106.200 578.800 ;
                RECT 666.880 578.480 674.320 578.800 ;
                RECT 0.160 579.840 83.080 580.160 ;
                RECT 95.680 579.840 106.200 580.160 ;
                RECT 666.880 579.840 674.320 580.160 ;
                RECT 0.160 581.200 83.080 581.520 ;
                RECT 95.680 581.200 106.200 581.520 ;
                RECT 666.880 581.200 674.320 581.520 ;
                RECT 0.160 582.560 83.080 582.880 ;
                RECT 95.680 582.560 106.200 582.880 ;
                RECT 666.880 582.560 674.320 582.880 ;
                RECT 0.160 583.920 106.200 584.240 ;
                RECT 666.880 583.920 674.320 584.240 ;
                RECT 0.160 585.280 83.080 585.600 ;
                RECT 95.680 585.280 106.200 585.600 ;
                RECT 666.880 585.280 674.320 585.600 ;
                RECT 0.160 586.640 83.080 586.960 ;
                RECT 95.680 586.640 106.200 586.960 ;
                RECT 666.880 586.640 674.320 586.960 ;
                RECT 0.160 588.000 88.520 588.320 ;
                RECT 95.680 588.000 106.200 588.320 ;
                RECT 666.880 588.000 674.320 588.320 ;
                RECT 0.160 589.360 83.080 589.680 ;
                RECT 95.680 589.360 106.200 589.680 ;
                RECT 666.880 589.360 674.320 589.680 ;
                RECT 0.160 590.720 83.080 591.040 ;
                RECT 95.680 590.720 106.200 591.040 ;
                RECT 666.880 590.720 674.320 591.040 ;
                RECT 0.160 592.080 106.200 592.400 ;
                RECT 666.880 592.080 674.320 592.400 ;
                RECT 0.160 593.440 83.080 593.760 ;
                RECT 95.680 593.440 106.200 593.760 ;
                RECT 666.880 593.440 674.320 593.760 ;
                RECT 0.160 594.800 83.080 595.120 ;
                RECT 95.680 594.800 106.200 595.120 ;
                RECT 666.880 594.800 674.320 595.120 ;
                RECT 0.160 596.160 83.080 596.480 ;
                RECT 95.680 596.160 106.200 596.480 ;
                RECT 666.880 596.160 674.320 596.480 ;
                RECT 0.160 597.520 91.240 597.840 ;
                RECT 95.680 597.520 106.200 597.840 ;
                RECT 666.880 597.520 674.320 597.840 ;
                RECT 0.160 598.880 83.080 599.200 ;
                RECT 95.680 598.880 106.200 599.200 ;
                RECT 666.880 598.880 674.320 599.200 ;
                RECT 0.160 600.240 106.200 600.560 ;
                RECT 666.880 600.240 674.320 600.560 ;
                RECT 0.160 601.600 83.080 601.920 ;
                RECT 95.680 601.600 106.200 601.920 ;
                RECT 666.880 601.600 674.320 601.920 ;
                RECT 0.160 602.960 83.080 603.280 ;
                RECT 95.680 602.960 106.200 603.280 ;
                RECT 666.880 602.960 674.320 603.280 ;
                RECT 0.160 604.320 83.080 604.640 ;
                RECT 95.680 604.320 106.200 604.640 ;
                RECT 666.880 604.320 674.320 604.640 ;
                RECT 0.160 605.680 83.080 606.000 ;
                RECT 95.680 605.680 106.200 606.000 ;
                RECT 666.880 605.680 674.320 606.000 ;
                RECT 0.160 607.040 106.200 607.360 ;
                RECT 666.880 607.040 674.320 607.360 ;
                RECT 0.160 608.400 85.800 608.720 ;
                RECT 95.680 608.400 106.200 608.720 ;
                RECT 666.880 608.400 674.320 608.720 ;
                RECT 0.160 609.760 83.760 610.080 ;
                RECT 95.680 609.760 106.200 610.080 ;
                RECT 666.880 609.760 674.320 610.080 ;
                RECT 0.160 611.120 83.760 611.440 ;
                RECT 95.680 611.120 106.200 611.440 ;
                RECT 666.880 611.120 674.320 611.440 ;
                RECT 0.160 612.480 83.760 612.800 ;
                RECT 95.680 612.480 106.200 612.800 ;
                RECT 666.880 612.480 674.320 612.800 ;
                RECT 0.160 613.840 83.760 614.160 ;
                RECT 95.680 613.840 106.200 614.160 ;
                RECT 666.880 613.840 674.320 614.160 ;
                RECT 0.160 615.200 106.200 615.520 ;
                RECT 666.880 615.200 674.320 615.520 ;
                RECT 0.160 616.560 87.840 616.880 ;
                RECT 95.680 616.560 106.200 616.880 ;
                RECT 666.880 616.560 674.320 616.880 ;
                RECT 0.160 617.920 88.520 618.240 ;
                RECT 95.680 617.920 106.200 618.240 ;
                RECT 666.880 617.920 674.320 618.240 ;
                RECT 0.160 619.280 83.760 619.600 ;
                RECT 95.680 619.280 106.200 619.600 ;
                RECT 666.880 619.280 674.320 619.600 ;
                RECT 0.160 620.640 83.760 620.960 ;
                RECT 95.680 620.640 106.200 620.960 ;
                RECT 666.880 620.640 674.320 620.960 ;
                RECT 0.160 622.000 83.760 622.320 ;
                RECT 95.680 622.000 106.200 622.320 ;
                RECT 666.880 622.000 674.320 622.320 ;
                RECT 0.160 623.360 106.200 623.680 ;
                RECT 666.880 623.360 674.320 623.680 ;
                RECT 0.160 624.720 83.760 625.040 ;
                RECT 95.680 624.720 106.200 625.040 ;
                RECT 666.880 624.720 674.320 625.040 ;
                RECT 0.160 626.080 83.760 626.400 ;
                RECT 95.680 626.080 106.200 626.400 ;
                RECT 666.880 626.080 674.320 626.400 ;
                RECT 0.160 627.440 90.560 627.760 ;
                RECT 95.680 627.440 106.200 627.760 ;
                RECT 666.880 627.440 674.320 627.760 ;
                RECT 0.160 628.800 83.760 629.120 ;
                RECT 95.680 628.800 106.200 629.120 ;
                RECT 666.880 628.800 674.320 629.120 ;
                RECT 0.160 630.160 83.760 630.480 ;
                RECT 95.680 630.160 106.200 630.480 ;
                RECT 666.880 630.160 674.320 630.480 ;
                RECT 0.160 631.520 106.200 631.840 ;
                RECT 666.880 631.520 674.320 631.840 ;
                RECT 0.160 632.880 83.760 633.200 ;
                RECT 95.680 632.880 106.200 633.200 ;
                RECT 666.880 632.880 674.320 633.200 ;
                RECT 0.160 634.240 83.760 634.560 ;
                RECT 95.680 634.240 106.200 634.560 ;
                RECT 666.880 634.240 674.320 634.560 ;
                RECT 0.160 635.600 83.760 635.920 ;
                RECT 95.680 635.600 106.200 635.920 ;
                RECT 666.880 635.600 674.320 635.920 ;
                RECT 0.160 636.960 93.280 637.280 ;
                RECT 95.680 636.960 106.200 637.280 ;
                RECT 666.880 636.960 674.320 637.280 ;
                RECT 0.160 638.320 83.760 638.640 ;
                RECT 95.680 638.320 106.200 638.640 ;
                RECT 666.880 638.320 674.320 638.640 ;
                RECT 0.160 639.680 106.200 640.000 ;
                RECT 666.880 639.680 674.320 640.000 ;
                RECT 0.160 641.040 83.760 641.360 ;
                RECT 95.680 641.040 106.200 641.360 ;
                RECT 666.880 641.040 674.320 641.360 ;
                RECT 0.160 642.400 83.760 642.720 ;
                RECT 95.680 642.400 106.200 642.720 ;
                RECT 666.880 642.400 674.320 642.720 ;
                RECT 0.160 643.760 83.760 644.080 ;
                RECT 95.680 643.760 106.200 644.080 ;
                RECT 666.880 643.760 674.320 644.080 ;
                RECT 0.160 645.120 83.760 645.440 ;
                RECT 95.680 645.120 106.200 645.440 ;
                RECT 666.880 645.120 674.320 645.440 ;
                RECT 0.160 646.480 106.200 646.800 ;
                RECT 666.880 646.480 674.320 646.800 ;
                RECT 0.160 647.840 87.840 648.160 ;
                RECT 95.680 647.840 106.200 648.160 ;
                RECT 666.880 647.840 674.320 648.160 ;
                RECT 0.160 649.200 83.760 649.520 ;
                RECT 95.680 649.200 106.200 649.520 ;
                RECT 666.880 649.200 674.320 649.520 ;
                RECT 0.160 650.560 83.760 650.880 ;
                RECT 95.680 650.560 106.200 650.880 ;
                RECT 666.880 650.560 674.320 650.880 ;
                RECT 0.160 651.920 83.760 652.240 ;
                RECT 95.680 651.920 106.200 652.240 ;
                RECT 666.880 651.920 674.320 652.240 ;
                RECT 0.160 653.280 83.760 653.600 ;
                RECT 95.680 653.280 106.200 653.600 ;
                RECT 666.880 653.280 674.320 653.600 ;
                RECT 0.160 654.640 106.200 654.960 ;
                RECT 666.880 654.640 674.320 654.960 ;
                RECT 0.160 656.000 89.880 656.320 ;
                RECT 95.680 656.000 106.200 656.320 ;
                RECT 666.880 656.000 674.320 656.320 ;
                RECT 0.160 657.360 83.760 657.680 ;
                RECT 95.680 657.360 106.200 657.680 ;
                RECT 666.880 657.360 674.320 657.680 ;
                RECT 0.160 658.720 83.760 659.040 ;
                RECT 95.680 658.720 106.200 659.040 ;
                RECT 666.880 658.720 674.320 659.040 ;
                RECT 0.160 660.080 83.760 660.400 ;
                RECT 95.680 660.080 106.200 660.400 ;
                RECT 666.880 660.080 674.320 660.400 ;
                RECT 0.160 661.440 83.760 661.760 ;
                RECT 95.680 661.440 106.200 661.760 ;
                RECT 666.880 661.440 674.320 661.760 ;
                RECT 0.160 662.800 106.200 663.120 ;
                RECT 666.880 662.800 674.320 663.120 ;
                RECT 0.160 664.160 83.760 664.480 ;
                RECT 95.680 664.160 106.200 664.480 ;
                RECT 666.880 664.160 674.320 664.480 ;
                RECT 0.160 665.520 91.920 665.840 ;
                RECT 95.680 665.520 106.200 665.840 ;
                RECT 666.880 665.520 674.320 665.840 ;
                RECT 0.160 666.880 92.600 667.200 ;
                RECT 95.680 666.880 106.200 667.200 ;
                RECT 666.880 666.880 674.320 667.200 ;
                RECT 0.160 668.240 83.760 668.560 ;
                RECT 95.680 668.240 106.200 668.560 ;
                RECT 666.880 668.240 674.320 668.560 ;
                RECT 0.160 669.600 83.760 669.920 ;
                RECT 95.680 669.600 106.200 669.920 ;
                RECT 666.880 669.600 674.320 669.920 ;
                RECT 0.160 670.960 106.200 671.280 ;
                RECT 666.880 670.960 674.320 671.280 ;
                RECT 0.160 672.320 84.440 672.640 ;
                RECT 95.680 672.320 106.200 672.640 ;
                RECT 666.880 672.320 674.320 672.640 ;
                RECT 0.160 673.680 84.440 674.000 ;
                RECT 95.680 673.680 106.200 674.000 ;
                RECT 666.880 673.680 674.320 674.000 ;
                RECT 0.160 675.040 84.440 675.360 ;
                RECT 95.680 675.040 106.200 675.360 ;
                RECT 666.880 675.040 674.320 675.360 ;
                RECT 0.160 676.400 87.160 676.720 ;
                RECT 95.680 676.400 106.200 676.720 ;
                RECT 666.880 676.400 674.320 676.720 ;
                RECT 0.160 677.760 84.440 678.080 ;
                RECT 95.680 677.760 106.200 678.080 ;
                RECT 666.880 677.760 674.320 678.080 ;
                RECT 0.160 679.120 106.200 679.440 ;
                RECT 666.880 679.120 674.320 679.440 ;
                RECT 0.160 680.480 84.440 680.800 ;
                RECT 95.680 680.480 106.200 680.800 ;
                RECT 666.880 680.480 674.320 680.800 ;
                RECT 0.160 681.840 84.440 682.160 ;
                RECT 95.680 681.840 106.200 682.160 ;
                RECT 666.880 681.840 674.320 682.160 ;
                RECT 0.160 683.200 84.440 683.520 ;
                RECT 95.680 683.200 106.200 683.520 ;
                RECT 666.880 683.200 674.320 683.520 ;
                RECT 0.160 684.560 84.440 684.880 ;
                RECT 95.680 684.560 106.200 684.880 ;
                RECT 666.880 684.560 674.320 684.880 ;
                RECT 0.160 685.920 106.200 686.240 ;
                RECT 666.880 685.920 674.320 686.240 ;
                RECT 0.160 687.280 89.880 687.600 ;
                RECT 95.680 687.280 106.200 687.600 ;
                RECT 666.880 687.280 674.320 687.600 ;
                RECT 0.160 688.640 84.440 688.960 ;
                RECT 95.680 688.640 106.200 688.960 ;
                RECT 666.880 688.640 674.320 688.960 ;
                RECT 0.160 690.000 84.440 690.320 ;
                RECT 95.680 690.000 106.200 690.320 ;
                RECT 666.880 690.000 674.320 690.320 ;
                RECT 0.160 691.360 84.440 691.680 ;
                RECT 95.680 691.360 106.200 691.680 ;
                RECT 666.880 691.360 674.320 691.680 ;
                RECT 0.160 692.720 84.440 693.040 ;
                RECT 95.680 692.720 106.200 693.040 ;
                RECT 666.880 692.720 674.320 693.040 ;
                RECT 0.160 694.080 106.200 694.400 ;
                RECT 666.880 694.080 674.320 694.400 ;
                RECT 0.160 695.440 91.920 695.760 ;
                RECT 95.680 695.440 106.200 695.760 ;
                RECT 666.880 695.440 674.320 695.760 ;
                RECT 0.160 696.800 84.440 697.120 ;
                RECT 95.680 696.800 106.200 697.120 ;
                RECT 666.880 696.800 674.320 697.120 ;
                RECT 0.160 698.160 84.440 698.480 ;
                RECT 95.680 698.160 106.200 698.480 ;
                RECT 666.880 698.160 674.320 698.480 ;
                RECT 0.160 699.520 84.440 699.840 ;
                RECT 95.680 699.520 106.200 699.840 ;
                RECT 666.880 699.520 674.320 699.840 ;
                RECT 0.160 700.880 84.440 701.200 ;
                RECT 95.680 700.880 106.200 701.200 ;
                RECT 666.880 700.880 674.320 701.200 ;
                RECT 0.160 702.240 106.200 702.560 ;
                RECT 666.880 702.240 674.320 702.560 ;
                RECT 0.160 703.600 85.120 703.920 ;
                RECT 95.680 703.600 106.200 703.920 ;
                RECT 666.880 703.600 674.320 703.920 ;
                RECT 0.160 704.960 86.480 705.280 ;
                RECT 95.680 704.960 106.200 705.280 ;
                RECT 666.880 704.960 674.320 705.280 ;
                RECT 0.160 706.320 85.120 706.640 ;
                RECT 95.680 706.320 106.200 706.640 ;
                RECT 666.880 706.320 674.320 706.640 ;
                RECT 0.160 707.680 85.120 708.000 ;
                RECT 95.680 707.680 106.200 708.000 ;
                RECT 666.880 707.680 674.320 708.000 ;
                RECT 0.160 709.040 85.120 709.360 ;
                RECT 95.680 709.040 106.200 709.360 ;
                RECT 666.880 709.040 674.320 709.360 ;
                RECT 0.160 710.400 106.200 710.720 ;
                RECT 666.880 710.400 674.320 710.720 ;
                RECT 0.160 711.760 85.120 712.080 ;
                RECT 95.680 711.760 106.200 712.080 ;
                RECT 666.880 711.760 674.320 712.080 ;
                RECT 0.160 713.120 85.120 713.440 ;
                RECT 95.680 713.120 106.200 713.440 ;
                RECT 666.880 713.120 674.320 713.440 ;
                RECT 0.160 714.480 88.520 714.800 ;
                RECT 95.680 714.480 106.200 714.800 ;
                RECT 666.880 714.480 674.320 714.800 ;
                RECT 0.160 715.840 89.200 716.160 ;
                RECT 95.680 715.840 106.200 716.160 ;
                RECT 666.880 715.840 674.320 716.160 ;
                RECT 0.160 717.200 85.120 717.520 ;
                RECT 95.680 717.200 106.200 717.520 ;
                RECT 666.880 717.200 674.320 717.520 ;
                RECT 0.160 718.560 106.200 718.880 ;
                RECT 666.880 718.560 674.320 718.880 ;
                RECT 0.160 719.920 85.120 720.240 ;
                RECT 95.680 719.920 106.200 720.240 ;
                RECT 666.880 719.920 674.320 720.240 ;
                RECT 0.160 721.280 85.120 721.600 ;
                RECT 95.680 721.280 106.200 721.600 ;
                RECT 666.880 721.280 674.320 721.600 ;
                RECT 0.160 722.640 85.120 722.960 ;
                RECT 95.680 722.640 106.200 722.960 ;
                RECT 666.880 722.640 674.320 722.960 ;
                RECT 0.160 724.000 91.240 724.320 ;
                RECT 95.680 724.000 106.200 724.320 ;
                RECT 666.880 724.000 674.320 724.320 ;
                RECT 0.160 725.360 106.200 725.680 ;
                RECT 666.880 725.360 674.320 725.680 ;
                RECT 0.160 726.720 91.920 727.040 ;
                RECT 95.680 726.720 106.200 727.040 ;
                RECT 666.880 726.720 674.320 727.040 ;
                RECT 0.160 728.080 85.120 728.400 ;
                RECT 95.680 728.080 106.200 728.400 ;
                RECT 666.880 728.080 674.320 728.400 ;
                RECT 0.160 729.440 85.120 729.760 ;
                RECT 95.680 729.440 106.200 729.760 ;
                RECT 666.880 729.440 674.320 729.760 ;
                RECT 0.160 730.800 85.120 731.120 ;
                RECT 95.680 730.800 106.200 731.120 ;
                RECT 666.880 730.800 674.320 731.120 ;
                RECT 0.160 732.160 85.120 732.480 ;
                RECT 95.680 732.160 106.200 732.480 ;
                RECT 666.880 732.160 674.320 732.480 ;
                RECT 0.160 733.520 106.200 733.840 ;
                RECT 666.880 733.520 674.320 733.840 ;
                RECT 0.160 734.880 85.800 735.200 ;
                RECT 95.680 734.880 106.200 735.200 ;
                RECT 666.880 734.880 674.320 735.200 ;
                RECT 0.160 736.240 85.800 736.560 ;
                RECT 95.680 736.240 106.200 736.560 ;
                RECT 666.880 736.240 674.320 736.560 ;
                RECT 0.160 737.600 85.800 737.920 ;
                RECT 95.680 737.600 106.200 737.920 ;
                RECT 666.880 737.600 674.320 737.920 ;
                RECT 0.160 738.960 85.800 739.280 ;
                RECT 95.680 738.960 106.200 739.280 ;
                RECT 666.880 738.960 674.320 739.280 ;
                RECT 0.160 740.320 85.800 740.640 ;
                RECT 95.680 740.320 106.200 740.640 ;
                RECT 666.880 740.320 674.320 740.640 ;
                RECT 0.160 741.680 106.200 742.000 ;
                RECT 666.880 741.680 674.320 742.000 ;
                RECT 0.160 743.040 85.800 743.360 ;
                RECT 95.680 743.040 106.200 743.360 ;
                RECT 666.880 743.040 674.320 743.360 ;
                RECT 0.160 744.400 88.520 744.720 ;
                RECT 95.680 744.400 106.200 744.720 ;
                RECT 666.880 744.400 674.320 744.720 ;
                RECT 0.160 745.760 85.800 746.080 ;
                RECT 95.680 745.760 106.200 746.080 ;
                RECT 666.880 745.760 674.320 746.080 ;
                RECT 0.160 747.120 85.800 747.440 ;
                RECT 95.680 747.120 106.200 747.440 ;
                RECT 666.880 747.120 674.320 747.440 ;
                RECT 0.160 748.480 85.800 748.800 ;
                RECT 95.680 748.480 106.200 748.800 ;
                RECT 666.880 748.480 674.320 748.800 ;
                RECT 0.160 749.840 106.200 750.160 ;
                RECT 666.880 749.840 674.320 750.160 ;
                RECT 0.160 751.200 85.800 751.520 ;
                RECT 95.680 751.200 106.200 751.520 ;
                RECT 666.880 751.200 674.320 751.520 ;
                RECT 0.160 752.560 85.800 752.880 ;
                RECT 95.680 752.560 106.200 752.880 ;
                RECT 666.880 752.560 674.320 752.880 ;
                RECT 0.160 753.920 90.560 754.240 ;
                RECT 95.680 753.920 106.200 754.240 ;
                RECT 666.880 753.920 674.320 754.240 ;
                RECT 0.160 755.280 85.800 755.600 ;
                RECT 95.680 755.280 106.200 755.600 ;
                RECT 666.880 755.280 674.320 755.600 ;
                RECT 0.160 756.640 85.800 756.960 ;
                RECT 95.680 756.640 106.200 756.960 ;
                RECT 666.880 756.640 674.320 756.960 ;
                RECT 0.160 758.000 106.200 758.320 ;
                RECT 666.880 758.000 674.320 758.320 ;
                RECT 0.160 759.360 85.800 759.680 ;
                RECT 95.680 759.360 106.200 759.680 ;
                RECT 666.880 759.360 674.320 759.680 ;
                RECT 0.160 760.720 85.800 761.040 ;
                RECT 95.680 760.720 106.200 761.040 ;
                RECT 666.880 760.720 674.320 761.040 ;
                RECT 0.160 762.080 85.800 762.400 ;
                RECT 95.680 762.080 106.200 762.400 ;
                RECT 666.880 762.080 674.320 762.400 ;
                RECT 0.160 763.440 93.280 763.760 ;
                RECT 95.680 763.440 106.200 763.760 ;
                RECT 666.880 763.440 674.320 763.760 ;
                RECT 0.160 764.800 85.800 765.120 ;
                RECT 95.680 764.800 106.200 765.120 ;
                RECT 666.880 764.800 674.320 765.120 ;
                RECT 0.160 766.160 106.200 766.480 ;
                RECT 666.880 766.160 674.320 766.480 ;
                RECT 0.160 767.520 298.640 767.840 ;
                RECT 666.880 767.520 674.320 767.840 ;
                RECT 0.160 768.880 298.640 769.200 ;
                RECT 666.880 768.880 674.320 769.200 ;
                RECT 0.160 770.240 298.640 770.560 ;
                RECT 666.880 770.240 674.320 770.560 ;
                RECT 0.160 771.600 674.320 771.920 ;
                RECT 0.160 772.960 674.320 773.280 ;
                RECT 0.160 774.320 674.320 774.640 ;
                RECT 0.160 775.680 674.320 776.000 ;
                RECT 0.160 0.160 674.320 1.520 ;
                RECT 0.160 780.400 674.320 781.760 ;
                RECT 302.780 50.590 308.580 51.960 ;
                RECT 657.080 50.590 662.880 51.960 ;
                RECT 302.780 55.845 308.580 57.395 ;
                RECT 657.080 55.845 662.880 57.395 ;
                RECT 302.780 61.700 308.580 63.500 ;
                RECT 657.080 61.700 662.880 63.500 ;
                RECT 302.780 67.230 308.580 68.480 ;
                RECT 657.080 67.230 662.880 68.480 ;
                RECT 302.780 71.990 308.580 73.280 ;
                RECT 657.080 71.990 662.880 73.280 ;
                RECT 302.780 76.810 308.580 78.100 ;
                RECT 657.080 76.810 662.880 78.100 ;
                RECT 302.780 121.930 662.880 125.530 ;
                RECT 302.780 99.240 662.880 100.040 ;
                RECT 302.780 170.625 662.880 172.425 ;
                RECT 302.780 96.230 662.880 97.030 ;
                RECT 302.780 84.760 662.880 86.560 ;
                RECT 302.780 104.130 662.880 104.930 ;
                RECT 302.780 235.165 662.880 238.765 ;
                RECT 302.780 131.735 662.880 132.025 ;
                RECT 302.780 34.835 662.880 36.635 ;
                RECT 110.570 259.275 112.490 766.455 ;
                RECT 114.410 259.275 116.330 766.455 ;
                RECT 126.605 259.275 128.525 766.455 ;
                RECT 130.445 259.275 132.365 766.455 ;
                RECT 134.285 259.275 136.205 766.455 ;
                RECT 138.125 259.275 140.045 766.455 ;
                RECT 159.440 259.275 161.360 766.455 ;
                RECT 163.280 259.275 165.200 766.455 ;
                RECT 167.120 259.275 169.040 766.455 ;
                RECT 170.960 259.275 172.880 766.455 ;
                RECT 174.800 259.275 176.720 766.455 ;
                RECT 178.640 259.275 180.560 766.455 ;
                RECT 182.480 259.275 184.400 766.455 ;
                RECT 186.320 259.275 188.240 766.455 ;
                RECT 224.845 259.275 226.765 766.455 ;
                RECT 228.685 259.275 230.605 766.455 ;
                RECT 232.525 259.275 234.445 766.455 ;
                RECT 236.365 259.275 238.285 766.455 ;
                RECT 240.205 259.275 242.125 766.455 ;
                RECT 244.045 259.275 245.965 766.455 ;
                RECT 247.885 259.275 249.805 766.455 ;
                RECT 251.725 259.275 253.645 766.455 ;
                RECT 255.565 259.275 257.485 766.455 ;
                RECT 259.405 259.275 261.325 766.455 ;
                RECT 263.245 259.275 265.165 766.455 ;
                RECT 267.085 259.275 269.005 766.455 ;
                RECT 270.925 259.275 272.845 766.455 ;
                RECT 274.765 259.275 276.685 766.455 ;
                RECT 278.605 259.275 280.525 766.455 ;
                RECT 282.445 259.275 284.365 766.455 ;
                RECT 286.285 259.275 288.205 766.455 ;
                RECT 290.125 259.275 292.045 766.455 ;
                RECT 293.965 259.275 295.885 766.455 ;
                RECT 175.050 55.735 176.970 142.735 ;
                RECT 182.025 55.735 183.945 142.735 ;
                RECT 190.720 55.735 192.640 142.735 ;
                RECT 204.390 55.735 206.310 142.735 ;
                RECT 208.230 55.735 210.150 142.735 ;
                RECT 212.070 55.735 213.990 142.735 ;
                RECT 235.750 55.735 237.670 142.735 ;
                RECT 239.590 55.735 241.510 142.735 ;
                RECT 243.430 55.735 245.350 142.735 ;
                RECT 247.270 55.735 249.190 142.735 ;
                RECT 251.110 55.735 253.030 142.735 ;
                RECT 254.950 55.735 256.870 142.735 ;
                RECT 258.790 55.735 260.710 142.735 ;
                RECT 262.630 55.735 264.550 142.735 ;
                RECT 266.470 55.735 268.390 142.735 ;
                RECT 208.355 203.560 210.275 252.640 ;
                RECT 215.845 203.560 217.595 252.640 ;
                RECT 222.065 203.560 223.605 252.640 ;
                RECT 231.645 203.560 233.565 252.640 ;
                RECT 248.585 203.560 250.505 252.640 ;
                RECT 252.425 203.560 254.345 252.640 ;
                RECT 256.265 203.560 258.185 252.640 ;
                RECT 260.105 203.560 262.025 252.640 ;
                RECT 263.945 203.560 265.865 252.640 ;
                RECT 267.785 203.560 269.705 252.640 ;
                RECT 222.520 192.400 224.440 197.560 ;
                RECT 231.660 192.400 233.580 197.560 ;
                RECT 235.500 192.400 237.420 197.560 ;
                RECT 251.150 192.400 253.070 197.560 ;
                RECT 254.990 192.400 256.910 197.560 ;
                RECT 258.830 192.400 260.750 197.560 ;
                RECT 262.670 192.400 264.590 197.560 ;
                RECT 266.510 192.400 268.430 197.560 ;
                RECT 267.665 46.155 269.585 49.735 ;
                RECT 27.350 261.545 36.510 262.295 ;
                RECT 27.350 266.945 36.510 268.865 ;
                RECT 111.790 247.555 127.830 249.205 ;
                RECT 90.190 247.685 109.830 251.285 ;
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 314.280 5.560 ;
                RECT 316.000 5.240 325.160 5.560 ;
                RECT 326.880 5.240 336.040 5.560 ;
                RECT 337.760 5.240 346.920 5.560 ;
                RECT 348.640 5.240 357.800 5.560 ;
                RECT 359.520 5.240 368.680 5.560 ;
                RECT 370.400 5.240 379.560 5.560 ;
                RECT 381.280 5.240 390.440 5.560 ;
                RECT 392.160 5.240 401.320 5.560 ;
                RECT 403.040 5.240 412.200 5.560 ;
                RECT 413.920 5.240 423.080 5.560 ;
                RECT 424.800 5.240 433.960 5.560 ;
                RECT 435.680 5.240 444.840 5.560 ;
                RECT 446.560 5.240 455.720 5.560 ;
                RECT 457.440 5.240 466.600 5.560 ;
                RECT 468.320 5.240 477.480 5.560 ;
                RECT 479.200 5.240 488.360 5.560 ;
                RECT 490.080 5.240 499.240 5.560 ;
                RECT 500.960 5.240 510.120 5.560 ;
                RECT 511.840 5.240 521.680 5.560 ;
                RECT 522.720 5.240 532.560 5.560 ;
                RECT 533.600 5.240 543.440 5.560 ;
                RECT 544.480 5.240 554.320 5.560 ;
                RECT 555.360 5.240 565.200 5.560 ;
                RECT 566.240 5.240 576.080 5.560 ;
                RECT 577.120 5.240 586.960 5.560 ;
                RECT 588.000 5.240 597.840 5.560 ;
                RECT 598.880 5.240 608.720 5.560 ;
                RECT 609.760 5.240 619.600 5.560 ;
                RECT 621.320 5.240 630.480 5.560 ;
                RECT 632.200 5.240 641.360 5.560 ;
                RECT 643.080 5.240 652.240 5.560 ;
                RECT 653.960 5.240 671.600 5.560 ;
                RECT 2.880 6.600 671.600 6.920 ;
                RECT 2.880 7.960 671.600 8.280 ;
                RECT 2.880 9.320 272.120 9.640 ;
                RECT 307.160 9.320 671.600 9.640 ;
                RECT 2.880 10.680 671.600 11.000 ;
                RECT 2.880 12.040 671.600 12.360 ;
                RECT 2.880 13.400 191.200 13.720 ;
                RECT 273.160 13.400 671.600 13.720 ;
                RECT 2.880 14.760 671.600 15.080 ;
                RECT 2.880 16.120 671.600 16.440 ;
                RECT 2.880 17.480 191.200 17.800 ;
                RECT 272.480 17.480 671.600 17.800 ;
                RECT 2.880 18.840 671.600 19.160 ;
                RECT 2.880 20.200 671.600 20.520 ;
                RECT 2.880 21.560 671.600 21.880 ;
                RECT 2.880 22.920 671.600 23.240 ;
                RECT 2.880 24.280 671.600 24.600 ;
                RECT 2.880 25.640 671.600 25.960 ;
                RECT 2.880 27.000 671.600 27.320 ;
                RECT 2.880 28.360 313.600 28.680 ;
                RECT 576.440 28.360 671.600 28.680 ;
                RECT 2.880 29.720 301.360 30.040 ;
                RECT 664.840 29.720 671.600 30.040 ;
                RECT 2.880 31.080 301.360 31.400 ;
                RECT 664.840 31.080 671.600 31.400 ;
                RECT 2.880 32.440 301.360 32.760 ;
                RECT 664.840 32.440 671.600 32.760 ;
                RECT 2.880 33.800 301.360 34.120 ;
                RECT 664.840 33.800 671.600 34.120 ;
                RECT 2.880 35.160 301.360 35.480 ;
                RECT 664.840 35.160 671.600 35.480 ;
                RECT 2.880 36.520 159.920 36.840 ;
                RECT 245.280 36.520 301.360 36.840 ;
                RECT 664.840 36.520 671.600 36.840 ;
                RECT 2.880 37.880 158.560 38.200 ;
                RECT 251.400 37.880 301.360 38.200 ;
                RECT 664.840 37.880 671.600 38.200 ;
                RECT 2.880 39.240 157.200 39.560 ;
                RECT 257.520 39.240 301.360 39.560 ;
                RECT 664.840 39.240 671.600 39.560 ;
                RECT 2.880 40.600 134.080 40.920 ;
                RECT 272.480 40.600 301.360 40.920 ;
                RECT 664.840 40.600 671.600 40.920 ;
                RECT 2.880 41.960 134.760 42.280 ;
                RECT 262.960 41.960 301.360 42.280 ;
                RECT 664.840 41.960 671.600 42.280 ;
                RECT 2.880 43.320 301.360 43.640 ;
                RECT 664.840 43.320 671.600 43.640 ;
                RECT 2.880 44.680 301.360 45.000 ;
                RECT 664.840 44.680 671.600 45.000 ;
                RECT 2.880 46.040 263.280 46.360 ;
                RECT 270.440 46.040 300.680 46.360 ;
                RECT 664.840 46.040 671.600 46.360 ;
                RECT 2.880 47.400 263.280 47.720 ;
                RECT 664.840 47.400 671.600 47.720 ;
                RECT 2.880 48.760 155.160 49.080 ;
                RECT 270.440 48.760 301.360 49.080 ;
                RECT 664.840 48.760 671.600 49.080 ;
                RECT 2.880 50.120 301.360 50.440 ;
                RECT 664.840 50.120 671.600 50.440 ;
                RECT 2.880 51.480 301.360 51.800 ;
                RECT 664.840 51.480 671.600 51.800 ;
                RECT 2.880 52.840 301.360 53.160 ;
                RECT 664.840 52.840 671.600 53.160 ;
                RECT 2.880 54.200 301.360 54.520 ;
                RECT 664.840 54.200 671.600 54.520 ;
                RECT 2.880 55.560 171.480 55.880 ;
                RECT 269.080 55.560 301.360 55.880 ;
                RECT 664.840 55.560 671.600 55.880 ;
                RECT 2.880 56.920 157.200 57.240 ;
                RECT 164.360 56.920 171.480 57.240 ;
                RECT 269.080 56.920 301.360 57.240 ;
                RECT 664.840 56.920 671.600 57.240 ;
                RECT 2.880 58.280 158.560 58.600 ;
                RECT 163.000 58.280 171.480 58.600 ;
                RECT 281.320 58.280 301.360 58.600 ;
                RECT 664.840 58.280 671.600 58.600 ;
                RECT 2.880 59.640 159.920 59.960 ;
                RECT 162.320 59.640 171.480 59.960 ;
                RECT 282.680 59.640 301.360 59.960 ;
                RECT 664.840 59.640 671.600 59.960 ;
                RECT 2.880 61.000 171.480 61.320 ;
                RECT 282.680 61.000 301.360 61.320 ;
                RECT 664.840 61.000 671.600 61.320 ;
                RECT 2.880 62.360 171.480 62.680 ;
                RECT 281.320 62.360 301.360 62.680 ;
                RECT 664.840 62.360 671.600 62.680 ;
                RECT 2.880 63.720 171.480 64.040 ;
                RECT 282.680 63.720 301.360 64.040 ;
                RECT 664.840 63.720 671.600 64.040 ;
                RECT 2.880 65.080 171.480 65.400 ;
                RECT 269.080 65.080 301.360 65.400 ;
                RECT 664.840 65.080 671.600 65.400 ;
                RECT 2.880 66.440 171.480 66.760 ;
                RECT 282.680 66.440 301.360 66.760 ;
                RECT 664.840 66.440 671.600 66.760 ;
                RECT 2.880 67.800 171.480 68.120 ;
                RECT 285.400 67.800 301.360 68.120 ;
                RECT 664.840 67.800 671.600 68.120 ;
                RECT 2.880 69.160 171.480 69.480 ;
                RECT 284.040 69.160 301.360 69.480 ;
                RECT 664.840 69.160 671.600 69.480 ;
                RECT 2.880 70.520 171.480 70.840 ;
                RECT 285.400 70.520 301.360 70.840 ;
                RECT 664.840 70.520 671.600 70.840 ;
                RECT 2.880 71.880 171.480 72.200 ;
                RECT 285.400 71.880 301.360 72.200 ;
                RECT 664.840 71.880 671.600 72.200 ;
                RECT 2.880 73.240 171.480 73.560 ;
                RECT 269.080 73.240 301.360 73.560 ;
                RECT 664.840 73.240 671.600 73.560 ;
                RECT 2.880 74.600 171.480 74.920 ;
                RECT 285.400 74.600 301.360 74.920 ;
                RECT 664.840 74.600 671.600 74.920 ;
                RECT 2.880 75.960 171.480 76.280 ;
                RECT 269.080 75.960 301.360 76.280 ;
                RECT 664.840 75.960 671.600 76.280 ;
                RECT 2.880 77.320 171.480 77.640 ;
                RECT 284.040 77.320 301.360 77.640 ;
                RECT 664.840 77.320 671.600 77.640 ;
                RECT 2.880 78.680 171.480 79.000 ;
                RECT 288.120 78.680 301.360 79.000 ;
                RECT 664.840 78.680 671.600 79.000 ;
                RECT 2.880 80.040 171.480 80.360 ;
                RECT 288.120 80.040 301.360 80.360 ;
                RECT 664.840 80.040 671.600 80.360 ;
                RECT 2.880 81.400 171.480 81.720 ;
                RECT 286.760 81.400 301.360 81.720 ;
                RECT 664.840 81.400 671.600 81.720 ;
                RECT 2.880 82.760 171.480 83.080 ;
                RECT 288.120 82.760 301.360 83.080 ;
                RECT 664.840 82.760 671.600 83.080 ;
                RECT 2.880 84.120 171.480 84.440 ;
                RECT 286.760 84.120 301.360 84.440 ;
                RECT 664.840 84.120 671.600 84.440 ;
                RECT 2.880 85.480 171.480 85.800 ;
                RECT 288.120 85.480 301.360 85.800 ;
                RECT 664.840 85.480 671.600 85.800 ;
                RECT 2.880 86.840 171.480 87.160 ;
                RECT 288.120 86.840 301.360 87.160 ;
                RECT 664.840 86.840 671.600 87.160 ;
                RECT 2.880 88.200 171.480 88.520 ;
                RECT 286.760 88.200 301.360 88.520 ;
                RECT 664.840 88.200 671.600 88.520 ;
                RECT 2.880 89.560 171.480 89.880 ;
                RECT 290.840 89.560 301.360 89.880 ;
                RECT 664.840 89.560 671.600 89.880 ;
                RECT 2.880 90.920 171.480 91.240 ;
                RECT 269.080 90.920 301.360 91.240 ;
                RECT 664.840 90.920 671.600 91.240 ;
                RECT 2.880 92.280 171.480 92.600 ;
                RECT 290.840 92.280 301.360 92.600 ;
                RECT 664.840 92.280 671.600 92.600 ;
                RECT 2.880 93.640 171.480 93.960 ;
                RECT 290.840 93.640 301.360 93.960 ;
                RECT 664.840 93.640 671.600 93.960 ;
                RECT 2.880 95.000 171.480 95.320 ;
                RECT 289.480 95.000 301.360 95.320 ;
                RECT 664.840 95.000 671.600 95.320 ;
                RECT 2.880 96.360 171.480 96.680 ;
                RECT 290.840 96.360 301.360 96.680 ;
                RECT 664.840 96.360 671.600 96.680 ;
                RECT 2.880 97.720 171.480 98.040 ;
                RECT 290.840 97.720 301.360 98.040 ;
                RECT 664.840 97.720 671.600 98.040 ;
                RECT 2.880 99.080 171.480 99.400 ;
                RECT 269.080 99.080 301.360 99.400 ;
                RECT 664.840 99.080 671.600 99.400 ;
                RECT 2.880 100.440 171.480 100.760 ;
                RECT 293.560 100.440 301.360 100.760 ;
                RECT 664.840 100.440 671.600 100.760 ;
                RECT 2.880 101.800 171.480 102.120 ;
                RECT 269.080 101.800 301.360 102.120 ;
                RECT 664.840 101.800 671.600 102.120 ;
                RECT 2.880 103.160 171.480 103.480 ;
                RECT 292.200 103.160 301.360 103.480 ;
                RECT 664.840 103.160 671.600 103.480 ;
                RECT 2.880 104.520 171.480 104.840 ;
                RECT 293.560 104.520 301.360 104.840 ;
                RECT 664.840 104.520 671.600 104.840 ;
                RECT 2.880 105.880 171.480 106.200 ;
                RECT 293.560 105.880 301.360 106.200 ;
                RECT 664.840 105.880 671.600 106.200 ;
                RECT 2.880 107.240 171.480 107.560 ;
                RECT 292.200 107.240 301.360 107.560 ;
                RECT 664.840 107.240 671.600 107.560 ;
                RECT 2.880 108.600 171.480 108.920 ;
                RECT 293.560 108.600 301.360 108.920 ;
                RECT 664.840 108.600 671.600 108.920 ;
                RECT 2.880 109.960 171.480 110.280 ;
                RECT 292.200 109.960 301.360 110.280 ;
                RECT 664.840 109.960 671.600 110.280 ;
                RECT 2.880 111.320 171.480 111.640 ;
                RECT 296.280 111.320 301.360 111.640 ;
                RECT 664.840 111.320 671.600 111.640 ;
                RECT 2.880 112.680 171.480 113.000 ;
                RECT 296.280 112.680 301.360 113.000 ;
                RECT 664.840 112.680 671.600 113.000 ;
                RECT 2.880 114.040 171.480 114.360 ;
                RECT 294.920 114.040 301.360 114.360 ;
                RECT 664.840 114.040 671.600 114.360 ;
                RECT 2.880 115.400 171.480 115.720 ;
                RECT 296.280 115.400 301.360 115.720 ;
                RECT 664.840 115.400 671.600 115.720 ;
                RECT 2.880 116.760 171.480 117.080 ;
                RECT 269.080 116.760 301.360 117.080 ;
                RECT 664.840 116.760 671.600 117.080 ;
                RECT 2.880 118.120 171.480 118.440 ;
                RECT 296.280 118.120 301.360 118.440 ;
                RECT 664.840 118.120 671.600 118.440 ;
                RECT 2.880 119.480 171.480 119.800 ;
                RECT 296.280 119.480 301.360 119.800 ;
                RECT 664.840 119.480 671.600 119.800 ;
                RECT 2.880 120.840 171.480 121.160 ;
                RECT 269.080 120.840 301.360 121.160 ;
                RECT 664.840 120.840 671.600 121.160 ;
                RECT 2.880 122.200 171.480 122.520 ;
                RECT 297.640 122.200 301.360 122.520 ;
                RECT 664.840 122.200 671.600 122.520 ;
                RECT 2.880 123.560 171.480 123.880 ;
                RECT 299.000 123.560 301.360 123.880 ;
                RECT 664.840 123.560 671.600 123.880 ;
                RECT 2.880 124.920 171.480 125.240 ;
                RECT 269.080 124.920 301.360 125.240 ;
                RECT 664.840 124.920 671.600 125.240 ;
                RECT 2.880 126.280 171.480 126.600 ;
                RECT 299.000 126.280 301.360 126.600 ;
                RECT 664.840 126.280 671.600 126.600 ;
                RECT 2.880 127.640 171.480 127.960 ;
                RECT 299.000 127.640 301.360 127.960 ;
                RECT 664.840 127.640 671.600 127.960 ;
                RECT 2.880 129.000 171.480 129.320 ;
                RECT 297.640 129.000 301.360 129.320 ;
                RECT 664.840 129.000 671.600 129.320 ;
                RECT 2.880 130.360 171.480 130.680 ;
                RECT 299.000 130.360 301.360 130.680 ;
                RECT 664.840 130.360 671.600 130.680 ;
                RECT 2.880 131.720 171.480 132.040 ;
                RECT 664.840 131.720 671.600 132.040 ;
                RECT 2.880 133.080 171.480 133.400 ;
                RECT 664.840 133.080 671.600 133.400 ;
                RECT 2.880 134.440 171.480 134.760 ;
                RECT 664.840 134.440 671.600 134.760 ;
                RECT 2.880 135.800 171.480 136.120 ;
                RECT 664.840 135.800 671.600 136.120 ;
                RECT 2.880 137.160 171.480 137.480 ;
                RECT 664.840 137.160 671.600 137.480 ;
                RECT 2.880 138.520 171.480 138.840 ;
                RECT 664.840 138.520 671.600 138.840 ;
                RECT 2.880 139.880 171.480 140.200 ;
                RECT 664.840 139.880 671.600 140.200 ;
                RECT 2.880 141.240 110.280 141.560 ;
                RECT 129.000 141.240 171.480 141.560 ;
                RECT 664.840 141.240 671.600 141.560 ;
                RECT 2.880 142.600 110.280 142.920 ;
                RECT 129.000 142.600 171.480 142.920 ;
                RECT 269.080 142.600 301.360 142.920 ;
                RECT 664.840 142.600 671.600 142.920 ;
                RECT 2.880 143.960 110.280 144.280 ;
                RECT 129.000 143.960 301.360 144.280 ;
                RECT 664.840 143.960 671.600 144.280 ;
                RECT 2.880 145.320 110.280 145.640 ;
                RECT 129.000 145.320 276.880 145.640 ;
                RECT 664.840 145.320 671.600 145.640 ;
                RECT 2.880 146.680 110.280 147.000 ;
                RECT 129.000 146.680 298.640 147.000 ;
                RECT 664.840 146.680 671.600 147.000 ;
                RECT 2.880 148.040 110.280 148.360 ;
                RECT 129.000 148.040 295.920 148.360 ;
                RECT 664.840 148.040 671.600 148.360 ;
                RECT 2.880 149.400 110.280 149.720 ;
                RECT 129.000 149.400 293.200 149.720 ;
                RECT 664.840 149.400 671.600 149.720 ;
                RECT 2.880 150.760 110.280 151.080 ;
                RECT 129.000 150.760 290.480 151.080 ;
                RECT 664.840 150.760 671.600 151.080 ;
                RECT 2.880 152.120 110.280 152.440 ;
                RECT 129.000 152.120 287.760 152.440 ;
                RECT 664.840 152.120 671.600 152.440 ;
                RECT 2.880 153.480 110.280 153.800 ;
                RECT 129.000 153.480 285.040 153.800 ;
                RECT 664.840 153.480 671.600 153.800 ;
                RECT 2.880 154.840 110.280 155.160 ;
                RECT 129.000 154.840 132.040 155.160 ;
                RECT 143.280 154.840 282.320 155.160 ;
                RECT 664.840 154.840 671.600 155.160 ;
                RECT 2.880 156.200 110.280 156.520 ;
                RECT 129.000 156.200 133.400 156.520 ;
                RECT 137.160 156.200 279.600 156.520 ;
                RECT 664.840 156.200 671.600 156.520 ;
                RECT 2.880 157.560 110.280 157.880 ;
                RECT 129.000 157.560 134.760 157.880 ;
                RECT 139.200 157.560 147.000 157.880 ;
                RECT 149.400 157.560 301.360 157.880 ;
                RECT 664.840 157.560 671.600 157.880 ;
                RECT 2.880 158.920 110.280 159.240 ;
                RECT 129.000 158.920 301.360 159.240 ;
                RECT 664.840 158.920 671.600 159.240 ;
                RECT 2.880 160.280 110.280 160.600 ;
                RECT 129.000 160.280 141.560 160.600 ;
                RECT 150.080 160.280 301.360 160.600 ;
                RECT 664.840 160.280 671.600 160.600 ;
                RECT 2.880 161.640 110.280 161.960 ;
                RECT 129.000 161.640 136.800 161.960 ;
                RECT 143.280 161.640 301.360 161.960 ;
                RECT 664.840 161.640 671.600 161.960 ;
                RECT 2.880 163.000 110.280 163.320 ;
                RECT 129.000 163.000 134.080 163.320 ;
                RECT 143.280 163.000 301.360 163.320 ;
                RECT 664.840 163.000 671.600 163.320 ;
                RECT 2.880 164.360 110.280 164.680 ;
                RECT 129.000 164.360 301.360 164.680 ;
                RECT 664.840 164.360 671.600 164.680 ;
                RECT 2.880 165.720 110.280 166.040 ;
                RECT 129.000 165.720 131.360 166.040 ;
                RECT 143.280 165.720 301.360 166.040 ;
                RECT 664.840 165.720 671.600 166.040 ;
                RECT 2.880 167.080 110.280 167.400 ;
                RECT 129.000 167.080 141.560 167.400 ;
                RECT 149.400 167.080 301.360 167.400 ;
                RECT 664.840 167.080 671.600 167.400 ;
                RECT 2.880 168.440 110.280 168.760 ;
                RECT 129.000 168.440 140.880 168.760 ;
                RECT 143.280 168.440 301.360 168.760 ;
                RECT 664.840 168.440 671.600 168.760 ;
                RECT 2.880 169.800 110.280 170.120 ;
                RECT 129.000 169.800 301.360 170.120 ;
                RECT 664.840 169.800 671.600 170.120 ;
                RECT 2.880 171.160 110.280 171.480 ;
                RECT 129.000 171.160 141.560 171.480 ;
                RECT 149.400 171.160 301.360 171.480 ;
                RECT 664.840 171.160 671.600 171.480 ;
                RECT 2.880 172.520 110.280 172.840 ;
                RECT 129.000 172.520 138.160 172.840 ;
                RECT 143.280 172.520 301.360 172.840 ;
                RECT 664.840 172.520 671.600 172.840 ;
                RECT 2.880 173.880 110.280 174.200 ;
                RECT 129.000 173.880 140.880 174.200 ;
                RECT 143.280 173.880 301.360 174.200 ;
                RECT 664.840 173.880 671.600 174.200 ;
                RECT 2.880 175.240 110.280 175.560 ;
                RECT 129.000 175.240 144.280 175.560 ;
                RECT 154.840 175.240 301.360 175.560 ;
                RECT 664.840 175.240 671.600 175.560 ;
                RECT 2.880 176.600 110.280 176.920 ;
                RECT 129.000 176.600 132.040 176.920 ;
                RECT 149.400 176.600 301.360 176.920 ;
                RECT 664.840 176.600 671.600 176.920 ;
                RECT 2.880 177.960 110.280 178.280 ;
                RECT 129.000 177.960 140.880 178.280 ;
                RECT 143.280 177.960 149.040 178.280 ;
                RECT 156.200 177.960 301.360 178.280 ;
                RECT 664.840 177.960 671.600 178.280 ;
                RECT 2.880 179.320 110.280 179.640 ;
                RECT 129.000 179.320 153.120 179.640 ;
                RECT 156.880 179.320 301.360 179.640 ;
                RECT 664.840 179.320 671.600 179.640 ;
                RECT 2.880 180.680 110.280 181.000 ;
                RECT 129.000 180.680 132.040 181.000 ;
                RECT 146.000 180.680 301.360 181.000 ;
                RECT 664.840 180.680 671.600 181.000 ;
                RECT 2.880 182.040 110.280 182.360 ;
                RECT 129.000 182.040 140.880 182.360 ;
                RECT 149.400 182.040 301.360 182.360 ;
                RECT 664.840 182.040 671.600 182.360 ;
                RECT 2.880 183.400 110.280 183.720 ;
                RECT 129.000 183.400 138.840 183.720 ;
                RECT 150.080 183.400 301.360 183.720 ;
                RECT 664.840 183.400 671.600 183.720 ;
                RECT 2.880 184.760 110.280 185.080 ;
                RECT 129.000 184.760 301.360 185.080 ;
                RECT 664.840 184.760 671.600 185.080 ;
                RECT 2.880 186.120 110.280 186.440 ;
                RECT 129.000 186.120 134.760 186.440 ;
                RECT 137.160 186.120 301.360 186.440 ;
                RECT 664.840 186.120 671.600 186.440 ;
                RECT 2.880 187.480 110.280 187.800 ;
                RECT 129.000 187.480 134.080 187.800 ;
                RECT 143.280 187.480 301.360 187.800 ;
                RECT 664.840 187.480 671.600 187.800 ;
                RECT 2.880 188.840 110.280 189.160 ;
                RECT 129.000 188.840 136.800 189.160 ;
                RECT 140.560 188.840 301.360 189.160 ;
                RECT 664.840 188.840 671.600 189.160 ;
                RECT 2.880 190.200 110.280 190.520 ;
                RECT 129.000 190.200 301.360 190.520 ;
                RECT 664.840 190.200 671.600 190.520 ;
                RECT 2.880 191.560 110.280 191.880 ;
                RECT 129.000 191.560 140.880 191.880 ;
                RECT 142.600 191.560 301.360 191.880 ;
                RECT 664.840 191.560 671.600 191.880 ;
                RECT 2.880 192.920 110.280 193.240 ;
                RECT 129.000 192.920 133.400 193.240 ;
                RECT 148.720 192.920 155.840 193.240 ;
                RECT 215.360 192.920 218.400 193.240 ;
                RECT 269.080 192.920 301.360 193.240 ;
                RECT 664.840 192.920 671.600 193.240 ;
                RECT 2.880 194.280 110.280 194.600 ;
                RECT 129.000 194.280 218.400 194.600 ;
                RECT 269.080 194.280 301.360 194.600 ;
                RECT 664.840 194.280 671.600 194.600 ;
                RECT 2.880 195.640 110.280 195.960 ;
                RECT 129.000 195.640 140.880 195.960 ;
                RECT 142.600 195.640 218.400 195.960 ;
                RECT 269.080 195.640 301.360 195.960 ;
                RECT 664.840 195.640 671.600 195.960 ;
                RECT 2.880 197.000 110.280 197.320 ;
                RECT 129.000 197.000 135.440 197.320 ;
                RECT 143.280 197.000 218.400 197.320 ;
                RECT 269.080 197.000 301.360 197.320 ;
                RECT 664.840 197.000 671.600 197.320 ;
                RECT 2.880 198.360 110.280 198.680 ;
                RECT 129.000 198.360 132.040 198.680 ;
                RECT 143.960 198.360 301.360 198.680 ;
                RECT 664.840 198.360 671.600 198.680 ;
                RECT 2.880 199.720 110.280 200.040 ;
                RECT 129.000 199.720 301.360 200.040 ;
                RECT 664.840 199.720 671.600 200.040 ;
                RECT 2.880 201.080 110.280 201.400 ;
                RECT 129.000 201.080 131.360 201.400 ;
                RECT 149.400 201.080 301.360 201.400 ;
                RECT 664.840 201.080 671.600 201.400 ;
                RECT 2.880 202.440 110.280 202.760 ;
                RECT 142.600 202.440 301.360 202.760 ;
                RECT 664.840 202.440 671.600 202.760 ;
                RECT 2.880 203.800 110.280 204.120 ;
                RECT 129.000 203.800 132.040 204.120 ;
                RECT 137.160 203.800 203.440 204.120 ;
                RECT 270.440 203.800 301.360 204.120 ;
                RECT 664.840 203.800 671.600 204.120 ;
                RECT 2.880 205.160 110.280 205.480 ;
                RECT 129.000 205.160 203.440 205.480 ;
                RECT 270.440 205.160 280.960 205.480 ;
                RECT 664.840 205.160 671.600 205.480 ;
                RECT 2.880 206.520 110.280 206.840 ;
                RECT 129.000 206.520 138.840 206.840 ;
                RECT 146.000 206.520 203.440 206.840 ;
                RECT 270.440 206.520 280.960 206.840 ;
                RECT 664.840 206.520 671.600 206.840 ;
                RECT 2.880 207.880 110.280 208.200 ;
                RECT 129.000 207.880 203.440 208.200 ;
                RECT 270.440 207.880 283.680 208.200 ;
                RECT 664.840 207.880 671.600 208.200 ;
                RECT 2.880 209.240 110.280 209.560 ;
                RECT 129.000 209.240 203.440 209.560 ;
                RECT 270.440 209.240 286.400 209.560 ;
                RECT 664.840 209.240 671.600 209.560 ;
                RECT 2.880 210.600 110.280 210.920 ;
                RECT 129.000 210.600 144.280 210.920 ;
                RECT 150.760 210.600 203.440 210.920 ;
                RECT 270.440 210.600 289.120 210.920 ;
                RECT 664.840 210.600 671.600 210.920 ;
                RECT 2.880 211.960 110.280 212.280 ;
                RECT 129.000 211.960 134.080 212.280 ;
                RECT 137.160 211.960 147.680 212.280 ;
                RECT 149.400 211.960 203.440 212.280 ;
                RECT 270.440 211.960 294.560 212.280 ;
                RECT 664.840 211.960 671.600 212.280 ;
                RECT 2.880 213.320 110.280 213.640 ;
                RECT 129.000 213.320 132.040 213.640 ;
                RECT 135.800 213.320 203.440 213.640 ;
                RECT 270.440 213.320 297.280 213.640 ;
                RECT 664.840 213.320 671.600 213.640 ;
                RECT 2.880 214.680 110.280 215.000 ;
                RECT 129.000 214.680 203.440 215.000 ;
                RECT 270.440 214.680 300.000 215.000 ;
                RECT 664.840 214.680 671.600 215.000 ;
                RECT 2.880 216.040 110.280 216.360 ;
                RECT 129.000 216.040 203.440 216.360 ;
                RECT 664.840 216.040 671.600 216.360 ;
                RECT 2.880 217.400 110.280 217.720 ;
                RECT 129.000 217.400 203.440 217.720 ;
                RECT 664.840 217.400 671.600 217.720 ;
                RECT 2.880 218.760 110.280 219.080 ;
                RECT 129.000 218.760 203.440 219.080 ;
                RECT 664.840 218.760 671.600 219.080 ;
                RECT 2.880 220.120 110.280 220.440 ;
                RECT 129.000 220.120 203.440 220.440 ;
                RECT 664.840 220.120 671.600 220.440 ;
                RECT 2.880 221.480 110.280 221.800 ;
                RECT 129.000 221.480 134.080 221.800 ;
                RECT 139.200 221.480 203.440 221.800 ;
                RECT 270.440 221.480 301.360 221.800 ;
                RECT 664.840 221.480 671.600 221.800 ;
                RECT 2.880 222.840 110.280 223.160 ;
                RECT 129.000 222.840 137.480 223.160 ;
                RECT 149.400 222.840 203.440 223.160 ;
                RECT 270.440 222.840 301.360 223.160 ;
                RECT 664.840 222.840 671.600 223.160 ;
                RECT 2.880 224.200 110.280 224.520 ;
                RECT 129.000 224.200 203.440 224.520 ;
                RECT 270.440 224.200 301.360 224.520 ;
                RECT 664.840 224.200 671.600 224.520 ;
                RECT 2.880 225.560 110.280 225.880 ;
                RECT 129.000 225.560 203.440 225.880 ;
                RECT 270.440 225.560 301.360 225.880 ;
                RECT 664.840 225.560 671.600 225.880 ;
                RECT 2.880 226.920 110.280 227.240 ;
                RECT 129.000 226.920 203.440 227.240 ;
                RECT 270.440 226.920 301.360 227.240 ;
                RECT 664.840 226.920 671.600 227.240 ;
                RECT 2.880 228.280 110.280 228.600 ;
                RECT 129.000 228.280 133.400 228.600 ;
                RECT 136.480 228.280 203.440 228.600 ;
                RECT 270.440 228.280 301.360 228.600 ;
                RECT 664.840 228.280 671.600 228.600 ;
                RECT 2.880 229.640 110.280 229.960 ;
                RECT 129.000 229.640 203.440 229.960 ;
                RECT 270.440 229.640 301.360 229.960 ;
                RECT 664.840 229.640 671.600 229.960 ;
                RECT 2.880 231.000 110.280 231.320 ;
                RECT 129.000 231.000 136.800 231.320 ;
                RECT 139.200 231.000 203.440 231.320 ;
                RECT 270.440 231.000 301.360 231.320 ;
                RECT 664.840 231.000 671.600 231.320 ;
                RECT 2.880 232.360 110.280 232.680 ;
                RECT 129.000 232.360 147.680 232.680 ;
                RECT 150.080 232.360 203.440 232.680 ;
                RECT 270.440 232.360 301.360 232.680 ;
                RECT 664.840 232.360 671.600 232.680 ;
                RECT 2.880 233.720 110.280 234.040 ;
                RECT 129.000 233.720 203.440 234.040 ;
                RECT 270.440 233.720 301.360 234.040 ;
                RECT 664.840 233.720 671.600 234.040 ;
                RECT 2.880 235.080 110.280 235.400 ;
                RECT 129.000 235.080 203.440 235.400 ;
                RECT 270.440 235.080 301.360 235.400 ;
                RECT 664.840 235.080 671.600 235.400 ;
                RECT 2.880 236.440 110.280 236.760 ;
                RECT 129.000 236.440 203.440 236.760 ;
                RECT 270.440 236.440 301.360 236.760 ;
                RECT 664.840 236.440 671.600 236.760 ;
                RECT 2.880 237.800 110.280 238.120 ;
                RECT 129.000 237.800 203.440 238.120 ;
                RECT 270.440 237.800 301.360 238.120 ;
                RECT 664.840 237.800 671.600 238.120 ;
                RECT 2.880 239.160 203.440 239.480 ;
                RECT 270.440 239.160 301.360 239.480 ;
                RECT 664.840 239.160 671.600 239.480 ;
                RECT 2.880 240.520 140.880 240.840 ;
                RECT 149.400 240.520 203.440 240.840 ;
                RECT 270.440 240.520 301.360 240.840 ;
                RECT 664.840 240.520 671.600 240.840 ;
                RECT 2.880 241.880 89.200 242.200 ;
                RECT 110.640 241.880 135.440 242.200 ;
                RECT 139.200 241.880 203.440 242.200 ;
                RECT 270.440 241.880 301.360 242.200 ;
                RECT 664.840 241.880 671.600 242.200 ;
                RECT 2.880 243.240 89.200 243.560 ;
                RECT 110.640 243.240 203.440 243.560 ;
                RECT 270.440 243.240 301.360 243.560 ;
                RECT 664.840 243.240 671.600 243.560 ;
                RECT 2.880 244.600 89.200 244.920 ;
                RECT 110.640 244.600 203.440 244.920 ;
                RECT 270.440 244.600 301.360 244.920 ;
                RECT 664.840 244.600 671.600 244.920 ;
                RECT 2.880 245.960 89.200 246.280 ;
                RECT 110.640 245.960 116.400 246.280 ;
                RECT 124.240 245.960 137.480 246.280 ;
                RECT 143.960 245.960 203.440 246.280 ;
                RECT 270.440 245.960 301.360 246.280 ;
                RECT 664.840 245.960 671.600 246.280 ;
                RECT 2.880 247.320 89.200 247.640 ;
                RECT 128.320 247.320 203.440 247.640 ;
                RECT 664.840 247.320 671.600 247.640 ;
                RECT 2.880 248.680 89.200 249.000 ;
                RECT 128.320 248.680 203.440 249.000 ;
                RECT 664.840 248.680 671.600 249.000 ;
                RECT 2.880 250.040 89.200 250.360 ;
                RECT 110.640 250.040 203.440 250.360 ;
                RECT 664.840 250.040 671.600 250.360 ;
                RECT 2.880 251.400 89.200 251.720 ;
                RECT 110.640 251.400 116.400 251.720 ;
                RECT 124.240 251.400 132.040 251.720 ;
                RECT 142.600 251.400 203.440 251.720 ;
                RECT 664.840 251.400 671.600 251.720 ;
                RECT 2.880 252.760 74.920 253.080 ;
                RECT 123.560 252.760 203.440 253.080 ;
                RECT 270.440 252.760 671.600 253.080 ;
                RECT 2.880 254.120 123.200 254.440 ;
                RECT 200.400 254.120 671.600 254.440 ;
                RECT 2.880 255.480 298.640 255.800 ;
                RECT 666.880 255.480 671.600 255.800 ;
                RECT 2.880 256.840 298.640 257.160 ;
                RECT 666.880 256.840 671.600 257.160 ;
                RECT 2.880 258.200 298.640 258.520 ;
                RECT 666.880 258.200 671.600 258.520 ;
                RECT 2.880 259.560 28.680 259.880 ;
                RECT 35.160 259.560 37.520 259.880 ;
                RECT 51.480 259.560 106.200 259.880 ;
                RECT 666.880 259.560 671.600 259.880 ;
                RECT 2.880 260.920 26.640 261.240 ;
                RECT 50.800 260.920 62.680 261.240 ;
                RECT 64.400 260.920 77.640 261.240 ;
                RECT 95.680 260.920 106.200 261.240 ;
                RECT 666.880 260.920 671.600 261.240 ;
                RECT 2.880 262.280 26.640 262.600 ;
                RECT 37.200 262.280 62.680 262.600 ;
                RECT 67.120 262.280 77.640 262.600 ;
                RECT 95.680 262.280 106.200 262.600 ;
                RECT 666.880 262.280 671.600 262.600 ;
                RECT 2.880 263.640 26.640 263.960 ;
                RECT 37.200 263.640 62.680 263.960 ;
                RECT 67.120 263.640 77.640 263.960 ;
                RECT 95.680 263.640 106.200 263.960 ;
                RECT 666.880 263.640 671.600 263.960 ;
                RECT 2.880 265.000 26.640 265.320 ;
                RECT 37.200 265.000 62.680 265.320 ;
                RECT 67.800 265.000 77.640 265.320 ;
                RECT 95.680 265.000 106.200 265.320 ;
                RECT 666.880 265.000 671.600 265.320 ;
                RECT 2.880 266.360 26.640 266.680 ;
                RECT 37.200 266.360 62.680 266.680 ;
                RECT 64.400 266.360 77.640 266.680 ;
                RECT 95.680 266.360 106.200 266.680 ;
                RECT 666.880 266.360 671.600 266.680 ;
                RECT 2.880 267.720 26.640 268.040 ;
                RECT 37.200 267.720 106.200 268.040 ;
                RECT 666.880 267.720 671.600 268.040 ;
                RECT 2.880 269.080 26.640 269.400 ;
                RECT 37.200 269.080 77.640 269.400 ;
                RECT 95.680 269.080 106.200 269.400 ;
                RECT 666.880 269.080 671.600 269.400 ;
                RECT 2.880 270.440 77.640 270.760 ;
                RECT 95.680 270.440 106.200 270.760 ;
                RECT 666.880 270.440 671.600 270.760 ;
                RECT 2.880 271.800 77.640 272.120 ;
                RECT 95.680 271.800 106.200 272.120 ;
                RECT 666.880 271.800 671.600 272.120 ;
                RECT 2.880 273.160 19.840 273.480 ;
                RECT 22.240 273.160 77.640 273.480 ;
                RECT 95.680 273.160 106.200 273.480 ;
                RECT 666.880 273.160 671.600 273.480 ;
                RECT 2.880 274.520 77.640 274.840 ;
                RECT 95.680 274.520 106.200 274.840 ;
                RECT 666.880 274.520 671.600 274.840 ;
                RECT 2.880 275.880 19.160 276.200 ;
                RECT 22.240 275.880 35.480 276.200 ;
                RECT 50.800 275.880 106.200 276.200 ;
                RECT 666.880 275.880 671.600 276.200 ;
                RECT 2.880 277.240 18.480 277.560 ;
                RECT 22.240 277.240 35.480 277.560 ;
                RECT 50.120 277.240 62.680 277.560 ;
                RECT 64.400 277.240 77.640 277.560 ;
                RECT 95.680 277.240 106.200 277.560 ;
                RECT 666.880 277.240 671.600 277.560 ;
                RECT 2.880 278.600 17.800 278.920 ;
                RECT 22.240 278.600 35.480 278.920 ;
                RECT 40.600 278.600 62.680 278.920 ;
                RECT 65.080 278.600 77.640 278.920 ;
                RECT 95.680 278.600 106.200 278.920 ;
                RECT 666.880 278.600 671.600 278.920 ;
                RECT 2.880 279.960 62.680 280.280 ;
                RECT 65.760 279.960 77.640 280.280 ;
                RECT 95.680 279.960 106.200 280.280 ;
                RECT 666.880 279.960 671.600 280.280 ;
                RECT 2.880 281.320 17.120 281.640 ;
                RECT 22.240 281.320 35.480 281.640 ;
                RECT 41.280 281.320 62.680 281.640 ;
                RECT 65.760 281.320 77.640 281.640 ;
                RECT 95.680 281.320 106.200 281.640 ;
                RECT 666.880 281.320 671.600 281.640 ;
                RECT 2.880 282.680 16.440 283.000 ;
                RECT 22.240 282.680 35.480 283.000 ;
                RECT 41.960 282.680 62.680 283.000 ;
                RECT 66.440 282.680 77.640 283.000 ;
                RECT 95.680 282.680 106.200 283.000 ;
                RECT 666.880 282.680 671.600 283.000 ;
                RECT 2.880 284.040 15.760 284.360 ;
                RECT 22.240 284.040 106.200 284.360 ;
                RECT 666.880 284.040 671.600 284.360 ;
                RECT 2.880 285.400 15.080 285.720 ;
                RECT 22.240 285.400 77.640 285.720 ;
                RECT 95.680 285.400 106.200 285.720 ;
                RECT 666.880 285.400 671.600 285.720 ;
                RECT 2.880 286.760 77.640 287.080 ;
                RECT 95.680 286.760 106.200 287.080 ;
                RECT 666.880 286.760 671.600 287.080 ;
                RECT 2.880 288.120 14.400 288.440 ;
                RECT 22.240 288.120 77.640 288.440 ;
                RECT 95.680 288.120 106.200 288.440 ;
                RECT 666.880 288.120 671.600 288.440 ;
                RECT 2.880 289.480 13.720 289.800 ;
                RECT 22.240 289.480 77.640 289.800 ;
                RECT 95.680 289.480 106.200 289.800 ;
                RECT 666.880 289.480 671.600 289.800 ;
                RECT 2.880 290.840 77.640 291.160 ;
                RECT 90.240 290.840 106.200 291.160 ;
                RECT 666.880 290.840 671.600 291.160 ;
                RECT 2.880 292.200 13.040 292.520 ;
                RECT 22.240 292.200 35.480 292.520 ;
                RECT 41.960 292.200 85.800 292.520 ;
                RECT 95.680 292.200 106.200 292.520 ;
                RECT 666.880 292.200 671.600 292.520 ;
                RECT 2.880 293.560 12.360 293.880 ;
                RECT 22.240 293.560 35.480 293.880 ;
                RECT 41.280 293.560 77.640 293.880 ;
                RECT 95.680 293.560 106.200 293.880 ;
                RECT 666.880 293.560 671.600 293.880 ;
                RECT 2.880 294.920 77.640 295.240 ;
                RECT 95.680 294.920 106.200 295.240 ;
                RECT 666.880 294.920 671.600 295.240 ;
                RECT 2.880 296.280 11.680 296.600 ;
                RECT 22.240 296.280 35.480 296.600 ;
                RECT 40.600 296.280 77.640 296.600 ;
                RECT 95.680 296.280 106.200 296.600 ;
                RECT 666.880 296.280 671.600 296.600 ;
                RECT 2.880 297.640 11.000 297.960 ;
                RECT 22.240 297.640 35.480 297.960 ;
                RECT 39.920 297.640 77.640 297.960 ;
                RECT 95.680 297.640 106.200 297.960 ;
                RECT 666.880 297.640 671.600 297.960 ;
                RECT 2.880 299.000 10.320 299.320 ;
                RECT 22.240 299.000 35.480 299.320 ;
                RECT 39.240 299.000 77.640 299.320 ;
                RECT 90.240 299.000 106.200 299.320 ;
                RECT 666.880 299.000 671.600 299.320 ;
                RECT 2.880 300.360 9.640 300.680 ;
                RECT 22.240 300.360 77.640 300.680 ;
                RECT 95.680 300.360 106.200 300.680 ;
                RECT 666.880 300.360 671.600 300.680 ;
                RECT 2.880 301.720 77.640 302.040 ;
                RECT 95.680 301.720 106.200 302.040 ;
                RECT 666.880 301.720 671.600 302.040 ;
                RECT 2.880 303.080 77.640 303.400 ;
                RECT 95.680 303.080 106.200 303.400 ;
                RECT 666.880 303.080 671.600 303.400 ;
                RECT 2.880 304.440 77.640 304.760 ;
                RECT 95.680 304.440 106.200 304.760 ;
                RECT 666.880 304.440 671.600 304.760 ;
                RECT 2.880 305.800 77.640 306.120 ;
                RECT 95.680 305.800 106.200 306.120 ;
                RECT 666.880 305.800 671.600 306.120 ;
                RECT 2.880 307.160 77.640 307.480 ;
                RECT 90.920 307.160 106.200 307.480 ;
                RECT 666.880 307.160 671.600 307.480 ;
                RECT 2.880 308.520 77.640 308.840 ;
                RECT 95.680 308.520 106.200 308.840 ;
                RECT 666.880 308.520 671.600 308.840 ;
                RECT 2.880 309.880 77.640 310.200 ;
                RECT 95.680 309.880 106.200 310.200 ;
                RECT 666.880 309.880 671.600 310.200 ;
                RECT 2.880 311.240 77.640 311.560 ;
                RECT 95.680 311.240 106.200 311.560 ;
                RECT 666.880 311.240 671.600 311.560 ;
                RECT 2.880 312.600 77.640 312.920 ;
                RECT 95.680 312.600 106.200 312.920 ;
                RECT 666.880 312.600 671.600 312.920 ;
                RECT 2.880 313.960 77.640 314.280 ;
                RECT 95.680 313.960 106.200 314.280 ;
                RECT 666.880 313.960 671.600 314.280 ;
                RECT 2.880 315.320 106.200 315.640 ;
                RECT 666.880 315.320 671.600 315.640 ;
                RECT 2.880 316.680 77.640 317.000 ;
                RECT 95.680 316.680 106.200 317.000 ;
                RECT 666.880 316.680 671.600 317.000 ;
                RECT 2.880 318.040 77.640 318.360 ;
                RECT 95.680 318.040 106.200 318.360 ;
                RECT 666.880 318.040 671.600 318.360 ;
                RECT 2.880 319.400 77.640 319.720 ;
                RECT 95.680 319.400 106.200 319.720 ;
                RECT 666.880 319.400 671.600 319.720 ;
                RECT 2.880 320.760 77.640 321.080 ;
                RECT 95.680 320.760 106.200 321.080 ;
                RECT 666.880 320.760 671.600 321.080 ;
                RECT 2.880 322.120 77.640 322.440 ;
                RECT 95.680 322.120 106.200 322.440 ;
                RECT 666.880 322.120 671.600 322.440 ;
                RECT 2.880 323.480 106.200 323.800 ;
                RECT 666.880 323.480 671.600 323.800 ;
                RECT 2.880 324.840 77.640 325.160 ;
                RECT 95.680 324.840 106.200 325.160 ;
                RECT 666.880 324.840 671.600 325.160 ;
                RECT 2.880 326.200 77.640 326.520 ;
                RECT 95.680 326.200 106.200 326.520 ;
                RECT 666.880 326.200 671.600 326.520 ;
                RECT 2.880 327.560 77.640 327.880 ;
                RECT 95.680 327.560 106.200 327.880 ;
                RECT 666.880 327.560 671.600 327.880 ;
                RECT 2.880 328.920 77.640 329.240 ;
                RECT 95.680 328.920 106.200 329.240 ;
                RECT 666.880 328.920 671.600 329.240 ;
                RECT 2.880 330.280 77.640 330.600 ;
                RECT 95.680 330.280 106.200 330.600 ;
                RECT 666.880 330.280 671.600 330.600 ;
                RECT 2.880 331.640 106.200 331.960 ;
                RECT 666.880 331.640 671.600 331.960 ;
                RECT 2.880 333.000 77.640 333.320 ;
                RECT 95.680 333.000 106.200 333.320 ;
                RECT 666.880 333.000 671.600 333.320 ;
                RECT 2.880 334.360 77.640 334.680 ;
                RECT 95.680 334.360 106.200 334.680 ;
                RECT 666.880 334.360 671.600 334.680 ;
                RECT 2.880 335.720 77.640 336.040 ;
                RECT 95.680 335.720 106.200 336.040 ;
                RECT 666.880 335.720 671.600 336.040 ;
                RECT 2.880 337.080 77.640 337.400 ;
                RECT 95.680 337.080 106.200 337.400 ;
                RECT 666.880 337.080 671.600 337.400 ;
                RECT 2.880 338.440 77.640 338.760 ;
                RECT 93.640 338.440 106.200 338.760 ;
                RECT 666.880 338.440 671.600 338.760 ;
                RECT 2.880 339.800 89.880 340.120 ;
                RECT 95.680 339.800 106.200 340.120 ;
                RECT 666.880 339.800 671.600 340.120 ;
                RECT 2.880 341.160 77.640 341.480 ;
                RECT 95.680 341.160 106.200 341.480 ;
                RECT 666.880 341.160 671.600 341.480 ;
                RECT 2.880 342.520 77.640 342.840 ;
                RECT 95.680 342.520 106.200 342.840 ;
                RECT 666.880 342.520 671.600 342.840 ;
                RECT 2.880 343.880 77.640 344.200 ;
                RECT 95.680 343.880 106.200 344.200 ;
                RECT 666.880 343.880 671.600 344.200 ;
                RECT 2.880 345.240 77.640 345.560 ;
                RECT 95.680 345.240 106.200 345.560 ;
                RECT 666.880 345.240 671.600 345.560 ;
                RECT 2.880 346.600 77.640 346.920 ;
                RECT 94.320 346.600 106.200 346.920 ;
                RECT 666.880 346.600 671.600 346.920 ;
                RECT 2.880 347.960 77.640 348.280 ;
                RECT 95.680 347.960 106.200 348.280 ;
                RECT 666.880 347.960 671.600 348.280 ;
                RECT 2.880 349.320 77.640 349.640 ;
                RECT 95.680 349.320 106.200 349.640 ;
                RECT 666.880 349.320 671.600 349.640 ;
                RECT 2.880 350.680 77.640 351.000 ;
                RECT 95.680 350.680 106.200 351.000 ;
                RECT 666.880 350.680 671.600 351.000 ;
                RECT 2.880 352.040 77.640 352.360 ;
                RECT 95.680 352.040 106.200 352.360 ;
                RECT 666.880 352.040 671.600 352.360 ;
                RECT 2.880 353.400 77.640 353.720 ;
                RECT 95.680 353.400 106.200 353.720 ;
                RECT 666.880 353.400 671.600 353.720 ;
                RECT 2.880 354.760 106.200 355.080 ;
                RECT 666.880 354.760 671.600 355.080 ;
                RECT 2.880 356.120 79.680 356.440 ;
                RECT 95.680 356.120 106.200 356.440 ;
                RECT 666.880 356.120 671.600 356.440 ;
                RECT 2.880 357.480 79.680 357.800 ;
                RECT 95.680 357.480 106.200 357.800 ;
                RECT 666.880 357.480 671.600 357.800 ;
                RECT 2.880 358.840 87.160 359.160 ;
                RECT 95.680 358.840 106.200 359.160 ;
                RECT 666.880 358.840 671.600 359.160 ;
                RECT 2.880 360.200 79.680 360.520 ;
                RECT 95.680 360.200 106.200 360.520 ;
                RECT 666.880 360.200 671.600 360.520 ;
                RECT 2.880 361.560 79.680 361.880 ;
                RECT 95.680 361.560 106.200 361.880 ;
                RECT 666.880 361.560 671.600 361.880 ;
                RECT 2.880 362.920 41.600 363.240 ;
                RECT 50.800 362.920 106.200 363.240 ;
                RECT 666.880 362.920 671.600 363.240 ;
                RECT 2.880 364.280 40.240 364.600 ;
                RECT 50.120 364.280 62.680 364.600 ;
                RECT 64.400 364.280 77.640 364.600 ;
                RECT 95.680 364.280 106.200 364.600 ;
                RECT 666.880 364.280 671.600 364.600 ;
                RECT 2.880 365.640 62.680 365.960 ;
                RECT 67.120 365.640 77.640 365.960 ;
                RECT 95.680 365.640 106.200 365.960 ;
                RECT 666.880 365.640 671.600 365.960 ;
                RECT 2.880 367.000 62.680 367.320 ;
                RECT 67.120 367.000 77.640 367.320 ;
                RECT 95.680 367.000 106.200 367.320 ;
                RECT 666.880 367.000 671.600 367.320 ;
                RECT 2.880 368.360 62.680 368.680 ;
                RECT 67.800 368.360 77.640 368.680 ;
                RECT 95.680 368.360 106.200 368.680 ;
                RECT 666.880 368.360 671.600 368.680 ;
                RECT 2.880 369.720 62.680 370.040 ;
                RECT 68.480 369.720 77.640 370.040 ;
                RECT 95.680 369.720 106.200 370.040 ;
                RECT 666.880 369.720 671.600 370.040 ;
                RECT 2.880 371.080 106.200 371.400 ;
                RECT 666.880 371.080 671.600 371.400 ;
                RECT 2.880 372.440 77.640 372.760 ;
                RECT 95.680 372.440 106.200 372.760 ;
                RECT 666.880 372.440 671.600 372.760 ;
                RECT 2.880 373.800 77.640 374.120 ;
                RECT 95.680 373.800 106.200 374.120 ;
                RECT 666.880 373.800 671.600 374.120 ;
                RECT 2.880 375.160 77.640 375.480 ;
                RECT 95.680 375.160 106.200 375.480 ;
                RECT 666.880 375.160 671.600 375.480 ;
                RECT 2.880 376.520 77.640 376.840 ;
                RECT 95.680 376.520 106.200 376.840 ;
                RECT 666.880 376.520 671.600 376.840 ;
                RECT 2.880 377.880 39.560 378.200 ;
                RECT 51.480 377.880 77.640 378.200 ;
                RECT 80.720 377.880 106.200 378.200 ;
                RECT 666.880 377.880 671.600 378.200 ;
                RECT 2.880 379.240 38.200 379.560 ;
                RECT 50.800 379.240 91.920 379.560 ;
                RECT 95.680 379.240 106.200 379.560 ;
                RECT 666.880 379.240 671.600 379.560 ;
                RECT 2.880 380.600 62.680 380.920 ;
                RECT 65.080 380.600 77.640 380.920 ;
                RECT 95.680 380.600 106.200 380.920 ;
                RECT 666.880 380.600 671.600 380.920 ;
                RECT 2.880 381.960 62.680 382.280 ;
                RECT 65.760 381.960 77.640 382.280 ;
                RECT 95.680 381.960 106.200 382.280 ;
                RECT 666.880 381.960 671.600 382.280 ;
                RECT 2.880 383.320 62.680 383.640 ;
                RECT 65.760 383.320 77.640 383.640 ;
                RECT 95.680 383.320 106.200 383.640 ;
                RECT 666.880 383.320 671.600 383.640 ;
                RECT 2.880 384.680 62.680 385.000 ;
                RECT 64.400 384.680 77.640 385.000 ;
                RECT 95.680 384.680 106.200 385.000 ;
                RECT 666.880 384.680 671.600 385.000 ;
                RECT 2.880 386.040 62.680 386.360 ;
                RECT 66.440 386.040 77.640 386.360 ;
                RECT 81.400 386.040 106.200 386.360 ;
                RECT 666.880 386.040 671.600 386.360 ;
                RECT 2.880 387.400 77.640 387.720 ;
                RECT 95.680 387.400 106.200 387.720 ;
                RECT 666.880 387.400 671.600 387.720 ;
                RECT 2.880 388.760 77.640 389.080 ;
                RECT 95.680 388.760 106.200 389.080 ;
                RECT 666.880 388.760 671.600 389.080 ;
                RECT 2.880 390.120 77.640 390.440 ;
                RECT 95.680 390.120 106.200 390.440 ;
                RECT 666.880 390.120 671.600 390.440 ;
                RECT 2.880 391.480 77.640 391.800 ;
                RECT 95.680 391.480 106.200 391.800 ;
                RECT 666.880 391.480 671.600 391.800 ;
                RECT 2.880 392.840 77.640 393.160 ;
                RECT 95.680 392.840 106.200 393.160 ;
                RECT 666.880 392.840 671.600 393.160 ;
                RECT 2.880 394.200 106.200 394.520 ;
                RECT 666.880 394.200 671.600 394.520 ;
                RECT 2.880 395.560 77.640 395.880 ;
                RECT 95.680 395.560 106.200 395.880 ;
                RECT 666.880 395.560 671.600 395.880 ;
                RECT 2.880 396.920 77.640 397.240 ;
                RECT 95.680 396.920 106.200 397.240 ;
                RECT 666.880 396.920 671.600 397.240 ;
                RECT 2.880 398.280 77.640 398.600 ;
                RECT 95.680 398.280 106.200 398.600 ;
                RECT 666.880 398.280 671.600 398.600 ;
                RECT 2.880 399.640 77.640 399.960 ;
                RECT 95.680 399.640 106.200 399.960 ;
                RECT 666.880 399.640 671.600 399.960 ;
                RECT 2.880 401.000 77.640 401.320 ;
                RECT 95.680 401.000 106.200 401.320 ;
                RECT 666.880 401.000 671.600 401.320 ;
                RECT 2.880 402.360 106.200 402.680 ;
                RECT 666.880 402.360 671.600 402.680 ;
                RECT 2.880 403.720 77.640 404.040 ;
                RECT 95.680 403.720 106.200 404.040 ;
                RECT 666.880 403.720 671.600 404.040 ;
                RECT 2.880 405.080 77.640 405.400 ;
                RECT 95.680 405.080 106.200 405.400 ;
                RECT 666.880 405.080 671.600 405.400 ;
                RECT 2.880 406.440 77.640 406.760 ;
                RECT 95.680 406.440 106.200 406.760 ;
                RECT 666.880 406.440 671.600 406.760 ;
                RECT 2.880 407.800 77.640 408.120 ;
                RECT 95.680 407.800 106.200 408.120 ;
                RECT 666.880 407.800 671.600 408.120 ;
                RECT 2.880 409.160 77.640 409.480 ;
                RECT 95.680 409.160 106.200 409.480 ;
                RECT 666.880 409.160 671.600 409.480 ;
                RECT 2.880 410.520 106.200 410.840 ;
                RECT 666.880 410.520 671.600 410.840 ;
                RECT 2.880 411.880 77.640 412.200 ;
                RECT 95.680 411.880 106.200 412.200 ;
                RECT 666.880 411.880 671.600 412.200 ;
                RECT 2.880 413.240 77.640 413.560 ;
                RECT 95.680 413.240 106.200 413.560 ;
                RECT 666.880 413.240 671.600 413.560 ;
                RECT 2.880 414.600 77.640 414.920 ;
                RECT 95.680 414.600 106.200 414.920 ;
                RECT 666.880 414.600 671.600 414.920 ;
                RECT 2.880 415.960 77.640 416.280 ;
                RECT 95.680 415.960 106.200 416.280 ;
                RECT 666.880 415.960 671.600 416.280 ;
                RECT 2.880 417.320 77.640 417.640 ;
                RECT 84.120 417.320 106.200 417.640 ;
                RECT 666.880 417.320 671.600 417.640 ;
                RECT 2.880 418.680 85.800 419.000 ;
                RECT 95.680 418.680 106.200 419.000 ;
                RECT 666.880 418.680 671.600 419.000 ;
                RECT 2.880 420.040 77.640 420.360 ;
                RECT 95.680 420.040 106.200 420.360 ;
                RECT 666.880 420.040 671.600 420.360 ;
                RECT 2.880 421.400 77.640 421.720 ;
                RECT 95.680 421.400 106.200 421.720 ;
                RECT 666.880 421.400 671.600 421.720 ;
                RECT 2.880 422.760 77.640 423.080 ;
                RECT 95.680 422.760 106.200 423.080 ;
                RECT 666.880 422.760 671.600 423.080 ;
                RECT 2.880 424.120 77.640 424.440 ;
                RECT 95.680 424.120 106.200 424.440 ;
                RECT 666.880 424.120 671.600 424.440 ;
                RECT 2.880 425.480 77.640 425.800 ;
                RECT 84.800 425.480 106.200 425.800 ;
                RECT 666.880 425.480 671.600 425.800 ;
                RECT 2.880 426.840 77.640 427.160 ;
                RECT 95.680 426.840 106.200 427.160 ;
                RECT 666.880 426.840 671.600 427.160 ;
                RECT 2.880 428.200 77.640 428.520 ;
                RECT 95.680 428.200 106.200 428.520 ;
                RECT 666.880 428.200 671.600 428.520 ;
                RECT 2.880 429.560 77.640 429.880 ;
                RECT 95.680 429.560 106.200 429.880 ;
                RECT 666.880 429.560 671.600 429.880 ;
                RECT 2.880 430.920 77.640 431.240 ;
                RECT 95.680 430.920 106.200 431.240 ;
                RECT 666.880 430.920 671.600 431.240 ;
                RECT 2.880 432.280 77.640 432.600 ;
                RECT 95.680 432.280 106.200 432.600 ;
                RECT 666.880 432.280 671.600 432.600 ;
                RECT 2.880 433.640 106.200 433.960 ;
                RECT 666.880 433.640 671.600 433.960 ;
                RECT 2.880 435.000 77.640 435.320 ;
                RECT 95.680 435.000 106.200 435.320 ;
                RECT 666.880 435.000 671.600 435.320 ;
                RECT 2.880 436.360 77.640 436.680 ;
                RECT 95.680 436.360 106.200 436.680 ;
                RECT 666.880 436.360 671.600 436.680 ;
                RECT 2.880 437.720 77.640 438.040 ;
                RECT 95.680 437.720 106.200 438.040 ;
                RECT 666.880 437.720 671.600 438.040 ;
                RECT 2.880 439.080 77.640 439.400 ;
                RECT 95.680 439.080 106.200 439.400 ;
                RECT 666.880 439.080 671.600 439.400 ;
                RECT 2.880 440.440 77.640 440.760 ;
                RECT 95.680 440.440 106.200 440.760 ;
                RECT 666.880 440.440 671.600 440.760 ;
                RECT 2.880 441.800 106.200 442.120 ;
                RECT 666.880 441.800 671.600 442.120 ;
                RECT 2.880 443.160 77.640 443.480 ;
                RECT 95.680 443.160 106.200 443.480 ;
                RECT 666.880 443.160 671.600 443.480 ;
                RECT 2.880 444.520 77.640 444.840 ;
                RECT 95.680 444.520 106.200 444.840 ;
                RECT 666.880 444.520 671.600 444.840 ;
                RECT 2.880 445.880 77.640 446.200 ;
                RECT 95.680 445.880 106.200 446.200 ;
                RECT 666.880 445.880 671.600 446.200 ;
                RECT 2.880 447.240 77.640 447.560 ;
                RECT 95.680 447.240 106.200 447.560 ;
                RECT 666.880 447.240 671.600 447.560 ;
                RECT 2.880 448.600 77.640 448.920 ;
                RECT 95.680 448.600 106.200 448.920 ;
                RECT 666.880 448.600 671.600 448.920 ;
                RECT 2.880 449.960 106.200 450.280 ;
                RECT 666.880 449.960 671.600 450.280 ;
                RECT 2.880 451.320 77.640 451.640 ;
                RECT 95.680 451.320 106.200 451.640 ;
                RECT 666.880 451.320 671.600 451.640 ;
                RECT 2.880 452.680 77.640 453.000 ;
                RECT 95.680 452.680 106.200 453.000 ;
                RECT 666.880 452.680 671.600 453.000 ;
                RECT 2.880 454.040 77.640 454.360 ;
                RECT 95.680 454.040 106.200 454.360 ;
                RECT 666.880 454.040 671.600 454.360 ;
                RECT 2.880 455.400 77.640 455.720 ;
                RECT 95.680 455.400 106.200 455.720 ;
                RECT 666.880 455.400 671.600 455.720 ;
                RECT 2.880 456.760 77.640 457.080 ;
                RECT 86.840 456.760 106.200 457.080 ;
                RECT 666.880 456.760 671.600 457.080 ;
                RECT 2.880 458.120 87.840 458.440 ;
                RECT 95.680 458.120 106.200 458.440 ;
                RECT 666.880 458.120 671.600 458.440 ;
                RECT 2.880 459.480 81.040 459.800 ;
                RECT 95.680 459.480 106.200 459.800 ;
                RECT 666.880 459.480 671.600 459.800 ;
                RECT 2.880 460.840 81.040 461.160 ;
                RECT 95.680 460.840 106.200 461.160 ;
                RECT 666.880 460.840 671.600 461.160 ;
                RECT 2.880 462.200 81.040 462.520 ;
                RECT 95.680 462.200 106.200 462.520 ;
                RECT 666.880 462.200 671.600 462.520 ;
                RECT 2.880 463.560 81.040 463.880 ;
                RECT 95.680 463.560 106.200 463.880 ;
                RECT 666.880 463.560 671.600 463.880 ;
                RECT 2.880 464.920 106.200 465.240 ;
                RECT 666.880 464.920 671.600 465.240 ;
                RECT 2.880 466.280 89.880 466.600 ;
                RECT 95.680 466.280 106.200 466.600 ;
                RECT 666.880 466.280 671.600 466.600 ;
                RECT 2.880 467.640 81.040 467.960 ;
                RECT 95.680 467.640 106.200 467.960 ;
                RECT 666.880 467.640 671.600 467.960 ;
                RECT 2.880 469.000 81.040 469.320 ;
                RECT 95.680 469.000 106.200 469.320 ;
                RECT 666.880 469.000 671.600 469.320 ;
                RECT 2.880 470.360 81.040 470.680 ;
                RECT 95.680 470.360 106.200 470.680 ;
                RECT 666.880 470.360 671.600 470.680 ;
                RECT 2.880 471.720 81.040 472.040 ;
                RECT 95.680 471.720 106.200 472.040 ;
                RECT 666.880 471.720 671.600 472.040 ;
                RECT 2.880 473.080 106.200 473.400 ;
                RECT 666.880 473.080 671.600 473.400 ;
                RECT 2.880 474.440 81.040 474.760 ;
                RECT 95.680 474.440 106.200 474.760 ;
                RECT 666.880 474.440 671.600 474.760 ;
                RECT 2.880 475.800 91.920 476.120 ;
                RECT 95.680 475.800 106.200 476.120 ;
                RECT 666.880 475.800 671.600 476.120 ;
                RECT 2.880 477.160 81.040 477.480 ;
                RECT 95.680 477.160 106.200 477.480 ;
                RECT 666.880 477.160 671.600 477.480 ;
                RECT 2.880 478.520 81.040 478.840 ;
                RECT 95.680 478.520 106.200 478.840 ;
                RECT 666.880 478.520 671.600 478.840 ;
                RECT 2.880 479.880 81.040 480.200 ;
                RECT 95.680 479.880 106.200 480.200 ;
                RECT 666.880 479.880 671.600 480.200 ;
                RECT 2.880 481.240 106.200 481.560 ;
                RECT 666.880 481.240 671.600 481.560 ;
                RECT 2.880 482.600 81.720 482.920 ;
                RECT 95.680 482.600 106.200 482.920 ;
                RECT 666.880 482.600 671.600 482.920 ;
                RECT 2.880 483.960 81.720 484.280 ;
                RECT 95.680 483.960 106.200 484.280 ;
                RECT 666.880 483.960 671.600 484.280 ;
                RECT 2.880 485.320 87.160 485.640 ;
                RECT 95.680 485.320 106.200 485.640 ;
                RECT 666.880 485.320 671.600 485.640 ;
                RECT 2.880 486.680 81.720 487.000 ;
                RECT 95.680 486.680 106.200 487.000 ;
                RECT 666.880 486.680 671.600 487.000 ;
                RECT 2.880 488.040 81.720 488.360 ;
                RECT 95.680 488.040 106.200 488.360 ;
                RECT 666.880 488.040 671.600 488.360 ;
                RECT 2.880 489.400 106.200 489.720 ;
                RECT 666.880 489.400 671.600 489.720 ;
                RECT 2.880 490.760 81.720 491.080 ;
                RECT 95.680 490.760 106.200 491.080 ;
                RECT 666.880 490.760 671.600 491.080 ;
                RECT 2.880 492.120 81.720 492.440 ;
                RECT 95.680 492.120 106.200 492.440 ;
                RECT 666.880 492.120 671.600 492.440 ;
                RECT 2.880 493.480 81.720 493.800 ;
                RECT 95.680 493.480 106.200 493.800 ;
                RECT 666.880 493.480 671.600 493.800 ;
                RECT 2.880 494.840 89.200 495.160 ;
                RECT 95.680 494.840 106.200 495.160 ;
                RECT 666.880 494.840 671.600 495.160 ;
                RECT 2.880 496.200 81.720 496.520 ;
                RECT 95.680 496.200 106.200 496.520 ;
                RECT 666.880 496.200 671.600 496.520 ;
                RECT 2.880 497.560 106.200 497.880 ;
                RECT 666.880 497.560 671.600 497.880 ;
                RECT 2.880 498.920 81.720 499.240 ;
                RECT 95.680 498.920 106.200 499.240 ;
                RECT 666.880 498.920 671.600 499.240 ;
                RECT 2.880 500.280 81.720 500.600 ;
                RECT 95.680 500.280 106.200 500.600 ;
                RECT 666.880 500.280 671.600 500.600 ;
                RECT 2.880 501.640 81.720 501.960 ;
                RECT 95.680 501.640 106.200 501.960 ;
                RECT 666.880 501.640 671.600 501.960 ;
                RECT 2.880 503.000 81.720 503.320 ;
                RECT 95.680 503.000 106.200 503.320 ;
                RECT 666.880 503.000 671.600 503.320 ;
                RECT 2.880 504.360 106.200 504.680 ;
                RECT 666.880 504.360 671.600 504.680 ;
                RECT 2.880 505.720 91.920 506.040 ;
                RECT 95.680 505.720 106.200 506.040 ;
                RECT 666.880 505.720 671.600 506.040 ;
                RECT 2.880 507.080 81.720 507.400 ;
                RECT 95.680 507.080 106.200 507.400 ;
                RECT 666.880 507.080 671.600 507.400 ;
                RECT 2.880 508.440 81.720 508.760 ;
                RECT 95.680 508.440 106.200 508.760 ;
                RECT 666.880 508.440 671.600 508.760 ;
                RECT 2.880 509.800 81.720 510.120 ;
                RECT 95.680 509.800 106.200 510.120 ;
                RECT 666.880 509.800 671.600 510.120 ;
                RECT 2.880 511.160 81.720 511.480 ;
                RECT 95.680 511.160 106.200 511.480 ;
                RECT 666.880 511.160 671.600 511.480 ;
                RECT 2.880 512.520 106.200 512.840 ;
                RECT 666.880 512.520 671.600 512.840 ;
                RECT 2.880 513.880 82.400 514.200 ;
                RECT 95.680 513.880 106.200 514.200 ;
                RECT 666.880 513.880 671.600 514.200 ;
                RECT 2.880 515.240 86.480 515.560 ;
                RECT 95.680 515.240 106.200 515.560 ;
                RECT 666.880 515.240 671.600 515.560 ;
                RECT 2.880 516.600 82.400 516.920 ;
                RECT 95.680 516.600 106.200 516.920 ;
                RECT 666.880 516.600 671.600 516.920 ;
                RECT 2.880 517.960 82.400 518.280 ;
                RECT 95.680 517.960 106.200 518.280 ;
                RECT 666.880 517.960 671.600 518.280 ;
                RECT 2.880 519.320 82.400 519.640 ;
                RECT 95.680 519.320 106.200 519.640 ;
                RECT 666.880 519.320 671.600 519.640 ;
                RECT 2.880 520.680 106.200 521.000 ;
                RECT 666.880 520.680 671.600 521.000 ;
                RECT 2.880 522.040 82.400 522.360 ;
                RECT 95.680 522.040 106.200 522.360 ;
                RECT 666.880 522.040 671.600 522.360 ;
                RECT 2.880 523.400 82.400 523.720 ;
                RECT 95.680 523.400 106.200 523.720 ;
                RECT 666.880 523.400 671.600 523.720 ;
                RECT 2.880 524.760 88.520 525.080 ;
                RECT 95.680 524.760 106.200 525.080 ;
                RECT 666.880 524.760 671.600 525.080 ;
                RECT 2.880 526.120 82.400 526.440 ;
                RECT 95.680 526.120 106.200 526.440 ;
                RECT 666.880 526.120 671.600 526.440 ;
                RECT 2.880 527.480 82.400 527.800 ;
                RECT 95.680 527.480 106.200 527.800 ;
                RECT 666.880 527.480 671.600 527.800 ;
                RECT 2.880 528.840 106.200 529.160 ;
                RECT 666.880 528.840 671.600 529.160 ;
                RECT 2.880 530.200 82.400 530.520 ;
                RECT 95.680 530.200 106.200 530.520 ;
                RECT 666.880 530.200 671.600 530.520 ;
                RECT 2.880 531.560 82.400 531.880 ;
                RECT 95.680 531.560 106.200 531.880 ;
                RECT 666.880 531.560 671.600 531.880 ;
                RECT 2.880 532.920 82.400 533.240 ;
                RECT 95.680 532.920 106.200 533.240 ;
                RECT 666.880 532.920 671.600 533.240 ;
                RECT 2.880 534.280 91.240 534.600 ;
                RECT 95.680 534.280 106.200 534.600 ;
                RECT 666.880 534.280 671.600 534.600 ;
                RECT 2.880 535.640 82.400 535.960 ;
                RECT 95.680 535.640 106.200 535.960 ;
                RECT 666.880 535.640 671.600 535.960 ;
                RECT 2.880 537.000 106.200 537.320 ;
                RECT 666.880 537.000 671.600 537.320 ;
                RECT 2.880 538.360 82.400 538.680 ;
                RECT 95.680 538.360 106.200 538.680 ;
                RECT 666.880 538.360 671.600 538.680 ;
                RECT 2.880 539.720 82.400 540.040 ;
                RECT 95.680 539.720 106.200 540.040 ;
                RECT 666.880 539.720 671.600 540.040 ;
                RECT 2.880 541.080 82.400 541.400 ;
                RECT 95.680 541.080 106.200 541.400 ;
                RECT 666.880 541.080 671.600 541.400 ;
                RECT 2.880 542.440 82.400 542.760 ;
                RECT 95.680 542.440 106.200 542.760 ;
                RECT 666.880 542.440 671.600 542.760 ;
                RECT 2.880 543.800 106.200 544.120 ;
                RECT 666.880 543.800 671.600 544.120 ;
                RECT 2.880 545.160 85.800 545.480 ;
                RECT 95.680 545.160 106.200 545.480 ;
                RECT 666.880 545.160 671.600 545.480 ;
                RECT 2.880 546.520 82.400 546.840 ;
                RECT 95.680 546.520 106.200 546.840 ;
                RECT 666.880 546.520 671.600 546.840 ;
                RECT 2.880 547.880 82.400 548.200 ;
                RECT 95.680 547.880 106.200 548.200 ;
                RECT 666.880 547.880 671.600 548.200 ;
                RECT 2.880 549.240 82.400 549.560 ;
                RECT 95.680 549.240 106.200 549.560 ;
                RECT 666.880 549.240 671.600 549.560 ;
                RECT 2.880 550.600 82.400 550.920 ;
                RECT 95.680 550.600 106.200 550.920 ;
                RECT 666.880 550.600 671.600 550.920 ;
                RECT 2.880 551.960 106.200 552.280 ;
                RECT 666.880 551.960 671.600 552.280 ;
                RECT 2.880 553.320 87.840 553.640 ;
                RECT 95.680 553.320 106.200 553.640 ;
                RECT 666.880 553.320 671.600 553.640 ;
                RECT 2.880 554.680 88.520 555.000 ;
                RECT 95.680 554.680 106.200 555.000 ;
                RECT 666.880 554.680 671.600 555.000 ;
                RECT 2.880 556.040 82.400 556.360 ;
                RECT 95.680 556.040 106.200 556.360 ;
                RECT 666.880 556.040 671.600 556.360 ;
                RECT 2.880 557.400 82.400 557.720 ;
                RECT 95.680 557.400 106.200 557.720 ;
                RECT 666.880 557.400 671.600 557.720 ;
                RECT 2.880 558.760 82.400 559.080 ;
                RECT 95.680 558.760 106.200 559.080 ;
                RECT 666.880 558.760 671.600 559.080 ;
                RECT 2.880 560.120 106.200 560.440 ;
                RECT 666.880 560.120 671.600 560.440 ;
                RECT 2.880 561.480 82.400 561.800 ;
                RECT 95.680 561.480 106.200 561.800 ;
                RECT 666.880 561.480 671.600 561.800 ;
                RECT 2.880 562.840 90.560 563.160 ;
                RECT 95.680 562.840 106.200 563.160 ;
                RECT 666.880 562.840 671.600 563.160 ;
                RECT 2.880 564.200 90.560 564.520 ;
                RECT 95.680 564.200 106.200 564.520 ;
                RECT 666.880 564.200 671.600 564.520 ;
                RECT 2.880 565.560 82.400 565.880 ;
                RECT 95.680 565.560 106.200 565.880 ;
                RECT 666.880 565.560 671.600 565.880 ;
                RECT 2.880 566.920 82.400 567.240 ;
                RECT 95.680 566.920 106.200 567.240 ;
                RECT 666.880 566.920 671.600 567.240 ;
                RECT 2.880 568.280 106.200 568.600 ;
                RECT 666.880 568.280 671.600 568.600 ;
                RECT 2.880 569.640 82.400 569.960 ;
                RECT 95.680 569.640 106.200 569.960 ;
                RECT 666.880 569.640 671.600 569.960 ;
                RECT 2.880 571.000 82.400 571.320 ;
                RECT 95.680 571.000 106.200 571.320 ;
                RECT 666.880 571.000 671.600 571.320 ;
                RECT 2.880 572.360 82.400 572.680 ;
                RECT 95.680 572.360 106.200 572.680 ;
                RECT 666.880 572.360 671.600 572.680 ;
                RECT 2.880 573.720 93.280 574.040 ;
                RECT 95.680 573.720 106.200 574.040 ;
                RECT 666.880 573.720 671.600 574.040 ;
                RECT 2.880 575.080 82.400 575.400 ;
                RECT 95.680 575.080 106.200 575.400 ;
                RECT 666.880 575.080 671.600 575.400 ;
                RECT 2.880 576.440 106.200 576.760 ;
                RECT 666.880 576.440 671.600 576.760 ;
                RECT 2.880 577.800 83.080 578.120 ;
                RECT 95.680 577.800 106.200 578.120 ;
                RECT 666.880 577.800 671.600 578.120 ;
                RECT 2.880 579.160 83.080 579.480 ;
                RECT 95.680 579.160 106.200 579.480 ;
                RECT 666.880 579.160 671.600 579.480 ;
                RECT 2.880 580.520 83.080 580.840 ;
                RECT 95.680 580.520 106.200 580.840 ;
                RECT 666.880 580.520 671.600 580.840 ;
                RECT 2.880 581.880 83.080 582.200 ;
                RECT 95.680 581.880 106.200 582.200 ;
                RECT 666.880 581.880 671.600 582.200 ;
                RECT 2.880 583.240 106.200 583.560 ;
                RECT 666.880 583.240 671.600 583.560 ;
                RECT 2.880 584.600 87.840 584.920 ;
                RECT 95.680 584.600 106.200 584.920 ;
                RECT 666.880 584.600 671.600 584.920 ;
                RECT 2.880 585.960 83.080 586.280 ;
                RECT 95.680 585.960 106.200 586.280 ;
                RECT 666.880 585.960 671.600 586.280 ;
                RECT 2.880 587.320 83.080 587.640 ;
                RECT 95.680 587.320 106.200 587.640 ;
                RECT 666.880 587.320 671.600 587.640 ;
                RECT 2.880 588.680 83.080 589.000 ;
                RECT 95.680 588.680 106.200 589.000 ;
                RECT 666.880 588.680 671.600 589.000 ;
                RECT 2.880 590.040 83.080 590.360 ;
                RECT 95.680 590.040 106.200 590.360 ;
                RECT 666.880 590.040 671.600 590.360 ;
                RECT 2.880 591.400 106.200 591.720 ;
                RECT 666.880 591.400 671.600 591.720 ;
                RECT 2.880 592.760 89.880 593.080 ;
                RECT 95.680 592.760 106.200 593.080 ;
                RECT 666.880 592.760 671.600 593.080 ;
                RECT 2.880 594.120 83.080 594.440 ;
                RECT 95.680 594.120 106.200 594.440 ;
                RECT 666.880 594.120 671.600 594.440 ;
                RECT 2.880 595.480 83.080 595.800 ;
                RECT 95.680 595.480 106.200 595.800 ;
                RECT 666.880 595.480 671.600 595.800 ;
                RECT 2.880 596.840 83.080 597.160 ;
                RECT 95.680 596.840 106.200 597.160 ;
                RECT 666.880 596.840 671.600 597.160 ;
                RECT 2.880 598.200 83.080 598.520 ;
                RECT 95.680 598.200 106.200 598.520 ;
                RECT 666.880 598.200 671.600 598.520 ;
                RECT 2.880 599.560 106.200 599.880 ;
                RECT 666.880 599.560 671.600 599.880 ;
                RECT 2.880 600.920 83.080 601.240 ;
                RECT 95.680 600.920 106.200 601.240 ;
                RECT 666.880 600.920 671.600 601.240 ;
                RECT 2.880 602.280 91.920 602.600 ;
                RECT 95.680 602.280 106.200 602.600 ;
                RECT 666.880 602.280 671.600 602.600 ;
                RECT 2.880 603.640 83.080 603.960 ;
                RECT 95.680 603.640 106.200 603.960 ;
                RECT 666.880 603.640 671.600 603.960 ;
                RECT 2.880 605.000 83.080 605.320 ;
                RECT 95.680 605.000 106.200 605.320 ;
                RECT 666.880 605.000 671.600 605.320 ;
                RECT 2.880 606.360 83.080 606.680 ;
                RECT 95.680 606.360 106.200 606.680 ;
                RECT 666.880 606.360 671.600 606.680 ;
                RECT 2.880 607.720 106.200 608.040 ;
                RECT 666.880 607.720 671.600 608.040 ;
                RECT 2.880 609.080 83.760 609.400 ;
                RECT 95.680 609.080 106.200 609.400 ;
                RECT 666.880 609.080 671.600 609.400 ;
                RECT 2.880 610.440 83.760 610.760 ;
                RECT 95.680 610.440 106.200 610.760 ;
                RECT 666.880 610.440 671.600 610.760 ;
                RECT 2.880 611.800 87.160 612.120 ;
                RECT 95.680 611.800 106.200 612.120 ;
                RECT 666.880 611.800 671.600 612.120 ;
                RECT 2.880 613.160 87.160 613.480 ;
                RECT 95.680 613.160 106.200 613.480 ;
                RECT 666.880 613.160 671.600 613.480 ;
                RECT 2.880 614.520 83.760 614.840 ;
                RECT 95.680 614.520 106.200 614.840 ;
                RECT 666.880 614.520 671.600 614.840 ;
                RECT 2.880 615.880 106.200 616.200 ;
                RECT 666.880 615.880 671.600 616.200 ;
                RECT 2.880 617.240 83.760 617.560 ;
                RECT 95.680 617.240 106.200 617.560 ;
                RECT 666.880 617.240 671.600 617.560 ;
                RECT 2.880 618.600 83.760 618.920 ;
                RECT 95.680 618.600 106.200 618.920 ;
                RECT 666.880 618.600 671.600 618.920 ;
                RECT 2.880 619.960 83.760 620.280 ;
                RECT 95.680 619.960 106.200 620.280 ;
                RECT 666.880 619.960 671.600 620.280 ;
                RECT 2.880 621.320 83.760 621.640 ;
                RECT 95.680 621.320 106.200 621.640 ;
                RECT 666.880 621.320 671.600 621.640 ;
                RECT 2.880 622.680 106.200 623.000 ;
                RECT 666.880 622.680 671.600 623.000 ;
                RECT 2.880 624.040 89.880 624.360 ;
                RECT 95.680 624.040 106.200 624.360 ;
                RECT 666.880 624.040 671.600 624.360 ;
                RECT 2.880 625.400 83.760 625.720 ;
                RECT 95.680 625.400 106.200 625.720 ;
                RECT 666.880 625.400 671.600 625.720 ;
                RECT 2.880 626.760 83.760 627.080 ;
                RECT 95.680 626.760 106.200 627.080 ;
                RECT 666.880 626.760 671.600 627.080 ;
                RECT 2.880 628.120 83.760 628.440 ;
                RECT 95.680 628.120 106.200 628.440 ;
                RECT 666.880 628.120 671.600 628.440 ;
                RECT 2.880 629.480 83.760 629.800 ;
                RECT 95.680 629.480 106.200 629.800 ;
                RECT 666.880 629.480 671.600 629.800 ;
                RECT 2.880 630.840 106.200 631.160 ;
                RECT 666.880 630.840 671.600 631.160 ;
                RECT 2.880 632.200 91.920 632.520 ;
                RECT 95.680 632.200 106.200 632.520 ;
                RECT 666.880 632.200 671.600 632.520 ;
                RECT 2.880 633.560 83.760 633.880 ;
                RECT 95.680 633.560 106.200 633.880 ;
                RECT 666.880 633.560 671.600 633.880 ;
                RECT 2.880 634.920 83.760 635.240 ;
                RECT 95.680 634.920 106.200 635.240 ;
                RECT 666.880 634.920 671.600 635.240 ;
                RECT 2.880 636.280 83.760 636.600 ;
                RECT 95.680 636.280 106.200 636.600 ;
                RECT 666.880 636.280 671.600 636.600 ;
                RECT 2.880 637.640 83.760 637.960 ;
                RECT 95.680 637.640 106.200 637.960 ;
                RECT 666.880 637.640 671.600 637.960 ;
                RECT 2.880 639.000 106.200 639.320 ;
                RECT 666.880 639.000 671.600 639.320 ;
                RECT 2.880 640.360 83.760 640.680 ;
                RECT 95.680 640.360 106.200 640.680 ;
                RECT 666.880 640.360 671.600 640.680 ;
                RECT 2.880 641.720 86.480 642.040 ;
                RECT 95.680 641.720 106.200 642.040 ;
                RECT 666.880 641.720 671.600 642.040 ;
                RECT 2.880 643.080 83.760 643.400 ;
                RECT 95.680 643.080 106.200 643.400 ;
                RECT 666.880 643.080 671.600 643.400 ;
                RECT 2.880 644.440 83.760 644.760 ;
                RECT 95.680 644.440 106.200 644.760 ;
                RECT 666.880 644.440 671.600 644.760 ;
                RECT 2.880 645.800 83.760 646.120 ;
                RECT 95.680 645.800 106.200 646.120 ;
                RECT 666.880 645.800 671.600 646.120 ;
                RECT 2.880 647.160 106.200 647.480 ;
                RECT 666.880 647.160 671.600 647.480 ;
                RECT 2.880 648.520 83.760 648.840 ;
                RECT 95.680 648.520 106.200 648.840 ;
                RECT 666.880 648.520 671.600 648.840 ;
                RECT 2.880 649.880 83.760 650.200 ;
                RECT 95.680 649.880 106.200 650.200 ;
                RECT 666.880 649.880 671.600 650.200 ;
                RECT 2.880 651.240 88.520 651.560 ;
                RECT 95.680 651.240 106.200 651.560 ;
                RECT 666.880 651.240 671.600 651.560 ;
                RECT 2.880 652.600 83.760 652.920 ;
                RECT 95.680 652.600 106.200 652.920 ;
                RECT 666.880 652.600 671.600 652.920 ;
                RECT 2.880 653.960 83.760 654.280 ;
                RECT 95.680 653.960 106.200 654.280 ;
                RECT 666.880 653.960 671.600 654.280 ;
                RECT 2.880 655.320 106.200 655.640 ;
                RECT 666.880 655.320 671.600 655.640 ;
                RECT 2.880 656.680 83.760 657.000 ;
                RECT 95.680 656.680 106.200 657.000 ;
                RECT 666.880 656.680 671.600 657.000 ;
                RECT 2.880 658.040 83.760 658.360 ;
                RECT 95.680 658.040 106.200 658.360 ;
                RECT 666.880 658.040 671.600 658.360 ;
                RECT 2.880 659.400 83.760 659.720 ;
                RECT 95.680 659.400 106.200 659.720 ;
                RECT 666.880 659.400 671.600 659.720 ;
                RECT 2.880 660.760 91.240 661.080 ;
                RECT 95.680 660.760 106.200 661.080 ;
                RECT 666.880 660.760 671.600 661.080 ;
                RECT 2.880 662.120 106.200 662.440 ;
                RECT 666.880 662.120 671.600 662.440 ;
                RECT 2.880 663.480 106.200 663.800 ;
                RECT 666.880 663.480 671.600 663.800 ;
                RECT 2.880 664.840 83.760 665.160 ;
                RECT 95.680 664.840 106.200 665.160 ;
                RECT 666.880 664.840 671.600 665.160 ;
                RECT 2.880 666.200 83.760 666.520 ;
                RECT 95.680 666.200 106.200 666.520 ;
                RECT 666.880 666.200 671.600 666.520 ;
                RECT 2.880 667.560 83.760 667.880 ;
                RECT 95.680 667.560 106.200 667.880 ;
                RECT 666.880 667.560 671.600 667.880 ;
                RECT 2.880 668.920 83.760 669.240 ;
                RECT 95.680 668.920 106.200 669.240 ;
                RECT 666.880 668.920 671.600 669.240 ;
                RECT 2.880 670.280 106.200 670.600 ;
                RECT 666.880 670.280 671.600 670.600 ;
                RECT 2.880 671.640 85.800 671.960 ;
                RECT 95.680 671.640 106.200 671.960 ;
                RECT 666.880 671.640 671.600 671.960 ;
                RECT 2.880 673.000 84.440 673.320 ;
                RECT 95.680 673.000 106.200 673.320 ;
                RECT 666.880 673.000 671.600 673.320 ;
                RECT 2.880 674.360 84.440 674.680 ;
                RECT 95.680 674.360 106.200 674.680 ;
                RECT 666.880 674.360 671.600 674.680 ;
                RECT 2.880 675.720 84.440 676.040 ;
                RECT 95.680 675.720 106.200 676.040 ;
                RECT 666.880 675.720 671.600 676.040 ;
                RECT 2.880 677.080 84.440 677.400 ;
                RECT 95.680 677.080 106.200 677.400 ;
                RECT 666.880 677.080 671.600 677.400 ;
                RECT 2.880 678.440 106.200 678.760 ;
                RECT 666.880 678.440 671.600 678.760 ;
                RECT 2.880 679.800 84.440 680.120 ;
                RECT 95.680 679.800 106.200 680.120 ;
                RECT 666.880 679.800 671.600 680.120 ;
                RECT 2.880 681.160 88.520 681.480 ;
                RECT 95.680 681.160 106.200 681.480 ;
                RECT 666.880 681.160 671.600 681.480 ;
                RECT 2.880 682.520 84.440 682.840 ;
                RECT 95.680 682.520 106.200 682.840 ;
                RECT 666.880 682.520 671.600 682.840 ;
                RECT 2.880 683.880 84.440 684.200 ;
                RECT 95.680 683.880 106.200 684.200 ;
                RECT 666.880 683.880 671.600 684.200 ;
                RECT 2.880 685.240 84.440 685.560 ;
                RECT 95.680 685.240 106.200 685.560 ;
                RECT 666.880 685.240 671.600 685.560 ;
                RECT 2.880 686.600 106.200 686.920 ;
                RECT 666.880 686.600 671.600 686.920 ;
                RECT 2.880 687.960 84.440 688.280 ;
                RECT 95.680 687.960 106.200 688.280 ;
                RECT 666.880 687.960 671.600 688.280 ;
                RECT 2.880 689.320 84.440 689.640 ;
                RECT 95.680 689.320 106.200 689.640 ;
                RECT 666.880 689.320 671.600 689.640 ;
                RECT 2.880 690.680 90.560 691.000 ;
                RECT 95.680 690.680 106.200 691.000 ;
                RECT 666.880 690.680 671.600 691.000 ;
                RECT 2.880 692.040 84.440 692.360 ;
                RECT 95.680 692.040 106.200 692.360 ;
                RECT 666.880 692.040 671.600 692.360 ;
                RECT 2.880 693.400 84.440 693.720 ;
                RECT 95.680 693.400 106.200 693.720 ;
                RECT 666.880 693.400 671.600 693.720 ;
                RECT 2.880 694.760 106.200 695.080 ;
                RECT 666.880 694.760 671.600 695.080 ;
                RECT 2.880 696.120 84.440 696.440 ;
                RECT 95.680 696.120 106.200 696.440 ;
                RECT 666.880 696.120 671.600 696.440 ;
                RECT 2.880 697.480 84.440 697.800 ;
                RECT 95.680 697.480 106.200 697.800 ;
                RECT 666.880 697.480 671.600 697.800 ;
                RECT 2.880 698.840 84.440 699.160 ;
                RECT 95.680 698.840 106.200 699.160 ;
                RECT 666.880 698.840 671.600 699.160 ;
                RECT 2.880 700.200 93.280 700.520 ;
                RECT 95.680 700.200 106.200 700.520 ;
                RECT 666.880 700.200 671.600 700.520 ;
                RECT 2.880 701.560 84.440 701.880 ;
                RECT 95.680 701.560 106.200 701.880 ;
                RECT 666.880 701.560 671.600 701.880 ;
                RECT 2.880 702.920 106.200 703.240 ;
                RECT 666.880 702.920 671.600 703.240 ;
                RECT 2.880 704.280 85.120 704.600 ;
                RECT 95.680 704.280 106.200 704.600 ;
                RECT 666.880 704.280 671.600 704.600 ;
                RECT 2.880 705.640 85.120 705.960 ;
                RECT 95.680 705.640 106.200 705.960 ;
                RECT 666.880 705.640 671.600 705.960 ;
                RECT 2.880 707.000 85.120 707.320 ;
                RECT 95.680 707.000 106.200 707.320 ;
                RECT 666.880 707.000 671.600 707.320 ;
                RECT 2.880 708.360 85.120 708.680 ;
                RECT 95.680 708.360 106.200 708.680 ;
                RECT 666.880 708.360 671.600 708.680 ;
                RECT 2.880 709.720 106.200 710.040 ;
                RECT 666.880 709.720 671.600 710.040 ;
                RECT 2.880 711.080 87.840 711.400 ;
                RECT 95.680 711.080 106.200 711.400 ;
                RECT 666.880 711.080 671.600 711.400 ;
                RECT 2.880 712.440 85.120 712.760 ;
                RECT 95.680 712.440 106.200 712.760 ;
                RECT 666.880 712.440 671.600 712.760 ;
                RECT 2.880 713.800 85.120 714.120 ;
                RECT 95.680 713.800 106.200 714.120 ;
                RECT 666.880 713.800 671.600 714.120 ;
                RECT 2.880 715.160 85.120 715.480 ;
                RECT 95.680 715.160 106.200 715.480 ;
                RECT 666.880 715.160 671.600 715.480 ;
                RECT 2.880 716.520 85.120 716.840 ;
                RECT 95.680 716.520 106.200 716.840 ;
                RECT 666.880 716.520 671.600 716.840 ;
                RECT 2.880 717.880 106.200 718.200 ;
                RECT 666.880 717.880 671.600 718.200 ;
                RECT 2.880 719.240 89.880 719.560 ;
                RECT 95.680 719.240 106.200 719.560 ;
                RECT 666.880 719.240 671.600 719.560 ;
                RECT 2.880 720.600 90.560 720.920 ;
                RECT 95.680 720.600 106.200 720.920 ;
                RECT 666.880 720.600 671.600 720.920 ;
                RECT 2.880 721.960 85.120 722.280 ;
                RECT 95.680 721.960 106.200 722.280 ;
                RECT 666.880 721.960 671.600 722.280 ;
                RECT 2.880 723.320 85.120 723.640 ;
                RECT 95.680 723.320 106.200 723.640 ;
                RECT 666.880 723.320 671.600 723.640 ;
                RECT 2.880 724.680 85.120 725.000 ;
                RECT 95.680 724.680 106.200 725.000 ;
                RECT 666.880 724.680 671.600 725.000 ;
                RECT 2.880 726.040 106.200 726.360 ;
                RECT 666.880 726.040 671.600 726.360 ;
                RECT 2.880 727.400 85.120 727.720 ;
                RECT 95.680 727.400 106.200 727.720 ;
                RECT 666.880 727.400 671.600 727.720 ;
                RECT 2.880 728.760 85.120 729.080 ;
                RECT 95.680 728.760 106.200 729.080 ;
                RECT 666.880 728.760 671.600 729.080 ;
                RECT 2.880 730.120 92.600 730.440 ;
                RECT 95.680 730.120 106.200 730.440 ;
                RECT 666.880 730.120 671.600 730.440 ;
                RECT 2.880 731.480 85.120 731.800 ;
                RECT 95.680 731.480 106.200 731.800 ;
                RECT 666.880 731.480 671.600 731.800 ;
                RECT 2.880 732.840 85.120 733.160 ;
                RECT 95.680 732.840 106.200 733.160 ;
                RECT 666.880 732.840 671.600 733.160 ;
                RECT 2.880 734.200 106.200 734.520 ;
                RECT 666.880 734.200 671.600 734.520 ;
                RECT 2.880 735.560 85.800 735.880 ;
                RECT 95.680 735.560 106.200 735.880 ;
                RECT 666.880 735.560 671.600 735.880 ;
                RECT 2.880 736.920 85.800 737.240 ;
                RECT 95.680 736.920 106.200 737.240 ;
                RECT 666.880 736.920 671.600 737.240 ;
                RECT 2.880 738.280 85.800 738.600 ;
                RECT 95.680 738.280 106.200 738.600 ;
                RECT 666.880 738.280 671.600 738.600 ;
                RECT 2.880 739.640 87.160 739.960 ;
                RECT 95.680 739.640 106.200 739.960 ;
                RECT 666.880 739.640 671.600 739.960 ;
                RECT 2.880 741.000 85.800 741.320 ;
                RECT 95.680 741.000 106.200 741.320 ;
                RECT 666.880 741.000 671.600 741.320 ;
                RECT 2.880 742.360 106.200 742.680 ;
                RECT 666.880 742.360 671.600 742.680 ;
                RECT 2.880 743.720 85.800 744.040 ;
                RECT 95.680 743.720 106.200 744.040 ;
                RECT 666.880 743.720 671.600 744.040 ;
                RECT 2.880 745.080 85.800 745.400 ;
                RECT 95.680 745.080 106.200 745.400 ;
                RECT 666.880 745.080 671.600 745.400 ;
                RECT 2.880 746.440 85.800 746.760 ;
                RECT 95.680 746.440 106.200 746.760 ;
                RECT 666.880 746.440 671.600 746.760 ;
                RECT 2.880 747.800 85.800 748.120 ;
                RECT 95.680 747.800 106.200 748.120 ;
                RECT 666.880 747.800 671.600 748.120 ;
                RECT 2.880 749.160 106.200 749.480 ;
                RECT 666.880 749.160 671.600 749.480 ;
                RECT 2.880 750.520 89.880 750.840 ;
                RECT 95.680 750.520 106.200 750.840 ;
                RECT 666.880 750.520 671.600 750.840 ;
                RECT 2.880 751.880 85.800 752.200 ;
                RECT 95.680 751.880 106.200 752.200 ;
                RECT 666.880 751.880 671.600 752.200 ;
                RECT 2.880 753.240 85.800 753.560 ;
                RECT 95.680 753.240 106.200 753.560 ;
                RECT 666.880 753.240 671.600 753.560 ;
                RECT 2.880 754.600 85.800 754.920 ;
                RECT 95.680 754.600 106.200 754.920 ;
                RECT 666.880 754.600 671.600 754.920 ;
                RECT 2.880 755.960 85.800 756.280 ;
                RECT 95.680 755.960 106.200 756.280 ;
                RECT 666.880 755.960 671.600 756.280 ;
                RECT 2.880 757.320 106.200 757.640 ;
                RECT 666.880 757.320 671.600 757.640 ;
                RECT 2.880 758.680 91.920 759.000 ;
                RECT 95.680 758.680 106.200 759.000 ;
                RECT 666.880 758.680 671.600 759.000 ;
                RECT 2.880 760.040 85.800 760.360 ;
                RECT 95.680 760.040 106.200 760.360 ;
                RECT 666.880 760.040 671.600 760.360 ;
                RECT 2.880 761.400 85.800 761.720 ;
                RECT 95.680 761.400 106.200 761.720 ;
                RECT 666.880 761.400 671.600 761.720 ;
                RECT 2.880 762.760 85.800 763.080 ;
                RECT 95.680 762.760 106.200 763.080 ;
                RECT 666.880 762.760 671.600 763.080 ;
                RECT 2.880 764.120 85.800 764.440 ;
                RECT 95.680 764.120 106.200 764.440 ;
                RECT 666.880 764.120 671.600 764.440 ;
                RECT 2.880 765.480 106.200 765.800 ;
                RECT 666.880 765.480 671.600 765.800 ;
                RECT 2.880 766.840 298.640 767.160 ;
                RECT 666.880 766.840 671.600 767.160 ;
                RECT 2.880 768.200 298.640 768.520 ;
                RECT 666.880 768.200 671.600 768.520 ;
                RECT 2.880 769.560 298.640 769.880 ;
                RECT 666.880 769.560 671.600 769.880 ;
                RECT 2.880 770.920 671.600 771.240 ;
                RECT 2.880 772.280 671.600 772.600 ;
                RECT 2.880 773.640 671.600 773.960 ;
                RECT 2.880 775.000 671.600 775.320 ;
                RECT 2.880 776.360 671.600 776.680 ;
                RECT 2.880 2.880 671.600 4.240 ;
                RECT 2.880 777.680 671.600 779.040 ;
                RECT 302.780 47.945 308.580 49.065 ;
                RECT 657.080 47.945 662.880 49.065 ;
                RECT 302.780 53.765 308.580 54.455 ;
                RECT 657.080 53.765 662.880 54.455 ;
                RECT 302.780 59.340 308.580 60.130 ;
                RECT 657.080 59.340 662.880 60.130 ;
                RECT 302.780 65.460 308.580 66.040 ;
                RECT 657.080 65.460 662.880 66.040 ;
                RECT 302.780 70.180 308.580 70.770 ;
                RECT 657.080 70.180 662.880 70.770 ;
                RECT 302.780 75.000 308.580 75.590 ;
                RECT 657.080 75.000 662.880 75.590 ;
                RECT 302.780 100.560 662.880 101.360 ;
                RECT 302.780 111.560 662.880 115.160 ;
                RECT 302.780 102.240 662.880 103.040 ;
                RECT 302.780 144.295 662.880 144.585 ;
                RECT 302.780 194.730 662.880 196.530 ;
                RECT 302.780 105.450 662.880 106.250 ;
                RECT 302.780 88.500 662.880 90.300 ;
                RECT 302.780 97.550 662.880 98.350 ;
                RECT 302.780 38.575 662.880 40.375 ;
                RECT 106.640 259.275 108.390 766.455 ;
                RECT 120.625 259.275 122.545 766.455 ;
                RECT 144.400 259.275 146.320 766.455 ;
                RECT 148.240 259.275 150.160 766.455 ;
                RECT 152.080 259.275 154.000 766.455 ;
                RECT 194.650 259.275 196.570 766.455 ;
                RECT 198.490 259.275 200.410 766.455 ;
                RECT 202.330 259.275 204.250 766.455 ;
                RECT 206.170 259.275 208.090 766.455 ;
                RECT 210.010 259.275 211.930 766.455 ;
                RECT 213.850 259.275 215.770 766.455 ;
                RECT 217.690 259.275 219.610 766.455 ;
                RECT 171.885 55.735 172.995 142.735 ;
                RECT 179.400 55.735 180.290 142.735 ;
                RECT 186.375 55.735 187.695 142.735 ;
                RECT 197.565 55.735 199.485 142.735 ;
                RECT 218.345 55.735 220.265 142.735 ;
                RECT 222.185 55.735 224.105 142.735 ;
                RECT 226.025 55.735 227.945 142.735 ;
                RECT 229.865 55.735 231.785 142.735 ;
                RECT 204.225 203.560 205.545 252.640 ;
                RECT 213.350 203.560 214.240 252.640 ;
                RECT 219.680 203.560 220.570 252.640 ;
                RECT 226.010 203.560 227.760 252.640 ;
                RECT 239.150 203.560 241.070 252.640 ;
                RECT 242.990 203.560 244.910 252.640 ;
                RECT 218.925 192.400 220.035 197.560 ;
                RECT 227.730 192.400 229.480 197.560 ;
                RECT 240.870 192.400 242.790 197.560 ;
                RECT 244.710 192.400 246.630 197.560 ;
                RECT 264.285 46.155 265.395 49.735 ;
                RECT 27.350 260.340 36.510 260.710 ;
                RECT 27.350 263.780 36.510 264.890 ;
                RECT 90.190 242.000 109.830 242.670 ;
                RECT 90.190 243.230 109.830 246.280 ;
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 674.480 781.920 ;
        LAYER met2 ;
            RECT 0.000 0.000 674.480 781.920 ;
    END 
END sram22_2048x32m8w8 
END LIBRARY 

