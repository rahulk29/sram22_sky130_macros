VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram22_256x32m4w8
  CLASS BLOCK ;
  ORIGIN 73.425 163.165 ;
  FOREIGN sram22_256x32m4w8 -73.425 -163.165 ;
  SIZE 286.25 BY 294.515 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 196.355 129.945 196.685 131.075 ;
        RECT 196.355 125.635 196.685 125.965 ;
        RECT 196.355 124.275 196.685 124.605 ;
        RECT 196.36 123.6 196.68 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -0.845 196.685 -0.515 ;
        RECT 196.355 -2.205 196.685 -1.875 ;
        RECT 196.355 -3.565 196.685 -3.235 ;
        RECT 196.36 -3.565 196.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -91.965 196.685 -91.635 ;
        RECT 196.355 -93.325 196.685 -92.995 ;
        RECT 196.355 -94.685 196.685 -94.355 ;
        RECT 196.355 -96.045 196.685 -95.715 ;
        RECT 196.355 -97.405 196.685 -97.075 ;
        RECT 196.355 -98.765 196.685 -98.435 ;
        RECT 196.355 -100.125 196.685 -99.795 ;
        RECT 196.355 -101.485 196.685 -101.155 ;
        RECT 196.355 -102.845 196.685 -102.515 ;
        RECT 196.355 -104.205 196.685 -103.875 ;
        RECT 196.355 -105.565 196.685 -105.235 ;
        RECT 196.355 -106.925 196.685 -106.595 ;
        RECT 196.355 -108.285 196.685 -107.955 ;
        RECT 196.355 -109.645 196.685 -109.315 ;
        RECT 196.355 -111.005 196.685 -110.675 ;
        RECT 196.355 -112.365 196.685 -112.035 ;
        RECT 196.355 -113.725 196.685 -113.395 ;
        RECT 196.355 -115.085 196.685 -114.755 ;
        RECT 196.355 -116.445 196.685 -116.115 ;
        RECT 196.355 -117.805 196.685 -117.475 ;
        RECT 196.355 -119.165 196.685 -118.835 ;
        RECT 196.355 -120.525 196.685 -120.195 ;
        RECT 196.355 -121.885 196.685 -121.555 ;
        RECT 196.355 -123.245 196.685 -122.915 ;
        RECT 196.355 -124.605 196.685 -124.275 ;
        RECT 196.355 -125.965 196.685 -125.635 ;
        RECT 196.355 -127.325 196.685 -126.995 ;
        RECT 196.355 -128.685 196.685 -128.355 ;
        RECT 196.355 -130.045 196.685 -129.715 ;
        RECT 196.355 -131.405 196.685 -131.075 ;
        RECT 196.355 -132.765 196.685 -132.435 ;
        RECT 196.355 -134.125 196.685 -133.795 ;
        RECT 196.355 -135.485 196.685 -135.155 ;
        RECT 196.355 -136.845 196.685 -136.515 ;
        RECT 196.355 -138.205 196.685 -137.875 ;
        RECT 196.355 -139.565 196.685 -139.235 ;
        RECT 196.355 -140.925 196.685 -140.595 ;
        RECT 196.355 -142.285 196.685 -141.955 ;
        RECT 196.355 -143.645 196.685 -143.315 ;
        RECT 196.355 -145.005 196.685 -144.675 ;
        RECT 196.355 -146.365 196.685 -146.035 ;
        RECT 196.355 -147.725 196.685 -147.395 ;
        RECT 196.355 -149.085 196.685 -148.755 ;
        RECT 196.355 -150.445 196.685 -150.115 ;
        RECT 196.355 -151.805 196.685 -151.475 ;
        RECT 196.355 -153.165 196.685 -152.835 ;
        RECT 196.355 -154.525 196.685 -154.195 ;
        RECT 196.355 -155.885 196.685 -155.555 ;
        RECT 196.355 -157.245 196.685 -156.915 ;
        RECT 196.355 -162.89 196.685 -161.76 ;
        RECT 196.36 -163.005 196.68 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 129.945 198.045 131.075 ;
        RECT 197.715 125.635 198.045 125.965 ;
        RECT 197.715 124.275 198.045 124.605 ;
        RECT 197.72 123.6 198.04 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 -96.045 198.045 -95.715 ;
        RECT 197.715 -97.405 198.045 -97.075 ;
        RECT 197.715 -98.765 198.045 -98.435 ;
        RECT 197.715 -100.125 198.045 -99.795 ;
        RECT 197.715 -101.485 198.045 -101.155 ;
        RECT 197.715 -102.845 198.045 -102.515 ;
        RECT 197.715 -104.205 198.045 -103.875 ;
        RECT 197.715 -105.565 198.045 -105.235 ;
        RECT 197.715 -106.925 198.045 -106.595 ;
        RECT 197.715 -108.285 198.045 -107.955 ;
        RECT 197.715 -109.645 198.045 -109.315 ;
        RECT 197.715 -111.005 198.045 -110.675 ;
        RECT 197.715 -112.365 198.045 -112.035 ;
        RECT 197.715 -113.725 198.045 -113.395 ;
        RECT 197.715 -115.085 198.045 -114.755 ;
        RECT 197.715 -116.445 198.045 -116.115 ;
        RECT 197.715 -117.805 198.045 -117.475 ;
        RECT 197.715 -119.165 198.045 -118.835 ;
        RECT 197.715 -120.525 198.045 -120.195 ;
        RECT 197.715 -121.885 198.045 -121.555 ;
        RECT 197.715 -123.245 198.045 -122.915 ;
        RECT 197.715 -124.605 198.045 -124.275 ;
        RECT 197.715 -125.965 198.045 -125.635 ;
        RECT 197.715 -127.325 198.045 -126.995 ;
        RECT 197.715 -128.685 198.045 -128.355 ;
        RECT 197.715 -130.045 198.045 -129.715 ;
        RECT 197.715 -131.405 198.045 -131.075 ;
        RECT 197.715 -132.765 198.045 -132.435 ;
        RECT 197.715 -134.125 198.045 -133.795 ;
        RECT 197.715 -135.485 198.045 -135.155 ;
        RECT 197.715 -136.845 198.045 -136.515 ;
        RECT 197.715 -138.205 198.045 -137.875 ;
        RECT 197.715 -139.565 198.045 -139.235 ;
        RECT 197.715 -140.925 198.045 -140.595 ;
        RECT 197.715 -142.285 198.045 -141.955 ;
        RECT 197.715 -143.645 198.045 -143.315 ;
        RECT 197.715 -145.005 198.045 -144.675 ;
        RECT 197.715 -146.365 198.045 -146.035 ;
        RECT 197.715 -147.725 198.045 -147.395 ;
        RECT 197.715 -149.085 198.045 -148.755 ;
        RECT 197.715 -150.445 198.045 -150.115 ;
        RECT 197.715 -151.805 198.045 -151.475 ;
        RECT 197.715 -153.165 198.045 -152.835 ;
        RECT 197.715 -154.525 198.045 -154.195 ;
        RECT 197.715 -155.885 198.045 -155.555 ;
        RECT 197.715 -157.245 198.045 -156.915 ;
        RECT 197.715 -162.89 198.045 -161.76 ;
        RECT 197.72 -163.005 198.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.51 -94.075 198.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 129.945 199.405 131.075 ;
        RECT 199.075 125.635 199.405 125.965 ;
        RECT 199.075 124.275 199.405 124.605 ;
        RECT 199.08 123.6 199.4 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 -96.045 199.405 -95.715 ;
        RECT 199.075 -97.405 199.405 -97.075 ;
        RECT 199.075 -98.765 199.405 -98.435 ;
        RECT 199.075 -100.125 199.405 -99.795 ;
        RECT 199.075 -101.485 199.405 -101.155 ;
        RECT 199.075 -102.845 199.405 -102.515 ;
        RECT 199.075 -104.205 199.405 -103.875 ;
        RECT 199.075 -105.565 199.405 -105.235 ;
        RECT 199.075 -106.925 199.405 -106.595 ;
        RECT 199.075 -108.285 199.405 -107.955 ;
        RECT 199.075 -109.645 199.405 -109.315 ;
        RECT 199.075 -111.005 199.405 -110.675 ;
        RECT 199.075 -112.365 199.405 -112.035 ;
        RECT 199.075 -113.725 199.405 -113.395 ;
        RECT 199.075 -115.085 199.405 -114.755 ;
        RECT 199.075 -116.445 199.405 -116.115 ;
        RECT 199.075 -117.805 199.405 -117.475 ;
        RECT 199.075 -119.165 199.405 -118.835 ;
        RECT 199.075 -120.525 199.405 -120.195 ;
        RECT 199.075 -121.885 199.405 -121.555 ;
        RECT 199.075 -123.245 199.405 -122.915 ;
        RECT 199.075 -124.605 199.405 -124.275 ;
        RECT 199.075 -125.965 199.405 -125.635 ;
        RECT 199.075 -127.325 199.405 -126.995 ;
        RECT 199.075 -128.685 199.405 -128.355 ;
        RECT 199.075 -130.045 199.405 -129.715 ;
        RECT 199.075 -131.405 199.405 -131.075 ;
        RECT 199.075 -132.765 199.405 -132.435 ;
        RECT 199.075 -134.125 199.405 -133.795 ;
        RECT 199.075 -135.485 199.405 -135.155 ;
        RECT 199.075 -136.845 199.405 -136.515 ;
        RECT 199.075 -138.205 199.405 -137.875 ;
        RECT 199.075 -139.565 199.405 -139.235 ;
        RECT 199.075 -140.925 199.405 -140.595 ;
        RECT 199.075 -142.285 199.405 -141.955 ;
        RECT 199.075 -143.645 199.405 -143.315 ;
        RECT 199.075 -145.005 199.405 -144.675 ;
        RECT 199.075 -146.365 199.405 -146.035 ;
        RECT 199.075 -147.725 199.405 -147.395 ;
        RECT 199.075 -149.085 199.405 -148.755 ;
        RECT 199.075 -150.445 199.405 -150.115 ;
        RECT 199.075 -151.805 199.405 -151.475 ;
        RECT 199.075 -153.165 199.405 -152.835 ;
        RECT 199.075 -154.525 199.405 -154.195 ;
        RECT 199.075 -155.885 199.405 -155.555 ;
        RECT 199.075 -157.245 199.405 -156.915 ;
        RECT 199.075 -162.89 199.405 -161.76 ;
        RECT 199.08 -163.005 199.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 129.945 200.765 131.075 ;
        RECT 200.435 125.635 200.765 125.965 ;
        RECT 200.435 124.275 200.765 124.605 ;
        RECT 200.44 123.6 200.76 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 -0.845 200.765 -0.515 ;
        RECT 200.435 -2.205 200.765 -1.875 ;
        RECT 200.435 -3.565 200.765 -3.235 ;
        RECT 200.44 -3.565 200.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 -91.965 200.765 -91.635 ;
        RECT 200.435 -93.325 200.765 -92.995 ;
        RECT 200.435 -94.685 200.765 -94.355 ;
        RECT 200.435 -96.045 200.765 -95.715 ;
        RECT 200.435 -97.405 200.765 -97.075 ;
        RECT 200.435 -98.765 200.765 -98.435 ;
        RECT 200.435 -100.125 200.765 -99.795 ;
        RECT 200.435 -101.485 200.765 -101.155 ;
        RECT 200.435 -102.845 200.765 -102.515 ;
        RECT 200.435 -104.205 200.765 -103.875 ;
        RECT 200.435 -105.565 200.765 -105.235 ;
        RECT 200.435 -106.925 200.765 -106.595 ;
        RECT 200.435 -108.285 200.765 -107.955 ;
        RECT 200.435 -109.645 200.765 -109.315 ;
        RECT 200.435 -111.005 200.765 -110.675 ;
        RECT 200.435 -112.365 200.765 -112.035 ;
        RECT 200.435 -113.725 200.765 -113.395 ;
        RECT 200.435 -115.085 200.765 -114.755 ;
        RECT 200.435 -116.445 200.765 -116.115 ;
        RECT 200.435 -117.805 200.765 -117.475 ;
        RECT 200.435 -119.165 200.765 -118.835 ;
        RECT 200.435 -120.525 200.765 -120.195 ;
        RECT 200.435 -121.885 200.765 -121.555 ;
        RECT 200.435 -123.245 200.765 -122.915 ;
        RECT 200.435 -124.605 200.765 -124.275 ;
        RECT 200.435 -125.965 200.765 -125.635 ;
        RECT 200.435 -127.325 200.765 -126.995 ;
        RECT 200.435 -128.685 200.765 -128.355 ;
        RECT 200.435 -130.045 200.765 -129.715 ;
        RECT 200.435 -131.405 200.765 -131.075 ;
        RECT 200.435 -132.765 200.765 -132.435 ;
        RECT 200.435 -134.125 200.765 -133.795 ;
        RECT 200.435 -135.485 200.765 -135.155 ;
        RECT 200.435 -136.845 200.765 -136.515 ;
        RECT 200.435 -138.205 200.765 -137.875 ;
        RECT 200.435 -139.565 200.765 -139.235 ;
        RECT 200.435 -140.925 200.765 -140.595 ;
        RECT 200.435 -142.285 200.765 -141.955 ;
        RECT 200.435 -143.645 200.765 -143.315 ;
        RECT 200.435 -145.005 200.765 -144.675 ;
        RECT 200.435 -146.365 200.765 -146.035 ;
        RECT 200.435 -147.725 200.765 -147.395 ;
        RECT 200.435 -149.085 200.765 -148.755 ;
        RECT 200.435 -150.445 200.765 -150.115 ;
        RECT 200.435 -151.805 200.765 -151.475 ;
        RECT 200.435 -153.165 200.765 -152.835 ;
        RECT 200.435 -154.525 200.765 -154.195 ;
        RECT 200.435 -155.885 200.765 -155.555 ;
        RECT 200.435 -157.245 200.765 -156.915 ;
        RECT 200.435 -162.89 200.765 -161.76 ;
        RECT 200.44 -163.005 200.76 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 129.945 202.125 131.075 ;
        RECT 201.795 125.635 202.125 125.965 ;
        RECT 201.795 124.275 202.125 124.605 ;
        RECT 201.8 123.6 202.12 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 -0.845 202.125 -0.515 ;
        RECT 201.795 -2.205 202.125 -1.875 ;
        RECT 201.795 -3.565 202.125 -3.235 ;
        RECT 201.8 -3.565 202.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 -91.965 202.125 -91.635 ;
        RECT 201.795 -93.325 202.125 -92.995 ;
        RECT 201.795 -94.685 202.125 -94.355 ;
        RECT 201.795 -96.045 202.125 -95.715 ;
        RECT 201.795 -97.405 202.125 -97.075 ;
        RECT 201.795 -98.765 202.125 -98.435 ;
        RECT 201.795 -100.125 202.125 -99.795 ;
        RECT 201.795 -101.485 202.125 -101.155 ;
        RECT 201.795 -102.845 202.125 -102.515 ;
        RECT 201.795 -104.205 202.125 -103.875 ;
        RECT 201.795 -105.565 202.125 -105.235 ;
        RECT 201.795 -106.925 202.125 -106.595 ;
        RECT 201.795 -108.285 202.125 -107.955 ;
        RECT 201.795 -109.645 202.125 -109.315 ;
        RECT 201.795 -111.005 202.125 -110.675 ;
        RECT 201.795 -112.365 202.125 -112.035 ;
        RECT 201.795 -113.725 202.125 -113.395 ;
        RECT 201.795 -115.085 202.125 -114.755 ;
        RECT 201.795 -116.445 202.125 -116.115 ;
        RECT 201.795 -117.805 202.125 -117.475 ;
        RECT 201.795 -119.165 202.125 -118.835 ;
        RECT 201.795 -120.525 202.125 -120.195 ;
        RECT 201.795 -121.885 202.125 -121.555 ;
        RECT 201.795 -123.245 202.125 -122.915 ;
        RECT 201.795 -124.605 202.125 -124.275 ;
        RECT 201.795 -125.965 202.125 -125.635 ;
        RECT 201.795 -127.325 202.125 -126.995 ;
        RECT 201.795 -128.685 202.125 -128.355 ;
        RECT 201.795 -130.045 202.125 -129.715 ;
        RECT 201.795 -131.405 202.125 -131.075 ;
        RECT 201.795 -132.765 202.125 -132.435 ;
        RECT 201.795 -134.125 202.125 -133.795 ;
        RECT 201.795 -135.485 202.125 -135.155 ;
        RECT 201.795 -136.845 202.125 -136.515 ;
        RECT 201.795 -138.205 202.125 -137.875 ;
        RECT 201.795 -139.565 202.125 -139.235 ;
        RECT 201.795 -140.925 202.125 -140.595 ;
        RECT 201.795 -142.285 202.125 -141.955 ;
        RECT 201.795 -143.645 202.125 -143.315 ;
        RECT 201.795 -145.005 202.125 -144.675 ;
        RECT 201.795 -146.365 202.125 -146.035 ;
        RECT 201.795 -147.725 202.125 -147.395 ;
        RECT 201.795 -149.085 202.125 -148.755 ;
        RECT 201.795 -150.445 202.125 -150.115 ;
        RECT 201.795 -151.805 202.125 -151.475 ;
        RECT 201.795 -153.165 202.125 -152.835 ;
        RECT 201.795 -154.525 202.125 -154.195 ;
        RECT 201.795 -155.885 202.125 -155.555 ;
        RECT 201.795 -157.245 202.125 -156.915 ;
        RECT 201.795 -162.89 202.125 -161.76 ;
        RECT 201.8 -163.005 202.12 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 129.945 203.485 131.075 ;
        RECT 203.155 125.635 203.485 125.965 ;
        RECT 203.155 124.275 203.485 124.605 ;
        RECT 203.155 121.41 203.485 121.74 ;
        RECT 203.155 119.235 203.485 119.565 ;
        RECT 203.155 117.655 203.485 117.985 ;
        RECT 203.155 116.805 203.485 117.135 ;
        RECT 203.155 114.495 203.485 114.825 ;
        RECT 203.155 113.645 203.485 113.975 ;
        RECT 203.155 111.335 203.485 111.665 ;
        RECT 203.155 110.485 203.485 110.815 ;
        RECT 203.155 108.175 203.485 108.505 ;
        RECT 203.155 107.325 203.485 107.655 ;
        RECT 203.155 105.015 203.485 105.345 ;
        RECT 203.155 103.435 203.485 103.765 ;
        RECT 203.155 102.585 203.485 102.915 ;
        RECT 203.155 100.275 203.485 100.605 ;
        RECT 203.155 99.425 203.485 99.755 ;
        RECT 203.155 97.115 203.485 97.445 ;
        RECT 203.155 96.265 203.485 96.595 ;
        RECT 203.155 93.955 203.485 94.285 ;
        RECT 203.155 93.105 203.485 93.435 ;
        RECT 203.155 90.795 203.485 91.125 ;
        RECT 203.155 89.215 203.485 89.545 ;
        RECT 203.155 88.365 203.485 88.695 ;
        RECT 203.155 86.055 203.485 86.385 ;
        RECT 203.155 85.205 203.485 85.535 ;
        RECT 203.155 82.895 203.485 83.225 ;
        RECT 203.155 82.045 203.485 82.375 ;
        RECT 203.155 79.735 203.485 80.065 ;
        RECT 203.155 78.885 203.485 79.215 ;
        RECT 203.155 76.575 203.485 76.905 ;
        RECT 203.155 74.995 203.485 75.325 ;
        RECT 203.155 74.145 203.485 74.475 ;
        RECT 203.155 71.835 203.485 72.165 ;
        RECT 203.155 70.985 203.485 71.315 ;
        RECT 203.155 68.675 203.485 69.005 ;
        RECT 203.155 67.825 203.485 68.155 ;
        RECT 203.155 65.515 203.485 65.845 ;
        RECT 203.155 64.665 203.485 64.995 ;
        RECT 203.155 62.355 203.485 62.685 ;
        RECT 203.155 60.775 203.485 61.105 ;
        RECT 203.155 59.925 203.485 60.255 ;
        RECT 203.155 57.615 203.485 57.945 ;
        RECT 203.155 56.765 203.485 57.095 ;
        RECT 203.155 54.455 203.485 54.785 ;
        RECT 203.155 53.605 203.485 53.935 ;
        RECT 203.155 51.295 203.485 51.625 ;
        RECT 203.155 50.445 203.485 50.775 ;
        RECT 203.155 48.135 203.485 48.465 ;
        RECT 203.155 46.555 203.485 46.885 ;
        RECT 203.155 45.705 203.485 46.035 ;
        RECT 203.155 43.395 203.485 43.725 ;
        RECT 203.155 42.545 203.485 42.875 ;
        RECT 203.155 40.235 203.485 40.565 ;
        RECT 203.155 39.385 203.485 39.715 ;
        RECT 203.155 37.075 203.485 37.405 ;
        RECT 203.155 36.225 203.485 36.555 ;
        RECT 203.155 33.915 203.485 34.245 ;
        RECT 203.155 32.335 203.485 32.665 ;
        RECT 203.155 31.485 203.485 31.815 ;
        RECT 203.155 29.175 203.485 29.505 ;
        RECT 203.155 28.325 203.485 28.655 ;
        RECT 203.155 26.015 203.485 26.345 ;
        RECT 203.155 25.165 203.485 25.495 ;
        RECT 203.155 22.855 203.485 23.185 ;
        RECT 203.155 22.005 203.485 22.335 ;
        RECT 203.155 19.695 203.485 20.025 ;
        RECT 203.155 18.115 203.485 18.445 ;
        RECT 203.155 17.265 203.485 17.595 ;
        RECT 203.155 14.955 203.485 15.285 ;
        RECT 203.155 14.105 203.485 14.435 ;
        RECT 203.155 11.795 203.485 12.125 ;
        RECT 203.155 10.945 203.485 11.275 ;
        RECT 203.155 8.635 203.485 8.965 ;
        RECT 203.155 7.785 203.485 8.115 ;
        RECT 203.155 5.475 203.485 5.805 ;
        RECT 203.155 3.895 203.485 4.225 ;
        RECT 203.155 3.045 203.485 3.375 ;
        RECT 203.155 0.87 203.485 1.2 ;
        RECT 203.155 -0.845 203.485 -0.515 ;
        RECT 203.155 -2.205 203.485 -1.875 ;
        RECT 203.155 -3.565 203.485 -3.235 ;
        RECT 203.155 -4.925 203.485 -4.595 ;
        RECT 203.155 -6.285 203.485 -5.955 ;
        RECT 203.155 -7.645 203.485 -7.315 ;
        RECT 203.155 -9.005 203.485 -8.675 ;
        RECT 203.155 -10.365 203.485 -10.035 ;
        RECT 203.155 -11.725 203.485 -11.395 ;
        RECT 203.155 -13.085 203.485 -12.755 ;
        RECT 203.155 -14.445 203.485 -14.115 ;
        RECT 203.155 -15.805 203.485 -15.475 ;
        RECT 203.155 -17.165 203.485 -16.835 ;
        RECT 203.155 -18.525 203.485 -18.195 ;
        RECT 203.155 -19.885 203.485 -19.555 ;
        RECT 203.155 -21.245 203.485 -20.915 ;
        RECT 203.155 -22.605 203.485 -22.275 ;
        RECT 203.155 -23.965 203.485 -23.635 ;
        RECT 203.155 -25.325 203.485 -24.995 ;
        RECT 203.155 -26.685 203.485 -26.355 ;
        RECT 203.155 -28.045 203.485 -27.715 ;
        RECT 203.155 -29.405 203.485 -29.075 ;
        RECT 203.155 -30.765 203.485 -30.435 ;
        RECT 203.155 -32.125 203.485 -31.795 ;
        RECT 203.155 -33.485 203.485 -33.155 ;
        RECT 203.155 -34.845 203.485 -34.515 ;
        RECT 203.155 -36.205 203.485 -35.875 ;
        RECT 203.155 -37.565 203.485 -37.235 ;
        RECT 203.155 -38.925 203.485 -38.595 ;
        RECT 203.155 -40.285 203.485 -39.955 ;
        RECT 203.155 -41.645 203.485 -41.315 ;
        RECT 203.155 -43.005 203.485 -42.675 ;
        RECT 203.155 -44.365 203.485 -44.035 ;
        RECT 203.155 -45.725 203.485 -45.395 ;
        RECT 203.155 -47.085 203.485 -46.755 ;
        RECT 203.155 -48.445 203.485 -48.115 ;
        RECT 203.155 -49.805 203.485 -49.475 ;
        RECT 203.155 -51.165 203.485 -50.835 ;
        RECT 203.155 -52.525 203.485 -52.195 ;
        RECT 203.155 -53.885 203.485 -53.555 ;
        RECT 203.155 -55.245 203.485 -54.915 ;
        RECT 203.155 -56.605 203.485 -56.275 ;
        RECT 203.155 -57.965 203.485 -57.635 ;
        RECT 203.155 -59.325 203.485 -58.995 ;
        RECT 203.155 -60.685 203.485 -60.355 ;
        RECT 203.155 -62.045 203.485 -61.715 ;
        RECT 203.155 -63.405 203.485 -63.075 ;
        RECT 203.155 -64.765 203.485 -64.435 ;
        RECT 203.155 -66.125 203.485 -65.795 ;
        RECT 203.155 -67.485 203.485 -67.155 ;
        RECT 203.155 -68.845 203.485 -68.515 ;
        RECT 203.155 -70.205 203.485 -69.875 ;
        RECT 203.155 -71.565 203.485 -71.235 ;
        RECT 203.155 -72.925 203.485 -72.595 ;
        RECT 203.155 -74.285 203.485 -73.955 ;
        RECT 203.155 -75.645 203.485 -75.315 ;
        RECT 203.155 -77.005 203.485 -76.675 ;
        RECT 203.155 -78.365 203.485 -78.035 ;
        RECT 203.155 -79.725 203.485 -79.395 ;
        RECT 203.155 -81.085 203.485 -80.755 ;
        RECT 203.155 -82.445 203.485 -82.115 ;
        RECT 203.155 -83.805 203.485 -83.475 ;
        RECT 203.155 -85.165 203.485 -84.835 ;
        RECT 203.155 -86.525 203.485 -86.195 ;
        RECT 203.155 -87.885 203.485 -87.555 ;
        RECT 203.155 -89.245 203.485 -88.915 ;
        RECT 203.155 -90.605 203.485 -90.275 ;
        RECT 203.155 -91.965 203.485 -91.635 ;
        RECT 203.155 -93.325 203.485 -92.995 ;
        RECT 203.155 -94.685 203.485 -94.355 ;
        RECT 203.155 -96.045 203.485 -95.715 ;
        RECT 203.155 -97.405 203.485 -97.075 ;
        RECT 203.155 -98.765 203.485 -98.435 ;
        RECT 203.155 -100.125 203.485 -99.795 ;
        RECT 203.155 -101.485 203.485 -101.155 ;
        RECT 203.155 -102.845 203.485 -102.515 ;
        RECT 203.155 -104.205 203.485 -103.875 ;
        RECT 203.155 -105.565 203.485 -105.235 ;
        RECT 203.155 -106.925 203.485 -106.595 ;
        RECT 203.155 -108.285 203.485 -107.955 ;
        RECT 203.155 -109.645 203.485 -109.315 ;
        RECT 203.155 -111.005 203.485 -110.675 ;
        RECT 203.155 -112.365 203.485 -112.035 ;
        RECT 203.155 -113.725 203.485 -113.395 ;
        RECT 203.155 -115.085 203.485 -114.755 ;
        RECT 203.155 -116.445 203.485 -116.115 ;
        RECT 203.155 -117.805 203.485 -117.475 ;
        RECT 203.155 -119.165 203.485 -118.835 ;
        RECT 203.155 -120.525 203.485 -120.195 ;
        RECT 203.155 -121.885 203.485 -121.555 ;
        RECT 203.155 -123.245 203.485 -122.915 ;
        RECT 203.155 -124.605 203.485 -124.275 ;
        RECT 203.155 -125.965 203.485 -125.635 ;
        RECT 203.155 -127.325 203.485 -126.995 ;
        RECT 203.155 -128.685 203.485 -128.355 ;
        RECT 203.155 -130.045 203.485 -129.715 ;
        RECT 203.155 -131.405 203.485 -131.075 ;
        RECT 203.155 -132.765 203.485 -132.435 ;
        RECT 203.155 -134.125 203.485 -133.795 ;
        RECT 203.155 -135.485 203.485 -135.155 ;
        RECT 203.155 -136.845 203.485 -136.515 ;
        RECT 203.155 -138.205 203.485 -137.875 ;
        RECT 203.155 -139.565 203.485 -139.235 ;
        RECT 203.155 -140.925 203.485 -140.595 ;
        RECT 203.155 -142.285 203.485 -141.955 ;
        RECT 203.155 -143.645 203.485 -143.315 ;
        RECT 203.155 -145.005 203.485 -144.675 ;
        RECT 203.155 -146.365 203.485 -146.035 ;
        RECT 203.155 -147.725 203.485 -147.395 ;
        RECT 203.155 -149.085 203.485 -148.755 ;
        RECT 203.155 -150.445 203.485 -150.115 ;
        RECT 203.155 -151.805 203.485 -151.475 ;
        RECT 203.155 -153.165 203.485 -152.835 ;
        RECT 203.155 -154.525 203.485 -154.195 ;
        RECT 203.155 -155.885 203.485 -155.555 ;
        RECT 203.155 -157.245 203.485 -156.915 ;
        RECT 203.155 -162.89 203.485 -161.76 ;
        RECT 203.16 -163.005 203.48 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 129.945 204.845 131.075 ;
        RECT 204.515 125.635 204.845 125.965 ;
        RECT 204.515 124.275 204.845 124.605 ;
        RECT 204.515 121.41 204.845 121.74 ;
        RECT 204.515 119.235 204.845 119.565 ;
        RECT 204.515 117.655 204.845 117.985 ;
        RECT 204.515 116.805 204.845 117.135 ;
        RECT 204.515 114.495 204.845 114.825 ;
        RECT 204.515 113.645 204.845 113.975 ;
        RECT 204.515 111.335 204.845 111.665 ;
        RECT 204.515 110.485 204.845 110.815 ;
        RECT 204.515 108.175 204.845 108.505 ;
        RECT 204.515 107.325 204.845 107.655 ;
        RECT 204.515 105.015 204.845 105.345 ;
        RECT 204.515 103.435 204.845 103.765 ;
        RECT 204.515 102.585 204.845 102.915 ;
        RECT 204.515 100.275 204.845 100.605 ;
        RECT 204.515 99.425 204.845 99.755 ;
        RECT 204.515 97.115 204.845 97.445 ;
        RECT 204.515 96.265 204.845 96.595 ;
        RECT 204.515 93.955 204.845 94.285 ;
        RECT 204.515 93.105 204.845 93.435 ;
        RECT 204.515 90.795 204.845 91.125 ;
        RECT 204.515 89.215 204.845 89.545 ;
        RECT 204.515 88.365 204.845 88.695 ;
        RECT 204.515 86.055 204.845 86.385 ;
        RECT 204.515 85.205 204.845 85.535 ;
        RECT 204.515 82.895 204.845 83.225 ;
        RECT 204.515 82.045 204.845 82.375 ;
        RECT 204.515 79.735 204.845 80.065 ;
        RECT 204.515 78.885 204.845 79.215 ;
        RECT 204.515 76.575 204.845 76.905 ;
        RECT 204.515 74.995 204.845 75.325 ;
        RECT 204.515 74.145 204.845 74.475 ;
        RECT 204.515 71.835 204.845 72.165 ;
        RECT 204.515 70.985 204.845 71.315 ;
        RECT 204.515 68.675 204.845 69.005 ;
        RECT 204.515 67.825 204.845 68.155 ;
        RECT 204.515 65.515 204.845 65.845 ;
        RECT 204.515 64.665 204.845 64.995 ;
        RECT 204.515 62.355 204.845 62.685 ;
        RECT 204.515 60.775 204.845 61.105 ;
        RECT 204.515 59.925 204.845 60.255 ;
        RECT 204.515 57.615 204.845 57.945 ;
        RECT 204.515 56.765 204.845 57.095 ;
        RECT 204.515 54.455 204.845 54.785 ;
        RECT 204.515 53.605 204.845 53.935 ;
        RECT 204.515 51.295 204.845 51.625 ;
        RECT 204.515 50.445 204.845 50.775 ;
        RECT 204.515 48.135 204.845 48.465 ;
        RECT 204.515 46.555 204.845 46.885 ;
        RECT 204.515 45.705 204.845 46.035 ;
        RECT 204.515 43.395 204.845 43.725 ;
        RECT 204.515 42.545 204.845 42.875 ;
        RECT 204.515 40.235 204.845 40.565 ;
        RECT 204.515 39.385 204.845 39.715 ;
        RECT 204.515 37.075 204.845 37.405 ;
        RECT 204.515 36.225 204.845 36.555 ;
        RECT 204.515 33.915 204.845 34.245 ;
        RECT 204.515 32.335 204.845 32.665 ;
        RECT 204.515 31.485 204.845 31.815 ;
        RECT 204.515 29.175 204.845 29.505 ;
        RECT 204.515 28.325 204.845 28.655 ;
        RECT 204.515 26.015 204.845 26.345 ;
        RECT 204.515 25.165 204.845 25.495 ;
        RECT 204.515 22.855 204.845 23.185 ;
        RECT 204.515 22.005 204.845 22.335 ;
        RECT 204.515 19.695 204.845 20.025 ;
        RECT 204.515 18.115 204.845 18.445 ;
        RECT 204.515 17.265 204.845 17.595 ;
        RECT 204.515 14.955 204.845 15.285 ;
        RECT 204.515 14.105 204.845 14.435 ;
        RECT 204.515 11.795 204.845 12.125 ;
        RECT 204.515 10.945 204.845 11.275 ;
        RECT 204.515 8.635 204.845 8.965 ;
        RECT 204.515 7.785 204.845 8.115 ;
        RECT 204.515 5.475 204.845 5.805 ;
        RECT 204.515 3.895 204.845 4.225 ;
        RECT 204.515 3.045 204.845 3.375 ;
        RECT 204.515 0.87 204.845 1.2 ;
        RECT 204.515 -0.845 204.845 -0.515 ;
        RECT 204.515 -2.205 204.845 -1.875 ;
        RECT 204.515 -3.565 204.845 -3.235 ;
        RECT 204.515 -4.925 204.845 -4.595 ;
        RECT 204.515 -6.285 204.845 -5.955 ;
        RECT 204.515 -7.645 204.845 -7.315 ;
        RECT 204.515 -9.005 204.845 -8.675 ;
        RECT 204.515 -10.365 204.845 -10.035 ;
        RECT 204.515 -11.725 204.845 -11.395 ;
        RECT 204.515 -13.085 204.845 -12.755 ;
        RECT 204.515 -14.445 204.845 -14.115 ;
        RECT 204.515 -15.805 204.845 -15.475 ;
        RECT 204.515 -17.165 204.845 -16.835 ;
        RECT 204.515 -18.525 204.845 -18.195 ;
        RECT 204.515 -19.885 204.845 -19.555 ;
        RECT 204.515 -21.245 204.845 -20.915 ;
        RECT 204.515 -22.605 204.845 -22.275 ;
        RECT 204.515 -23.965 204.845 -23.635 ;
        RECT 204.515 -25.325 204.845 -24.995 ;
        RECT 204.515 -26.685 204.845 -26.355 ;
        RECT 204.515 -28.045 204.845 -27.715 ;
        RECT 204.515 -29.405 204.845 -29.075 ;
        RECT 204.515 -30.765 204.845 -30.435 ;
        RECT 204.515 -32.125 204.845 -31.795 ;
        RECT 204.515 -33.485 204.845 -33.155 ;
        RECT 204.515 -34.845 204.845 -34.515 ;
        RECT 204.515 -36.205 204.845 -35.875 ;
        RECT 204.515 -37.565 204.845 -37.235 ;
        RECT 204.515 -38.925 204.845 -38.595 ;
        RECT 204.515 -40.285 204.845 -39.955 ;
        RECT 204.515 -41.645 204.845 -41.315 ;
        RECT 204.515 -43.005 204.845 -42.675 ;
        RECT 204.515 -44.365 204.845 -44.035 ;
        RECT 204.515 -45.725 204.845 -45.395 ;
        RECT 204.515 -47.085 204.845 -46.755 ;
        RECT 204.515 -48.445 204.845 -48.115 ;
        RECT 204.515 -49.805 204.845 -49.475 ;
        RECT 204.515 -51.165 204.845 -50.835 ;
        RECT 204.515 -52.525 204.845 -52.195 ;
        RECT 204.515 -53.885 204.845 -53.555 ;
        RECT 204.515 -55.245 204.845 -54.915 ;
        RECT 204.515 -56.605 204.845 -56.275 ;
        RECT 204.515 -57.965 204.845 -57.635 ;
        RECT 204.515 -59.325 204.845 -58.995 ;
        RECT 204.515 -60.685 204.845 -60.355 ;
        RECT 204.515 -62.045 204.845 -61.715 ;
        RECT 204.515 -63.405 204.845 -63.075 ;
        RECT 204.515 -64.765 204.845 -64.435 ;
        RECT 204.515 -66.125 204.845 -65.795 ;
        RECT 204.515 -67.485 204.845 -67.155 ;
        RECT 204.515 -68.845 204.845 -68.515 ;
        RECT 204.515 -70.205 204.845 -69.875 ;
        RECT 204.515 -71.565 204.845 -71.235 ;
        RECT 204.515 -72.925 204.845 -72.595 ;
        RECT 204.515 -74.285 204.845 -73.955 ;
        RECT 204.515 -75.645 204.845 -75.315 ;
        RECT 204.515 -77.005 204.845 -76.675 ;
        RECT 204.515 -78.365 204.845 -78.035 ;
        RECT 204.515 -79.725 204.845 -79.395 ;
        RECT 204.515 -81.085 204.845 -80.755 ;
        RECT 204.515 -82.445 204.845 -82.115 ;
        RECT 204.515 -83.805 204.845 -83.475 ;
        RECT 204.515 -85.165 204.845 -84.835 ;
        RECT 204.515 -86.525 204.845 -86.195 ;
        RECT 204.515 -87.885 204.845 -87.555 ;
        RECT 204.515 -89.245 204.845 -88.915 ;
        RECT 204.515 -90.605 204.845 -90.275 ;
        RECT 204.515 -91.965 204.845 -91.635 ;
        RECT 204.515 -93.325 204.845 -92.995 ;
        RECT 204.515 -94.685 204.845 -94.355 ;
        RECT 204.515 -96.045 204.845 -95.715 ;
        RECT 204.515 -97.405 204.845 -97.075 ;
        RECT 204.515 -98.765 204.845 -98.435 ;
        RECT 204.515 -100.125 204.845 -99.795 ;
        RECT 204.515 -101.485 204.845 -101.155 ;
        RECT 204.515 -102.845 204.845 -102.515 ;
        RECT 204.515 -104.205 204.845 -103.875 ;
        RECT 204.515 -105.565 204.845 -105.235 ;
        RECT 204.515 -106.925 204.845 -106.595 ;
        RECT 204.515 -108.285 204.845 -107.955 ;
        RECT 204.515 -109.645 204.845 -109.315 ;
        RECT 204.515 -111.005 204.845 -110.675 ;
        RECT 204.515 -112.365 204.845 -112.035 ;
        RECT 204.515 -113.725 204.845 -113.395 ;
        RECT 204.515 -115.085 204.845 -114.755 ;
        RECT 204.515 -116.445 204.845 -116.115 ;
        RECT 204.515 -117.805 204.845 -117.475 ;
        RECT 204.515 -119.165 204.845 -118.835 ;
        RECT 204.515 -120.525 204.845 -120.195 ;
        RECT 204.515 -121.885 204.845 -121.555 ;
        RECT 204.515 -123.245 204.845 -122.915 ;
        RECT 204.515 -124.605 204.845 -124.275 ;
        RECT 204.515 -125.965 204.845 -125.635 ;
        RECT 204.515 -127.325 204.845 -126.995 ;
        RECT 204.515 -128.685 204.845 -128.355 ;
        RECT 204.515 -130.045 204.845 -129.715 ;
        RECT 204.515 -131.405 204.845 -131.075 ;
        RECT 204.515 -132.765 204.845 -132.435 ;
        RECT 204.515 -134.125 204.845 -133.795 ;
        RECT 204.515 -135.485 204.845 -135.155 ;
        RECT 204.515 -136.845 204.845 -136.515 ;
        RECT 204.515 -138.205 204.845 -137.875 ;
        RECT 204.515 -139.565 204.845 -139.235 ;
        RECT 204.515 -140.925 204.845 -140.595 ;
        RECT 204.515 -142.285 204.845 -141.955 ;
        RECT 204.515 -143.645 204.845 -143.315 ;
        RECT 204.515 -145.005 204.845 -144.675 ;
        RECT 204.515 -146.365 204.845 -146.035 ;
        RECT 204.515 -147.725 204.845 -147.395 ;
        RECT 204.515 -149.085 204.845 -148.755 ;
        RECT 204.515 -150.445 204.845 -150.115 ;
        RECT 204.515 -151.805 204.845 -151.475 ;
        RECT 204.515 -153.165 204.845 -152.835 ;
        RECT 204.515 -154.525 204.845 -154.195 ;
        RECT 204.515 -155.885 204.845 -155.555 ;
        RECT 204.515 -157.245 204.845 -156.915 ;
        RECT 204.515 -162.89 204.845 -161.76 ;
        RECT 204.52 -163.005 204.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 129.945 206.205 131.075 ;
        RECT 205.875 125.635 206.205 125.965 ;
        RECT 205.875 124.275 206.205 124.605 ;
        RECT 205.875 121.41 206.205 121.74 ;
        RECT 205.875 119.235 206.205 119.565 ;
        RECT 205.875 117.655 206.205 117.985 ;
        RECT 205.875 116.805 206.205 117.135 ;
        RECT 205.875 114.495 206.205 114.825 ;
        RECT 205.875 113.645 206.205 113.975 ;
        RECT 205.875 111.335 206.205 111.665 ;
        RECT 205.875 110.485 206.205 110.815 ;
        RECT 205.875 108.175 206.205 108.505 ;
        RECT 205.875 107.325 206.205 107.655 ;
        RECT 205.875 105.015 206.205 105.345 ;
        RECT 205.875 103.435 206.205 103.765 ;
        RECT 205.875 102.585 206.205 102.915 ;
        RECT 205.875 100.275 206.205 100.605 ;
        RECT 205.875 99.425 206.205 99.755 ;
        RECT 205.875 97.115 206.205 97.445 ;
        RECT 205.875 96.265 206.205 96.595 ;
        RECT 205.875 93.955 206.205 94.285 ;
        RECT 205.875 93.105 206.205 93.435 ;
        RECT 205.875 90.795 206.205 91.125 ;
        RECT 205.875 89.215 206.205 89.545 ;
        RECT 205.875 88.365 206.205 88.695 ;
        RECT 205.875 86.055 206.205 86.385 ;
        RECT 205.875 85.205 206.205 85.535 ;
        RECT 205.875 82.895 206.205 83.225 ;
        RECT 205.875 82.045 206.205 82.375 ;
        RECT 205.875 79.735 206.205 80.065 ;
        RECT 205.875 78.885 206.205 79.215 ;
        RECT 205.875 76.575 206.205 76.905 ;
        RECT 205.875 74.995 206.205 75.325 ;
        RECT 205.875 74.145 206.205 74.475 ;
        RECT 205.875 71.835 206.205 72.165 ;
        RECT 205.875 70.985 206.205 71.315 ;
        RECT 205.875 68.675 206.205 69.005 ;
        RECT 205.875 67.825 206.205 68.155 ;
        RECT 205.875 65.515 206.205 65.845 ;
        RECT 205.875 64.665 206.205 64.995 ;
        RECT 205.875 62.355 206.205 62.685 ;
        RECT 205.875 60.775 206.205 61.105 ;
        RECT 205.875 59.925 206.205 60.255 ;
        RECT 205.875 57.615 206.205 57.945 ;
        RECT 205.875 56.765 206.205 57.095 ;
        RECT 205.875 54.455 206.205 54.785 ;
        RECT 205.875 53.605 206.205 53.935 ;
        RECT 205.875 51.295 206.205 51.625 ;
        RECT 205.875 50.445 206.205 50.775 ;
        RECT 205.875 48.135 206.205 48.465 ;
        RECT 205.875 46.555 206.205 46.885 ;
        RECT 205.875 45.705 206.205 46.035 ;
        RECT 205.875 43.395 206.205 43.725 ;
        RECT 205.875 42.545 206.205 42.875 ;
        RECT 205.875 40.235 206.205 40.565 ;
        RECT 205.875 39.385 206.205 39.715 ;
        RECT 205.875 37.075 206.205 37.405 ;
        RECT 205.875 36.225 206.205 36.555 ;
        RECT 205.875 33.915 206.205 34.245 ;
        RECT 205.875 32.335 206.205 32.665 ;
        RECT 205.875 31.485 206.205 31.815 ;
        RECT 205.875 29.175 206.205 29.505 ;
        RECT 205.875 28.325 206.205 28.655 ;
        RECT 205.875 26.015 206.205 26.345 ;
        RECT 205.875 25.165 206.205 25.495 ;
        RECT 205.875 22.855 206.205 23.185 ;
        RECT 205.875 22.005 206.205 22.335 ;
        RECT 205.875 19.695 206.205 20.025 ;
        RECT 205.875 18.115 206.205 18.445 ;
        RECT 205.875 17.265 206.205 17.595 ;
        RECT 205.875 14.955 206.205 15.285 ;
        RECT 205.875 14.105 206.205 14.435 ;
        RECT 205.875 11.795 206.205 12.125 ;
        RECT 205.875 10.945 206.205 11.275 ;
        RECT 205.875 8.635 206.205 8.965 ;
        RECT 205.875 7.785 206.205 8.115 ;
        RECT 205.875 5.475 206.205 5.805 ;
        RECT 205.875 3.895 206.205 4.225 ;
        RECT 205.875 3.045 206.205 3.375 ;
        RECT 205.875 0.87 206.205 1.2 ;
        RECT 205.875 -0.845 206.205 -0.515 ;
        RECT 205.875 -2.205 206.205 -1.875 ;
        RECT 205.875 -3.565 206.205 -3.235 ;
        RECT 205.875 -4.925 206.205 -4.595 ;
        RECT 205.875 -6.285 206.205 -5.955 ;
        RECT 205.875 -7.645 206.205 -7.315 ;
        RECT 205.875 -9.005 206.205 -8.675 ;
        RECT 205.875 -10.365 206.205 -10.035 ;
        RECT 205.875 -11.725 206.205 -11.395 ;
        RECT 205.875 -13.085 206.205 -12.755 ;
        RECT 205.875 -14.445 206.205 -14.115 ;
        RECT 205.875 -15.805 206.205 -15.475 ;
        RECT 205.875 -17.165 206.205 -16.835 ;
        RECT 205.875 -18.525 206.205 -18.195 ;
        RECT 205.875 -19.885 206.205 -19.555 ;
        RECT 205.875 -21.245 206.205 -20.915 ;
        RECT 205.875 -22.605 206.205 -22.275 ;
        RECT 205.875 -23.965 206.205 -23.635 ;
        RECT 205.875 -25.325 206.205 -24.995 ;
        RECT 205.875 -26.685 206.205 -26.355 ;
        RECT 205.875 -28.045 206.205 -27.715 ;
        RECT 205.875 -29.405 206.205 -29.075 ;
        RECT 205.875 -30.765 206.205 -30.435 ;
        RECT 205.875 -32.125 206.205 -31.795 ;
        RECT 205.875 -33.485 206.205 -33.155 ;
        RECT 205.875 -34.845 206.205 -34.515 ;
        RECT 205.875 -36.205 206.205 -35.875 ;
        RECT 205.875 -37.565 206.205 -37.235 ;
        RECT 205.875 -38.925 206.205 -38.595 ;
        RECT 205.875 -40.285 206.205 -39.955 ;
        RECT 205.875 -41.645 206.205 -41.315 ;
        RECT 205.875 -43.005 206.205 -42.675 ;
        RECT 205.875 -44.365 206.205 -44.035 ;
        RECT 205.875 -45.725 206.205 -45.395 ;
        RECT 205.875 -47.085 206.205 -46.755 ;
        RECT 205.875 -48.445 206.205 -48.115 ;
        RECT 205.875 -49.805 206.205 -49.475 ;
        RECT 205.875 -51.165 206.205 -50.835 ;
        RECT 205.875 -52.525 206.205 -52.195 ;
        RECT 205.875 -53.885 206.205 -53.555 ;
        RECT 205.875 -55.245 206.205 -54.915 ;
        RECT 205.875 -56.605 206.205 -56.275 ;
        RECT 205.875 -57.965 206.205 -57.635 ;
        RECT 205.875 -59.325 206.205 -58.995 ;
        RECT 205.875 -60.685 206.205 -60.355 ;
        RECT 205.875 -62.045 206.205 -61.715 ;
        RECT 205.875 -63.405 206.205 -63.075 ;
        RECT 205.875 -64.765 206.205 -64.435 ;
        RECT 205.875 -66.125 206.205 -65.795 ;
        RECT 205.875 -67.485 206.205 -67.155 ;
        RECT 205.875 -68.845 206.205 -68.515 ;
        RECT 205.875 -70.205 206.205 -69.875 ;
        RECT 205.875 -71.565 206.205 -71.235 ;
        RECT 205.875 -72.925 206.205 -72.595 ;
        RECT 205.875 -74.285 206.205 -73.955 ;
        RECT 205.875 -75.645 206.205 -75.315 ;
        RECT 205.875 -77.005 206.205 -76.675 ;
        RECT 205.875 -78.365 206.205 -78.035 ;
        RECT 205.875 -79.725 206.205 -79.395 ;
        RECT 205.875 -81.085 206.205 -80.755 ;
        RECT 205.875 -82.445 206.205 -82.115 ;
        RECT 205.875 -83.805 206.205 -83.475 ;
        RECT 205.875 -85.165 206.205 -84.835 ;
        RECT 205.875 -86.525 206.205 -86.195 ;
        RECT 205.875 -87.885 206.205 -87.555 ;
        RECT 205.875 -89.245 206.205 -88.915 ;
        RECT 205.875 -90.605 206.205 -90.275 ;
        RECT 205.875 -91.965 206.205 -91.635 ;
        RECT 205.875 -93.325 206.205 -92.995 ;
        RECT 205.875 -94.685 206.205 -94.355 ;
        RECT 205.875 -96.045 206.205 -95.715 ;
        RECT 205.875 -97.405 206.205 -97.075 ;
        RECT 205.875 -98.765 206.205 -98.435 ;
        RECT 205.875 -100.125 206.205 -99.795 ;
        RECT 205.875 -101.485 206.205 -101.155 ;
        RECT 205.875 -102.845 206.205 -102.515 ;
        RECT 205.875 -104.205 206.205 -103.875 ;
        RECT 205.875 -105.565 206.205 -105.235 ;
        RECT 205.875 -106.925 206.205 -106.595 ;
        RECT 205.875 -108.285 206.205 -107.955 ;
        RECT 205.875 -109.645 206.205 -109.315 ;
        RECT 205.875 -111.005 206.205 -110.675 ;
        RECT 205.875 -112.365 206.205 -112.035 ;
        RECT 205.875 -113.725 206.205 -113.395 ;
        RECT 205.875 -115.085 206.205 -114.755 ;
        RECT 205.875 -116.445 206.205 -116.115 ;
        RECT 205.875 -117.805 206.205 -117.475 ;
        RECT 205.875 -119.165 206.205 -118.835 ;
        RECT 205.875 -120.525 206.205 -120.195 ;
        RECT 205.875 -121.885 206.205 -121.555 ;
        RECT 205.875 -123.245 206.205 -122.915 ;
        RECT 205.875 -124.605 206.205 -124.275 ;
        RECT 205.875 -125.965 206.205 -125.635 ;
        RECT 205.875 -127.325 206.205 -126.995 ;
        RECT 205.875 -128.685 206.205 -128.355 ;
        RECT 205.875 -130.045 206.205 -129.715 ;
        RECT 205.875 -131.405 206.205 -131.075 ;
        RECT 205.875 -132.765 206.205 -132.435 ;
        RECT 205.875 -134.125 206.205 -133.795 ;
        RECT 205.875 -135.485 206.205 -135.155 ;
        RECT 205.875 -136.845 206.205 -136.515 ;
        RECT 205.875 -138.205 206.205 -137.875 ;
        RECT 205.875 -139.565 206.205 -139.235 ;
        RECT 205.875 -140.925 206.205 -140.595 ;
        RECT 205.875 -142.285 206.205 -141.955 ;
        RECT 205.875 -143.645 206.205 -143.315 ;
        RECT 205.875 -145.005 206.205 -144.675 ;
        RECT 205.875 -146.365 206.205 -146.035 ;
        RECT 205.875 -147.725 206.205 -147.395 ;
        RECT 205.875 -149.085 206.205 -148.755 ;
        RECT 205.875 -150.445 206.205 -150.115 ;
        RECT 205.875 -151.805 206.205 -151.475 ;
        RECT 205.875 -153.165 206.205 -152.835 ;
        RECT 205.875 -154.525 206.205 -154.195 ;
        RECT 205.875 -155.885 206.205 -155.555 ;
        RECT 205.875 -157.245 206.205 -156.915 ;
        RECT 205.875 -162.89 206.205 -161.76 ;
        RECT 205.88 -163.005 206.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 129.945 207.565 131.075 ;
        RECT 207.235 125.635 207.565 125.965 ;
        RECT 207.235 124.275 207.565 124.605 ;
        RECT 207.235 -0.845 207.565 -0.515 ;
        RECT 207.235 -2.205 207.565 -1.875 ;
        RECT 207.235 -3.565 207.565 -3.235 ;
        RECT 207.235 -4.925 207.565 -4.595 ;
        RECT 207.235 -6.285 207.565 -5.955 ;
        RECT 207.235 -7.645 207.565 -7.315 ;
        RECT 207.235 -9.005 207.565 -8.675 ;
        RECT 207.235 -10.365 207.565 -10.035 ;
        RECT 207.235 -11.725 207.565 -11.395 ;
        RECT 207.235 -13.085 207.565 -12.755 ;
        RECT 207.235 -14.445 207.565 -14.115 ;
        RECT 207.235 -15.805 207.565 -15.475 ;
        RECT 207.235 -17.165 207.565 -16.835 ;
        RECT 207.235 -18.525 207.565 -18.195 ;
        RECT 207.235 -19.885 207.565 -19.555 ;
        RECT 207.235 -21.245 207.565 -20.915 ;
        RECT 207.235 -22.605 207.565 -22.275 ;
        RECT 207.235 -23.965 207.565 -23.635 ;
        RECT 207.235 -25.325 207.565 -24.995 ;
        RECT 207.235 -26.685 207.565 -26.355 ;
        RECT 207.235 -28.045 207.565 -27.715 ;
        RECT 207.235 -29.405 207.565 -29.075 ;
        RECT 207.235 -30.765 207.565 -30.435 ;
        RECT 207.235 -32.125 207.565 -31.795 ;
        RECT 207.235 -33.485 207.565 -33.155 ;
        RECT 207.235 -34.845 207.565 -34.515 ;
        RECT 207.235 -36.205 207.565 -35.875 ;
        RECT 207.235 -37.565 207.565 -37.235 ;
        RECT 207.235 -38.925 207.565 -38.595 ;
        RECT 207.235 -40.285 207.565 -39.955 ;
        RECT 207.235 -41.645 207.565 -41.315 ;
        RECT 207.235 -43.005 207.565 -42.675 ;
        RECT 207.235 -44.365 207.565 -44.035 ;
        RECT 207.235 -45.725 207.565 -45.395 ;
        RECT 207.235 -47.085 207.565 -46.755 ;
        RECT 207.235 -48.445 207.565 -48.115 ;
        RECT 207.235 -49.805 207.565 -49.475 ;
        RECT 207.235 -51.165 207.565 -50.835 ;
        RECT 207.235 -52.525 207.565 -52.195 ;
        RECT 207.235 -53.885 207.565 -53.555 ;
        RECT 207.235 -55.245 207.565 -54.915 ;
        RECT 207.235 -56.605 207.565 -56.275 ;
        RECT 207.235 -57.965 207.565 -57.635 ;
        RECT 207.235 -59.325 207.565 -58.995 ;
        RECT 207.235 -60.685 207.565 -60.355 ;
        RECT 207.235 -62.045 207.565 -61.715 ;
        RECT 207.235 -63.405 207.565 -63.075 ;
        RECT 207.235 -64.765 207.565 -64.435 ;
        RECT 207.235 -66.125 207.565 -65.795 ;
        RECT 207.235 -67.485 207.565 -67.155 ;
        RECT 207.235 -68.845 207.565 -68.515 ;
        RECT 207.235 -70.205 207.565 -69.875 ;
        RECT 207.235 -71.565 207.565 -71.235 ;
        RECT 207.235 -72.925 207.565 -72.595 ;
        RECT 207.235 -74.285 207.565 -73.955 ;
        RECT 207.235 -75.645 207.565 -75.315 ;
        RECT 207.235 -77.005 207.565 -76.675 ;
        RECT 207.235 -78.365 207.565 -78.035 ;
        RECT 207.235 -79.725 207.565 -79.395 ;
        RECT 207.235 -81.085 207.565 -80.755 ;
        RECT 207.235 -82.445 207.565 -82.115 ;
        RECT 207.235 -83.805 207.565 -83.475 ;
        RECT 207.235 -85.165 207.565 -84.835 ;
        RECT 207.235 -86.525 207.565 -86.195 ;
        RECT 207.235 -87.885 207.565 -87.555 ;
        RECT 207.235 -89.245 207.565 -88.915 ;
        RECT 207.235 -90.605 207.565 -90.275 ;
        RECT 207.235 -91.965 207.565 -91.635 ;
        RECT 207.235 -93.325 207.565 -92.995 ;
        RECT 207.235 -94.685 207.565 -94.355 ;
        RECT 207.235 -96.045 207.565 -95.715 ;
        RECT 207.235 -97.405 207.565 -97.075 ;
        RECT 207.235 -98.765 207.565 -98.435 ;
        RECT 207.235 -100.125 207.565 -99.795 ;
        RECT 207.235 -101.485 207.565 -101.155 ;
        RECT 207.235 -102.845 207.565 -102.515 ;
        RECT 207.235 -104.205 207.565 -103.875 ;
        RECT 207.235 -105.565 207.565 -105.235 ;
        RECT 207.235 -106.925 207.565 -106.595 ;
        RECT 207.235 -108.285 207.565 -107.955 ;
        RECT 207.235 -109.645 207.565 -109.315 ;
        RECT 207.235 -111.005 207.565 -110.675 ;
        RECT 207.235 -112.365 207.565 -112.035 ;
        RECT 207.235 -113.725 207.565 -113.395 ;
        RECT 207.235 -115.085 207.565 -114.755 ;
        RECT 207.235 -116.445 207.565 -116.115 ;
        RECT 207.235 -117.805 207.565 -117.475 ;
        RECT 207.235 -119.165 207.565 -118.835 ;
        RECT 207.235 -120.525 207.565 -120.195 ;
        RECT 207.235 -121.885 207.565 -121.555 ;
        RECT 207.235 -123.245 207.565 -122.915 ;
        RECT 207.235 -124.605 207.565 -124.275 ;
        RECT 207.235 -125.965 207.565 -125.635 ;
        RECT 207.235 -127.325 207.565 -126.995 ;
        RECT 207.235 -128.685 207.565 -128.355 ;
        RECT 207.235 -130.045 207.565 -129.715 ;
        RECT 207.235 -131.405 207.565 -131.075 ;
        RECT 207.235 -132.765 207.565 -132.435 ;
        RECT 207.235 -134.125 207.565 -133.795 ;
        RECT 207.235 -135.485 207.565 -135.155 ;
        RECT 207.235 -136.845 207.565 -136.515 ;
        RECT 207.235 -138.205 207.565 -137.875 ;
        RECT 207.235 -139.565 207.565 -139.235 ;
        RECT 207.235 -140.925 207.565 -140.595 ;
        RECT 207.235 -142.285 207.565 -141.955 ;
        RECT 207.235 -143.645 207.565 -143.315 ;
        RECT 207.235 -145.005 207.565 -144.675 ;
        RECT 207.235 -146.365 207.565 -146.035 ;
        RECT 207.235 -147.725 207.565 -147.395 ;
        RECT 207.235 -149.085 207.565 -148.755 ;
        RECT 207.235 -150.445 207.565 -150.115 ;
        RECT 207.235 -151.805 207.565 -151.475 ;
        RECT 207.235 -153.165 207.565 -152.835 ;
        RECT 207.235 -154.525 207.565 -154.195 ;
        RECT 207.235 -155.885 207.565 -155.555 ;
        RECT 207.235 -157.245 207.565 -156.915 ;
        RECT 207.235 -162.89 207.565 -161.76 ;
        RECT 207.24 -163.005 207.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.16 -94.075 155.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 129.945 155.885 131.075 ;
        RECT 155.555 125.635 155.885 125.965 ;
        RECT 155.555 124.275 155.885 124.605 ;
        RECT 155.56 123.6 155.88 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 -96.045 155.885 -95.715 ;
        RECT 155.555 -97.405 155.885 -97.075 ;
        RECT 155.555 -98.765 155.885 -98.435 ;
        RECT 155.555 -100.125 155.885 -99.795 ;
        RECT 155.555 -101.485 155.885 -101.155 ;
        RECT 155.555 -102.845 155.885 -102.515 ;
        RECT 155.555 -104.205 155.885 -103.875 ;
        RECT 155.555 -105.565 155.885 -105.235 ;
        RECT 155.555 -106.925 155.885 -106.595 ;
        RECT 155.555 -108.285 155.885 -107.955 ;
        RECT 155.555 -109.645 155.885 -109.315 ;
        RECT 155.555 -111.005 155.885 -110.675 ;
        RECT 155.555 -112.365 155.885 -112.035 ;
        RECT 155.555 -113.725 155.885 -113.395 ;
        RECT 155.555 -115.085 155.885 -114.755 ;
        RECT 155.555 -116.445 155.885 -116.115 ;
        RECT 155.555 -117.805 155.885 -117.475 ;
        RECT 155.555 -119.165 155.885 -118.835 ;
        RECT 155.555 -120.525 155.885 -120.195 ;
        RECT 155.555 -121.885 155.885 -121.555 ;
        RECT 155.555 -123.245 155.885 -122.915 ;
        RECT 155.555 -124.605 155.885 -124.275 ;
        RECT 155.555 -125.965 155.885 -125.635 ;
        RECT 155.555 -127.325 155.885 -126.995 ;
        RECT 155.555 -128.685 155.885 -128.355 ;
        RECT 155.555 -130.045 155.885 -129.715 ;
        RECT 155.555 -131.405 155.885 -131.075 ;
        RECT 155.555 -132.765 155.885 -132.435 ;
        RECT 155.555 -134.125 155.885 -133.795 ;
        RECT 155.555 -135.485 155.885 -135.155 ;
        RECT 155.555 -136.845 155.885 -136.515 ;
        RECT 155.555 -138.205 155.885 -137.875 ;
        RECT 155.555 -139.565 155.885 -139.235 ;
        RECT 155.555 -140.925 155.885 -140.595 ;
        RECT 155.555 -142.285 155.885 -141.955 ;
        RECT 155.555 -143.645 155.885 -143.315 ;
        RECT 155.555 -145.005 155.885 -144.675 ;
        RECT 155.555 -146.365 155.885 -146.035 ;
        RECT 155.555 -147.725 155.885 -147.395 ;
        RECT 155.555 -149.085 155.885 -148.755 ;
        RECT 155.555 -150.445 155.885 -150.115 ;
        RECT 155.555 -151.805 155.885 -151.475 ;
        RECT 155.555 -153.165 155.885 -152.835 ;
        RECT 155.555 -154.525 155.885 -154.195 ;
        RECT 155.555 -155.885 155.885 -155.555 ;
        RECT 155.555 -157.245 155.885 -156.915 ;
        RECT 155.555 -162.89 155.885 -161.76 ;
        RECT 155.56 -163.005 155.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 129.945 157.245 131.075 ;
        RECT 156.915 125.635 157.245 125.965 ;
        RECT 156.915 124.275 157.245 124.605 ;
        RECT 156.92 123.6 157.24 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 -0.845 157.245 -0.515 ;
        RECT 156.915 -2.205 157.245 -1.875 ;
        RECT 156.915 -3.565 157.245 -3.235 ;
        RECT 156.92 -3.565 157.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 129.945 158.605 131.075 ;
        RECT 158.275 125.635 158.605 125.965 ;
        RECT 158.275 124.275 158.605 124.605 ;
        RECT 158.28 123.6 158.6 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 -0.845 158.605 -0.515 ;
        RECT 158.275 -2.205 158.605 -1.875 ;
        RECT 158.275 -3.565 158.605 -3.235 ;
        RECT 158.28 -3.565 158.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 129.945 159.965 131.075 ;
        RECT 159.635 125.635 159.965 125.965 ;
        RECT 159.635 124.275 159.965 124.605 ;
        RECT 159.64 123.6 159.96 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -0.845 159.965 -0.515 ;
        RECT 159.635 -2.205 159.965 -1.875 ;
        RECT 159.635 -3.565 159.965 -3.235 ;
        RECT 159.64 -3.565 159.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -91.965 159.965 -91.635 ;
        RECT 159.635 -93.325 159.965 -92.995 ;
        RECT 159.635 -94.685 159.965 -94.355 ;
        RECT 159.635 -96.045 159.965 -95.715 ;
        RECT 159.635 -97.405 159.965 -97.075 ;
        RECT 159.635 -98.765 159.965 -98.435 ;
        RECT 159.635 -100.125 159.965 -99.795 ;
        RECT 159.635 -101.485 159.965 -101.155 ;
        RECT 159.635 -102.845 159.965 -102.515 ;
        RECT 159.635 -104.205 159.965 -103.875 ;
        RECT 159.635 -105.565 159.965 -105.235 ;
        RECT 159.635 -106.925 159.965 -106.595 ;
        RECT 159.635 -108.285 159.965 -107.955 ;
        RECT 159.635 -109.645 159.965 -109.315 ;
        RECT 159.635 -111.005 159.965 -110.675 ;
        RECT 159.635 -112.365 159.965 -112.035 ;
        RECT 159.635 -113.725 159.965 -113.395 ;
        RECT 159.635 -115.085 159.965 -114.755 ;
        RECT 159.635 -116.445 159.965 -116.115 ;
        RECT 159.635 -117.805 159.965 -117.475 ;
        RECT 159.635 -119.165 159.965 -118.835 ;
        RECT 159.635 -120.525 159.965 -120.195 ;
        RECT 159.635 -121.885 159.965 -121.555 ;
        RECT 159.635 -123.245 159.965 -122.915 ;
        RECT 159.635 -124.605 159.965 -124.275 ;
        RECT 159.635 -125.965 159.965 -125.635 ;
        RECT 159.635 -127.325 159.965 -126.995 ;
        RECT 159.635 -128.685 159.965 -128.355 ;
        RECT 159.635 -130.045 159.965 -129.715 ;
        RECT 159.635 -131.405 159.965 -131.075 ;
        RECT 159.635 -132.765 159.965 -132.435 ;
        RECT 159.635 -134.125 159.965 -133.795 ;
        RECT 159.635 -135.485 159.965 -135.155 ;
        RECT 159.635 -136.845 159.965 -136.515 ;
        RECT 159.635 -138.205 159.965 -137.875 ;
        RECT 159.635 -139.565 159.965 -139.235 ;
        RECT 159.635 -140.925 159.965 -140.595 ;
        RECT 159.635 -142.285 159.965 -141.955 ;
        RECT 159.635 -143.645 159.965 -143.315 ;
        RECT 159.635 -145.005 159.965 -144.675 ;
        RECT 159.635 -146.365 159.965 -146.035 ;
        RECT 159.635 -147.725 159.965 -147.395 ;
        RECT 159.635 -149.085 159.965 -148.755 ;
        RECT 159.635 -150.445 159.965 -150.115 ;
        RECT 159.635 -151.805 159.965 -151.475 ;
        RECT 159.635 -153.165 159.965 -152.835 ;
        RECT 159.635 -154.525 159.965 -154.195 ;
        RECT 159.635 -155.885 159.965 -155.555 ;
        RECT 159.635 -157.245 159.965 -156.915 ;
        RECT 159.635 -162.89 159.965 -161.76 ;
        RECT 159.64 -163.005 159.96 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 129.945 161.325 131.075 ;
        RECT 160.995 125.635 161.325 125.965 ;
        RECT 160.995 124.275 161.325 124.605 ;
        RECT 161 123.6 161.32 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 -96.045 161.325 -95.715 ;
        RECT 160.995 -97.405 161.325 -97.075 ;
        RECT 160.995 -98.765 161.325 -98.435 ;
        RECT 160.995 -100.125 161.325 -99.795 ;
        RECT 160.995 -101.485 161.325 -101.155 ;
        RECT 160.995 -102.845 161.325 -102.515 ;
        RECT 160.995 -104.205 161.325 -103.875 ;
        RECT 160.995 -105.565 161.325 -105.235 ;
        RECT 160.995 -106.925 161.325 -106.595 ;
        RECT 160.995 -108.285 161.325 -107.955 ;
        RECT 160.995 -109.645 161.325 -109.315 ;
        RECT 160.995 -111.005 161.325 -110.675 ;
        RECT 160.995 -112.365 161.325 -112.035 ;
        RECT 160.995 -113.725 161.325 -113.395 ;
        RECT 160.995 -115.085 161.325 -114.755 ;
        RECT 160.995 -116.445 161.325 -116.115 ;
        RECT 160.995 -117.805 161.325 -117.475 ;
        RECT 160.995 -119.165 161.325 -118.835 ;
        RECT 160.995 -120.525 161.325 -120.195 ;
        RECT 160.995 -121.885 161.325 -121.555 ;
        RECT 160.995 -123.245 161.325 -122.915 ;
        RECT 160.995 -124.605 161.325 -124.275 ;
        RECT 160.995 -125.965 161.325 -125.635 ;
        RECT 160.995 -127.325 161.325 -126.995 ;
        RECT 160.995 -128.685 161.325 -128.355 ;
        RECT 160.995 -130.045 161.325 -129.715 ;
        RECT 160.995 -131.405 161.325 -131.075 ;
        RECT 160.995 -132.765 161.325 -132.435 ;
        RECT 160.995 -134.125 161.325 -133.795 ;
        RECT 160.995 -135.485 161.325 -135.155 ;
        RECT 160.995 -136.845 161.325 -136.515 ;
        RECT 160.995 -138.205 161.325 -137.875 ;
        RECT 160.995 -139.565 161.325 -139.235 ;
        RECT 160.995 -140.925 161.325 -140.595 ;
        RECT 160.995 -142.285 161.325 -141.955 ;
        RECT 160.995 -143.645 161.325 -143.315 ;
        RECT 160.995 -145.005 161.325 -144.675 ;
        RECT 160.995 -146.365 161.325 -146.035 ;
        RECT 160.995 -147.725 161.325 -147.395 ;
        RECT 160.995 -149.085 161.325 -148.755 ;
        RECT 160.995 -150.445 161.325 -150.115 ;
        RECT 160.995 -151.805 161.325 -151.475 ;
        RECT 160.995 -153.165 161.325 -152.835 ;
        RECT 160.995 -154.525 161.325 -154.195 ;
        RECT 160.995 -155.885 161.325 -155.555 ;
        RECT 160.995 -157.245 161.325 -156.915 ;
        RECT 160.995 -162.89 161.325 -161.76 ;
        RECT 161 -163.005 161.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.26 -94.075 161.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 129.945 162.685 131.075 ;
        RECT 162.355 125.635 162.685 125.965 ;
        RECT 162.355 124.275 162.685 124.605 ;
        RECT 162.36 123.6 162.68 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 129.945 164.045 131.075 ;
        RECT 163.715 125.635 164.045 125.965 ;
        RECT 163.715 124.275 164.045 124.605 ;
        RECT 163.72 123.6 164.04 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 -0.845 164.045 -0.515 ;
        RECT 163.715 -2.205 164.045 -1.875 ;
        RECT 163.715 -3.565 164.045 -3.235 ;
        RECT 163.72 -3.565 164.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 129.945 165.405 131.075 ;
        RECT 165.075 125.635 165.405 125.965 ;
        RECT 165.075 124.275 165.405 124.605 ;
        RECT 165.08 123.6 165.4 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -0.845 165.405 -0.515 ;
        RECT 165.075 -2.205 165.405 -1.875 ;
        RECT 165.075 -3.565 165.405 -3.235 ;
        RECT 165.08 -3.565 165.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -91.965 165.405 -91.635 ;
        RECT 165.075 -93.325 165.405 -92.995 ;
        RECT 165.075 -94.685 165.405 -94.355 ;
        RECT 165.075 -96.045 165.405 -95.715 ;
        RECT 165.075 -97.405 165.405 -97.075 ;
        RECT 165.075 -98.765 165.405 -98.435 ;
        RECT 165.075 -100.125 165.405 -99.795 ;
        RECT 165.075 -101.485 165.405 -101.155 ;
        RECT 165.075 -102.845 165.405 -102.515 ;
        RECT 165.075 -104.205 165.405 -103.875 ;
        RECT 165.075 -105.565 165.405 -105.235 ;
        RECT 165.075 -106.925 165.405 -106.595 ;
        RECT 165.075 -108.285 165.405 -107.955 ;
        RECT 165.075 -109.645 165.405 -109.315 ;
        RECT 165.075 -111.005 165.405 -110.675 ;
        RECT 165.075 -112.365 165.405 -112.035 ;
        RECT 165.075 -113.725 165.405 -113.395 ;
        RECT 165.075 -115.085 165.405 -114.755 ;
        RECT 165.075 -116.445 165.405 -116.115 ;
        RECT 165.075 -117.805 165.405 -117.475 ;
        RECT 165.075 -119.165 165.405 -118.835 ;
        RECT 165.075 -120.525 165.405 -120.195 ;
        RECT 165.075 -121.885 165.405 -121.555 ;
        RECT 165.075 -123.245 165.405 -122.915 ;
        RECT 165.075 -124.605 165.405 -124.275 ;
        RECT 165.075 -125.965 165.405 -125.635 ;
        RECT 165.075 -127.325 165.405 -126.995 ;
        RECT 165.075 -128.685 165.405 -128.355 ;
        RECT 165.075 -130.045 165.405 -129.715 ;
        RECT 165.075 -131.405 165.405 -131.075 ;
        RECT 165.075 -132.765 165.405 -132.435 ;
        RECT 165.075 -134.125 165.405 -133.795 ;
        RECT 165.075 -135.485 165.405 -135.155 ;
        RECT 165.075 -136.845 165.405 -136.515 ;
        RECT 165.075 -138.205 165.405 -137.875 ;
        RECT 165.075 -139.565 165.405 -139.235 ;
        RECT 165.075 -140.925 165.405 -140.595 ;
        RECT 165.075 -142.285 165.405 -141.955 ;
        RECT 165.075 -143.645 165.405 -143.315 ;
        RECT 165.075 -145.005 165.405 -144.675 ;
        RECT 165.075 -146.365 165.405 -146.035 ;
        RECT 165.075 -147.725 165.405 -147.395 ;
        RECT 165.075 -149.085 165.405 -148.755 ;
        RECT 165.075 -150.445 165.405 -150.115 ;
        RECT 165.075 -151.805 165.405 -151.475 ;
        RECT 165.075 -153.165 165.405 -152.835 ;
        RECT 165.075 -154.525 165.405 -154.195 ;
        RECT 165.075 -155.885 165.405 -155.555 ;
        RECT 165.075 -157.245 165.405 -156.915 ;
        RECT 165.075 -162.89 165.405 -161.76 ;
        RECT 165.08 -163.005 165.4 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 129.945 166.765 131.075 ;
        RECT 166.435 125.635 166.765 125.965 ;
        RECT 166.435 124.275 166.765 124.605 ;
        RECT 166.44 123.6 166.76 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -0.845 166.765 -0.515 ;
        RECT 166.435 -2.205 166.765 -1.875 ;
        RECT 166.435 -3.565 166.765 -3.235 ;
        RECT 166.44 -3.565 166.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -91.965 166.765 -91.635 ;
        RECT 166.435 -93.325 166.765 -92.995 ;
        RECT 166.435 -94.685 166.765 -94.355 ;
        RECT 166.435 -96.045 166.765 -95.715 ;
        RECT 166.435 -97.405 166.765 -97.075 ;
        RECT 166.435 -98.765 166.765 -98.435 ;
        RECT 166.435 -100.125 166.765 -99.795 ;
        RECT 166.435 -101.485 166.765 -101.155 ;
        RECT 166.435 -102.845 166.765 -102.515 ;
        RECT 166.435 -104.205 166.765 -103.875 ;
        RECT 166.435 -105.565 166.765 -105.235 ;
        RECT 166.435 -106.925 166.765 -106.595 ;
        RECT 166.435 -108.285 166.765 -107.955 ;
        RECT 166.435 -109.645 166.765 -109.315 ;
        RECT 166.435 -111.005 166.765 -110.675 ;
        RECT 166.435 -112.365 166.765 -112.035 ;
        RECT 166.435 -113.725 166.765 -113.395 ;
        RECT 166.435 -115.085 166.765 -114.755 ;
        RECT 166.435 -116.445 166.765 -116.115 ;
        RECT 166.435 -117.805 166.765 -117.475 ;
        RECT 166.435 -119.165 166.765 -118.835 ;
        RECT 166.435 -120.525 166.765 -120.195 ;
        RECT 166.435 -121.885 166.765 -121.555 ;
        RECT 166.435 -123.245 166.765 -122.915 ;
        RECT 166.435 -124.605 166.765 -124.275 ;
        RECT 166.435 -125.965 166.765 -125.635 ;
        RECT 166.435 -127.325 166.765 -126.995 ;
        RECT 166.435 -128.685 166.765 -128.355 ;
        RECT 166.435 -130.045 166.765 -129.715 ;
        RECT 166.435 -131.405 166.765 -131.075 ;
        RECT 166.435 -132.765 166.765 -132.435 ;
        RECT 166.435 -134.125 166.765 -133.795 ;
        RECT 166.435 -135.485 166.765 -135.155 ;
        RECT 166.435 -136.845 166.765 -136.515 ;
        RECT 166.435 -138.205 166.765 -137.875 ;
        RECT 166.435 -139.565 166.765 -139.235 ;
        RECT 166.435 -140.925 166.765 -140.595 ;
        RECT 166.435 -142.285 166.765 -141.955 ;
        RECT 166.435 -143.645 166.765 -143.315 ;
        RECT 166.435 -145.005 166.765 -144.675 ;
        RECT 166.435 -146.365 166.765 -146.035 ;
        RECT 166.435 -147.725 166.765 -147.395 ;
        RECT 166.435 -149.085 166.765 -148.755 ;
        RECT 166.435 -150.445 166.765 -150.115 ;
        RECT 166.435 -151.805 166.765 -151.475 ;
        RECT 166.435 -153.165 166.765 -152.835 ;
        RECT 166.435 -154.525 166.765 -154.195 ;
        RECT 166.435 -155.885 166.765 -155.555 ;
        RECT 166.435 -157.245 166.765 -156.915 ;
        RECT 166.435 -162.89 166.765 -161.76 ;
        RECT 166.44 -163.005 166.76 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.36 -94.075 167.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 129.945 168.125 131.075 ;
        RECT 167.795 125.635 168.125 125.965 ;
        RECT 167.795 124.275 168.125 124.605 ;
        RECT 167.8 123.6 168.12 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 -96.045 168.125 -95.715 ;
        RECT 167.795 -97.405 168.125 -97.075 ;
        RECT 167.795 -98.765 168.125 -98.435 ;
        RECT 167.795 -100.125 168.125 -99.795 ;
        RECT 167.795 -101.485 168.125 -101.155 ;
        RECT 167.795 -102.845 168.125 -102.515 ;
        RECT 167.795 -104.205 168.125 -103.875 ;
        RECT 167.795 -105.565 168.125 -105.235 ;
        RECT 167.795 -106.925 168.125 -106.595 ;
        RECT 167.795 -108.285 168.125 -107.955 ;
        RECT 167.795 -109.645 168.125 -109.315 ;
        RECT 167.795 -111.005 168.125 -110.675 ;
        RECT 167.795 -112.365 168.125 -112.035 ;
        RECT 167.795 -113.725 168.125 -113.395 ;
        RECT 167.795 -115.085 168.125 -114.755 ;
        RECT 167.795 -116.445 168.125 -116.115 ;
        RECT 167.795 -117.805 168.125 -117.475 ;
        RECT 167.795 -119.165 168.125 -118.835 ;
        RECT 167.795 -120.525 168.125 -120.195 ;
        RECT 167.795 -121.885 168.125 -121.555 ;
        RECT 167.795 -123.245 168.125 -122.915 ;
        RECT 167.795 -124.605 168.125 -124.275 ;
        RECT 167.795 -125.965 168.125 -125.635 ;
        RECT 167.795 -127.325 168.125 -126.995 ;
        RECT 167.795 -128.685 168.125 -128.355 ;
        RECT 167.795 -130.045 168.125 -129.715 ;
        RECT 167.795 -131.405 168.125 -131.075 ;
        RECT 167.795 -132.765 168.125 -132.435 ;
        RECT 167.795 -134.125 168.125 -133.795 ;
        RECT 167.795 -135.485 168.125 -135.155 ;
        RECT 167.795 -136.845 168.125 -136.515 ;
        RECT 167.795 -138.205 168.125 -137.875 ;
        RECT 167.795 -139.565 168.125 -139.235 ;
        RECT 167.795 -140.925 168.125 -140.595 ;
        RECT 167.795 -142.285 168.125 -141.955 ;
        RECT 167.795 -143.645 168.125 -143.315 ;
        RECT 167.795 -145.005 168.125 -144.675 ;
        RECT 167.795 -146.365 168.125 -146.035 ;
        RECT 167.795 -147.725 168.125 -147.395 ;
        RECT 167.795 -149.085 168.125 -148.755 ;
        RECT 167.795 -150.445 168.125 -150.115 ;
        RECT 167.795 -151.805 168.125 -151.475 ;
        RECT 167.795 -153.165 168.125 -152.835 ;
        RECT 167.795 -154.525 168.125 -154.195 ;
        RECT 167.795 -155.885 168.125 -155.555 ;
        RECT 167.795 -157.245 168.125 -156.915 ;
        RECT 167.795 -162.89 168.125 -161.76 ;
        RECT 167.8 -163.005 168.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 129.945 169.485 131.075 ;
        RECT 169.155 125.635 169.485 125.965 ;
        RECT 169.155 124.275 169.485 124.605 ;
        RECT 169.16 123.6 169.48 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 -0.845 169.485 -0.515 ;
        RECT 169.155 -2.205 169.485 -1.875 ;
        RECT 169.155 -3.565 169.485 -3.235 ;
        RECT 169.16 -3.565 169.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 129.945 170.845 131.075 ;
        RECT 170.515 125.635 170.845 125.965 ;
        RECT 170.515 124.275 170.845 124.605 ;
        RECT 170.52 123.6 170.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 -0.845 170.845 -0.515 ;
        RECT 170.515 -2.205 170.845 -1.875 ;
        RECT 170.515 -3.565 170.845 -3.235 ;
        RECT 170.52 -3.565 170.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 129.945 172.205 131.075 ;
        RECT 171.875 125.635 172.205 125.965 ;
        RECT 171.875 124.275 172.205 124.605 ;
        RECT 171.88 123.6 172.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -0.845 172.205 -0.515 ;
        RECT 171.875 -2.205 172.205 -1.875 ;
        RECT 171.875 -3.565 172.205 -3.235 ;
        RECT 171.88 -3.565 172.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -91.965 172.205 -91.635 ;
        RECT 171.875 -93.325 172.205 -92.995 ;
        RECT 171.875 -94.685 172.205 -94.355 ;
        RECT 171.875 -96.045 172.205 -95.715 ;
        RECT 171.875 -97.405 172.205 -97.075 ;
        RECT 171.875 -98.765 172.205 -98.435 ;
        RECT 171.875 -100.125 172.205 -99.795 ;
        RECT 171.875 -101.485 172.205 -101.155 ;
        RECT 171.875 -102.845 172.205 -102.515 ;
        RECT 171.875 -104.205 172.205 -103.875 ;
        RECT 171.875 -105.565 172.205 -105.235 ;
        RECT 171.875 -106.925 172.205 -106.595 ;
        RECT 171.875 -108.285 172.205 -107.955 ;
        RECT 171.875 -109.645 172.205 -109.315 ;
        RECT 171.875 -111.005 172.205 -110.675 ;
        RECT 171.875 -112.365 172.205 -112.035 ;
        RECT 171.875 -113.725 172.205 -113.395 ;
        RECT 171.875 -115.085 172.205 -114.755 ;
        RECT 171.875 -116.445 172.205 -116.115 ;
        RECT 171.875 -117.805 172.205 -117.475 ;
        RECT 171.875 -119.165 172.205 -118.835 ;
        RECT 171.875 -120.525 172.205 -120.195 ;
        RECT 171.875 -121.885 172.205 -121.555 ;
        RECT 171.875 -123.245 172.205 -122.915 ;
        RECT 171.875 -124.605 172.205 -124.275 ;
        RECT 171.875 -125.965 172.205 -125.635 ;
        RECT 171.875 -127.325 172.205 -126.995 ;
        RECT 171.875 -128.685 172.205 -128.355 ;
        RECT 171.875 -130.045 172.205 -129.715 ;
        RECT 171.875 -131.405 172.205 -131.075 ;
        RECT 171.875 -132.765 172.205 -132.435 ;
        RECT 171.875 -134.125 172.205 -133.795 ;
        RECT 171.875 -135.485 172.205 -135.155 ;
        RECT 171.875 -136.845 172.205 -136.515 ;
        RECT 171.875 -138.205 172.205 -137.875 ;
        RECT 171.875 -139.565 172.205 -139.235 ;
        RECT 171.875 -140.925 172.205 -140.595 ;
        RECT 171.875 -142.285 172.205 -141.955 ;
        RECT 171.875 -143.645 172.205 -143.315 ;
        RECT 171.875 -145.005 172.205 -144.675 ;
        RECT 171.875 -146.365 172.205 -146.035 ;
        RECT 171.875 -147.725 172.205 -147.395 ;
        RECT 171.875 -149.085 172.205 -148.755 ;
        RECT 171.875 -150.445 172.205 -150.115 ;
        RECT 171.875 -151.805 172.205 -151.475 ;
        RECT 171.875 -153.165 172.205 -152.835 ;
        RECT 171.875 -154.525 172.205 -154.195 ;
        RECT 171.875 -155.885 172.205 -155.555 ;
        RECT 171.875 -157.245 172.205 -156.915 ;
        RECT 171.875 -162.89 172.205 -161.76 ;
        RECT 171.88 -163.005 172.2 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 129.945 173.565 131.075 ;
        RECT 173.235 125.635 173.565 125.965 ;
        RECT 173.235 124.275 173.565 124.605 ;
        RECT 173.24 123.6 173.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 -96.045 173.565 -95.715 ;
        RECT 173.235 -97.405 173.565 -97.075 ;
        RECT 173.235 -98.765 173.565 -98.435 ;
        RECT 173.235 -100.125 173.565 -99.795 ;
        RECT 173.235 -101.485 173.565 -101.155 ;
        RECT 173.235 -102.845 173.565 -102.515 ;
        RECT 173.235 -104.205 173.565 -103.875 ;
        RECT 173.235 -105.565 173.565 -105.235 ;
        RECT 173.235 -106.925 173.565 -106.595 ;
        RECT 173.235 -108.285 173.565 -107.955 ;
        RECT 173.235 -109.645 173.565 -109.315 ;
        RECT 173.235 -111.005 173.565 -110.675 ;
        RECT 173.235 -112.365 173.565 -112.035 ;
        RECT 173.235 -113.725 173.565 -113.395 ;
        RECT 173.235 -115.085 173.565 -114.755 ;
        RECT 173.235 -116.445 173.565 -116.115 ;
        RECT 173.235 -117.805 173.565 -117.475 ;
        RECT 173.235 -119.165 173.565 -118.835 ;
        RECT 173.235 -120.525 173.565 -120.195 ;
        RECT 173.235 -121.885 173.565 -121.555 ;
        RECT 173.235 -123.245 173.565 -122.915 ;
        RECT 173.235 -124.605 173.565 -124.275 ;
        RECT 173.235 -125.965 173.565 -125.635 ;
        RECT 173.235 -127.325 173.565 -126.995 ;
        RECT 173.235 -128.685 173.565 -128.355 ;
        RECT 173.235 -130.045 173.565 -129.715 ;
        RECT 173.235 -131.405 173.565 -131.075 ;
        RECT 173.235 -132.765 173.565 -132.435 ;
        RECT 173.235 -134.125 173.565 -133.795 ;
        RECT 173.235 -135.485 173.565 -135.155 ;
        RECT 173.235 -136.845 173.565 -136.515 ;
        RECT 173.235 -138.205 173.565 -137.875 ;
        RECT 173.235 -139.565 173.565 -139.235 ;
        RECT 173.235 -140.925 173.565 -140.595 ;
        RECT 173.235 -142.285 173.565 -141.955 ;
        RECT 173.235 -143.645 173.565 -143.315 ;
        RECT 173.235 -145.005 173.565 -144.675 ;
        RECT 173.235 -146.365 173.565 -146.035 ;
        RECT 173.235 -147.725 173.565 -147.395 ;
        RECT 173.235 -149.085 173.565 -148.755 ;
        RECT 173.235 -150.445 173.565 -150.115 ;
        RECT 173.235 -151.805 173.565 -151.475 ;
        RECT 173.235 -153.165 173.565 -152.835 ;
        RECT 173.235 -154.525 173.565 -154.195 ;
        RECT 173.235 -155.885 173.565 -155.555 ;
        RECT 173.235 -157.245 173.565 -156.915 ;
        RECT 173.235 -162.89 173.565 -161.76 ;
        RECT 173.24 -163.005 173.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.46 -94.075 173.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 129.945 174.925 131.075 ;
        RECT 174.595 125.635 174.925 125.965 ;
        RECT 174.595 124.275 174.925 124.605 ;
        RECT 174.6 123.6 174.92 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 129.945 176.285 131.075 ;
        RECT 175.955 125.635 176.285 125.965 ;
        RECT 175.955 124.275 176.285 124.605 ;
        RECT 175.96 123.6 176.28 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 -0.845 176.285 -0.515 ;
        RECT 175.955 -2.205 176.285 -1.875 ;
        RECT 175.955 -3.565 176.285 -3.235 ;
        RECT 175.96 -3.565 176.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 129.945 177.645 131.075 ;
        RECT 177.315 125.635 177.645 125.965 ;
        RECT 177.315 124.275 177.645 124.605 ;
        RECT 177.32 123.6 177.64 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 -0.845 177.645 -0.515 ;
        RECT 177.315 -2.205 177.645 -1.875 ;
        RECT 177.315 -3.565 177.645 -3.235 ;
        RECT 177.32 -3.565 177.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 -91.965 177.645 -91.635 ;
        RECT 177.315 -93.325 177.645 -92.995 ;
        RECT 177.315 -94.685 177.645 -94.355 ;
        RECT 177.315 -96.045 177.645 -95.715 ;
        RECT 177.315 -97.405 177.645 -97.075 ;
        RECT 177.315 -98.765 177.645 -98.435 ;
        RECT 177.315 -100.125 177.645 -99.795 ;
        RECT 177.315 -101.485 177.645 -101.155 ;
        RECT 177.315 -102.845 177.645 -102.515 ;
        RECT 177.315 -104.205 177.645 -103.875 ;
        RECT 177.315 -105.565 177.645 -105.235 ;
        RECT 177.315 -106.925 177.645 -106.595 ;
        RECT 177.315 -108.285 177.645 -107.955 ;
        RECT 177.315 -109.645 177.645 -109.315 ;
        RECT 177.315 -111.005 177.645 -110.675 ;
        RECT 177.315 -112.365 177.645 -112.035 ;
        RECT 177.315 -113.725 177.645 -113.395 ;
        RECT 177.315 -115.085 177.645 -114.755 ;
        RECT 177.315 -116.445 177.645 -116.115 ;
        RECT 177.315 -117.805 177.645 -117.475 ;
        RECT 177.315 -119.165 177.645 -118.835 ;
        RECT 177.315 -120.525 177.645 -120.195 ;
        RECT 177.315 -121.885 177.645 -121.555 ;
        RECT 177.315 -123.245 177.645 -122.915 ;
        RECT 177.315 -124.605 177.645 -124.275 ;
        RECT 177.315 -125.965 177.645 -125.635 ;
        RECT 177.315 -127.325 177.645 -126.995 ;
        RECT 177.315 -128.685 177.645 -128.355 ;
        RECT 177.315 -130.045 177.645 -129.715 ;
        RECT 177.315 -131.405 177.645 -131.075 ;
        RECT 177.315 -132.765 177.645 -132.435 ;
        RECT 177.315 -134.125 177.645 -133.795 ;
        RECT 177.315 -135.485 177.645 -135.155 ;
        RECT 177.315 -136.845 177.645 -136.515 ;
        RECT 177.315 -138.205 177.645 -137.875 ;
        RECT 177.315 -139.565 177.645 -139.235 ;
        RECT 177.315 -140.925 177.645 -140.595 ;
        RECT 177.315 -142.285 177.645 -141.955 ;
        RECT 177.315 -143.645 177.645 -143.315 ;
        RECT 177.315 -145.005 177.645 -144.675 ;
        RECT 177.315 -146.365 177.645 -146.035 ;
        RECT 177.315 -147.725 177.645 -147.395 ;
        RECT 177.315 -149.085 177.645 -148.755 ;
        RECT 177.315 -150.445 177.645 -150.115 ;
        RECT 177.315 -151.805 177.645 -151.475 ;
        RECT 177.315 -153.165 177.645 -152.835 ;
        RECT 177.315 -154.525 177.645 -154.195 ;
        RECT 177.315 -155.885 177.645 -155.555 ;
        RECT 177.315 -157.245 177.645 -156.915 ;
        RECT 177.315 -162.89 177.645 -161.76 ;
        RECT 177.32 -163.005 177.64 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 129.945 179.005 131.075 ;
        RECT 178.675 125.635 179.005 125.965 ;
        RECT 178.675 124.275 179.005 124.605 ;
        RECT 178.68 123.6 179 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 -0.845 179.005 -0.515 ;
        RECT 178.675 -2.205 179.005 -1.875 ;
        RECT 178.675 -3.565 179.005 -3.235 ;
        RECT 178.68 -3.565 179 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 -91.965 179.005 -91.635 ;
        RECT 178.675 -93.325 179.005 -92.995 ;
        RECT 178.675 -94.685 179.005 -94.355 ;
        RECT 178.675 -96.045 179.005 -95.715 ;
        RECT 178.675 -97.405 179.005 -97.075 ;
        RECT 178.675 -98.765 179.005 -98.435 ;
        RECT 178.675 -100.125 179.005 -99.795 ;
        RECT 178.675 -101.485 179.005 -101.155 ;
        RECT 178.675 -102.845 179.005 -102.515 ;
        RECT 178.675 -104.205 179.005 -103.875 ;
        RECT 178.675 -105.565 179.005 -105.235 ;
        RECT 178.675 -106.925 179.005 -106.595 ;
        RECT 178.675 -108.285 179.005 -107.955 ;
        RECT 178.675 -109.645 179.005 -109.315 ;
        RECT 178.675 -111.005 179.005 -110.675 ;
        RECT 178.675 -112.365 179.005 -112.035 ;
        RECT 178.675 -113.725 179.005 -113.395 ;
        RECT 178.675 -115.085 179.005 -114.755 ;
        RECT 178.675 -116.445 179.005 -116.115 ;
        RECT 178.675 -117.805 179.005 -117.475 ;
        RECT 178.675 -119.165 179.005 -118.835 ;
        RECT 178.675 -120.525 179.005 -120.195 ;
        RECT 178.675 -121.885 179.005 -121.555 ;
        RECT 178.675 -123.245 179.005 -122.915 ;
        RECT 178.675 -124.605 179.005 -124.275 ;
        RECT 178.675 -125.965 179.005 -125.635 ;
        RECT 178.675 -127.325 179.005 -126.995 ;
        RECT 178.675 -128.685 179.005 -128.355 ;
        RECT 178.675 -130.045 179.005 -129.715 ;
        RECT 178.675 -131.405 179.005 -131.075 ;
        RECT 178.675 -132.765 179.005 -132.435 ;
        RECT 178.675 -134.125 179.005 -133.795 ;
        RECT 178.675 -135.485 179.005 -135.155 ;
        RECT 178.675 -136.845 179.005 -136.515 ;
        RECT 178.675 -138.205 179.005 -137.875 ;
        RECT 178.675 -139.565 179.005 -139.235 ;
        RECT 178.675 -140.925 179.005 -140.595 ;
        RECT 178.675 -142.285 179.005 -141.955 ;
        RECT 178.675 -143.645 179.005 -143.315 ;
        RECT 178.675 -145.005 179.005 -144.675 ;
        RECT 178.675 -146.365 179.005 -146.035 ;
        RECT 178.675 -147.725 179.005 -147.395 ;
        RECT 178.675 -149.085 179.005 -148.755 ;
        RECT 178.675 -150.445 179.005 -150.115 ;
        RECT 178.675 -151.805 179.005 -151.475 ;
        RECT 178.675 -153.165 179.005 -152.835 ;
        RECT 178.675 -154.525 179.005 -154.195 ;
        RECT 178.675 -155.885 179.005 -155.555 ;
        RECT 178.675 -157.245 179.005 -156.915 ;
        RECT 178.675 -162.89 179.005 -161.76 ;
        RECT 178.68 -163.005 179 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.56 -94.075 179.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 129.945 180.365 131.075 ;
        RECT 180.035 125.635 180.365 125.965 ;
        RECT 180.035 124.275 180.365 124.605 ;
        RECT 180.04 123.6 180.36 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 -96.045 180.365 -95.715 ;
        RECT 180.035 -97.405 180.365 -97.075 ;
        RECT 180.035 -98.765 180.365 -98.435 ;
        RECT 180.035 -100.125 180.365 -99.795 ;
        RECT 180.035 -101.485 180.365 -101.155 ;
        RECT 180.035 -102.845 180.365 -102.515 ;
        RECT 180.035 -104.205 180.365 -103.875 ;
        RECT 180.035 -105.565 180.365 -105.235 ;
        RECT 180.035 -106.925 180.365 -106.595 ;
        RECT 180.035 -108.285 180.365 -107.955 ;
        RECT 180.035 -109.645 180.365 -109.315 ;
        RECT 180.035 -111.005 180.365 -110.675 ;
        RECT 180.035 -112.365 180.365 -112.035 ;
        RECT 180.035 -113.725 180.365 -113.395 ;
        RECT 180.035 -115.085 180.365 -114.755 ;
        RECT 180.035 -116.445 180.365 -116.115 ;
        RECT 180.035 -117.805 180.365 -117.475 ;
        RECT 180.035 -119.165 180.365 -118.835 ;
        RECT 180.035 -120.525 180.365 -120.195 ;
        RECT 180.035 -121.885 180.365 -121.555 ;
        RECT 180.035 -123.245 180.365 -122.915 ;
        RECT 180.035 -124.605 180.365 -124.275 ;
        RECT 180.035 -125.965 180.365 -125.635 ;
        RECT 180.035 -127.325 180.365 -126.995 ;
        RECT 180.035 -128.685 180.365 -128.355 ;
        RECT 180.035 -130.045 180.365 -129.715 ;
        RECT 180.035 -131.405 180.365 -131.075 ;
        RECT 180.035 -132.765 180.365 -132.435 ;
        RECT 180.035 -134.125 180.365 -133.795 ;
        RECT 180.035 -135.485 180.365 -135.155 ;
        RECT 180.035 -136.845 180.365 -136.515 ;
        RECT 180.035 -138.205 180.365 -137.875 ;
        RECT 180.035 -139.565 180.365 -139.235 ;
        RECT 180.035 -140.925 180.365 -140.595 ;
        RECT 180.035 -142.285 180.365 -141.955 ;
        RECT 180.035 -143.645 180.365 -143.315 ;
        RECT 180.035 -145.005 180.365 -144.675 ;
        RECT 180.035 -146.365 180.365 -146.035 ;
        RECT 180.035 -147.725 180.365 -147.395 ;
        RECT 180.035 -149.085 180.365 -148.755 ;
        RECT 180.035 -150.445 180.365 -150.115 ;
        RECT 180.035 -151.805 180.365 -151.475 ;
        RECT 180.035 -153.165 180.365 -152.835 ;
        RECT 180.035 -154.525 180.365 -154.195 ;
        RECT 180.035 -155.885 180.365 -155.555 ;
        RECT 180.035 -157.245 180.365 -156.915 ;
        RECT 180.035 -162.89 180.365 -161.76 ;
        RECT 180.04 -163.005 180.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 129.945 181.725 131.075 ;
        RECT 181.395 125.635 181.725 125.965 ;
        RECT 181.395 124.275 181.725 124.605 ;
        RECT 181.4 123.6 181.72 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 -0.845 181.725 -0.515 ;
        RECT 181.395 -2.205 181.725 -1.875 ;
        RECT 181.395 -3.565 181.725 -3.235 ;
        RECT 181.4 -3.565 181.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 129.945 183.085 131.075 ;
        RECT 182.755 125.635 183.085 125.965 ;
        RECT 182.755 124.275 183.085 124.605 ;
        RECT 182.76 123.6 183.08 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 -0.845 183.085 -0.515 ;
        RECT 182.755 -2.205 183.085 -1.875 ;
        RECT 182.755 -3.565 183.085 -3.235 ;
        RECT 182.76 -3.565 183.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 129.945 184.445 131.075 ;
        RECT 184.115 125.635 184.445 125.965 ;
        RECT 184.115 124.275 184.445 124.605 ;
        RECT 184.12 123.6 184.44 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -0.845 184.445 -0.515 ;
        RECT 184.115 -2.205 184.445 -1.875 ;
        RECT 184.115 -3.565 184.445 -3.235 ;
        RECT 184.12 -3.565 184.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -91.965 184.445 -91.635 ;
        RECT 184.115 -93.325 184.445 -92.995 ;
        RECT 184.115 -94.685 184.445 -94.355 ;
        RECT 184.115 -96.045 184.445 -95.715 ;
        RECT 184.115 -97.405 184.445 -97.075 ;
        RECT 184.115 -98.765 184.445 -98.435 ;
        RECT 184.115 -100.125 184.445 -99.795 ;
        RECT 184.115 -101.485 184.445 -101.155 ;
        RECT 184.115 -102.845 184.445 -102.515 ;
        RECT 184.115 -104.205 184.445 -103.875 ;
        RECT 184.115 -105.565 184.445 -105.235 ;
        RECT 184.115 -106.925 184.445 -106.595 ;
        RECT 184.115 -108.285 184.445 -107.955 ;
        RECT 184.115 -109.645 184.445 -109.315 ;
        RECT 184.115 -111.005 184.445 -110.675 ;
        RECT 184.115 -112.365 184.445 -112.035 ;
        RECT 184.115 -113.725 184.445 -113.395 ;
        RECT 184.115 -115.085 184.445 -114.755 ;
        RECT 184.115 -116.445 184.445 -116.115 ;
        RECT 184.115 -117.805 184.445 -117.475 ;
        RECT 184.115 -119.165 184.445 -118.835 ;
        RECT 184.115 -120.525 184.445 -120.195 ;
        RECT 184.115 -121.885 184.445 -121.555 ;
        RECT 184.115 -123.245 184.445 -122.915 ;
        RECT 184.115 -124.605 184.445 -124.275 ;
        RECT 184.115 -125.965 184.445 -125.635 ;
        RECT 184.115 -127.325 184.445 -126.995 ;
        RECT 184.115 -128.685 184.445 -128.355 ;
        RECT 184.115 -130.045 184.445 -129.715 ;
        RECT 184.115 -131.405 184.445 -131.075 ;
        RECT 184.115 -132.765 184.445 -132.435 ;
        RECT 184.115 -134.125 184.445 -133.795 ;
        RECT 184.115 -135.485 184.445 -135.155 ;
        RECT 184.115 -136.845 184.445 -136.515 ;
        RECT 184.115 -138.205 184.445 -137.875 ;
        RECT 184.115 -139.565 184.445 -139.235 ;
        RECT 184.115 -140.925 184.445 -140.595 ;
        RECT 184.115 -142.285 184.445 -141.955 ;
        RECT 184.115 -143.645 184.445 -143.315 ;
        RECT 184.115 -145.005 184.445 -144.675 ;
        RECT 184.115 -146.365 184.445 -146.035 ;
        RECT 184.115 -147.725 184.445 -147.395 ;
        RECT 184.115 -149.085 184.445 -148.755 ;
        RECT 184.115 -150.445 184.445 -150.115 ;
        RECT 184.115 -151.805 184.445 -151.475 ;
        RECT 184.115 -153.165 184.445 -152.835 ;
        RECT 184.115 -154.525 184.445 -154.195 ;
        RECT 184.115 -155.885 184.445 -155.555 ;
        RECT 184.115 -157.245 184.445 -156.915 ;
        RECT 184.115 -162.89 184.445 -161.76 ;
        RECT 184.12 -163.005 184.44 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 129.945 185.805 131.075 ;
        RECT 185.475 125.635 185.805 125.965 ;
        RECT 185.475 124.275 185.805 124.605 ;
        RECT 185.48 123.6 185.8 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 -96.045 185.805 -95.715 ;
        RECT 185.475 -97.405 185.805 -97.075 ;
        RECT 185.475 -98.765 185.805 -98.435 ;
        RECT 185.475 -100.125 185.805 -99.795 ;
        RECT 185.475 -101.485 185.805 -101.155 ;
        RECT 185.475 -102.845 185.805 -102.515 ;
        RECT 185.475 -104.205 185.805 -103.875 ;
        RECT 185.475 -105.565 185.805 -105.235 ;
        RECT 185.475 -106.925 185.805 -106.595 ;
        RECT 185.475 -108.285 185.805 -107.955 ;
        RECT 185.475 -109.645 185.805 -109.315 ;
        RECT 185.475 -111.005 185.805 -110.675 ;
        RECT 185.475 -112.365 185.805 -112.035 ;
        RECT 185.475 -113.725 185.805 -113.395 ;
        RECT 185.475 -115.085 185.805 -114.755 ;
        RECT 185.475 -116.445 185.805 -116.115 ;
        RECT 185.475 -117.805 185.805 -117.475 ;
        RECT 185.475 -119.165 185.805 -118.835 ;
        RECT 185.475 -120.525 185.805 -120.195 ;
        RECT 185.475 -121.885 185.805 -121.555 ;
        RECT 185.475 -123.245 185.805 -122.915 ;
        RECT 185.475 -124.605 185.805 -124.275 ;
        RECT 185.475 -125.965 185.805 -125.635 ;
        RECT 185.475 -127.325 185.805 -126.995 ;
        RECT 185.475 -128.685 185.805 -128.355 ;
        RECT 185.475 -130.045 185.805 -129.715 ;
        RECT 185.475 -131.405 185.805 -131.075 ;
        RECT 185.475 -132.765 185.805 -132.435 ;
        RECT 185.475 -134.125 185.805 -133.795 ;
        RECT 185.475 -135.485 185.805 -135.155 ;
        RECT 185.475 -136.845 185.805 -136.515 ;
        RECT 185.475 -138.205 185.805 -137.875 ;
        RECT 185.475 -139.565 185.805 -139.235 ;
        RECT 185.475 -140.925 185.805 -140.595 ;
        RECT 185.475 -142.285 185.805 -141.955 ;
        RECT 185.475 -143.645 185.805 -143.315 ;
        RECT 185.475 -145.005 185.805 -144.675 ;
        RECT 185.475 -146.365 185.805 -146.035 ;
        RECT 185.475 -147.725 185.805 -147.395 ;
        RECT 185.475 -149.085 185.805 -148.755 ;
        RECT 185.475 -150.445 185.805 -150.115 ;
        RECT 185.475 -151.805 185.805 -151.475 ;
        RECT 185.475 -153.165 185.805 -152.835 ;
        RECT 185.475 -154.525 185.805 -154.195 ;
        RECT 185.475 -155.885 185.805 -155.555 ;
        RECT 185.475 -157.245 185.805 -156.915 ;
        RECT 185.475 -162.89 185.805 -161.76 ;
        RECT 185.48 -163.005 185.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.66 -94.075 185.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 129.945 187.165 131.075 ;
        RECT 186.835 125.635 187.165 125.965 ;
        RECT 186.835 124.275 187.165 124.605 ;
        RECT 186.84 123.6 187.16 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 129.945 188.525 131.075 ;
        RECT 188.195 125.635 188.525 125.965 ;
        RECT 188.195 124.275 188.525 124.605 ;
        RECT 188.2 123.6 188.52 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 -0.845 188.525 -0.515 ;
        RECT 188.195 -2.205 188.525 -1.875 ;
        RECT 188.195 -3.565 188.525 -3.235 ;
        RECT 188.2 -3.565 188.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 129.945 189.885 131.075 ;
        RECT 189.555 125.635 189.885 125.965 ;
        RECT 189.555 124.275 189.885 124.605 ;
        RECT 189.56 123.6 189.88 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 -0.845 189.885 -0.515 ;
        RECT 189.555 -2.205 189.885 -1.875 ;
        RECT 189.555 -3.565 189.885 -3.235 ;
        RECT 189.56 -3.565 189.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 -91.965 189.885 -91.635 ;
        RECT 189.555 -93.325 189.885 -92.995 ;
        RECT 189.555 -94.685 189.885 -94.355 ;
        RECT 189.555 -96.045 189.885 -95.715 ;
        RECT 189.555 -97.405 189.885 -97.075 ;
        RECT 189.555 -98.765 189.885 -98.435 ;
        RECT 189.555 -100.125 189.885 -99.795 ;
        RECT 189.555 -101.485 189.885 -101.155 ;
        RECT 189.555 -102.845 189.885 -102.515 ;
        RECT 189.555 -104.205 189.885 -103.875 ;
        RECT 189.555 -105.565 189.885 -105.235 ;
        RECT 189.555 -106.925 189.885 -106.595 ;
        RECT 189.555 -108.285 189.885 -107.955 ;
        RECT 189.555 -109.645 189.885 -109.315 ;
        RECT 189.555 -111.005 189.885 -110.675 ;
        RECT 189.555 -112.365 189.885 -112.035 ;
        RECT 189.555 -113.725 189.885 -113.395 ;
        RECT 189.555 -115.085 189.885 -114.755 ;
        RECT 189.555 -116.445 189.885 -116.115 ;
        RECT 189.555 -117.805 189.885 -117.475 ;
        RECT 189.555 -119.165 189.885 -118.835 ;
        RECT 189.555 -120.525 189.885 -120.195 ;
        RECT 189.555 -121.885 189.885 -121.555 ;
        RECT 189.555 -123.245 189.885 -122.915 ;
        RECT 189.555 -124.605 189.885 -124.275 ;
        RECT 189.555 -125.965 189.885 -125.635 ;
        RECT 189.555 -127.325 189.885 -126.995 ;
        RECT 189.555 -128.685 189.885 -128.355 ;
        RECT 189.555 -130.045 189.885 -129.715 ;
        RECT 189.555 -131.405 189.885 -131.075 ;
        RECT 189.555 -132.765 189.885 -132.435 ;
        RECT 189.555 -134.125 189.885 -133.795 ;
        RECT 189.555 -135.485 189.885 -135.155 ;
        RECT 189.555 -136.845 189.885 -136.515 ;
        RECT 189.555 -138.205 189.885 -137.875 ;
        RECT 189.555 -139.565 189.885 -139.235 ;
        RECT 189.555 -140.925 189.885 -140.595 ;
        RECT 189.555 -142.285 189.885 -141.955 ;
        RECT 189.555 -143.645 189.885 -143.315 ;
        RECT 189.555 -145.005 189.885 -144.675 ;
        RECT 189.555 -146.365 189.885 -146.035 ;
        RECT 189.555 -147.725 189.885 -147.395 ;
        RECT 189.555 -149.085 189.885 -148.755 ;
        RECT 189.555 -150.445 189.885 -150.115 ;
        RECT 189.555 -151.805 189.885 -151.475 ;
        RECT 189.555 -153.165 189.885 -152.835 ;
        RECT 189.555 -154.525 189.885 -154.195 ;
        RECT 189.555 -155.885 189.885 -155.555 ;
        RECT 189.555 -157.245 189.885 -156.915 ;
        RECT 189.555 -162.89 189.885 -161.76 ;
        RECT 189.56 -163.005 189.88 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 129.945 191.245 131.075 ;
        RECT 190.915 125.635 191.245 125.965 ;
        RECT 190.915 124.275 191.245 124.605 ;
        RECT 190.92 123.6 191.24 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 -0.845 191.245 -0.515 ;
        RECT 190.915 -2.205 191.245 -1.875 ;
        RECT 190.915 -3.565 191.245 -3.235 ;
        RECT 190.92 -3.565 191.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 -91.965 191.245 -91.635 ;
        RECT 190.915 -93.325 191.245 -92.995 ;
        RECT 190.915 -94.685 191.245 -94.355 ;
        RECT 190.915 -96.045 191.245 -95.715 ;
        RECT 190.915 -97.405 191.245 -97.075 ;
        RECT 190.915 -98.765 191.245 -98.435 ;
        RECT 190.915 -100.125 191.245 -99.795 ;
        RECT 190.915 -101.485 191.245 -101.155 ;
        RECT 190.915 -102.845 191.245 -102.515 ;
        RECT 190.915 -104.205 191.245 -103.875 ;
        RECT 190.915 -105.565 191.245 -105.235 ;
        RECT 190.915 -106.925 191.245 -106.595 ;
        RECT 190.915 -108.285 191.245 -107.955 ;
        RECT 190.915 -109.645 191.245 -109.315 ;
        RECT 190.915 -111.005 191.245 -110.675 ;
        RECT 190.915 -112.365 191.245 -112.035 ;
        RECT 190.915 -113.725 191.245 -113.395 ;
        RECT 190.915 -115.085 191.245 -114.755 ;
        RECT 190.915 -116.445 191.245 -116.115 ;
        RECT 190.915 -117.805 191.245 -117.475 ;
        RECT 190.915 -119.165 191.245 -118.835 ;
        RECT 190.915 -120.525 191.245 -120.195 ;
        RECT 190.915 -121.885 191.245 -121.555 ;
        RECT 190.915 -123.245 191.245 -122.915 ;
        RECT 190.915 -124.605 191.245 -124.275 ;
        RECT 190.915 -125.965 191.245 -125.635 ;
        RECT 190.915 -127.325 191.245 -126.995 ;
        RECT 190.915 -128.685 191.245 -128.355 ;
        RECT 190.915 -130.045 191.245 -129.715 ;
        RECT 190.915 -131.405 191.245 -131.075 ;
        RECT 190.915 -132.765 191.245 -132.435 ;
        RECT 190.915 -134.125 191.245 -133.795 ;
        RECT 190.915 -135.485 191.245 -135.155 ;
        RECT 190.915 -136.845 191.245 -136.515 ;
        RECT 190.915 -138.205 191.245 -137.875 ;
        RECT 190.915 -139.565 191.245 -139.235 ;
        RECT 190.915 -140.925 191.245 -140.595 ;
        RECT 190.915 -142.285 191.245 -141.955 ;
        RECT 190.915 -143.645 191.245 -143.315 ;
        RECT 190.915 -145.005 191.245 -144.675 ;
        RECT 190.915 -146.365 191.245 -146.035 ;
        RECT 190.915 -147.725 191.245 -147.395 ;
        RECT 190.915 -149.085 191.245 -148.755 ;
        RECT 190.915 -150.445 191.245 -150.115 ;
        RECT 190.915 -151.805 191.245 -151.475 ;
        RECT 190.915 -153.165 191.245 -152.835 ;
        RECT 190.915 -154.525 191.245 -154.195 ;
        RECT 190.915 -155.885 191.245 -155.555 ;
        RECT 190.915 -157.245 191.245 -156.915 ;
        RECT 190.915 -162.89 191.245 -161.76 ;
        RECT 190.92 -163.005 191.24 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.76 -94.075 192.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 129.945 192.605 131.075 ;
        RECT 192.275 125.635 192.605 125.965 ;
        RECT 192.275 124.275 192.605 124.605 ;
        RECT 192.28 123.6 192.6 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 -96.045 192.605 -95.715 ;
        RECT 192.275 -97.405 192.605 -97.075 ;
        RECT 192.275 -98.765 192.605 -98.435 ;
        RECT 192.275 -100.125 192.605 -99.795 ;
        RECT 192.275 -101.485 192.605 -101.155 ;
        RECT 192.275 -102.845 192.605 -102.515 ;
        RECT 192.275 -104.205 192.605 -103.875 ;
        RECT 192.275 -105.565 192.605 -105.235 ;
        RECT 192.275 -106.925 192.605 -106.595 ;
        RECT 192.275 -108.285 192.605 -107.955 ;
        RECT 192.275 -109.645 192.605 -109.315 ;
        RECT 192.275 -111.005 192.605 -110.675 ;
        RECT 192.275 -112.365 192.605 -112.035 ;
        RECT 192.275 -113.725 192.605 -113.395 ;
        RECT 192.275 -115.085 192.605 -114.755 ;
        RECT 192.275 -116.445 192.605 -116.115 ;
        RECT 192.275 -117.805 192.605 -117.475 ;
        RECT 192.275 -119.165 192.605 -118.835 ;
        RECT 192.275 -120.525 192.605 -120.195 ;
        RECT 192.275 -121.885 192.605 -121.555 ;
        RECT 192.275 -123.245 192.605 -122.915 ;
        RECT 192.275 -124.605 192.605 -124.275 ;
        RECT 192.275 -125.965 192.605 -125.635 ;
        RECT 192.275 -127.325 192.605 -126.995 ;
        RECT 192.275 -128.685 192.605 -128.355 ;
        RECT 192.275 -130.045 192.605 -129.715 ;
        RECT 192.275 -131.405 192.605 -131.075 ;
        RECT 192.275 -132.765 192.605 -132.435 ;
        RECT 192.275 -134.125 192.605 -133.795 ;
        RECT 192.275 -135.485 192.605 -135.155 ;
        RECT 192.275 -136.845 192.605 -136.515 ;
        RECT 192.275 -138.205 192.605 -137.875 ;
        RECT 192.275 -139.565 192.605 -139.235 ;
        RECT 192.275 -140.925 192.605 -140.595 ;
        RECT 192.275 -142.285 192.605 -141.955 ;
        RECT 192.275 -143.645 192.605 -143.315 ;
        RECT 192.275 -145.005 192.605 -144.675 ;
        RECT 192.275 -146.365 192.605 -146.035 ;
        RECT 192.275 -147.725 192.605 -147.395 ;
        RECT 192.275 -149.085 192.605 -148.755 ;
        RECT 192.275 -150.445 192.605 -150.115 ;
        RECT 192.275 -151.805 192.605 -151.475 ;
        RECT 192.275 -153.165 192.605 -152.835 ;
        RECT 192.275 -154.525 192.605 -154.195 ;
        RECT 192.275 -155.885 192.605 -155.555 ;
        RECT 192.275 -157.245 192.605 -156.915 ;
        RECT 192.275 -162.89 192.605 -161.76 ;
        RECT 192.28 -163.005 192.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 129.945 193.965 131.075 ;
        RECT 193.635 125.635 193.965 125.965 ;
        RECT 193.635 124.275 193.965 124.605 ;
        RECT 193.64 123.6 193.96 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 -0.845 193.965 -0.515 ;
        RECT 193.635 -2.205 193.965 -1.875 ;
        RECT 193.635 -3.565 193.965 -3.235 ;
        RECT 193.64 -3.565 193.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 129.945 195.325 131.075 ;
        RECT 194.995 125.635 195.325 125.965 ;
        RECT 194.995 124.275 195.325 124.605 ;
        RECT 195 123.6 195.32 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -3.565 195.32 -0.515 ;
        RECT 194.995 -0.845 195.325 -0.515 ;
        RECT 194.995 -2.205 195.325 -1.875 ;
        RECT 194.995 -3.565 195.325 -3.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.46 -94.075 112.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 129.945 113.725 131.075 ;
        RECT 113.395 125.635 113.725 125.965 ;
        RECT 113.395 124.275 113.725 124.605 ;
        RECT 113.4 123.6 113.72 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 129.945 115.085 131.075 ;
        RECT 114.755 125.635 115.085 125.965 ;
        RECT 114.755 124.275 115.085 124.605 ;
        RECT 114.76 123.6 115.08 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 -0.845 115.085 -0.515 ;
        RECT 114.755 -2.205 115.085 -1.875 ;
        RECT 114.755 -3.565 115.085 -3.235 ;
        RECT 114.76 -3.565 115.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 129.945 116.445 131.075 ;
        RECT 116.115 125.635 116.445 125.965 ;
        RECT 116.115 124.275 116.445 124.605 ;
        RECT 116.12 123.6 116.44 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 -0.845 116.445 -0.515 ;
        RECT 116.115 -2.205 116.445 -1.875 ;
        RECT 116.115 -3.565 116.445 -3.235 ;
        RECT 116.12 -3.565 116.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 129.945 117.805 131.075 ;
        RECT 117.475 125.635 117.805 125.965 ;
        RECT 117.475 124.275 117.805 124.605 ;
        RECT 117.48 123.6 117.8 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -0.845 117.805 -0.515 ;
        RECT 117.475 -2.205 117.805 -1.875 ;
        RECT 117.475 -3.565 117.805 -3.235 ;
        RECT 117.48 -3.565 117.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -91.965 117.805 -91.635 ;
        RECT 117.475 -93.325 117.805 -92.995 ;
        RECT 117.475 -94.685 117.805 -94.355 ;
        RECT 117.475 -96.045 117.805 -95.715 ;
        RECT 117.475 -97.405 117.805 -97.075 ;
        RECT 117.475 -98.765 117.805 -98.435 ;
        RECT 117.475 -100.125 117.805 -99.795 ;
        RECT 117.475 -101.485 117.805 -101.155 ;
        RECT 117.475 -102.845 117.805 -102.515 ;
        RECT 117.475 -104.205 117.805 -103.875 ;
        RECT 117.475 -105.565 117.805 -105.235 ;
        RECT 117.475 -106.925 117.805 -106.595 ;
        RECT 117.475 -108.285 117.805 -107.955 ;
        RECT 117.475 -109.645 117.805 -109.315 ;
        RECT 117.475 -111.005 117.805 -110.675 ;
        RECT 117.475 -112.365 117.805 -112.035 ;
        RECT 117.475 -113.725 117.805 -113.395 ;
        RECT 117.475 -115.085 117.805 -114.755 ;
        RECT 117.475 -116.445 117.805 -116.115 ;
        RECT 117.475 -117.805 117.805 -117.475 ;
        RECT 117.475 -119.165 117.805 -118.835 ;
        RECT 117.475 -120.525 117.805 -120.195 ;
        RECT 117.475 -121.885 117.805 -121.555 ;
        RECT 117.475 -123.245 117.805 -122.915 ;
        RECT 117.475 -124.605 117.805 -124.275 ;
        RECT 117.475 -125.965 117.805 -125.635 ;
        RECT 117.475 -127.325 117.805 -126.995 ;
        RECT 117.475 -128.685 117.805 -128.355 ;
        RECT 117.475 -130.045 117.805 -129.715 ;
        RECT 117.475 -131.405 117.805 -131.075 ;
        RECT 117.475 -132.765 117.805 -132.435 ;
        RECT 117.475 -134.125 117.805 -133.795 ;
        RECT 117.475 -135.485 117.805 -135.155 ;
        RECT 117.475 -136.845 117.805 -136.515 ;
        RECT 117.475 -138.205 117.805 -137.875 ;
        RECT 117.475 -139.565 117.805 -139.235 ;
        RECT 117.475 -140.925 117.805 -140.595 ;
        RECT 117.475 -142.285 117.805 -141.955 ;
        RECT 117.475 -143.645 117.805 -143.315 ;
        RECT 117.475 -145.005 117.805 -144.675 ;
        RECT 117.475 -146.365 117.805 -146.035 ;
        RECT 117.475 -147.725 117.805 -147.395 ;
        RECT 117.475 -149.085 117.805 -148.755 ;
        RECT 117.475 -150.445 117.805 -150.115 ;
        RECT 117.475 -151.805 117.805 -151.475 ;
        RECT 117.475 -153.165 117.805 -152.835 ;
        RECT 117.475 -154.525 117.805 -154.195 ;
        RECT 117.475 -155.885 117.805 -155.555 ;
        RECT 117.475 -157.245 117.805 -156.915 ;
        RECT 117.475 -162.89 117.805 -161.76 ;
        RECT 117.48 -163.005 117.8 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.56 -94.075 118.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 129.945 119.165 131.075 ;
        RECT 118.835 125.635 119.165 125.965 ;
        RECT 118.835 124.275 119.165 124.605 ;
        RECT 118.84 123.6 119.16 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 -96.045 119.165 -95.715 ;
        RECT 118.835 -97.405 119.165 -97.075 ;
        RECT 118.835 -98.765 119.165 -98.435 ;
        RECT 118.835 -100.125 119.165 -99.795 ;
        RECT 118.835 -101.485 119.165 -101.155 ;
        RECT 118.835 -102.845 119.165 -102.515 ;
        RECT 118.835 -104.205 119.165 -103.875 ;
        RECT 118.835 -105.565 119.165 -105.235 ;
        RECT 118.835 -106.925 119.165 -106.595 ;
        RECT 118.835 -108.285 119.165 -107.955 ;
        RECT 118.835 -109.645 119.165 -109.315 ;
        RECT 118.835 -111.005 119.165 -110.675 ;
        RECT 118.835 -112.365 119.165 -112.035 ;
        RECT 118.835 -113.725 119.165 -113.395 ;
        RECT 118.835 -115.085 119.165 -114.755 ;
        RECT 118.835 -116.445 119.165 -116.115 ;
        RECT 118.835 -117.805 119.165 -117.475 ;
        RECT 118.835 -119.165 119.165 -118.835 ;
        RECT 118.835 -120.525 119.165 -120.195 ;
        RECT 118.835 -121.885 119.165 -121.555 ;
        RECT 118.835 -123.245 119.165 -122.915 ;
        RECT 118.835 -124.605 119.165 -124.275 ;
        RECT 118.835 -125.965 119.165 -125.635 ;
        RECT 118.835 -127.325 119.165 -126.995 ;
        RECT 118.835 -128.685 119.165 -128.355 ;
        RECT 118.835 -130.045 119.165 -129.715 ;
        RECT 118.835 -131.405 119.165 -131.075 ;
        RECT 118.835 -132.765 119.165 -132.435 ;
        RECT 118.835 -134.125 119.165 -133.795 ;
        RECT 118.835 -135.485 119.165 -135.155 ;
        RECT 118.835 -136.845 119.165 -136.515 ;
        RECT 118.835 -138.205 119.165 -137.875 ;
        RECT 118.835 -139.565 119.165 -139.235 ;
        RECT 118.835 -140.925 119.165 -140.595 ;
        RECT 118.835 -142.285 119.165 -141.955 ;
        RECT 118.835 -143.645 119.165 -143.315 ;
        RECT 118.835 -145.005 119.165 -144.675 ;
        RECT 118.835 -146.365 119.165 -146.035 ;
        RECT 118.835 -147.725 119.165 -147.395 ;
        RECT 118.835 -149.085 119.165 -148.755 ;
        RECT 118.835 -150.445 119.165 -150.115 ;
        RECT 118.835 -151.805 119.165 -151.475 ;
        RECT 118.835 -153.165 119.165 -152.835 ;
        RECT 118.835 -154.525 119.165 -154.195 ;
        RECT 118.835 -155.885 119.165 -155.555 ;
        RECT 118.835 -157.245 119.165 -156.915 ;
        RECT 118.835 -162.89 119.165 -161.76 ;
        RECT 118.84 -163.005 119.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 129.945 120.525 131.075 ;
        RECT 120.195 125.635 120.525 125.965 ;
        RECT 120.195 124.275 120.525 124.605 ;
        RECT 120.2 123.6 120.52 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 -0.845 120.525 -0.515 ;
        RECT 120.195 -2.205 120.525 -1.875 ;
        RECT 120.195 -3.565 120.525 -3.235 ;
        RECT 120.2 -3.565 120.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 129.945 121.885 131.075 ;
        RECT 121.555 125.635 121.885 125.965 ;
        RECT 121.555 124.275 121.885 124.605 ;
        RECT 121.56 123.6 121.88 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 -0.845 121.885 -0.515 ;
        RECT 121.555 -2.205 121.885 -1.875 ;
        RECT 121.555 -3.565 121.885 -3.235 ;
        RECT 121.56 -3.565 121.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 129.945 123.245 131.075 ;
        RECT 122.915 125.635 123.245 125.965 ;
        RECT 122.915 124.275 123.245 124.605 ;
        RECT 122.92 123.6 123.24 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -0.845 123.245 -0.515 ;
        RECT 122.915 -2.205 123.245 -1.875 ;
        RECT 122.915 -3.565 123.245 -3.235 ;
        RECT 122.92 -3.565 123.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -91.965 123.245 -91.635 ;
        RECT 122.915 -93.325 123.245 -92.995 ;
        RECT 122.915 -94.685 123.245 -94.355 ;
        RECT 122.915 -96.045 123.245 -95.715 ;
        RECT 122.915 -97.405 123.245 -97.075 ;
        RECT 122.915 -98.765 123.245 -98.435 ;
        RECT 122.915 -100.125 123.245 -99.795 ;
        RECT 122.915 -101.485 123.245 -101.155 ;
        RECT 122.915 -102.845 123.245 -102.515 ;
        RECT 122.915 -104.205 123.245 -103.875 ;
        RECT 122.915 -105.565 123.245 -105.235 ;
        RECT 122.915 -106.925 123.245 -106.595 ;
        RECT 122.915 -108.285 123.245 -107.955 ;
        RECT 122.915 -109.645 123.245 -109.315 ;
        RECT 122.915 -111.005 123.245 -110.675 ;
        RECT 122.915 -112.365 123.245 -112.035 ;
        RECT 122.915 -113.725 123.245 -113.395 ;
        RECT 122.915 -115.085 123.245 -114.755 ;
        RECT 122.915 -116.445 123.245 -116.115 ;
        RECT 122.915 -117.805 123.245 -117.475 ;
        RECT 122.915 -119.165 123.245 -118.835 ;
        RECT 122.915 -120.525 123.245 -120.195 ;
        RECT 122.915 -121.885 123.245 -121.555 ;
        RECT 122.915 -123.245 123.245 -122.915 ;
        RECT 122.915 -124.605 123.245 -124.275 ;
        RECT 122.915 -125.965 123.245 -125.635 ;
        RECT 122.915 -127.325 123.245 -126.995 ;
        RECT 122.915 -128.685 123.245 -128.355 ;
        RECT 122.915 -130.045 123.245 -129.715 ;
        RECT 122.915 -131.405 123.245 -131.075 ;
        RECT 122.915 -132.765 123.245 -132.435 ;
        RECT 122.915 -134.125 123.245 -133.795 ;
        RECT 122.915 -135.485 123.245 -135.155 ;
        RECT 122.915 -136.845 123.245 -136.515 ;
        RECT 122.915 -138.205 123.245 -137.875 ;
        RECT 122.915 -139.565 123.245 -139.235 ;
        RECT 122.915 -140.925 123.245 -140.595 ;
        RECT 122.915 -142.285 123.245 -141.955 ;
        RECT 122.915 -143.645 123.245 -143.315 ;
        RECT 122.915 -145.005 123.245 -144.675 ;
        RECT 122.915 -146.365 123.245 -146.035 ;
        RECT 122.915 -147.725 123.245 -147.395 ;
        RECT 122.915 -149.085 123.245 -148.755 ;
        RECT 122.915 -150.445 123.245 -150.115 ;
        RECT 122.915 -151.805 123.245 -151.475 ;
        RECT 122.915 -153.165 123.245 -152.835 ;
        RECT 122.915 -154.525 123.245 -154.195 ;
        RECT 122.915 -155.885 123.245 -155.555 ;
        RECT 122.915 -157.245 123.245 -156.915 ;
        RECT 122.915 -162.89 123.245 -161.76 ;
        RECT 122.92 -163.005 123.24 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 129.945 124.605 131.075 ;
        RECT 124.275 125.635 124.605 125.965 ;
        RECT 124.275 124.275 124.605 124.605 ;
        RECT 124.28 123.6 124.6 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 -96.045 124.605 -95.715 ;
        RECT 124.275 -97.405 124.605 -97.075 ;
        RECT 124.275 -98.765 124.605 -98.435 ;
        RECT 124.275 -100.125 124.605 -99.795 ;
        RECT 124.275 -101.485 124.605 -101.155 ;
        RECT 124.275 -102.845 124.605 -102.515 ;
        RECT 124.275 -104.205 124.605 -103.875 ;
        RECT 124.275 -105.565 124.605 -105.235 ;
        RECT 124.275 -106.925 124.605 -106.595 ;
        RECT 124.275 -108.285 124.605 -107.955 ;
        RECT 124.275 -109.645 124.605 -109.315 ;
        RECT 124.275 -111.005 124.605 -110.675 ;
        RECT 124.275 -112.365 124.605 -112.035 ;
        RECT 124.275 -113.725 124.605 -113.395 ;
        RECT 124.275 -115.085 124.605 -114.755 ;
        RECT 124.275 -116.445 124.605 -116.115 ;
        RECT 124.275 -117.805 124.605 -117.475 ;
        RECT 124.275 -119.165 124.605 -118.835 ;
        RECT 124.275 -120.525 124.605 -120.195 ;
        RECT 124.275 -121.885 124.605 -121.555 ;
        RECT 124.275 -123.245 124.605 -122.915 ;
        RECT 124.275 -124.605 124.605 -124.275 ;
        RECT 124.275 -125.965 124.605 -125.635 ;
        RECT 124.275 -127.325 124.605 -126.995 ;
        RECT 124.275 -128.685 124.605 -128.355 ;
        RECT 124.275 -130.045 124.605 -129.715 ;
        RECT 124.275 -131.405 124.605 -131.075 ;
        RECT 124.275 -132.765 124.605 -132.435 ;
        RECT 124.275 -134.125 124.605 -133.795 ;
        RECT 124.275 -135.485 124.605 -135.155 ;
        RECT 124.275 -136.845 124.605 -136.515 ;
        RECT 124.275 -138.205 124.605 -137.875 ;
        RECT 124.275 -139.565 124.605 -139.235 ;
        RECT 124.275 -140.925 124.605 -140.595 ;
        RECT 124.275 -142.285 124.605 -141.955 ;
        RECT 124.275 -143.645 124.605 -143.315 ;
        RECT 124.275 -145.005 124.605 -144.675 ;
        RECT 124.275 -146.365 124.605 -146.035 ;
        RECT 124.275 -147.725 124.605 -147.395 ;
        RECT 124.275 -149.085 124.605 -148.755 ;
        RECT 124.275 -150.445 124.605 -150.115 ;
        RECT 124.275 -151.805 124.605 -151.475 ;
        RECT 124.275 -153.165 124.605 -152.835 ;
        RECT 124.275 -154.525 124.605 -154.195 ;
        RECT 124.275 -155.885 124.605 -155.555 ;
        RECT 124.275 -157.245 124.605 -156.915 ;
        RECT 124.275 -162.89 124.605 -161.76 ;
        RECT 124.28 -163.005 124.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.66 -94.075 124.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 129.945 125.965 131.075 ;
        RECT 125.635 125.635 125.965 125.965 ;
        RECT 125.635 124.275 125.965 124.605 ;
        RECT 125.64 123.6 125.96 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 129.945 127.325 131.075 ;
        RECT 126.995 125.635 127.325 125.965 ;
        RECT 126.995 124.275 127.325 124.605 ;
        RECT 127 123.6 127.32 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 -0.845 127.325 -0.515 ;
        RECT 126.995 -2.205 127.325 -1.875 ;
        RECT 126.995 -3.565 127.325 -3.235 ;
        RECT 127 -3.565 127.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 129.945 128.685 131.075 ;
        RECT 128.355 125.635 128.685 125.965 ;
        RECT 128.355 124.275 128.685 124.605 ;
        RECT 128.36 123.6 128.68 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -0.845 128.685 -0.515 ;
        RECT 128.355 -2.205 128.685 -1.875 ;
        RECT 128.355 -3.565 128.685 -3.235 ;
        RECT 128.36 -3.565 128.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -91.965 128.685 -91.635 ;
        RECT 128.355 -93.325 128.685 -92.995 ;
        RECT 128.355 -94.685 128.685 -94.355 ;
        RECT 128.355 -96.045 128.685 -95.715 ;
        RECT 128.355 -97.405 128.685 -97.075 ;
        RECT 128.355 -98.765 128.685 -98.435 ;
        RECT 128.355 -100.125 128.685 -99.795 ;
        RECT 128.355 -101.485 128.685 -101.155 ;
        RECT 128.355 -102.845 128.685 -102.515 ;
        RECT 128.355 -104.205 128.685 -103.875 ;
        RECT 128.355 -105.565 128.685 -105.235 ;
        RECT 128.355 -106.925 128.685 -106.595 ;
        RECT 128.355 -108.285 128.685 -107.955 ;
        RECT 128.355 -109.645 128.685 -109.315 ;
        RECT 128.355 -111.005 128.685 -110.675 ;
        RECT 128.355 -112.365 128.685 -112.035 ;
        RECT 128.355 -113.725 128.685 -113.395 ;
        RECT 128.355 -115.085 128.685 -114.755 ;
        RECT 128.355 -116.445 128.685 -116.115 ;
        RECT 128.355 -117.805 128.685 -117.475 ;
        RECT 128.355 -119.165 128.685 -118.835 ;
        RECT 128.355 -120.525 128.685 -120.195 ;
        RECT 128.355 -121.885 128.685 -121.555 ;
        RECT 128.355 -123.245 128.685 -122.915 ;
        RECT 128.355 -124.605 128.685 -124.275 ;
        RECT 128.355 -125.965 128.685 -125.635 ;
        RECT 128.355 -127.325 128.685 -126.995 ;
        RECT 128.355 -128.685 128.685 -128.355 ;
        RECT 128.355 -130.045 128.685 -129.715 ;
        RECT 128.355 -131.405 128.685 -131.075 ;
        RECT 128.355 -132.765 128.685 -132.435 ;
        RECT 128.355 -134.125 128.685 -133.795 ;
        RECT 128.355 -135.485 128.685 -135.155 ;
        RECT 128.355 -136.845 128.685 -136.515 ;
        RECT 128.355 -138.205 128.685 -137.875 ;
        RECT 128.355 -139.565 128.685 -139.235 ;
        RECT 128.355 -140.925 128.685 -140.595 ;
        RECT 128.355 -142.285 128.685 -141.955 ;
        RECT 128.355 -143.645 128.685 -143.315 ;
        RECT 128.355 -145.005 128.685 -144.675 ;
        RECT 128.355 -146.365 128.685 -146.035 ;
        RECT 128.355 -147.725 128.685 -147.395 ;
        RECT 128.355 -149.085 128.685 -148.755 ;
        RECT 128.355 -150.445 128.685 -150.115 ;
        RECT 128.355 -151.805 128.685 -151.475 ;
        RECT 128.355 -153.165 128.685 -152.835 ;
        RECT 128.355 -154.525 128.685 -154.195 ;
        RECT 128.355 -155.885 128.685 -155.555 ;
        RECT 128.355 -157.245 128.685 -156.915 ;
        RECT 128.355 -162.89 128.685 -161.76 ;
        RECT 128.36 -163.005 128.68 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 129.945 130.045 131.075 ;
        RECT 129.715 125.635 130.045 125.965 ;
        RECT 129.715 124.275 130.045 124.605 ;
        RECT 129.72 123.6 130.04 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -0.845 130.045 -0.515 ;
        RECT 129.715 -2.205 130.045 -1.875 ;
        RECT 129.715 -3.565 130.045 -3.235 ;
        RECT 129.72 -3.565 130.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -91.965 130.045 -91.635 ;
        RECT 129.715 -93.325 130.045 -92.995 ;
        RECT 129.715 -94.685 130.045 -94.355 ;
        RECT 129.715 -96.045 130.045 -95.715 ;
        RECT 129.715 -97.405 130.045 -97.075 ;
        RECT 129.715 -98.765 130.045 -98.435 ;
        RECT 129.715 -100.125 130.045 -99.795 ;
        RECT 129.715 -101.485 130.045 -101.155 ;
        RECT 129.715 -102.845 130.045 -102.515 ;
        RECT 129.715 -104.205 130.045 -103.875 ;
        RECT 129.715 -105.565 130.045 -105.235 ;
        RECT 129.715 -106.925 130.045 -106.595 ;
        RECT 129.715 -108.285 130.045 -107.955 ;
        RECT 129.715 -109.645 130.045 -109.315 ;
        RECT 129.715 -111.005 130.045 -110.675 ;
        RECT 129.715 -112.365 130.045 -112.035 ;
        RECT 129.715 -113.725 130.045 -113.395 ;
        RECT 129.715 -115.085 130.045 -114.755 ;
        RECT 129.715 -116.445 130.045 -116.115 ;
        RECT 129.715 -117.805 130.045 -117.475 ;
        RECT 129.715 -119.165 130.045 -118.835 ;
        RECT 129.715 -120.525 130.045 -120.195 ;
        RECT 129.715 -121.885 130.045 -121.555 ;
        RECT 129.715 -123.245 130.045 -122.915 ;
        RECT 129.715 -124.605 130.045 -124.275 ;
        RECT 129.715 -125.965 130.045 -125.635 ;
        RECT 129.715 -127.325 130.045 -126.995 ;
        RECT 129.715 -128.685 130.045 -128.355 ;
        RECT 129.715 -130.045 130.045 -129.715 ;
        RECT 129.715 -131.405 130.045 -131.075 ;
        RECT 129.715 -132.765 130.045 -132.435 ;
        RECT 129.715 -134.125 130.045 -133.795 ;
        RECT 129.715 -135.485 130.045 -135.155 ;
        RECT 129.715 -136.845 130.045 -136.515 ;
        RECT 129.715 -138.205 130.045 -137.875 ;
        RECT 129.715 -139.565 130.045 -139.235 ;
        RECT 129.715 -140.925 130.045 -140.595 ;
        RECT 129.715 -142.285 130.045 -141.955 ;
        RECT 129.715 -143.645 130.045 -143.315 ;
        RECT 129.715 -145.005 130.045 -144.675 ;
        RECT 129.715 -146.365 130.045 -146.035 ;
        RECT 129.715 -147.725 130.045 -147.395 ;
        RECT 129.715 -149.085 130.045 -148.755 ;
        RECT 129.715 -150.445 130.045 -150.115 ;
        RECT 129.715 -151.805 130.045 -151.475 ;
        RECT 129.715 -153.165 130.045 -152.835 ;
        RECT 129.715 -154.525 130.045 -154.195 ;
        RECT 129.715 -155.885 130.045 -155.555 ;
        RECT 129.715 -157.245 130.045 -156.915 ;
        RECT 129.715 -162.89 130.045 -161.76 ;
        RECT 129.72 -163.005 130.04 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.76 -94.075 131.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 129.945 131.405 131.075 ;
        RECT 131.075 125.635 131.405 125.965 ;
        RECT 131.075 124.275 131.405 124.605 ;
        RECT 131.08 123.6 131.4 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 -96.045 131.405 -95.715 ;
        RECT 131.075 -97.405 131.405 -97.075 ;
        RECT 131.075 -98.765 131.405 -98.435 ;
        RECT 131.075 -100.125 131.405 -99.795 ;
        RECT 131.075 -101.485 131.405 -101.155 ;
        RECT 131.075 -102.845 131.405 -102.515 ;
        RECT 131.075 -104.205 131.405 -103.875 ;
        RECT 131.075 -105.565 131.405 -105.235 ;
        RECT 131.075 -106.925 131.405 -106.595 ;
        RECT 131.075 -108.285 131.405 -107.955 ;
        RECT 131.075 -109.645 131.405 -109.315 ;
        RECT 131.075 -111.005 131.405 -110.675 ;
        RECT 131.075 -112.365 131.405 -112.035 ;
        RECT 131.075 -113.725 131.405 -113.395 ;
        RECT 131.075 -115.085 131.405 -114.755 ;
        RECT 131.075 -116.445 131.405 -116.115 ;
        RECT 131.075 -117.805 131.405 -117.475 ;
        RECT 131.075 -119.165 131.405 -118.835 ;
        RECT 131.075 -120.525 131.405 -120.195 ;
        RECT 131.075 -121.885 131.405 -121.555 ;
        RECT 131.075 -123.245 131.405 -122.915 ;
        RECT 131.075 -124.605 131.405 -124.275 ;
        RECT 131.075 -125.965 131.405 -125.635 ;
        RECT 131.075 -127.325 131.405 -126.995 ;
        RECT 131.075 -128.685 131.405 -128.355 ;
        RECT 131.075 -130.045 131.405 -129.715 ;
        RECT 131.075 -131.405 131.405 -131.075 ;
        RECT 131.075 -132.765 131.405 -132.435 ;
        RECT 131.075 -134.125 131.405 -133.795 ;
        RECT 131.075 -135.485 131.405 -135.155 ;
        RECT 131.075 -136.845 131.405 -136.515 ;
        RECT 131.075 -138.205 131.405 -137.875 ;
        RECT 131.075 -139.565 131.405 -139.235 ;
        RECT 131.075 -140.925 131.405 -140.595 ;
        RECT 131.075 -142.285 131.405 -141.955 ;
        RECT 131.075 -143.645 131.405 -143.315 ;
        RECT 131.075 -145.005 131.405 -144.675 ;
        RECT 131.075 -146.365 131.405 -146.035 ;
        RECT 131.075 -147.725 131.405 -147.395 ;
        RECT 131.075 -149.085 131.405 -148.755 ;
        RECT 131.075 -150.445 131.405 -150.115 ;
        RECT 131.075 -151.805 131.405 -151.475 ;
        RECT 131.075 -153.165 131.405 -152.835 ;
        RECT 131.075 -154.525 131.405 -154.195 ;
        RECT 131.075 -155.885 131.405 -155.555 ;
        RECT 131.075 -157.245 131.405 -156.915 ;
        RECT 131.075 -162.89 131.405 -161.76 ;
        RECT 131.08 -163.005 131.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 129.945 132.765 131.075 ;
        RECT 132.435 125.635 132.765 125.965 ;
        RECT 132.435 124.275 132.765 124.605 ;
        RECT 132.44 123.6 132.76 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 -0.845 132.765 -0.515 ;
        RECT 132.435 -2.205 132.765 -1.875 ;
        RECT 132.435 -3.565 132.765 -3.235 ;
        RECT 132.44 -3.565 132.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 129.945 134.125 131.075 ;
        RECT 133.795 125.635 134.125 125.965 ;
        RECT 133.795 124.275 134.125 124.605 ;
        RECT 133.8 123.6 134.12 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 -0.845 134.125 -0.515 ;
        RECT 133.795 -2.205 134.125 -1.875 ;
        RECT 133.795 -3.565 134.125 -3.235 ;
        RECT 133.8 -3.565 134.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 129.945 135.485 131.075 ;
        RECT 135.155 125.635 135.485 125.965 ;
        RECT 135.155 124.275 135.485 124.605 ;
        RECT 135.16 123.6 135.48 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 -0.845 135.485 -0.515 ;
        RECT 135.155 -2.205 135.485 -1.875 ;
        RECT 135.155 -3.565 135.485 -3.235 ;
        RECT 135.16 -3.565 135.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 -91.965 135.485 -91.635 ;
        RECT 135.155 -93.325 135.485 -92.995 ;
        RECT 135.155 -94.685 135.485 -94.355 ;
        RECT 135.155 -96.045 135.485 -95.715 ;
        RECT 135.155 -97.405 135.485 -97.075 ;
        RECT 135.155 -98.765 135.485 -98.435 ;
        RECT 135.155 -100.125 135.485 -99.795 ;
        RECT 135.155 -101.485 135.485 -101.155 ;
        RECT 135.155 -102.845 135.485 -102.515 ;
        RECT 135.155 -104.205 135.485 -103.875 ;
        RECT 135.155 -105.565 135.485 -105.235 ;
        RECT 135.155 -106.925 135.485 -106.595 ;
        RECT 135.155 -108.285 135.485 -107.955 ;
        RECT 135.155 -109.645 135.485 -109.315 ;
        RECT 135.155 -111.005 135.485 -110.675 ;
        RECT 135.155 -112.365 135.485 -112.035 ;
        RECT 135.155 -113.725 135.485 -113.395 ;
        RECT 135.155 -115.085 135.485 -114.755 ;
        RECT 135.155 -116.445 135.485 -116.115 ;
        RECT 135.155 -117.805 135.485 -117.475 ;
        RECT 135.155 -119.165 135.485 -118.835 ;
        RECT 135.155 -120.525 135.485 -120.195 ;
        RECT 135.155 -121.885 135.485 -121.555 ;
        RECT 135.155 -123.245 135.485 -122.915 ;
        RECT 135.155 -124.605 135.485 -124.275 ;
        RECT 135.155 -125.965 135.485 -125.635 ;
        RECT 135.155 -127.325 135.485 -126.995 ;
        RECT 135.155 -128.685 135.485 -128.355 ;
        RECT 135.155 -130.045 135.485 -129.715 ;
        RECT 135.155 -131.405 135.485 -131.075 ;
        RECT 135.155 -132.765 135.485 -132.435 ;
        RECT 135.155 -134.125 135.485 -133.795 ;
        RECT 135.155 -135.485 135.485 -135.155 ;
        RECT 135.155 -136.845 135.485 -136.515 ;
        RECT 135.155 -138.205 135.485 -137.875 ;
        RECT 135.155 -139.565 135.485 -139.235 ;
        RECT 135.155 -140.925 135.485 -140.595 ;
        RECT 135.155 -142.285 135.485 -141.955 ;
        RECT 135.155 -143.645 135.485 -143.315 ;
        RECT 135.155 -145.005 135.485 -144.675 ;
        RECT 135.155 -146.365 135.485 -146.035 ;
        RECT 135.155 -147.725 135.485 -147.395 ;
        RECT 135.155 -149.085 135.485 -148.755 ;
        RECT 135.155 -150.445 135.485 -150.115 ;
        RECT 135.155 -151.805 135.485 -151.475 ;
        RECT 135.155 -153.165 135.485 -152.835 ;
        RECT 135.155 -154.525 135.485 -154.195 ;
        RECT 135.155 -155.885 135.485 -155.555 ;
        RECT 135.155 -157.245 135.485 -156.915 ;
        RECT 135.155 -162.89 135.485 -161.76 ;
        RECT 135.16 -163.005 135.48 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 129.945 136.845 131.075 ;
        RECT 136.515 125.635 136.845 125.965 ;
        RECT 136.515 124.275 136.845 124.605 ;
        RECT 136.52 123.6 136.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 -96.045 136.845 -95.715 ;
        RECT 136.515 -97.405 136.845 -97.075 ;
        RECT 136.515 -98.765 136.845 -98.435 ;
        RECT 136.515 -100.125 136.845 -99.795 ;
        RECT 136.515 -101.485 136.845 -101.155 ;
        RECT 136.515 -102.845 136.845 -102.515 ;
        RECT 136.515 -104.205 136.845 -103.875 ;
        RECT 136.515 -105.565 136.845 -105.235 ;
        RECT 136.515 -106.925 136.845 -106.595 ;
        RECT 136.515 -108.285 136.845 -107.955 ;
        RECT 136.515 -109.645 136.845 -109.315 ;
        RECT 136.515 -111.005 136.845 -110.675 ;
        RECT 136.515 -112.365 136.845 -112.035 ;
        RECT 136.515 -113.725 136.845 -113.395 ;
        RECT 136.515 -115.085 136.845 -114.755 ;
        RECT 136.515 -116.445 136.845 -116.115 ;
        RECT 136.515 -117.805 136.845 -117.475 ;
        RECT 136.515 -119.165 136.845 -118.835 ;
        RECT 136.515 -120.525 136.845 -120.195 ;
        RECT 136.515 -121.885 136.845 -121.555 ;
        RECT 136.515 -123.245 136.845 -122.915 ;
        RECT 136.515 -124.605 136.845 -124.275 ;
        RECT 136.515 -125.965 136.845 -125.635 ;
        RECT 136.515 -127.325 136.845 -126.995 ;
        RECT 136.515 -128.685 136.845 -128.355 ;
        RECT 136.515 -130.045 136.845 -129.715 ;
        RECT 136.515 -131.405 136.845 -131.075 ;
        RECT 136.515 -132.765 136.845 -132.435 ;
        RECT 136.515 -134.125 136.845 -133.795 ;
        RECT 136.515 -135.485 136.845 -135.155 ;
        RECT 136.515 -136.845 136.845 -136.515 ;
        RECT 136.515 -138.205 136.845 -137.875 ;
        RECT 136.515 -139.565 136.845 -139.235 ;
        RECT 136.515 -140.925 136.845 -140.595 ;
        RECT 136.515 -142.285 136.845 -141.955 ;
        RECT 136.515 -143.645 136.845 -143.315 ;
        RECT 136.515 -145.005 136.845 -144.675 ;
        RECT 136.515 -146.365 136.845 -146.035 ;
        RECT 136.515 -147.725 136.845 -147.395 ;
        RECT 136.515 -149.085 136.845 -148.755 ;
        RECT 136.515 -150.445 136.845 -150.115 ;
        RECT 136.515 -151.805 136.845 -151.475 ;
        RECT 136.515 -153.165 136.845 -152.835 ;
        RECT 136.515 -154.525 136.845 -154.195 ;
        RECT 136.515 -155.885 136.845 -155.555 ;
        RECT 136.515 -157.245 136.845 -156.915 ;
        RECT 136.515 -162.89 136.845 -161.76 ;
        RECT 136.52 -163.005 136.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.86 -94.075 137.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 129.945 138.205 131.075 ;
        RECT 137.875 125.635 138.205 125.965 ;
        RECT 137.875 124.275 138.205 124.605 ;
        RECT 137.88 123.6 138.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 129.945 139.565 131.075 ;
        RECT 139.235 125.635 139.565 125.965 ;
        RECT 139.235 124.275 139.565 124.605 ;
        RECT 139.24 123.6 139.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 -0.845 139.565 -0.515 ;
        RECT 139.235 -2.205 139.565 -1.875 ;
        RECT 139.235 -3.565 139.565 -3.235 ;
        RECT 139.24 -3.565 139.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 129.945 140.925 131.075 ;
        RECT 140.595 125.635 140.925 125.965 ;
        RECT 140.595 124.275 140.925 124.605 ;
        RECT 140.6 123.6 140.92 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -0.845 140.925 -0.515 ;
        RECT 140.595 -2.205 140.925 -1.875 ;
        RECT 140.595 -3.565 140.925 -3.235 ;
        RECT 140.6 -3.565 140.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -91.965 140.925 -91.635 ;
        RECT 140.595 -93.325 140.925 -92.995 ;
        RECT 140.595 -94.685 140.925 -94.355 ;
        RECT 140.595 -96.045 140.925 -95.715 ;
        RECT 140.595 -97.405 140.925 -97.075 ;
        RECT 140.595 -98.765 140.925 -98.435 ;
        RECT 140.595 -100.125 140.925 -99.795 ;
        RECT 140.595 -101.485 140.925 -101.155 ;
        RECT 140.595 -102.845 140.925 -102.515 ;
        RECT 140.595 -104.205 140.925 -103.875 ;
        RECT 140.595 -105.565 140.925 -105.235 ;
        RECT 140.595 -106.925 140.925 -106.595 ;
        RECT 140.595 -108.285 140.925 -107.955 ;
        RECT 140.595 -109.645 140.925 -109.315 ;
        RECT 140.595 -111.005 140.925 -110.675 ;
        RECT 140.595 -112.365 140.925 -112.035 ;
        RECT 140.595 -113.725 140.925 -113.395 ;
        RECT 140.595 -115.085 140.925 -114.755 ;
        RECT 140.595 -116.445 140.925 -116.115 ;
        RECT 140.595 -117.805 140.925 -117.475 ;
        RECT 140.595 -119.165 140.925 -118.835 ;
        RECT 140.595 -120.525 140.925 -120.195 ;
        RECT 140.595 -121.885 140.925 -121.555 ;
        RECT 140.595 -123.245 140.925 -122.915 ;
        RECT 140.595 -124.605 140.925 -124.275 ;
        RECT 140.595 -125.965 140.925 -125.635 ;
        RECT 140.595 -127.325 140.925 -126.995 ;
        RECT 140.595 -128.685 140.925 -128.355 ;
        RECT 140.595 -130.045 140.925 -129.715 ;
        RECT 140.595 -131.405 140.925 -131.075 ;
        RECT 140.595 -132.765 140.925 -132.435 ;
        RECT 140.595 -134.125 140.925 -133.795 ;
        RECT 140.595 -135.485 140.925 -135.155 ;
        RECT 140.595 -136.845 140.925 -136.515 ;
        RECT 140.595 -138.205 140.925 -137.875 ;
        RECT 140.595 -139.565 140.925 -139.235 ;
        RECT 140.595 -140.925 140.925 -140.595 ;
        RECT 140.595 -142.285 140.925 -141.955 ;
        RECT 140.595 -143.645 140.925 -143.315 ;
        RECT 140.595 -145.005 140.925 -144.675 ;
        RECT 140.595 -146.365 140.925 -146.035 ;
        RECT 140.595 -147.725 140.925 -147.395 ;
        RECT 140.595 -149.085 140.925 -148.755 ;
        RECT 140.595 -150.445 140.925 -150.115 ;
        RECT 140.595 -151.805 140.925 -151.475 ;
        RECT 140.595 -153.165 140.925 -152.835 ;
        RECT 140.595 -154.525 140.925 -154.195 ;
        RECT 140.595 -155.885 140.925 -155.555 ;
        RECT 140.595 -157.245 140.925 -156.915 ;
        RECT 140.595 -162.89 140.925 -161.76 ;
        RECT 140.6 -163.005 140.92 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 129.945 142.285 131.075 ;
        RECT 141.955 125.635 142.285 125.965 ;
        RECT 141.955 124.275 142.285 124.605 ;
        RECT 141.96 123.6 142.28 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -0.845 142.285 -0.515 ;
        RECT 141.955 -2.205 142.285 -1.875 ;
        RECT 141.955 -3.565 142.285 -3.235 ;
        RECT 141.96 -3.565 142.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -91.965 142.285 -91.635 ;
        RECT 141.955 -93.325 142.285 -92.995 ;
        RECT 141.955 -94.685 142.285 -94.355 ;
        RECT 141.955 -96.045 142.285 -95.715 ;
        RECT 141.955 -97.405 142.285 -97.075 ;
        RECT 141.955 -98.765 142.285 -98.435 ;
        RECT 141.955 -100.125 142.285 -99.795 ;
        RECT 141.955 -101.485 142.285 -101.155 ;
        RECT 141.955 -102.845 142.285 -102.515 ;
        RECT 141.955 -104.205 142.285 -103.875 ;
        RECT 141.955 -105.565 142.285 -105.235 ;
        RECT 141.955 -106.925 142.285 -106.595 ;
        RECT 141.955 -108.285 142.285 -107.955 ;
        RECT 141.955 -109.645 142.285 -109.315 ;
        RECT 141.955 -111.005 142.285 -110.675 ;
        RECT 141.955 -112.365 142.285 -112.035 ;
        RECT 141.955 -113.725 142.285 -113.395 ;
        RECT 141.955 -115.085 142.285 -114.755 ;
        RECT 141.955 -116.445 142.285 -116.115 ;
        RECT 141.955 -117.805 142.285 -117.475 ;
        RECT 141.955 -119.165 142.285 -118.835 ;
        RECT 141.955 -120.525 142.285 -120.195 ;
        RECT 141.955 -121.885 142.285 -121.555 ;
        RECT 141.955 -123.245 142.285 -122.915 ;
        RECT 141.955 -124.605 142.285 -124.275 ;
        RECT 141.955 -125.965 142.285 -125.635 ;
        RECT 141.955 -127.325 142.285 -126.995 ;
        RECT 141.955 -128.685 142.285 -128.355 ;
        RECT 141.955 -130.045 142.285 -129.715 ;
        RECT 141.955 -131.405 142.285 -131.075 ;
        RECT 141.955 -132.765 142.285 -132.435 ;
        RECT 141.955 -134.125 142.285 -133.795 ;
        RECT 141.955 -135.485 142.285 -135.155 ;
        RECT 141.955 -136.845 142.285 -136.515 ;
        RECT 141.955 -138.205 142.285 -137.875 ;
        RECT 141.955 -139.565 142.285 -139.235 ;
        RECT 141.955 -140.925 142.285 -140.595 ;
        RECT 141.955 -142.285 142.285 -141.955 ;
        RECT 141.955 -143.645 142.285 -143.315 ;
        RECT 141.955 -145.005 142.285 -144.675 ;
        RECT 141.955 -146.365 142.285 -146.035 ;
        RECT 141.955 -147.725 142.285 -147.395 ;
        RECT 141.955 -149.085 142.285 -148.755 ;
        RECT 141.955 -150.445 142.285 -150.115 ;
        RECT 141.955 -151.805 142.285 -151.475 ;
        RECT 141.955 -153.165 142.285 -152.835 ;
        RECT 141.955 -154.525 142.285 -154.195 ;
        RECT 141.955 -155.885 142.285 -155.555 ;
        RECT 141.955 -157.245 142.285 -156.915 ;
        RECT 141.955 -162.89 142.285 -161.76 ;
        RECT 141.96 -163.005 142.28 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.96 -94.075 143.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 129.945 143.645 131.075 ;
        RECT 143.315 125.635 143.645 125.965 ;
        RECT 143.315 124.275 143.645 124.605 ;
        RECT 143.32 123.6 143.64 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 -96.045 143.645 -95.715 ;
        RECT 143.315 -97.405 143.645 -97.075 ;
        RECT 143.315 -98.765 143.645 -98.435 ;
        RECT 143.315 -100.125 143.645 -99.795 ;
        RECT 143.315 -101.485 143.645 -101.155 ;
        RECT 143.315 -102.845 143.645 -102.515 ;
        RECT 143.315 -104.205 143.645 -103.875 ;
        RECT 143.315 -105.565 143.645 -105.235 ;
        RECT 143.315 -106.925 143.645 -106.595 ;
        RECT 143.315 -108.285 143.645 -107.955 ;
        RECT 143.315 -109.645 143.645 -109.315 ;
        RECT 143.315 -111.005 143.645 -110.675 ;
        RECT 143.315 -112.365 143.645 -112.035 ;
        RECT 143.315 -113.725 143.645 -113.395 ;
        RECT 143.315 -115.085 143.645 -114.755 ;
        RECT 143.315 -116.445 143.645 -116.115 ;
        RECT 143.315 -117.805 143.645 -117.475 ;
        RECT 143.315 -119.165 143.645 -118.835 ;
        RECT 143.315 -120.525 143.645 -120.195 ;
        RECT 143.315 -121.885 143.645 -121.555 ;
        RECT 143.315 -123.245 143.645 -122.915 ;
        RECT 143.315 -124.605 143.645 -124.275 ;
        RECT 143.315 -125.965 143.645 -125.635 ;
        RECT 143.315 -127.325 143.645 -126.995 ;
        RECT 143.315 -128.685 143.645 -128.355 ;
        RECT 143.315 -130.045 143.645 -129.715 ;
        RECT 143.315 -131.405 143.645 -131.075 ;
        RECT 143.315 -132.765 143.645 -132.435 ;
        RECT 143.315 -134.125 143.645 -133.795 ;
        RECT 143.315 -135.485 143.645 -135.155 ;
        RECT 143.315 -136.845 143.645 -136.515 ;
        RECT 143.315 -138.205 143.645 -137.875 ;
        RECT 143.315 -139.565 143.645 -139.235 ;
        RECT 143.315 -140.925 143.645 -140.595 ;
        RECT 143.315 -142.285 143.645 -141.955 ;
        RECT 143.315 -143.645 143.645 -143.315 ;
        RECT 143.315 -145.005 143.645 -144.675 ;
        RECT 143.315 -146.365 143.645 -146.035 ;
        RECT 143.315 -147.725 143.645 -147.395 ;
        RECT 143.315 -149.085 143.645 -148.755 ;
        RECT 143.315 -150.445 143.645 -150.115 ;
        RECT 143.315 -151.805 143.645 -151.475 ;
        RECT 143.315 -153.165 143.645 -152.835 ;
        RECT 143.315 -154.525 143.645 -154.195 ;
        RECT 143.315 -155.885 143.645 -155.555 ;
        RECT 143.315 -157.245 143.645 -156.915 ;
        RECT 143.315 -162.89 143.645 -161.76 ;
        RECT 143.32 -163.005 143.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 129.945 145.005 131.075 ;
        RECT 144.675 125.635 145.005 125.965 ;
        RECT 144.675 124.275 145.005 124.605 ;
        RECT 144.68 123.6 145 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 -0.845 145.005 -0.515 ;
        RECT 144.675 -2.205 145.005 -1.875 ;
        RECT 144.675 -3.565 145.005 -3.235 ;
        RECT 144.68 -3.565 145 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 129.945 146.365 131.075 ;
        RECT 146.035 125.635 146.365 125.965 ;
        RECT 146.035 124.275 146.365 124.605 ;
        RECT 146.04 123.6 146.36 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 -0.845 146.365 -0.515 ;
        RECT 146.035 -2.205 146.365 -1.875 ;
        RECT 146.035 -3.565 146.365 -3.235 ;
        RECT 146.04 -3.565 146.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 129.945 147.725 131.075 ;
        RECT 147.395 125.635 147.725 125.965 ;
        RECT 147.395 124.275 147.725 124.605 ;
        RECT 147.4 123.6 147.72 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 -0.845 147.725 -0.515 ;
        RECT 147.395 -2.205 147.725 -1.875 ;
        RECT 147.395 -3.565 147.725 -3.235 ;
        RECT 147.4 -3.565 147.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 -91.965 147.725 -91.635 ;
        RECT 147.395 -93.325 147.725 -92.995 ;
        RECT 147.395 -94.685 147.725 -94.355 ;
        RECT 147.395 -96.045 147.725 -95.715 ;
        RECT 147.395 -97.405 147.725 -97.075 ;
        RECT 147.395 -98.765 147.725 -98.435 ;
        RECT 147.395 -100.125 147.725 -99.795 ;
        RECT 147.395 -101.485 147.725 -101.155 ;
        RECT 147.395 -102.845 147.725 -102.515 ;
        RECT 147.395 -104.205 147.725 -103.875 ;
        RECT 147.395 -105.565 147.725 -105.235 ;
        RECT 147.395 -106.925 147.725 -106.595 ;
        RECT 147.395 -108.285 147.725 -107.955 ;
        RECT 147.395 -109.645 147.725 -109.315 ;
        RECT 147.395 -111.005 147.725 -110.675 ;
        RECT 147.395 -112.365 147.725 -112.035 ;
        RECT 147.395 -113.725 147.725 -113.395 ;
        RECT 147.395 -115.085 147.725 -114.755 ;
        RECT 147.395 -116.445 147.725 -116.115 ;
        RECT 147.395 -117.805 147.725 -117.475 ;
        RECT 147.395 -119.165 147.725 -118.835 ;
        RECT 147.395 -120.525 147.725 -120.195 ;
        RECT 147.395 -121.885 147.725 -121.555 ;
        RECT 147.395 -123.245 147.725 -122.915 ;
        RECT 147.395 -124.605 147.725 -124.275 ;
        RECT 147.395 -125.965 147.725 -125.635 ;
        RECT 147.395 -127.325 147.725 -126.995 ;
        RECT 147.395 -128.685 147.725 -128.355 ;
        RECT 147.395 -130.045 147.725 -129.715 ;
        RECT 147.395 -131.405 147.725 -131.075 ;
        RECT 147.395 -132.765 147.725 -132.435 ;
        RECT 147.395 -134.125 147.725 -133.795 ;
        RECT 147.395 -135.485 147.725 -135.155 ;
        RECT 147.395 -136.845 147.725 -136.515 ;
        RECT 147.395 -138.205 147.725 -137.875 ;
        RECT 147.395 -139.565 147.725 -139.235 ;
        RECT 147.395 -140.925 147.725 -140.595 ;
        RECT 147.395 -142.285 147.725 -141.955 ;
        RECT 147.395 -143.645 147.725 -143.315 ;
        RECT 147.395 -145.005 147.725 -144.675 ;
        RECT 147.395 -146.365 147.725 -146.035 ;
        RECT 147.395 -147.725 147.725 -147.395 ;
        RECT 147.395 -149.085 147.725 -148.755 ;
        RECT 147.395 -150.445 147.725 -150.115 ;
        RECT 147.395 -151.805 147.725 -151.475 ;
        RECT 147.395 -153.165 147.725 -152.835 ;
        RECT 147.395 -154.525 147.725 -154.195 ;
        RECT 147.395 -155.885 147.725 -155.555 ;
        RECT 147.395 -157.245 147.725 -156.915 ;
        RECT 147.395 -162.89 147.725 -161.76 ;
        RECT 147.4 -163.005 147.72 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 129.945 149.085 131.075 ;
        RECT 148.755 125.635 149.085 125.965 ;
        RECT 148.755 124.275 149.085 124.605 ;
        RECT 148.76 123.6 149.08 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 -96.045 149.085 -95.715 ;
        RECT 148.755 -97.405 149.085 -97.075 ;
        RECT 148.755 -98.765 149.085 -98.435 ;
        RECT 148.755 -100.125 149.085 -99.795 ;
        RECT 148.755 -101.485 149.085 -101.155 ;
        RECT 148.755 -102.845 149.085 -102.515 ;
        RECT 148.755 -104.205 149.085 -103.875 ;
        RECT 148.755 -105.565 149.085 -105.235 ;
        RECT 148.755 -106.925 149.085 -106.595 ;
        RECT 148.755 -108.285 149.085 -107.955 ;
        RECT 148.755 -109.645 149.085 -109.315 ;
        RECT 148.755 -111.005 149.085 -110.675 ;
        RECT 148.755 -112.365 149.085 -112.035 ;
        RECT 148.755 -113.725 149.085 -113.395 ;
        RECT 148.755 -115.085 149.085 -114.755 ;
        RECT 148.755 -116.445 149.085 -116.115 ;
        RECT 148.755 -117.805 149.085 -117.475 ;
        RECT 148.755 -119.165 149.085 -118.835 ;
        RECT 148.755 -120.525 149.085 -120.195 ;
        RECT 148.755 -121.885 149.085 -121.555 ;
        RECT 148.755 -123.245 149.085 -122.915 ;
        RECT 148.755 -124.605 149.085 -124.275 ;
        RECT 148.755 -125.965 149.085 -125.635 ;
        RECT 148.755 -127.325 149.085 -126.995 ;
        RECT 148.755 -128.685 149.085 -128.355 ;
        RECT 148.755 -130.045 149.085 -129.715 ;
        RECT 148.755 -131.405 149.085 -131.075 ;
        RECT 148.755 -132.765 149.085 -132.435 ;
        RECT 148.755 -134.125 149.085 -133.795 ;
        RECT 148.755 -135.485 149.085 -135.155 ;
        RECT 148.755 -136.845 149.085 -136.515 ;
        RECT 148.755 -138.205 149.085 -137.875 ;
        RECT 148.755 -139.565 149.085 -139.235 ;
        RECT 148.755 -140.925 149.085 -140.595 ;
        RECT 148.755 -142.285 149.085 -141.955 ;
        RECT 148.755 -143.645 149.085 -143.315 ;
        RECT 148.755 -145.005 149.085 -144.675 ;
        RECT 148.755 -146.365 149.085 -146.035 ;
        RECT 148.755 -147.725 149.085 -147.395 ;
        RECT 148.755 -149.085 149.085 -148.755 ;
        RECT 148.755 -150.445 149.085 -150.115 ;
        RECT 148.755 -151.805 149.085 -151.475 ;
        RECT 148.755 -153.165 149.085 -152.835 ;
        RECT 148.755 -154.525 149.085 -154.195 ;
        RECT 148.755 -155.885 149.085 -155.555 ;
        RECT 148.755 -157.245 149.085 -156.915 ;
        RECT 148.755 -162.89 149.085 -161.76 ;
        RECT 148.76 -163.005 149.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.06 -94.075 149.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 129.945 150.445 131.075 ;
        RECT 150.115 125.635 150.445 125.965 ;
        RECT 150.115 124.275 150.445 124.605 ;
        RECT 150.12 123.6 150.44 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 129.945 151.805 131.075 ;
        RECT 151.475 125.635 151.805 125.965 ;
        RECT 151.475 124.275 151.805 124.605 ;
        RECT 151.48 123.6 151.8 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 -0.845 151.805 -0.515 ;
        RECT 151.475 -2.205 151.805 -1.875 ;
        RECT 151.475 -3.565 151.805 -3.235 ;
        RECT 151.48 -3.565 151.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 129.945 153.165 131.075 ;
        RECT 152.835 125.635 153.165 125.965 ;
        RECT 152.835 124.275 153.165 124.605 ;
        RECT 152.84 123.6 153.16 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 -0.845 153.165 -0.515 ;
        RECT 152.835 -2.205 153.165 -1.875 ;
        RECT 152.835 -3.565 153.165 -3.235 ;
        RECT 152.84 -3.565 153.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 129.945 154.525 131.075 ;
        RECT 154.195 125.635 154.525 125.965 ;
        RECT 154.195 124.275 154.525 124.605 ;
        RECT 154.2 123.6 154.52 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -0.845 154.525 -0.515 ;
        RECT 154.195 -2.205 154.525 -1.875 ;
        RECT 154.195 -3.565 154.525 -3.235 ;
        RECT 154.2 -3.565 154.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -93.325 154.525 -92.995 ;
        RECT 154.195 -94.685 154.525 -94.355 ;
        RECT 154.195 -96.045 154.525 -95.715 ;
        RECT 154.195 -97.405 154.525 -97.075 ;
        RECT 154.195 -98.765 154.525 -98.435 ;
        RECT 154.195 -100.125 154.525 -99.795 ;
        RECT 154.195 -101.485 154.525 -101.155 ;
        RECT 154.195 -102.845 154.525 -102.515 ;
        RECT 154.195 -104.205 154.525 -103.875 ;
        RECT 154.195 -105.565 154.525 -105.235 ;
        RECT 154.195 -106.925 154.525 -106.595 ;
        RECT 154.195 -108.285 154.525 -107.955 ;
        RECT 154.195 -109.645 154.525 -109.315 ;
        RECT 154.195 -111.005 154.525 -110.675 ;
        RECT 154.195 -112.365 154.525 -112.035 ;
        RECT 154.195 -113.725 154.525 -113.395 ;
        RECT 154.195 -115.085 154.525 -114.755 ;
        RECT 154.195 -116.445 154.525 -116.115 ;
        RECT 154.195 -117.805 154.525 -117.475 ;
        RECT 154.195 -119.165 154.525 -118.835 ;
        RECT 154.195 -120.525 154.525 -120.195 ;
        RECT 154.195 -121.885 154.525 -121.555 ;
        RECT 154.195 -123.245 154.525 -122.915 ;
        RECT 154.195 -124.605 154.525 -124.275 ;
        RECT 154.195 -125.965 154.525 -125.635 ;
        RECT 154.195 -127.325 154.525 -126.995 ;
        RECT 154.195 -128.685 154.525 -128.355 ;
        RECT 154.195 -130.045 154.525 -129.715 ;
        RECT 154.195 -131.405 154.525 -131.075 ;
        RECT 154.195 -132.765 154.525 -132.435 ;
        RECT 154.195 -134.125 154.525 -133.795 ;
        RECT 154.195 -135.485 154.525 -135.155 ;
        RECT 154.195 -136.845 154.525 -136.515 ;
        RECT 154.195 -138.205 154.525 -137.875 ;
        RECT 154.195 -139.565 154.525 -139.235 ;
        RECT 154.195 -140.925 154.525 -140.595 ;
        RECT 154.195 -142.285 154.525 -141.955 ;
        RECT 154.195 -143.645 154.525 -143.315 ;
        RECT 154.195 -145.005 154.525 -144.675 ;
        RECT 154.195 -146.365 154.525 -146.035 ;
        RECT 154.195 -147.725 154.525 -147.395 ;
        RECT 154.195 -149.085 154.525 -148.755 ;
        RECT 154.195 -150.445 154.525 -150.115 ;
        RECT 154.195 -151.805 154.525 -151.475 ;
        RECT 154.195 -153.165 154.525 -152.835 ;
        RECT 154.195 -154.525 154.525 -154.195 ;
        RECT 154.195 -155.885 154.525 -155.555 ;
        RECT 154.195 -157.245 154.525 -156.915 ;
        RECT 154.195 -162.89 154.525 -161.76 ;
        RECT 154.2 -163.005 154.52 -90.96 ;
        RECT 154.195 -91.965 154.525 -91.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -91.965 74.285 -91.635 ;
        RECT 73.955 -93.325 74.285 -92.995 ;
        RECT 73.955 -94.685 74.285 -94.355 ;
        RECT 73.955 -96.045 74.285 -95.715 ;
        RECT 73.955 -97.405 74.285 -97.075 ;
        RECT 73.955 -98.765 74.285 -98.435 ;
        RECT 73.955 -100.125 74.285 -99.795 ;
        RECT 73.955 -101.485 74.285 -101.155 ;
        RECT 73.955 -102.845 74.285 -102.515 ;
        RECT 73.955 -104.205 74.285 -103.875 ;
        RECT 73.955 -105.565 74.285 -105.235 ;
        RECT 73.955 -106.925 74.285 -106.595 ;
        RECT 73.955 -108.285 74.285 -107.955 ;
        RECT 73.955 -109.645 74.285 -109.315 ;
        RECT 73.955 -111.005 74.285 -110.675 ;
        RECT 73.955 -112.365 74.285 -112.035 ;
        RECT 73.955 -113.725 74.285 -113.395 ;
        RECT 73.955 -115.085 74.285 -114.755 ;
        RECT 73.955 -116.445 74.285 -116.115 ;
        RECT 73.955 -117.805 74.285 -117.475 ;
        RECT 73.955 -119.165 74.285 -118.835 ;
        RECT 73.955 -120.525 74.285 -120.195 ;
        RECT 73.955 -121.885 74.285 -121.555 ;
        RECT 73.955 -123.245 74.285 -122.915 ;
        RECT 73.955 -124.605 74.285 -124.275 ;
        RECT 73.955 -125.965 74.285 -125.635 ;
        RECT 73.955 -127.325 74.285 -126.995 ;
        RECT 73.955 -128.685 74.285 -128.355 ;
        RECT 73.955 -130.045 74.285 -129.715 ;
        RECT 73.955 -131.405 74.285 -131.075 ;
        RECT 73.955 -132.765 74.285 -132.435 ;
        RECT 73.955 -134.125 74.285 -133.795 ;
        RECT 73.955 -135.485 74.285 -135.155 ;
        RECT 73.955 -136.845 74.285 -136.515 ;
        RECT 73.955 -138.205 74.285 -137.875 ;
        RECT 73.955 -139.565 74.285 -139.235 ;
        RECT 73.955 -140.925 74.285 -140.595 ;
        RECT 73.955 -142.285 74.285 -141.955 ;
        RECT 73.955 -143.645 74.285 -143.315 ;
        RECT 73.955 -145.005 74.285 -144.675 ;
        RECT 73.955 -146.365 74.285 -146.035 ;
        RECT 73.955 -147.725 74.285 -147.395 ;
        RECT 73.955 -149.085 74.285 -148.755 ;
        RECT 73.955 -150.445 74.285 -150.115 ;
        RECT 73.955 -151.805 74.285 -151.475 ;
        RECT 73.955 -153.165 74.285 -152.835 ;
        RECT 73.955 -154.525 74.285 -154.195 ;
        RECT 73.955 -155.885 74.285 -155.555 ;
        RECT 73.955 -157.245 74.285 -156.915 ;
        RECT 73.955 -162.89 74.285 -161.76 ;
        RECT 73.96 -163.005 74.28 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 129.945 75.645 131.075 ;
        RECT 75.315 125.635 75.645 125.965 ;
        RECT 75.315 124.275 75.645 124.605 ;
        RECT 75.32 123.6 75.64 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 -96.045 75.645 -95.715 ;
        RECT 75.315 -97.405 75.645 -97.075 ;
        RECT 75.315 -98.765 75.645 -98.435 ;
        RECT 75.315 -100.125 75.645 -99.795 ;
        RECT 75.315 -101.485 75.645 -101.155 ;
        RECT 75.315 -102.845 75.645 -102.515 ;
        RECT 75.315 -104.205 75.645 -103.875 ;
        RECT 75.315 -105.565 75.645 -105.235 ;
        RECT 75.315 -106.925 75.645 -106.595 ;
        RECT 75.315 -108.285 75.645 -107.955 ;
        RECT 75.315 -109.645 75.645 -109.315 ;
        RECT 75.315 -111.005 75.645 -110.675 ;
        RECT 75.315 -112.365 75.645 -112.035 ;
        RECT 75.315 -113.725 75.645 -113.395 ;
        RECT 75.315 -115.085 75.645 -114.755 ;
        RECT 75.315 -116.445 75.645 -116.115 ;
        RECT 75.315 -117.805 75.645 -117.475 ;
        RECT 75.315 -119.165 75.645 -118.835 ;
        RECT 75.315 -120.525 75.645 -120.195 ;
        RECT 75.315 -121.885 75.645 -121.555 ;
        RECT 75.315 -123.245 75.645 -122.915 ;
        RECT 75.315 -124.605 75.645 -124.275 ;
        RECT 75.315 -125.965 75.645 -125.635 ;
        RECT 75.315 -127.325 75.645 -126.995 ;
        RECT 75.315 -128.685 75.645 -128.355 ;
        RECT 75.315 -130.045 75.645 -129.715 ;
        RECT 75.315 -131.405 75.645 -131.075 ;
        RECT 75.315 -132.765 75.645 -132.435 ;
        RECT 75.315 -134.125 75.645 -133.795 ;
        RECT 75.315 -135.485 75.645 -135.155 ;
        RECT 75.315 -136.845 75.645 -136.515 ;
        RECT 75.315 -138.205 75.645 -137.875 ;
        RECT 75.315 -139.565 75.645 -139.235 ;
        RECT 75.315 -140.925 75.645 -140.595 ;
        RECT 75.315 -142.285 75.645 -141.955 ;
        RECT 75.315 -143.645 75.645 -143.315 ;
        RECT 75.315 -145.005 75.645 -144.675 ;
        RECT 75.315 -146.365 75.645 -146.035 ;
        RECT 75.315 -147.725 75.645 -147.395 ;
        RECT 75.315 -149.085 75.645 -148.755 ;
        RECT 75.315 -150.445 75.645 -150.115 ;
        RECT 75.315 -151.805 75.645 -151.475 ;
        RECT 75.315 -153.165 75.645 -152.835 ;
        RECT 75.315 -154.525 75.645 -154.195 ;
        RECT 75.315 -155.885 75.645 -155.555 ;
        RECT 75.315 -157.245 75.645 -156.915 ;
        RECT 75.315 -162.89 75.645 -161.76 ;
        RECT 75.32 -163.005 75.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.86 -94.075 76.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 129.945 77.005 131.075 ;
        RECT 76.675 125.635 77.005 125.965 ;
        RECT 76.675 124.275 77.005 124.605 ;
        RECT 76.68 123.6 77 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 129.945 78.365 131.075 ;
        RECT 78.035 125.635 78.365 125.965 ;
        RECT 78.035 124.275 78.365 124.605 ;
        RECT 78.04 123.6 78.36 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -0.845 78.365 -0.515 ;
        RECT 78.035 -2.205 78.365 -1.875 ;
        RECT 78.035 -3.565 78.365 -3.235 ;
        RECT 78.04 -3.565 78.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -91.965 78.365 -91.635 ;
        RECT 78.035 -93.325 78.365 -92.995 ;
        RECT 78.035 -94.685 78.365 -94.355 ;
        RECT 78.035 -96.045 78.365 -95.715 ;
        RECT 78.035 -97.405 78.365 -97.075 ;
        RECT 78.035 -98.765 78.365 -98.435 ;
        RECT 78.035 -100.125 78.365 -99.795 ;
        RECT 78.035 -101.485 78.365 -101.155 ;
        RECT 78.035 -102.845 78.365 -102.515 ;
        RECT 78.035 -104.205 78.365 -103.875 ;
        RECT 78.035 -105.565 78.365 -105.235 ;
        RECT 78.035 -106.925 78.365 -106.595 ;
        RECT 78.035 -108.285 78.365 -107.955 ;
        RECT 78.035 -109.645 78.365 -109.315 ;
        RECT 78.035 -111.005 78.365 -110.675 ;
        RECT 78.035 -112.365 78.365 -112.035 ;
        RECT 78.035 -113.725 78.365 -113.395 ;
        RECT 78.035 -115.085 78.365 -114.755 ;
        RECT 78.035 -116.445 78.365 -116.115 ;
        RECT 78.035 -117.805 78.365 -117.475 ;
        RECT 78.035 -119.165 78.365 -118.835 ;
        RECT 78.035 -120.525 78.365 -120.195 ;
        RECT 78.035 -121.885 78.365 -121.555 ;
        RECT 78.035 -123.245 78.365 -122.915 ;
        RECT 78.035 -124.605 78.365 -124.275 ;
        RECT 78.035 -125.965 78.365 -125.635 ;
        RECT 78.035 -127.325 78.365 -126.995 ;
        RECT 78.035 -128.685 78.365 -128.355 ;
        RECT 78.035 -130.045 78.365 -129.715 ;
        RECT 78.035 -131.405 78.365 -131.075 ;
        RECT 78.035 -132.765 78.365 -132.435 ;
        RECT 78.035 -134.125 78.365 -133.795 ;
        RECT 78.035 -135.485 78.365 -135.155 ;
        RECT 78.035 -136.845 78.365 -136.515 ;
        RECT 78.035 -138.205 78.365 -137.875 ;
        RECT 78.035 -139.565 78.365 -139.235 ;
        RECT 78.035 -140.925 78.365 -140.595 ;
        RECT 78.035 -142.285 78.365 -141.955 ;
        RECT 78.035 -143.645 78.365 -143.315 ;
        RECT 78.035 -145.005 78.365 -144.675 ;
        RECT 78.035 -146.365 78.365 -146.035 ;
        RECT 78.035 -147.725 78.365 -147.395 ;
        RECT 78.035 -149.085 78.365 -148.755 ;
        RECT 78.035 -150.445 78.365 -150.115 ;
        RECT 78.035 -151.805 78.365 -151.475 ;
        RECT 78.035 -153.165 78.365 -152.835 ;
        RECT 78.035 -154.525 78.365 -154.195 ;
        RECT 78.035 -155.885 78.365 -155.555 ;
        RECT 78.035 -157.245 78.365 -156.915 ;
        RECT 78.035 -162.89 78.365 -161.76 ;
        RECT 78.04 -163.005 78.36 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 129.945 79.725 131.075 ;
        RECT 79.395 125.635 79.725 125.965 ;
        RECT 79.395 124.275 79.725 124.605 ;
        RECT 79.4 123.6 79.72 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 -0.845 79.725 -0.515 ;
        RECT 79.395 -2.205 79.725 -1.875 ;
        RECT 79.395 -3.565 79.725 -3.235 ;
        RECT 79.4 -3.565 79.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 129.945 81.085 131.075 ;
        RECT 80.755 125.635 81.085 125.965 ;
        RECT 80.755 124.275 81.085 124.605 ;
        RECT 80.76 123.6 81.08 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 -0.845 81.085 -0.515 ;
        RECT 80.755 -2.205 81.085 -1.875 ;
        RECT 80.755 -3.565 81.085 -3.235 ;
        RECT 80.76 -3.565 81.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 -91.965 81.085 -91.635 ;
        RECT 80.755 -93.325 81.085 -92.995 ;
        RECT 80.755 -94.685 81.085 -94.355 ;
        RECT 80.755 -96.045 81.085 -95.715 ;
        RECT 80.755 -97.405 81.085 -97.075 ;
        RECT 80.755 -98.765 81.085 -98.435 ;
        RECT 80.755 -100.125 81.085 -99.795 ;
        RECT 80.755 -101.485 81.085 -101.155 ;
        RECT 80.755 -102.845 81.085 -102.515 ;
        RECT 80.755 -104.205 81.085 -103.875 ;
        RECT 80.755 -105.565 81.085 -105.235 ;
        RECT 80.755 -106.925 81.085 -106.595 ;
        RECT 80.755 -108.285 81.085 -107.955 ;
        RECT 80.755 -109.645 81.085 -109.315 ;
        RECT 80.755 -111.005 81.085 -110.675 ;
        RECT 80.755 -112.365 81.085 -112.035 ;
        RECT 80.755 -113.725 81.085 -113.395 ;
        RECT 80.755 -115.085 81.085 -114.755 ;
        RECT 80.755 -116.445 81.085 -116.115 ;
        RECT 80.755 -117.805 81.085 -117.475 ;
        RECT 80.755 -119.165 81.085 -118.835 ;
        RECT 80.755 -120.525 81.085 -120.195 ;
        RECT 80.755 -121.885 81.085 -121.555 ;
        RECT 80.755 -123.245 81.085 -122.915 ;
        RECT 80.755 -124.605 81.085 -124.275 ;
        RECT 80.755 -125.965 81.085 -125.635 ;
        RECT 80.755 -127.325 81.085 -126.995 ;
        RECT 80.755 -128.685 81.085 -128.355 ;
        RECT 80.755 -130.045 81.085 -129.715 ;
        RECT 80.755 -131.405 81.085 -131.075 ;
        RECT 80.755 -132.765 81.085 -132.435 ;
        RECT 80.755 -134.125 81.085 -133.795 ;
        RECT 80.755 -135.485 81.085 -135.155 ;
        RECT 80.755 -136.845 81.085 -136.515 ;
        RECT 80.755 -138.205 81.085 -137.875 ;
        RECT 80.755 -139.565 81.085 -139.235 ;
        RECT 80.755 -140.925 81.085 -140.595 ;
        RECT 80.755 -142.285 81.085 -141.955 ;
        RECT 80.755 -143.645 81.085 -143.315 ;
        RECT 80.755 -145.005 81.085 -144.675 ;
        RECT 80.755 -146.365 81.085 -146.035 ;
        RECT 80.755 -147.725 81.085 -147.395 ;
        RECT 80.755 -149.085 81.085 -148.755 ;
        RECT 80.755 -150.445 81.085 -150.115 ;
        RECT 80.755 -151.805 81.085 -151.475 ;
        RECT 80.755 -153.165 81.085 -152.835 ;
        RECT 80.755 -154.525 81.085 -154.195 ;
        RECT 80.755 -155.885 81.085 -155.555 ;
        RECT 80.755 -157.245 81.085 -156.915 ;
        RECT 80.755 -162.89 81.085 -161.76 ;
        RECT 80.76 -163.005 81.08 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.96 -94.075 82.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 129.945 82.445 131.075 ;
        RECT 82.115 125.635 82.445 125.965 ;
        RECT 82.115 124.275 82.445 124.605 ;
        RECT 82.12 123.6 82.44 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 -96.045 82.445 -95.715 ;
        RECT 82.115 -97.405 82.445 -97.075 ;
        RECT 82.115 -98.765 82.445 -98.435 ;
        RECT 82.115 -100.125 82.445 -99.795 ;
        RECT 82.115 -101.485 82.445 -101.155 ;
        RECT 82.115 -102.845 82.445 -102.515 ;
        RECT 82.115 -104.205 82.445 -103.875 ;
        RECT 82.115 -105.565 82.445 -105.235 ;
        RECT 82.115 -106.925 82.445 -106.595 ;
        RECT 82.115 -108.285 82.445 -107.955 ;
        RECT 82.115 -109.645 82.445 -109.315 ;
        RECT 82.115 -111.005 82.445 -110.675 ;
        RECT 82.115 -112.365 82.445 -112.035 ;
        RECT 82.115 -113.725 82.445 -113.395 ;
        RECT 82.115 -115.085 82.445 -114.755 ;
        RECT 82.115 -116.445 82.445 -116.115 ;
        RECT 82.115 -117.805 82.445 -117.475 ;
        RECT 82.115 -119.165 82.445 -118.835 ;
        RECT 82.115 -120.525 82.445 -120.195 ;
        RECT 82.115 -121.885 82.445 -121.555 ;
        RECT 82.115 -123.245 82.445 -122.915 ;
        RECT 82.115 -124.605 82.445 -124.275 ;
        RECT 82.115 -125.965 82.445 -125.635 ;
        RECT 82.115 -127.325 82.445 -126.995 ;
        RECT 82.115 -128.685 82.445 -128.355 ;
        RECT 82.115 -130.045 82.445 -129.715 ;
        RECT 82.115 -131.405 82.445 -131.075 ;
        RECT 82.115 -132.765 82.445 -132.435 ;
        RECT 82.115 -134.125 82.445 -133.795 ;
        RECT 82.115 -135.485 82.445 -135.155 ;
        RECT 82.115 -136.845 82.445 -136.515 ;
        RECT 82.115 -138.205 82.445 -137.875 ;
        RECT 82.115 -139.565 82.445 -139.235 ;
        RECT 82.115 -140.925 82.445 -140.595 ;
        RECT 82.115 -142.285 82.445 -141.955 ;
        RECT 82.115 -143.645 82.445 -143.315 ;
        RECT 82.115 -145.005 82.445 -144.675 ;
        RECT 82.115 -146.365 82.445 -146.035 ;
        RECT 82.115 -147.725 82.445 -147.395 ;
        RECT 82.115 -149.085 82.445 -148.755 ;
        RECT 82.115 -150.445 82.445 -150.115 ;
        RECT 82.115 -151.805 82.445 -151.475 ;
        RECT 82.115 -153.165 82.445 -152.835 ;
        RECT 82.115 -154.525 82.445 -154.195 ;
        RECT 82.115 -155.885 82.445 -155.555 ;
        RECT 82.115 -157.245 82.445 -156.915 ;
        RECT 82.115 -162.89 82.445 -161.76 ;
        RECT 82.12 -163.005 82.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 129.945 83.805 131.075 ;
        RECT 83.475 125.635 83.805 125.965 ;
        RECT 83.475 124.275 83.805 124.605 ;
        RECT 83.48 123.6 83.8 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 -0.845 83.805 -0.515 ;
        RECT 83.475 -2.205 83.805 -1.875 ;
        RECT 83.475 -3.565 83.805 -3.235 ;
        RECT 83.48 -3.565 83.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 129.945 85.165 131.075 ;
        RECT 84.835 125.635 85.165 125.965 ;
        RECT 84.835 124.275 85.165 124.605 ;
        RECT 84.84 123.6 85.16 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 -0.845 85.165 -0.515 ;
        RECT 84.835 -2.205 85.165 -1.875 ;
        RECT 84.835 -3.565 85.165 -3.235 ;
        RECT 84.84 -3.565 85.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 129.945 86.525 131.075 ;
        RECT 86.195 125.635 86.525 125.965 ;
        RECT 86.195 124.275 86.525 124.605 ;
        RECT 86.2 123.6 86.52 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -0.845 86.525 -0.515 ;
        RECT 86.195 -2.205 86.525 -1.875 ;
        RECT 86.195 -3.565 86.525 -3.235 ;
        RECT 86.2 -3.565 86.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -91.965 86.525 -91.635 ;
        RECT 86.195 -93.325 86.525 -92.995 ;
        RECT 86.195 -94.685 86.525 -94.355 ;
        RECT 86.195 -96.045 86.525 -95.715 ;
        RECT 86.195 -97.405 86.525 -97.075 ;
        RECT 86.195 -98.765 86.525 -98.435 ;
        RECT 86.195 -100.125 86.525 -99.795 ;
        RECT 86.195 -101.485 86.525 -101.155 ;
        RECT 86.195 -102.845 86.525 -102.515 ;
        RECT 86.195 -104.205 86.525 -103.875 ;
        RECT 86.195 -105.565 86.525 -105.235 ;
        RECT 86.195 -106.925 86.525 -106.595 ;
        RECT 86.195 -108.285 86.525 -107.955 ;
        RECT 86.195 -109.645 86.525 -109.315 ;
        RECT 86.195 -111.005 86.525 -110.675 ;
        RECT 86.195 -112.365 86.525 -112.035 ;
        RECT 86.195 -113.725 86.525 -113.395 ;
        RECT 86.195 -115.085 86.525 -114.755 ;
        RECT 86.195 -116.445 86.525 -116.115 ;
        RECT 86.195 -117.805 86.525 -117.475 ;
        RECT 86.195 -119.165 86.525 -118.835 ;
        RECT 86.195 -120.525 86.525 -120.195 ;
        RECT 86.195 -121.885 86.525 -121.555 ;
        RECT 86.195 -123.245 86.525 -122.915 ;
        RECT 86.195 -124.605 86.525 -124.275 ;
        RECT 86.195 -125.965 86.525 -125.635 ;
        RECT 86.195 -127.325 86.525 -126.995 ;
        RECT 86.195 -128.685 86.525 -128.355 ;
        RECT 86.195 -130.045 86.525 -129.715 ;
        RECT 86.195 -131.405 86.525 -131.075 ;
        RECT 86.195 -132.765 86.525 -132.435 ;
        RECT 86.195 -134.125 86.525 -133.795 ;
        RECT 86.195 -135.485 86.525 -135.155 ;
        RECT 86.195 -136.845 86.525 -136.515 ;
        RECT 86.195 -138.205 86.525 -137.875 ;
        RECT 86.195 -139.565 86.525 -139.235 ;
        RECT 86.195 -140.925 86.525 -140.595 ;
        RECT 86.195 -142.285 86.525 -141.955 ;
        RECT 86.195 -143.645 86.525 -143.315 ;
        RECT 86.195 -145.005 86.525 -144.675 ;
        RECT 86.195 -146.365 86.525 -146.035 ;
        RECT 86.195 -147.725 86.525 -147.395 ;
        RECT 86.195 -149.085 86.525 -148.755 ;
        RECT 86.195 -150.445 86.525 -150.115 ;
        RECT 86.195 -151.805 86.525 -151.475 ;
        RECT 86.195 -153.165 86.525 -152.835 ;
        RECT 86.195 -154.525 86.525 -154.195 ;
        RECT 86.195 -155.885 86.525 -155.555 ;
        RECT 86.195 -157.245 86.525 -156.915 ;
        RECT 86.195 -162.89 86.525 -161.76 ;
        RECT 86.2 -163.005 86.52 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 129.945 87.885 131.075 ;
        RECT 87.555 125.635 87.885 125.965 ;
        RECT 87.555 124.275 87.885 124.605 ;
        RECT 87.56 123.6 87.88 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 -96.045 87.885 -95.715 ;
        RECT 87.555 -97.405 87.885 -97.075 ;
        RECT 87.555 -98.765 87.885 -98.435 ;
        RECT 87.555 -100.125 87.885 -99.795 ;
        RECT 87.555 -101.485 87.885 -101.155 ;
        RECT 87.555 -102.845 87.885 -102.515 ;
        RECT 87.555 -104.205 87.885 -103.875 ;
        RECT 87.555 -105.565 87.885 -105.235 ;
        RECT 87.555 -106.925 87.885 -106.595 ;
        RECT 87.555 -108.285 87.885 -107.955 ;
        RECT 87.555 -109.645 87.885 -109.315 ;
        RECT 87.555 -111.005 87.885 -110.675 ;
        RECT 87.555 -112.365 87.885 -112.035 ;
        RECT 87.555 -113.725 87.885 -113.395 ;
        RECT 87.555 -115.085 87.885 -114.755 ;
        RECT 87.555 -116.445 87.885 -116.115 ;
        RECT 87.555 -117.805 87.885 -117.475 ;
        RECT 87.555 -119.165 87.885 -118.835 ;
        RECT 87.555 -120.525 87.885 -120.195 ;
        RECT 87.555 -121.885 87.885 -121.555 ;
        RECT 87.555 -123.245 87.885 -122.915 ;
        RECT 87.555 -124.605 87.885 -124.275 ;
        RECT 87.555 -125.965 87.885 -125.635 ;
        RECT 87.555 -127.325 87.885 -126.995 ;
        RECT 87.555 -128.685 87.885 -128.355 ;
        RECT 87.555 -130.045 87.885 -129.715 ;
        RECT 87.555 -131.405 87.885 -131.075 ;
        RECT 87.555 -132.765 87.885 -132.435 ;
        RECT 87.555 -134.125 87.885 -133.795 ;
        RECT 87.555 -135.485 87.885 -135.155 ;
        RECT 87.555 -136.845 87.885 -136.515 ;
        RECT 87.555 -138.205 87.885 -137.875 ;
        RECT 87.555 -139.565 87.885 -139.235 ;
        RECT 87.555 -140.925 87.885 -140.595 ;
        RECT 87.555 -142.285 87.885 -141.955 ;
        RECT 87.555 -143.645 87.885 -143.315 ;
        RECT 87.555 -145.005 87.885 -144.675 ;
        RECT 87.555 -146.365 87.885 -146.035 ;
        RECT 87.555 -147.725 87.885 -147.395 ;
        RECT 87.555 -149.085 87.885 -148.755 ;
        RECT 87.555 -150.445 87.885 -150.115 ;
        RECT 87.555 -151.805 87.885 -151.475 ;
        RECT 87.555 -153.165 87.885 -152.835 ;
        RECT 87.555 -154.525 87.885 -154.195 ;
        RECT 87.555 -155.885 87.885 -155.555 ;
        RECT 87.555 -157.245 87.885 -156.915 ;
        RECT 87.555 -162.89 87.885 -161.76 ;
        RECT 87.56 -163.005 87.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.06 -94.075 88.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 129.945 89.245 131.075 ;
        RECT 88.915 125.635 89.245 125.965 ;
        RECT 88.915 124.275 89.245 124.605 ;
        RECT 88.92 123.6 89.24 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 129.945 90.605 131.075 ;
        RECT 90.275 125.635 90.605 125.965 ;
        RECT 90.275 124.275 90.605 124.605 ;
        RECT 90.28 123.6 90.6 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 -0.845 90.605 -0.515 ;
        RECT 90.275 -2.205 90.605 -1.875 ;
        RECT 90.275 -3.565 90.605 -3.235 ;
        RECT 90.28 -3.565 90.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 -91.965 90.605 -91.635 ;
        RECT 90.275 -93.325 90.605 -92.995 ;
        RECT 90.275 -94.685 90.605 -94.355 ;
        RECT 90.275 -96.045 90.605 -95.715 ;
        RECT 90.275 -97.405 90.605 -97.075 ;
        RECT 90.275 -98.765 90.605 -98.435 ;
        RECT 90.275 -100.125 90.605 -99.795 ;
        RECT 90.275 -101.485 90.605 -101.155 ;
        RECT 90.275 -102.845 90.605 -102.515 ;
        RECT 90.275 -104.205 90.605 -103.875 ;
        RECT 90.275 -105.565 90.605 -105.235 ;
        RECT 90.275 -106.925 90.605 -106.595 ;
        RECT 90.275 -108.285 90.605 -107.955 ;
        RECT 90.275 -109.645 90.605 -109.315 ;
        RECT 90.275 -111.005 90.605 -110.675 ;
        RECT 90.275 -112.365 90.605 -112.035 ;
        RECT 90.275 -113.725 90.605 -113.395 ;
        RECT 90.275 -115.085 90.605 -114.755 ;
        RECT 90.275 -116.445 90.605 -116.115 ;
        RECT 90.275 -117.805 90.605 -117.475 ;
        RECT 90.275 -119.165 90.605 -118.835 ;
        RECT 90.275 -120.525 90.605 -120.195 ;
        RECT 90.275 -121.885 90.605 -121.555 ;
        RECT 90.275 -123.245 90.605 -122.915 ;
        RECT 90.275 -124.605 90.605 -124.275 ;
        RECT 90.275 -125.965 90.605 -125.635 ;
        RECT 90.275 -127.325 90.605 -126.995 ;
        RECT 90.275 -128.685 90.605 -128.355 ;
        RECT 90.275 -130.045 90.605 -129.715 ;
        RECT 90.275 -131.405 90.605 -131.075 ;
        RECT 90.275 -132.765 90.605 -132.435 ;
        RECT 90.275 -134.125 90.605 -133.795 ;
        RECT 90.275 -135.485 90.605 -135.155 ;
        RECT 90.275 -136.845 90.605 -136.515 ;
        RECT 90.275 -138.205 90.605 -137.875 ;
        RECT 90.275 -139.565 90.605 -139.235 ;
        RECT 90.275 -140.925 90.605 -140.595 ;
        RECT 90.275 -142.285 90.605 -141.955 ;
        RECT 90.275 -143.645 90.605 -143.315 ;
        RECT 90.275 -145.005 90.605 -144.675 ;
        RECT 90.275 -146.365 90.605 -146.035 ;
        RECT 90.275 -147.725 90.605 -147.395 ;
        RECT 90.275 -149.085 90.605 -148.755 ;
        RECT 90.275 -150.445 90.605 -150.115 ;
        RECT 90.275 -151.805 90.605 -151.475 ;
        RECT 90.275 -153.165 90.605 -152.835 ;
        RECT 90.275 -154.525 90.605 -154.195 ;
        RECT 90.275 -155.885 90.605 -155.555 ;
        RECT 90.275 -157.245 90.605 -156.915 ;
        RECT 90.275 -162.89 90.605 -161.76 ;
        RECT 90.28 -163.005 90.6 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 129.945 91.965 131.075 ;
        RECT 91.635 125.635 91.965 125.965 ;
        RECT 91.635 124.275 91.965 124.605 ;
        RECT 91.64 123.6 91.96 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 -0.845 91.965 -0.515 ;
        RECT 91.635 -2.205 91.965 -1.875 ;
        RECT 91.635 -3.565 91.965 -3.235 ;
        RECT 91.64 -3.565 91.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 129.945 93.325 131.075 ;
        RECT 92.995 125.635 93.325 125.965 ;
        RECT 92.995 124.275 93.325 124.605 ;
        RECT 93 123.6 93.32 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 -0.845 93.325 -0.515 ;
        RECT 92.995 -2.205 93.325 -1.875 ;
        RECT 92.995 -3.565 93.325 -3.235 ;
        RECT 93 -3.565 93.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 -91.965 93.325 -91.635 ;
        RECT 92.995 -93.325 93.325 -92.995 ;
        RECT 92.995 -94.685 93.325 -94.355 ;
        RECT 92.995 -96.045 93.325 -95.715 ;
        RECT 92.995 -97.405 93.325 -97.075 ;
        RECT 92.995 -98.765 93.325 -98.435 ;
        RECT 92.995 -100.125 93.325 -99.795 ;
        RECT 92.995 -101.485 93.325 -101.155 ;
        RECT 92.995 -102.845 93.325 -102.515 ;
        RECT 92.995 -104.205 93.325 -103.875 ;
        RECT 92.995 -105.565 93.325 -105.235 ;
        RECT 92.995 -106.925 93.325 -106.595 ;
        RECT 92.995 -108.285 93.325 -107.955 ;
        RECT 92.995 -109.645 93.325 -109.315 ;
        RECT 92.995 -111.005 93.325 -110.675 ;
        RECT 92.995 -112.365 93.325 -112.035 ;
        RECT 92.995 -113.725 93.325 -113.395 ;
        RECT 92.995 -115.085 93.325 -114.755 ;
        RECT 92.995 -116.445 93.325 -116.115 ;
        RECT 92.995 -117.805 93.325 -117.475 ;
        RECT 92.995 -119.165 93.325 -118.835 ;
        RECT 92.995 -120.525 93.325 -120.195 ;
        RECT 92.995 -121.885 93.325 -121.555 ;
        RECT 92.995 -123.245 93.325 -122.915 ;
        RECT 92.995 -124.605 93.325 -124.275 ;
        RECT 92.995 -125.965 93.325 -125.635 ;
        RECT 92.995 -127.325 93.325 -126.995 ;
        RECT 92.995 -128.685 93.325 -128.355 ;
        RECT 92.995 -130.045 93.325 -129.715 ;
        RECT 92.995 -131.405 93.325 -131.075 ;
        RECT 92.995 -132.765 93.325 -132.435 ;
        RECT 92.995 -134.125 93.325 -133.795 ;
        RECT 92.995 -135.485 93.325 -135.155 ;
        RECT 92.995 -136.845 93.325 -136.515 ;
        RECT 92.995 -138.205 93.325 -137.875 ;
        RECT 92.995 -139.565 93.325 -139.235 ;
        RECT 92.995 -140.925 93.325 -140.595 ;
        RECT 92.995 -142.285 93.325 -141.955 ;
        RECT 92.995 -143.645 93.325 -143.315 ;
        RECT 92.995 -145.005 93.325 -144.675 ;
        RECT 92.995 -146.365 93.325 -146.035 ;
        RECT 92.995 -147.725 93.325 -147.395 ;
        RECT 92.995 -149.085 93.325 -148.755 ;
        RECT 92.995 -150.445 93.325 -150.115 ;
        RECT 92.995 -151.805 93.325 -151.475 ;
        RECT 92.995 -153.165 93.325 -152.835 ;
        RECT 92.995 -154.525 93.325 -154.195 ;
        RECT 92.995 -155.885 93.325 -155.555 ;
        RECT 92.995 -157.245 93.325 -156.915 ;
        RECT 92.995 -162.89 93.325 -161.76 ;
        RECT 93 -163.005 93.32 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.16 -94.075 94.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 129.945 94.685 131.075 ;
        RECT 94.355 125.635 94.685 125.965 ;
        RECT 94.355 124.275 94.685 124.605 ;
        RECT 94.36 123.6 94.68 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 -96.045 94.685 -95.715 ;
        RECT 94.355 -97.405 94.685 -97.075 ;
        RECT 94.355 -98.765 94.685 -98.435 ;
        RECT 94.355 -100.125 94.685 -99.795 ;
        RECT 94.355 -101.485 94.685 -101.155 ;
        RECT 94.355 -102.845 94.685 -102.515 ;
        RECT 94.355 -104.205 94.685 -103.875 ;
        RECT 94.355 -105.565 94.685 -105.235 ;
        RECT 94.355 -106.925 94.685 -106.595 ;
        RECT 94.355 -108.285 94.685 -107.955 ;
        RECT 94.355 -109.645 94.685 -109.315 ;
        RECT 94.355 -111.005 94.685 -110.675 ;
        RECT 94.355 -112.365 94.685 -112.035 ;
        RECT 94.355 -113.725 94.685 -113.395 ;
        RECT 94.355 -115.085 94.685 -114.755 ;
        RECT 94.355 -116.445 94.685 -116.115 ;
        RECT 94.355 -117.805 94.685 -117.475 ;
        RECT 94.355 -119.165 94.685 -118.835 ;
        RECT 94.355 -120.525 94.685 -120.195 ;
        RECT 94.355 -121.885 94.685 -121.555 ;
        RECT 94.355 -123.245 94.685 -122.915 ;
        RECT 94.355 -124.605 94.685 -124.275 ;
        RECT 94.355 -125.965 94.685 -125.635 ;
        RECT 94.355 -127.325 94.685 -126.995 ;
        RECT 94.355 -128.685 94.685 -128.355 ;
        RECT 94.355 -130.045 94.685 -129.715 ;
        RECT 94.355 -131.405 94.685 -131.075 ;
        RECT 94.355 -132.765 94.685 -132.435 ;
        RECT 94.355 -134.125 94.685 -133.795 ;
        RECT 94.355 -135.485 94.685 -135.155 ;
        RECT 94.355 -136.845 94.685 -136.515 ;
        RECT 94.355 -138.205 94.685 -137.875 ;
        RECT 94.355 -139.565 94.685 -139.235 ;
        RECT 94.355 -140.925 94.685 -140.595 ;
        RECT 94.355 -142.285 94.685 -141.955 ;
        RECT 94.355 -143.645 94.685 -143.315 ;
        RECT 94.355 -145.005 94.685 -144.675 ;
        RECT 94.355 -146.365 94.685 -146.035 ;
        RECT 94.355 -147.725 94.685 -147.395 ;
        RECT 94.355 -149.085 94.685 -148.755 ;
        RECT 94.355 -150.445 94.685 -150.115 ;
        RECT 94.355 -151.805 94.685 -151.475 ;
        RECT 94.355 -153.165 94.685 -152.835 ;
        RECT 94.355 -154.525 94.685 -154.195 ;
        RECT 94.355 -155.885 94.685 -155.555 ;
        RECT 94.355 -157.245 94.685 -156.915 ;
        RECT 94.355 -162.89 94.685 -161.76 ;
        RECT 94.36 -163.005 94.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 129.945 96.045 131.075 ;
        RECT 95.715 125.635 96.045 125.965 ;
        RECT 95.715 124.275 96.045 124.605 ;
        RECT 95.72 123.6 96.04 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 -0.845 96.045 -0.515 ;
        RECT 95.715 -2.205 96.045 -1.875 ;
        RECT 95.715 -3.565 96.045 -3.235 ;
        RECT 95.72 -3.565 96.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 129.945 97.405 131.075 ;
        RECT 97.075 125.635 97.405 125.965 ;
        RECT 97.075 124.275 97.405 124.605 ;
        RECT 97.08 123.6 97.4 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 -0.845 97.405 -0.515 ;
        RECT 97.075 -2.205 97.405 -1.875 ;
        RECT 97.075 -3.565 97.405 -3.235 ;
        RECT 97.08 -3.565 97.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 129.945 98.765 131.075 ;
        RECT 98.435 125.635 98.765 125.965 ;
        RECT 98.435 124.275 98.765 124.605 ;
        RECT 98.44 123.6 98.76 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -0.845 98.765 -0.515 ;
        RECT 98.435 -2.205 98.765 -1.875 ;
        RECT 98.435 -3.565 98.765 -3.235 ;
        RECT 98.44 -3.565 98.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -91.965 98.765 -91.635 ;
        RECT 98.435 -93.325 98.765 -92.995 ;
        RECT 98.435 -94.685 98.765 -94.355 ;
        RECT 98.435 -96.045 98.765 -95.715 ;
        RECT 98.435 -97.405 98.765 -97.075 ;
        RECT 98.435 -98.765 98.765 -98.435 ;
        RECT 98.435 -100.125 98.765 -99.795 ;
        RECT 98.435 -101.485 98.765 -101.155 ;
        RECT 98.435 -102.845 98.765 -102.515 ;
        RECT 98.435 -104.205 98.765 -103.875 ;
        RECT 98.435 -105.565 98.765 -105.235 ;
        RECT 98.435 -106.925 98.765 -106.595 ;
        RECT 98.435 -108.285 98.765 -107.955 ;
        RECT 98.435 -109.645 98.765 -109.315 ;
        RECT 98.435 -111.005 98.765 -110.675 ;
        RECT 98.435 -112.365 98.765 -112.035 ;
        RECT 98.435 -113.725 98.765 -113.395 ;
        RECT 98.435 -115.085 98.765 -114.755 ;
        RECT 98.435 -116.445 98.765 -116.115 ;
        RECT 98.435 -117.805 98.765 -117.475 ;
        RECT 98.435 -119.165 98.765 -118.835 ;
        RECT 98.435 -120.525 98.765 -120.195 ;
        RECT 98.435 -121.885 98.765 -121.555 ;
        RECT 98.435 -123.245 98.765 -122.915 ;
        RECT 98.435 -124.605 98.765 -124.275 ;
        RECT 98.435 -125.965 98.765 -125.635 ;
        RECT 98.435 -127.325 98.765 -126.995 ;
        RECT 98.435 -128.685 98.765 -128.355 ;
        RECT 98.435 -130.045 98.765 -129.715 ;
        RECT 98.435 -131.405 98.765 -131.075 ;
        RECT 98.435 -132.765 98.765 -132.435 ;
        RECT 98.435 -134.125 98.765 -133.795 ;
        RECT 98.435 -135.485 98.765 -135.155 ;
        RECT 98.435 -136.845 98.765 -136.515 ;
        RECT 98.435 -138.205 98.765 -137.875 ;
        RECT 98.435 -139.565 98.765 -139.235 ;
        RECT 98.435 -140.925 98.765 -140.595 ;
        RECT 98.435 -142.285 98.765 -141.955 ;
        RECT 98.435 -143.645 98.765 -143.315 ;
        RECT 98.435 -145.005 98.765 -144.675 ;
        RECT 98.435 -146.365 98.765 -146.035 ;
        RECT 98.435 -147.725 98.765 -147.395 ;
        RECT 98.435 -149.085 98.765 -148.755 ;
        RECT 98.435 -150.445 98.765 -150.115 ;
        RECT 98.435 -151.805 98.765 -151.475 ;
        RECT 98.435 -153.165 98.765 -152.835 ;
        RECT 98.435 -154.525 98.765 -154.195 ;
        RECT 98.435 -155.885 98.765 -155.555 ;
        RECT 98.435 -157.245 98.765 -156.915 ;
        RECT 98.435 -162.89 98.765 -161.76 ;
        RECT 98.44 -163.005 98.76 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 129.945 100.125 131.075 ;
        RECT 99.795 125.635 100.125 125.965 ;
        RECT 99.795 124.275 100.125 124.605 ;
        RECT 99.8 123.6 100.12 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 -96.045 100.125 -95.715 ;
        RECT 99.795 -97.405 100.125 -97.075 ;
        RECT 99.795 -98.765 100.125 -98.435 ;
        RECT 99.795 -100.125 100.125 -99.795 ;
        RECT 99.795 -101.485 100.125 -101.155 ;
        RECT 99.795 -102.845 100.125 -102.515 ;
        RECT 99.795 -104.205 100.125 -103.875 ;
        RECT 99.795 -105.565 100.125 -105.235 ;
        RECT 99.795 -106.925 100.125 -106.595 ;
        RECT 99.795 -108.285 100.125 -107.955 ;
        RECT 99.795 -109.645 100.125 -109.315 ;
        RECT 99.795 -111.005 100.125 -110.675 ;
        RECT 99.795 -112.365 100.125 -112.035 ;
        RECT 99.795 -113.725 100.125 -113.395 ;
        RECT 99.795 -115.085 100.125 -114.755 ;
        RECT 99.795 -116.445 100.125 -116.115 ;
        RECT 99.795 -117.805 100.125 -117.475 ;
        RECT 99.795 -119.165 100.125 -118.835 ;
        RECT 99.795 -120.525 100.125 -120.195 ;
        RECT 99.795 -121.885 100.125 -121.555 ;
        RECT 99.795 -123.245 100.125 -122.915 ;
        RECT 99.795 -124.605 100.125 -124.275 ;
        RECT 99.795 -125.965 100.125 -125.635 ;
        RECT 99.795 -127.325 100.125 -126.995 ;
        RECT 99.795 -128.685 100.125 -128.355 ;
        RECT 99.795 -130.045 100.125 -129.715 ;
        RECT 99.795 -131.405 100.125 -131.075 ;
        RECT 99.795 -132.765 100.125 -132.435 ;
        RECT 99.795 -134.125 100.125 -133.795 ;
        RECT 99.795 -135.485 100.125 -135.155 ;
        RECT 99.795 -136.845 100.125 -136.515 ;
        RECT 99.795 -138.205 100.125 -137.875 ;
        RECT 99.795 -139.565 100.125 -139.235 ;
        RECT 99.795 -140.925 100.125 -140.595 ;
        RECT 99.795 -142.285 100.125 -141.955 ;
        RECT 99.795 -143.645 100.125 -143.315 ;
        RECT 99.795 -145.005 100.125 -144.675 ;
        RECT 99.795 -146.365 100.125 -146.035 ;
        RECT 99.795 -147.725 100.125 -147.395 ;
        RECT 99.795 -149.085 100.125 -148.755 ;
        RECT 99.795 -150.445 100.125 -150.115 ;
        RECT 99.795 -151.805 100.125 -151.475 ;
        RECT 99.795 -153.165 100.125 -152.835 ;
        RECT 99.795 -154.525 100.125 -154.195 ;
        RECT 99.795 -155.885 100.125 -155.555 ;
        RECT 99.795 -157.245 100.125 -156.915 ;
        RECT 99.795 -162.89 100.125 -161.76 ;
        RECT 99.8 -163.005 100.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.26 -94.075 100.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 129.945 101.485 131.075 ;
        RECT 101.155 125.635 101.485 125.965 ;
        RECT 101.155 124.275 101.485 124.605 ;
        RECT 101.16 123.6 101.48 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 129.945 102.845 131.075 ;
        RECT 102.515 125.635 102.845 125.965 ;
        RECT 102.515 124.275 102.845 124.605 ;
        RECT 102.52 123.6 102.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 -0.845 102.845 -0.515 ;
        RECT 102.515 -2.205 102.845 -1.875 ;
        RECT 102.515 -3.565 102.845 -3.235 ;
        RECT 102.52 -3.565 102.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 -91.965 102.845 -91.635 ;
        RECT 102.515 -93.325 102.845 -92.995 ;
        RECT 102.515 -94.685 102.845 -94.355 ;
        RECT 102.515 -96.045 102.845 -95.715 ;
        RECT 102.515 -97.405 102.845 -97.075 ;
        RECT 102.515 -98.765 102.845 -98.435 ;
        RECT 102.515 -100.125 102.845 -99.795 ;
        RECT 102.515 -101.485 102.845 -101.155 ;
        RECT 102.515 -102.845 102.845 -102.515 ;
        RECT 102.515 -104.205 102.845 -103.875 ;
        RECT 102.515 -105.565 102.845 -105.235 ;
        RECT 102.515 -106.925 102.845 -106.595 ;
        RECT 102.515 -108.285 102.845 -107.955 ;
        RECT 102.515 -109.645 102.845 -109.315 ;
        RECT 102.515 -111.005 102.845 -110.675 ;
        RECT 102.515 -112.365 102.845 -112.035 ;
        RECT 102.515 -113.725 102.845 -113.395 ;
        RECT 102.515 -115.085 102.845 -114.755 ;
        RECT 102.515 -116.445 102.845 -116.115 ;
        RECT 102.515 -117.805 102.845 -117.475 ;
        RECT 102.515 -119.165 102.845 -118.835 ;
        RECT 102.515 -120.525 102.845 -120.195 ;
        RECT 102.515 -121.885 102.845 -121.555 ;
        RECT 102.515 -123.245 102.845 -122.915 ;
        RECT 102.515 -124.605 102.845 -124.275 ;
        RECT 102.515 -125.965 102.845 -125.635 ;
        RECT 102.515 -127.325 102.845 -126.995 ;
        RECT 102.515 -128.685 102.845 -128.355 ;
        RECT 102.515 -130.045 102.845 -129.715 ;
        RECT 102.515 -131.405 102.845 -131.075 ;
        RECT 102.515 -132.765 102.845 -132.435 ;
        RECT 102.515 -134.125 102.845 -133.795 ;
        RECT 102.515 -135.485 102.845 -135.155 ;
        RECT 102.515 -136.845 102.845 -136.515 ;
        RECT 102.515 -138.205 102.845 -137.875 ;
        RECT 102.515 -139.565 102.845 -139.235 ;
        RECT 102.515 -140.925 102.845 -140.595 ;
        RECT 102.515 -142.285 102.845 -141.955 ;
        RECT 102.515 -143.645 102.845 -143.315 ;
        RECT 102.515 -145.005 102.845 -144.675 ;
        RECT 102.515 -146.365 102.845 -146.035 ;
        RECT 102.515 -147.725 102.845 -147.395 ;
        RECT 102.515 -149.085 102.845 -148.755 ;
        RECT 102.515 -150.445 102.845 -150.115 ;
        RECT 102.515 -151.805 102.845 -151.475 ;
        RECT 102.515 -153.165 102.845 -152.835 ;
        RECT 102.515 -154.525 102.845 -154.195 ;
        RECT 102.515 -155.885 102.845 -155.555 ;
        RECT 102.515 -157.245 102.845 -156.915 ;
        RECT 102.515 -162.89 102.845 -161.76 ;
        RECT 102.52 -163.005 102.84 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 129.945 104.205 131.075 ;
        RECT 103.875 125.635 104.205 125.965 ;
        RECT 103.875 124.275 104.205 124.605 ;
        RECT 103.88 123.6 104.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 -0.845 104.205 -0.515 ;
        RECT 103.875 -2.205 104.205 -1.875 ;
        RECT 103.875 -3.565 104.205 -3.235 ;
        RECT 103.88 -3.565 104.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 129.945 105.565 131.075 ;
        RECT 105.235 125.635 105.565 125.965 ;
        RECT 105.235 124.275 105.565 124.605 ;
        RECT 105.24 123.6 105.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -0.845 105.565 -0.515 ;
        RECT 105.235 -2.205 105.565 -1.875 ;
        RECT 105.235 -3.565 105.565 -3.235 ;
        RECT 105.24 -3.565 105.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -91.965 105.565 -91.635 ;
        RECT 105.235 -93.325 105.565 -92.995 ;
        RECT 105.235 -94.685 105.565 -94.355 ;
        RECT 105.235 -96.045 105.565 -95.715 ;
        RECT 105.235 -97.405 105.565 -97.075 ;
        RECT 105.235 -98.765 105.565 -98.435 ;
        RECT 105.235 -100.125 105.565 -99.795 ;
        RECT 105.235 -101.485 105.565 -101.155 ;
        RECT 105.235 -102.845 105.565 -102.515 ;
        RECT 105.235 -104.205 105.565 -103.875 ;
        RECT 105.235 -105.565 105.565 -105.235 ;
        RECT 105.235 -106.925 105.565 -106.595 ;
        RECT 105.235 -108.285 105.565 -107.955 ;
        RECT 105.235 -109.645 105.565 -109.315 ;
        RECT 105.235 -111.005 105.565 -110.675 ;
        RECT 105.235 -112.365 105.565 -112.035 ;
        RECT 105.235 -113.725 105.565 -113.395 ;
        RECT 105.235 -115.085 105.565 -114.755 ;
        RECT 105.235 -116.445 105.565 -116.115 ;
        RECT 105.235 -117.805 105.565 -117.475 ;
        RECT 105.235 -119.165 105.565 -118.835 ;
        RECT 105.235 -120.525 105.565 -120.195 ;
        RECT 105.235 -121.885 105.565 -121.555 ;
        RECT 105.235 -123.245 105.565 -122.915 ;
        RECT 105.235 -124.605 105.565 -124.275 ;
        RECT 105.235 -125.965 105.565 -125.635 ;
        RECT 105.235 -127.325 105.565 -126.995 ;
        RECT 105.235 -128.685 105.565 -128.355 ;
        RECT 105.235 -130.045 105.565 -129.715 ;
        RECT 105.235 -131.405 105.565 -131.075 ;
        RECT 105.235 -132.765 105.565 -132.435 ;
        RECT 105.235 -134.125 105.565 -133.795 ;
        RECT 105.235 -135.485 105.565 -135.155 ;
        RECT 105.235 -136.845 105.565 -136.515 ;
        RECT 105.235 -138.205 105.565 -137.875 ;
        RECT 105.235 -139.565 105.565 -139.235 ;
        RECT 105.235 -140.925 105.565 -140.595 ;
        RECT 105.235 -142.285 105.565 -141.955 ;
        RECT 105.235 -143.645 105.565 -143.315 ;
        RECT 105.235 -145.005 105.565 -144.675 ;
        RECT 105.235 -146.365 105.565 -146.035 ;
        RECT 105.235 -147.725 105.565 -147.395 ;
        RECT 105.235 -149.085 105.565 -148.755 ;
        RECT 105.235 -150.445 105.565 -150.115 ;
        RECT 105.235 -151.805 105.565 -151.475 ;
        RECT 105.235 -153.165 105.565 -152.835 ;
        RECT 105.235 -154.525 105.565 -154.195 ;
        RECT 105.235 -155.885 105.565 -155.555 ;
        RECT 105.235 -157.245 105.565 -156.915 ;
        RECT 105.235 -162.89 105.565 -161.76 ;
        RECT 105.24 -163.005 105.56 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.36 -94.075 106.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 129.945 106.925 131.075 ;
        RECT 106.595 125.635 106.925 125.965 ;
        RECT 106.595 124.275 106.925 124.605 ;
        RECT 106.6 123.6 106.92 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 -96.045 106.925 -95.715 ;
        RECT 106.595 -97.405 106.925 -97.075 ;
        RECT 106.595 -98.765 106.925 -98.435 ;
        RECT 106.595 -100.125 106.925 -99.795 ;
        RECT 106.595 -101.485 106.925 -101.155 ;
        RECT 106.595 -102.845 106.925 -102.515 ;
        RECT 106.595 -104.205 106.925 -103.875 ;
        RECT 106.595 -105.565 106.925 -105.235 ;
        RECT 106.595 -106.925 106.925 -106.595 ;
        RECT 106.595 -108.285 106.925 -107.955 ;
        RECT 106.595 -109.645 106.925 -109.315 ;
        RECT 106.595 -111.005 106.925 -110.675 ;
        RECT 106.595 -112.365 106.925 -112.035 ;
        RECT 106.595 -113.725 106.925 -113.395 ;
        RECT 106.595 -115.085 106.925 -114.755 ;
        RECT 106.595 -116.445 106.925 -116.115 ;
        RECT 106.595 -117.805 106.925 -117.475 ;
        RECT 106.595 -119.165 106.925 -118.835 ;
        RECT 106.595 -120.525 106.925 -120.195 ;
        RECT 106.595 -121.885 106.925 -121.555 ;
        RECT 106.595 -123.245 106.925 -122.915 ;
        RECT 106.595 -124.605 106.925 -124.275 ;
        RECT 106.595 -125.965 106.925 -125.635 ;
        RECT 106.595 -127.325 106.925 -126.995 ;
        RECT 106.595 -128.685 106.925 -128.355 ;
        RECT 106.595 -130.045 106.925 -129.715 ;
        RECT 106.595 -131.405 106.925 -131.075 ;
        RECT 106.595 -132.765 106.925 -132.435 ;
        RECT 106.595 -134.125 106.925 -133.795 ;
        RECT 106.595 -135.485 106.925 -135.155 ;
        RECT 106.595 -136.845 106.925 -136.515 ;
        RECT 106.595 -138.205 106.925 -137.875 ;
        RECT 106.595 -139.565 106.925 -139.235 ;
        RECT 106.595 -140.925 106.925 -140.595 ;
        RECT 106.595 -142.285 106.925 -141.955 ;
        RECT 106.595 -143.645 106.925 -143.315 ;
        RECT 106.595 -145.005 106.925 -144.675 ;
        RECT 106.595 -146.365 106.925 -146.035 ;
        RECT 106.595 -147.725 106.925 -147.395 ;
        RECT 106.595 -149.085 106.925 -148.755 ;
        RECT 106.595 -150.445 106.925 -150.115 ;
        RECT 106.595 -151.805 106.925 -151.475 ;
        RECT 106.595 -153.165 106.925 -152.835 ;
        RECT 106.595 -154.525 106.925 -154.195 ;
        RECT 106.595 -155.885 106.925 -155.555 ;
        RECT 106.595 -157.245 106.925 -156.915 ;
        RECT 106.595 -162.89 106.925 -161.76 ;
        RECT 106.6 -163.005 106.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 129.945 108.285 131.075 ;
        RECT 107.955 125.635 108.285 125.965 ;
        RECT 107.955 124.275 108.285 124.605 ;
        RECT 107.96 123.6 108.28 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 -0.845 108.285 -0.515 ;
        RECT 107.955 -2.205 108.285 -1.875 ;
        RECT 107.955 -3.565 108.285 -3.235 ;
        RECT 107.96 -3.565 108.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 129.945 109.645 131.075 ;
        RECT 109.315 125.635 109.645 125.965 ;
        RECT 109.315 124.275 109.645 124.605 ;
        RECT 109.32 123.6 109.64 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 -0.845 109.645 -0.515 ;
        RECT 109.315 -2.205 109.645 -1.875 ;
        RECT 109.315 -3.565 109.645 -3.235 ;
        RECT 109.32 -3.565 109.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 129.945 111.005 131.075 ;
        RECT 110.675 125.635 111.005 125.965 ;
        RECT 110.675 124.275 111.005 124.605 ;
        RECT 110.68 123.6 111 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -0.845 111.005 -0.515 ;
        RECT 110.675 -2.205 111.005 -1.875 ;
        RECT 110.675 -3.565 111.005 -3.235 ;
        RECT 110.68 -3.565 111 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -91.965 111.005 -91.635 ;
        RECT 110.675 -93.325 111.005 -92.995 ;
        RECT 110.675 -94.685 111.005 -94.355 ;
        RECT 110.675 -96.045 111.005 -95.715 ;
        RECT 110.675 -97.405 111.005 -97.075 ;
        RECT 110.675 -98.765 111.005 -98.435 ;
        RECT 110.675 -100.125 111.005 -99.795 ;
        RECT 110.675 -101.485 111.005 -101.155 ;
        RECT 110.675 -102.845 111.005 -102.515 ;
        RECT 110.675 -104.205 111.005 -103.875 ;
        RECT 110.675 -105.565 111.005 -105.235 ;
        RECT 110.675 -106.925 111.005 -106.595 ;
        RECT 110.675 -108.285 111.005 -107.955 ;
        RECT 110.675 -109.645 111.005 -109.315 ;
        RECT 110.675 -111.005 111.005 -110.675 ;
        RECT 110.675 -112.365 111.005 -112.035 ;
        RECT 110.675 -113.725 111.005 -113.395 ;
        RECT 110.675 -115.085 111.005 -114.755 ;
        RECT 110.675 -116.445 111.005 -116.115 ;
        RECT 110.675 -117.805 111.005 -117.475 ;
        RECT 110.675 -119.165 111.005 -118.835 ;
        RECT 110.675 -120.525 111.005 -120.195 ;
        RECT 110.675 -121.885 111.005 -121.555 ;
        RECT 110.675 -123.245 111.005 -122.915 ;
        RECT 110.675 -124.605 111.005 -124.275 ;
        RECT 110.675 -125.965 111.005 -125.635 ;
        RECT 110.675 -127.325 111.005 -126.995 ;
        RECT 110.675 -128.685 111.005 -128.355 ;
        RECT 110.675 -130.045 111.005 -129.715 ;
        RECT 110.675 -131.405 111.005 -131.075 ;
        RECT 110.675 -132.765 111.005 -132.435 ;
        RECT 110.675 -134.125 111.005 -133.795 ;
        RECT 110.675 -135.485 111.005 -135.155 ;
        RECT 110.675 -136.845 111.005 -136.515 ;
        RECT 110.675 -138.205 111.005 -137.875 ;
        RECT 110.675 -139.565 111.005 -139.235 ;
        RECT 110.675 -140.925 111.005 -140.595 ;
        RECT 110.675 -142.285 111.005 -141.955 ;
        RECT 110.675 -143.645 111.005 -143.315 ;
        RECT 110.675 -145.005 111.005 -144.675 ;
        RECT 110.675 -146.365 111.005 -146.035 ;
        RECT 110.675 -147.725 111.005 -147.395 ;
        RECT 110.675 -149.085 111.005 -148.755 ;
        RECT 110.675 -150.445 111.005 -150.115 ;
        RECT 110.675 -151.805 111.005 -151.475 ;
        RECT 110.675 -153.165 111.005 -152.835 ;
        RECT 110.675 -154.525 111.005 -154.195 ;
        RECT 110.675 -155.885 111.005 -155.555 ;
        RECT 110.675 -157.245 111.005 -156.915 ;
        RECT 110.675 -162.89 111.005 -161.76 ;
        RECT 110.68 -163.005 111 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 129.945 112.365 131.075 ;
        RECT 112.035 125.635 112.365 125.965 ;
        RECT 112.035 124.275 112.365 124.605 ;
        RECT 112.04 123.6 112.36 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 -149.085 112.365 -148.755 ;
        RECT 112.035 -150.445 112.365 -150.115 ;
        RECT 112.035 -151.805 112.365 -151.475 ;
        RECT 112.035 -153.165 112.365 -152.835 ;
        RECT 112.035 -154.525 112.365 -154.195 ;
        RECT 112.035 -155.885 112.365 -155.555 ;
        RECT 112.035 -157.245 112.365 -156.915 ;
        RECT 112.035 -162.89 112.365 -161.76 ;
        RECT 112.04 -163.005 112.36 -95.04 ;
        RECT 112.035 -96.045 112.365 -95.715 ;
        RECT 112.035 -97.405 112.365 -97.075 ;
        RECT 112.035 -98.765 112.365 -98.435 ;
        RECT 112.035 -100.125 112.365 -99.795 ;
        RECT 112.035 -101.485 112.365 -101.155 ;
        RECT 112.035 -102.845 112.365 -102.515 ;
        RECT 112.035 -104.205 112.365 -103.875 ;
        RECT 112.035 -105.565 112.365 -105.235 ;
        RECT 112.035 -106.925 112.365 -106.595 ;
        RECT 112.035 -108.285 112.365 -107.955 ;
        RECT 112.035 -109.645 112.365 -109.315 ;
        RECT 112.035 -111.005 112.365 -110.675 ;
        RECT 112.035 -112.365 112.365 -112.035 ;
        RECT 112.035 -113.725 112.365 -113.395 ;
        RECT 112.035 -115.085 112.365 -114.755 ;
        RECT 112.035 -116.445 112.365 -116.115 ;
        RECT 112.035 -117.805 112.365 -117.475 ;
        RECT 112.035 -119.165 112.365 -118.835 ;
        RECT 112.035 -120.525 112.365 -120.195 ;
        RECT 112.035 -121.885 112.365 -121.555 ;
        RECT 112.035 -123.245 112.365 -122.915 ;
        RECT 112.035 -124.605 112.365 -124.275 ;
        RECT 112.035 -125.965 112.365 -125.635 ;
        RECT 112.035 -127.325 112.365 -126.995 ;
        RECT 112.035 -128.685 112.365 -128.355 ;
        RECT 112.035 -130.045 112.365 -129.715 ;
        RECT 112.035 -131.405 112.365 -131.075 ;
        RECT 112.035 -132.765 112.365 -132.435 ;
        RECT 112.035 -134.125 112.365 -133.795 ;
        RECT 112.035 -135.485 112.365 -135.155 ;
        RECT 112.035 -136.845 112.365 -136.515 ;
        RECT 112.035 -138.205 112.365 -137.875 ;
        RECT 112.035 -139.565 112.365 -139.235 ;
        RECT 112.035 -140.925 112.365 -140.595 ;
        RECT 112.035 -142.285 112.365 -141.955 ;
        RECT 112.035 -143.645 112.365 -143.315 ;
        RECT 112.035 -145.005 112.365 -144.675 ;
        RECT 112.035 -146.365 112.365 -146.035 ;
        RECT 112.035 -147.725 112.365 -147.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 129.945 33.485 131.075 ;
        RECT 33.155 125.635 33.485 125.965 ;
        RECT 33.155 124.275 33.485 124.605 ;
        RECT 33.16 123.6 33.48 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 -96.045 33.485 -95.715 ;
        RECT 33.155 -97.405 33.485 -97.075 ;
        RECT 33.155 -98.765 33.485 -98.435 ;
        RECT 33.155 -100.125 33.485 -99.795 ;
        RECT 33.155 -101.485 33.485 -101.155 ;
        RECT 33.155 -102.845 33.485 -102.515 ;
        RECT 33.155 -104.205 33.485 -103.875 ;
        RECT 33.155 -105.565 33.485 -105.235 ;
        RECT 33.155 -106.925 33.485 -106.595 ;
        RECT 33.155 -108.285 33.485 -107.955 ;
        RECT 33.155 -109.645 33.485 -109.315 ;
        RECT 33.155 -111.005 33.485 -110.675 ;
        RECT 33.155 -112.365 33.485 -112.035 ;
        RECT 33.155 -113.725 33.485 -113.395 ;
        RECT 33.155 -115.085 33.485 -114.755 ;
        RECT 33.155 -116.445 33.485 -116.115 ;
        RECT 33.155 -117.805 33.485 -117.475 ;
        RECT 33.155 -119.165 33.485 -118.835 ;
        RECT 33.155 -120.525 33.485 -120.195 ;
        RECT 33.155 -121.885 33.485 -121.555 ;
        RECT 33.155 -123.245 33.485 -122.915 ;
        RECT 33.155 -124.605 33.485 -124.275 ;
        RECT 33.155 -125.965 33.485 -125.635 ;
        RECT 33.155 -127.325 33.485 -126.995 ;
        RECT 33.155 -128.685 33.485 -128.355 ;
        RECT 33.155 -130.045 33.485 -129.715 ;
        RECT 33.155 -131.405 33.485 -131.075 ;
        RECT 33.155 -132.765 33.485 -132.435 ;
        RECT 33.155 -134.125 33.485 -133.795 ;
        RECT 33.155 -135.485 33.485 -135.155 ;
        RECT 33.155 -136.845 33.485 -136.515 ;
        RECT 33.155 -138.205 33.485 -137.875 ;
        RECT 33.155 -139.565 33.485 -139.235 ;
        RECT 33.155 -140.925 33.485 -140.595 ;
        RECT 33.155 -142.285 33.485 -141.955 ;
        RECT 33.155 -143.645 33.485 -143.315 ;
        RECT 33.155 -145.005 33.485 -144.675 ;
        RECT 33.155 -146.365 33.485 -146.035 ;
        RECT 33.155 -147.725 33.485 -147.395 ;
        RECT 33.155 -149.085 33.485 -148.755 ;
        RECT 33.155 -150.445 33.485 -150.115 ;
        RECT 33.155 -151.805 33.485 -151.475 ;
        RECT 33.155 -153.165 33.485 -152.835 ;
        RECT 33.155 -154.525 33.485 -154.195 ;
        RECT 33.155 -155.885 33.485 -155.555 ;
        RECT 33.155 -157.245 33.485 -156.915 ;
        RECT 33.155 -162.89 33.485 -161.76 ;
        RECT 33.16 -163.005 33.48 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.16 -94.075 33.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 129.945 34.845 131.075 ;
        RECT 34.515 125.635 34.845 125.965 ;
        RECT 34.515 124.275 34.845 124.605 ;
        RECT 34.52 123.6 34.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 -0.845 34.845 -0.515 ;
        RECT 34.515 -2.205 34.845 -1.875 ;
        RECT 34.515 -3.565 34.845 -3.235 ;
        RECT 34.52 -3.565 34.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 129.945 36.205 131.075 ;
        RECT 35.875 125.635 36.205 125.965 ;
        RECT 35.875 124.275 36.205 124.605 ;
        RECT 35.88 123.6 36.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 -0.845 36.205 -0.515 ;
        RECT 35.875 -2.205 36.205 -1.875 ;
        RECT 35.875 -3.565 36.205 -3.235 ;
        RECT 35.88 -3.565 36.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 129.945 37.565 131.075 ;
        RECT 37.235 125.635 37.565 125.965 ;
        RECT 37.235 124.275 37.565 124.605 ;
        RECT 37.24 123.6 37.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 -0.845 37.565 -0.515 ;
        RECT 37.235 -2.205 37.565 -1.875 ;
        RECT 37.235 -3.565 37.565 -3.235 ;
        RECT 37.24 -3.565 37.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 -91.965 37.565 -91.635 ;
        RECT 37.235 -93.325 37.565 -92.995 ;
        RECT 37.235 -94.685 37.565 -94.355 ;
        RECT 37.235 -96.045 37.565 -95.715 ;
        RECT 37.235 -97.405 37.565 -97.075 ;
        RECT 37.235 -98.765 37.565 -98.435 ;
        RECT 37.235 -100.125 37.565 -99.795 ;
        RECT 37.235 -101.485 37.565 -101.155 ;
        RECT 37.235 -102.845 37.565 -102.515 ;
        RECT 37.235 -104.205 37.565 -103.875 ;
        RECT 37.235 -105.565 37.565 -105.235 ;
        RECT 37.235 -106.925 37.565 -106.595 ;
        RECT 37.235 -108.285 37.565 -107.955 ;
        RECT 37.235 -109.645 37.565 -109.315 ;
        RECT 37.235 -111.005 37.565 -110.675 ;
        RECT 37.235 -112.365 37.565 -112.035 ;
        RECT 37.235 -113.725 37.565 -113.395 ;
        RECT 37.235 -115.085 37.565 -114.755 ;
        RECT 37.235 -116.445 37.565 -116.115 ;
        RECT 37.235 -117.805 37.565 -117.475 ;
        RECT 37.235 -119.165 37.565 -118.835 ;
        RECT 37.235 -120.525 37.565 -120.195 ;
        RECT 37.235 -121.885 37.565 -121.555 ;
        RECT 37.235 -123.245 37.565 -122.915 ;
        RECT 37.235 -124.605 37.565 -124.275 ;
        RECT 37.235 -125.965 37.565 -125.635 ;
        RECT 37.235 -127.325 37.565 -126.995 ;
        RECT 37.235 -128.685 37.565 -128.355 ;
        RECT 37.235 -130.045 37.565 -129.715 ;
        RECT 37.235 -131.405 37.565 -131.075 ;
        RECT 37.235 -132.765 37.565 -132.435 ;
        RECT 37.235 -134.125 37.565 -133.795 ;
        RECT 37.235 -135.485 37.565 -135.155 ;
        RECT 37.235 -136.845 37.565 -136.515 ;
        RECT 37.235 -138.205 37.565 -137.875 ;
        RECT 37.235 -139.565 37.565 -139.235 ;
        RECT 37.235 -140.925 37.565 -140.595 ;
        RECT 37.235 -142.285 37.565 -141.955 ;
        RECT 37.235 -143.645 37.565 -143.315 ;
        RECT 37.235 -145.005 37.565 -144.675 ;
        RECT 37.235 -146.365 37.565 -146.035 ;
        RECT 37.235 -147.725 37.565 -147.395 ;
        RECT 37.235 -149.085 37.565 -148.755 ;
        RECT 37.235 -150.445 37.565 -150.115 ;
        RECT 37.235 -151.805 37.565 -151.475 ;
        RECT 37.235 -153.165 37.565 -152.835 ;
        RECT 37.235 -154.525 37.565 -154.195 ;
        RECT 37.235 -155.885 37.565 -155.555 ;
        RECT 37.235 -157.245 37.565 -156.915 ;
        RECT 37.235 -162.89 37.565 -161.76 ;
        RECT 37.24 -163.005 37.56 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 129.945 38.925 131.075 ;
        RECT 38.595 125.635 38.925 125.965 ;
        RECT 38.595 124.275 38.925 124.605 ;
        RECT 38.6 123.6 38.92 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 -96.045 38.925 -95.715 ;
        RECT 38.595 -97.405 38.925 -97.075 ;
        RECT 38.595 -98.765 38.925 -98.435 ;
        RECT 38.595 -100.125 38.925 -99.795 ;
        RECT 38.595 -101.485 38.925 -101.155 ;
        RECT 38.595 -102.845 38.925 -102.515 ;
        RECT 38.595 -104.205 38.925 -103.875 ;
        RECT 38.595 -105.565 38.925 -105.235 ;
        RECT 38.595 -106.925 38.925 -106.595 ;
        RECT 38.595 -108.285 38.925 -107.955 ;
        RECT 38.595 -109.645 38.925 -109.315 ;
        RECT 38.595 -111.005 38.925 -110.675 ;
        RECT 38.595 -112.365 38.925 -112.035 ;
        RECT 38.595 -113.725 38.925 -113.395 ;
        RECT 38.595 -115.085 38.925 -114.755 ;
        RECT 38.595 -116.445 38.925 -116.115 ;
        RECT 38.595 -117.805 38.925 -117.475 ;
        RECT 38.595 -119.165 38.925 -118.835 ;
        RECT 38.595 -120.525 38.925 -120.195 ;
        RECT 38.595 -121.885 38.925 -121.555 ;
        RECT 38.595 -123.245 38.925 -122.915 ;
        RECT 38.595 -124.605 38.925 -124.275 ;
        RECT 38.595 -125.965 38.925 -125.635 ;
        RECT 38.595 -127.325 38.925 -126.995 ;
        RECT 38.595 -128.685 38.925 -128.355 ;
        RECT 38.595 -130.045 38.925 -129.715 ;
        RECT 38.595 -131.405 38.925 -131.075 ;
        RECT 38.595 -132.765 38.925 -132.435 ;
        RECT 38.595 -134.125 38.925 -133.795 ;
        RECT 38.595 -135.485 38.925 -135.155 ;
        RECT 38.595 -136.845 38.925 -136.515 ;
        RECT 38.595 -138.205 38.925 -137.875 ;
        RECT 38.595 -139.565 38.925 -139.235 ;
        RECT 38.595 -140.925 38.925 -140.595 ;
        RECT 38.595 -142.285 38.925 -141.955 ;
        RECT 38.595 -143.645 38.925 -143.315 ;
        RECT 38.595 -145.005 38.925 -144.675 ;
        RECT 38.595 -146.365 38.925 -146.035 ;
        RECT 38.595 -147.725 38.925 -147.395 ;
        RECT 38.595 -149.085 38.925 -148.755 ;
        RECT 38.595 -150.445 38.925 -150.115 ;
        RECT 38.595 -151.805 38.925 -151.475 ;
        RECT 38.595 -153.165 38.925 -152.835 ;
        RECT 38.595 -154.525 38.925 -154.195 ;
        RECT 38.595 -155.885 38.925 -155.555 ;
        RECT 38.595 -157.245 38.925 -156.915 ;
        RECT 38.595 -162.89 38.925 -161.76 ;
        RECT 38.6 -163.005 38.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.26 -94.075 39.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 129.945 40.285 131.075 ;
        RECT 39.955 125.635 40.285 125.965 ;
        RECT 39.955 124.275 40.285 124.605 ;
        RECT 39.96 123.6 40.28 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 129.945 41.645 131.075 ;
        RECT 41.315 125.635 41.645 125.965 ;
        RECT 41.315 124.275 41.645 124.605 ;
        RECT 41.32 123.6 41.64 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 -0.845 41.645 -0.515 ;
        RECT 41.315 -2.205 41.645 -1.875 ;
        RECT 41.315 -3.565 41.645 -3.235 ;
        RECT 41.32 -3.565 41.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 129.945 43.005 131.075 ;
        RECT 42.675 125.635 43.005 125.965 ;
        RECT 42.675 124.275 43.005 124.605 ;
        RECT 42.68 123.6 43 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 -0.845 43.005 -0.515 ;
        RECT 42.675 -2.205 43.005 -1.875 ;
        RECT 42.675 -3.565 43.005 -3.235 ;
        RECT 42.68 -3.565 43 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 129.945 44.365 131.075 ;
        RECT 44.035 125.635 44.365 125.965 ;
        RECT 44.035 124.275 44.365 124.605 ;
        RECT 44.04 123.6 44.36 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -0.845 44.365 -0.515 ;
        RECT 44.035 -2.205 44.365 -1.875 ;
        RECT 44.035 -3.565 44.365 -3.235 ;
        RECT 44.04 -3.565 44.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -91.965 44.365 -91.635 ;
        RECT 44.035 -93.325 44.365 -92.995 ;
        RECT 44.035 -94.685 44.365 -94.355 ;
        RECT 44.035 -96.045 44.365 -95.715 ;
        RECT 44.035 -97.405 44.365 -97.075 ;
        RECT 44.035 -98.765 44.365 -98.435 ;
        RECT 44.035 -100.125 44.365 -99.795 ;
        RECT 44.035 -101.485 44.365 -101.155 ;
        RECT 44.035 -102.845 44.365 -102.515 ;
        RECT 44.035 -104.205 44.365 -103.875 ;
        RECT 44.035 -105.565 44.365 -105.235 ;
        RECT 44.035 -106.925 44.365 -106.595 ;
        RECT 44.035 -108.285 44.365 -107.955 ;
        RECT 44.035 -109.645 44.365 -109.315 ;
        RECT 44.035 -111.005 44.365 -110.675 ;
        RECT 44.035 -112.365 44.365 -112.035 ;
        RECT 44.035 -113.725 44.365 -113.395 ;
        RECT 44.035 -115.085 44.365 -114.755 ;
        RECT 44.035 -116.445 44.365 -116.115 ;
        RECT 44.035 -117.805 44.365 -117.475 ;
        RECT 44.035 -119.165 44.365 -118.835 ;
        RECT 44.035 -120.525 44.365 -120.195 ;
        RECT 44.035 -121.885 44.365 -121.555 ;
        RECT 44.035 -123.245 44.365 -122.915 ;
        RECT 44.035 -124.605 44.365 -124.275 ;
        RECT 44.035 -125.965 44.365 -125.635 ;
        RECT 44.035 -127.325 44.365 -126.995 ;
        RECT 44.035 -128.685 44.365 -128.355 ;
        RECT 44.035 -130.045 44.365 -129.715 ;
        RECT 44.035 -131.405 44.365 -131.075 ;
        RECT 44.035 -132.765 44.365 -132.435 ;
        RECT 44.035 -134.125 44.365 -133.795 ;
        RECT 44.035 -135.485 44.365 -135.155 ;
        RECT 44.035 -136.845 44.365 -136.515 ;
        RECT 44.035 -138.205 44.365 -137.875 ;
        RECT 44.035 -139.565 44.365 -139.235 ;
        RECT 44.035 -140.925 44.365 -140.595 ;
        RECT 44.035 -142.285 44.365 -141.955 ;
        RECT 44.035 -143.645 44.365 -143.315 ;
        RECT 44.035 -145.005 44.365 -144.675 ;
        RECT 44.035 -146.365 44.365 -146.035 ;
        RECT 44.035 -147.725 44.365 -147.395 ;
        RECT 44.035 -149.085 44.365 -148.755 ;
        RECT 44.035 -150.445 44.365 -150.115 ;
        RECT 44.035 -151.805 44.365 -151.475 ;
        RECT 44.035 -153.165 44.365 -152.835 ;
        RECT 44.035 -154.525 44.365 -154.195 ;
        RECT 44.035 -155.885 44.365 -155.555 ;
        RECT 44.035 -157.245 44.365 -156.915 ;
        RECT 44.035 -162.89 44.365 -161.76 ;
        RECT 44.04 -163.005 44.36 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.36 -94.075 45.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 129.945 45.725 131.075 ;
        RECT 45.395 125.635 45.725 125.965 ;
        RECT 45.395 124.275 45.725 124.605 ;
        RECT 45.4 123.6 45.72 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 -96.045 45.725 -95.715 ;
        RECT 45.395 -97.405 45.725 -97.075 ;
        RECT 45.395 -98.765 45.725 -98.435 ;
        RECT 45.395 -100.125 45.725 -99.795 ;
        RECT 45.395 -101.485 45.725 -101.155 ;
        RECT 45.395 -102.845 45.725 -102.515 ;
        RECT 45.395 -104.205 45.725 -103.875 ;
        RECT 45.395 -105.565 45.725 -105.235 ;
        RECT 45.395 -106.925 45.725 -106.595 ;
        RECT 45.395 -108.285 45.725 -107.955 ;
        RECT 45.395 -109.645 45.725 -109.315 ;
        RECT 45.395 -111.005 45.725 -110.675 ;
        RECT 45.395 -112.365 45.725 -112.035 ;
        RECT 45.395 -113.725 45.725 -113.395 ;
        RECT 45.395 -115.085 45.725 -114.755 ;
        RECT 45.395 -116.445 45.725 -116.115 ;
        RECT 45.395 -117.805 45.725 -117.475 ;
        RECT 45.395 -119.165 45.725 -118.835 ;
        RECT 45.395 -120.525 45.725 -120.195 ;
        RECT 45.395 -121.885 45.725 -121.555 ;
        RECT 45.395 -123.245 45.725 -122.915 ;
        RECT 45.395 -124.605 45.725 -124.275 ;
        RECT 45.395 -125.965 45.725 -125.635 ;
        RECT 45.395 -127.325 45.725 -126.995 ;
        RECT 45.395 -128.685 45.725 -128.355 ;
        RECT 45.395 -130.045 45.725 -129.715 ;
        RECT 45.395 -131.405 45.725 -131.075 ;
        RECT 45.395 -132.765 45.725 -132.435 ;
        RECT 45.395 -134.125 45.725 -133.795 ;
        RECT 45.395 -135.485 45.725 -135.155 ;
        RECT 45.395 -136.845 45.725 -136.515 ;
        RECT 45.395 -138.205 45.725 -137.875 ;
        RECT 45.395 -139.565 45.725 -139.235 ;
        RECT 45.395 -140.925 45.725 -140.595 ;
        RECT 45.395 -142.285 45.725 -141.955 ;
        RECT 45.395 -143.645 45.725 -143.315 ;
        RECT 45.395 -145.005 45.725 -144.675 ;
        RECT 45.395 -146.365 45.725 -146.035 ;
        RECT 45.395 -147.725 45.725 -147.395 ;
        RECT 45.395 -149.085 45.725 -148.755 ;
        RECT 45.395 -150.445 45.725 -150.115 ;
        RECT 45.395 -151.805 45.725 -151.475 ;
        RECT 45.395 -153.165 45.725 -152.835 ;
        RECT 45.395 -154.525 45.725 -154.195 ;
        RECT 45.395 -155.885 45.725 -155.555 ;
        RECT 45.395 -157.245 45.725 -156.915 ;
        RECT 45.395 -162.89 45.725 -161.76 ;
        RECT 45.4 -163.005 45.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 129.945 47.085 131.075 ;
        RECT 46.755 125.635 47.085 125.965 ;
        RECT 46.755 124.275 47.085 124.605 ;
        RECT 46.76 123.6 47.08 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 -0.845 47.085 -0.515 ;
        RECT 46.755 -2.205 47.085 -1.875 ;
        RECT 46.755 -3.565 47.085 -3.235 ;
        RECT 46.76 -3.565 47.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 129.945 48.445 131.075 ;
        RECT 48.115 125.635 48.445 125.965 ;
        RECT 48.115 124.275 48.445 124.605 ;
        RECT 48.12 123.6 48.44 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 -0.845 48.445 -0.515 ;
        RECT 48.115 -2.205 48.445 -1.875 ;
        RECT 48.115 -3.565 48.445 -3.235 ;
        RECT 48.12 -3.565 48.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 129.945 49.805 131.075 ;
        RECT 49.475 125.635 49.805 125.965 ;
        RECT 49.475 124.275 49.805 124.605 ;
        RECT 49.48 123.6 49.8 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 -0.845 49.805 -0.515 ;
        RECT 49.475 -2.205 49.805 -1.875 ;
        RECT 49.475 -3.565 49.805 -3.235 ;
        RECT 49.48 -3.565 49.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 -91.965 49.805 -91.635 ;
        RECT 49.475 -93.325 49.805 -92.995 ;
        RECT 49.475 -94.685 49.805 -94.355 ;
        RECT 49.475 -96.045 49.805 -95.715 ;
        RECT 49.475 -97.405 49.805 -97.075 ;
        RECT 49.475 -98.765 49.805 -98.435 ;
        RECT 49.475 -100.125 49.805 -99.795 ;
        RECT 49.475 -101.485 49.805 -101.155 ;
        RECT 49.475 -102.845 49.805 -102.515 ;
        RECT 49.475 -104.205 49.805 -103.875 ;
        RECT 49.475 -105.565 49.805 -105.235 ;
        RECT 49.475 -106.925 49.805 -106.595 ;
        RECT 49.475 -108.285 49.805 -107.955 ;
        RECT 49.475 -109.645 49.805 -109.315 ;
        RECT 49.475 -111.005 49.805 -110.675 ;
        RECT 49.475 -112.365 49.805 -112.035 ;
        RECT 49.475 -113.725 49.805 -113.395 ;
        RECT 49.475 -115.085 49.805 -114.755 ;
        RECT 49.475 -116.445 49.805 -116.115 ;
        RECT 49.475 -117.805 49.805 -117.475 ;
        RECT 49.475 -119.165 49.805 -118.835 ;
        RECT 49.475 -120.525 49.805 -120.195 ;
        RECT 49.475 -121.885 49.805 -121.555 ;
        RECT 49.475 -123.245 49.805 -122.915 ;
        RECT 49.475 -124.605 49.805 -124.275 ;
        RECT 49.475 -125.965 49.805 -125.635 ;
        RECT 49.475 -127.325 49.805 -126.995 ;
        RECT 49.475 -128.685 49.805 -128.355 ;
        RECT 49.475 -130.045 49.805 -129.715 ;
        RECT 49.475 -131.405 49.805 -131.075 ;
        RECT 49.475 -132.765 49.805 -132.435 ;
        RECT 49.475 -134.125 49.805 -133.795 ;
        RECT 49.475 -135.485 49.805 -135.155 ;
        RECT 49.475 -136.845 49.805 -136.515 ;
        RECT 49.475 -138.205 49.805 -137.875 ;
        RECT 49.475 -139.565 49.805 -139.235 ;
        RECT 49.475 -140.925 49.805 -140.595 ;
        RECT 49.475 -142.285 49.805 -141.955 ;
        RECT 49.475 -143.645 49.805 -143.315 ;
        RECT 49.475 -145.005 49.805 -144.675 ;
        RECT 49.475 -146.365 49.805 -146.035 ;
        RECT 49.475 -147.725 49.805 -147.395 ;
        RECT 49.475 -149.085 49.805 -148.755 ;
        RECT 49.475 -150.445 49.805 -150.115 ;
        RECT 49.475 -151.805 49.805 -151.475 ;
        RECT 49.475 -153.165 49.805 -152.835 ;
        RECT 49.475 -154.525 49.805 -154.195 ;
        RECT 49.475 -155.885 49.805 -155.555 ;
        RECT 49.475 -157.245 49.805 -156.915 ;
        RECT 49.475 -162.89 49.805 -161.76 ;
        RECT 49.48 -163.005 49.8 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 129.945 51.165 131.075 ;
        RECT 50.835 125.635 51.165 125.965 ;
        RECT 50.835 124.275 51.165 124.605 ;
        RECT 50.84 123.6 51.16 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 -96.045 51.165 -95.715 ;
        RECT 50.835 -97.405 51.165 -97.075 ;
        RECT 50.835 -98.765 51.165 -98.435 ;
        RECT 50.835 -100.125 51.165 -99.795 ;
        RECT 50.835 -101.485 51.165 -101.155 ;
        RECT 50.835 -102.845 51.165 -102.515 ;
        RECT 50.835 -104.205 51.165 -103.875 ;
        RECT 50.835 -105.565 51.165 -105.235 ;
        RECT 50.835 -106.925 51.165 -106.595 ;
        RECT 50.835 -108.285 51.165 -107.955 ;
        RECT 50.835 -109.645 51.165 -109.315 ;
        RECT 50.835 -111.005 51.165 -110.675 ;
        RECT 50.835 -112.365 51.165 -112.035 ;
        RECT 50.835 -113.725 51.165 -113.395 ;
        RECT 50.835 -115.085 51.165 -114.755 ;
        RECT 50.835 -116.445 51.165 -116.115 ;
        RECT 50.835 -117.805 51.165 -117.475 ;
        RECT 50.835 -119.165 51.165 -118.835 ;
        RECT 50.835 -120.525 51.165 -120.195 ;
        RECT 50.835 -121.885 51.165 -121.555 ;
        RECT 50.835 -123.245 51.165 -122.915 ;
        RECT 50.835 -124.605 51.165 -124.275 ;
        RECT 50.835 -125.965 51.165 -125.635 ;
        RECT 50.835 -127.325 51.165 -126.995 ;
        RECT 50.835 -128.685 51.165 -128.355 ;
        RECT 50.835 -130.045 51.165 -129.715 ;
        RECT 50.835 -131.405 51.165 -131.075 ;
        RECT 50.835 -132.765 51.165 -132.435 ;
        RECT 50.835 -134.125 51.165 -133.795 ;
        RECT 50.835 -135.485 51.165 -135.155 ;
        RECT 50.835 -136.845 51.165 -136.515 ;
        RECT 50.835 -138.205 51.165 -137.875 ;
        RECT 50.835 -139.565 51.165 -139.235 ;
        RECT 50.835 -140.925 51.165 -140.595 ;
        RECT 50.835 -142.285 51.165 -141.955 ;
        RECT 50.835 -143.645 51.165 -143.315 ;
        RECT 50.835 -145.005 51.165 -144.675 ;
        RECT 50.835 -146.365 51.165 -146.035 ;
        RECT 50.835 -147.725 51.165 -147.395 ;
        RECT 50.835 -149.085 51.165 -148.755 ;
        RECT 50.835 -150.445 51.165 -150.115 ;
        RECT 50.835 -151.805 51.165 -151.475 ;
        RECT 50.835 -153.165 51.165 -152.835 ;
        RECT 50.835 -154.525 51.165 -154.195 ;
        RECT 50.835 -155.885 51.165 -155.555 ;
        RECT 50.835 -157.245 51.165 -156.915 ;
        RECT 50.835 -162.89 51.165 -161.76 ;
        RECT 50.84 -163.005 51.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.46 -94.075 51.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 129.945 52.525 131.075 ;
        RECT 52.195 125.635 52.525 125.965 ;
        RECT 52.195 124.275 52.525 124.605 ;
        RECT 52.2 123.6 52.52 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 129.945 53.885 131.075 ;
        RECT 53.555 125.635 53.885 125.965 ;
        RECT 53.555 124.275 53.885 124.605 ;
        RECT 53.56 123.6 53.88 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -0.845 53.885 -0.515 ;
        RECT 53.555 -2.205 53.885 -1.875 ;
        RECT 53.555 -3.565 53.885 -3.235 ;
        RECT 53.56 -3.565 53.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -91.965 53.885 -91.635 ;
        RECT 53.555 -93.325 53.885 -92.995 ;
        RECT 53.555 -94.685 53.885 -94.355 ;
        RECT 53.555 -96.045 53.885 -95.715 ;
        RECT 53.555 -97.405 53.885 -97.075 ;
        RECT 53.555 -98.765 53.885 -98.435 ;
        RECT 53.555 -100.125 53.885 -99.795 ;
        RECT 53.555 -101.485 53.885 -101.155 ;
        RECT 53.555 -102.845 53.885 -102.515 ;
        RECT 53.555 -104.205 53.885 -103.875 ;
        RECT 53.555 -105.565 53.885 -105.235 ;
        RECT 53.555 -106.925 53.885 -106.595 ;
        RECT 53.555 -108.285 53.885 -107.955 ;
        RECT 53.555 -109.645 53.885 -109.315 ;
        RECT 53.555 -111.005 53.885 -110.675 ;
        RECT 53.555 -112.365 53.885 -112.035 ;
        RECT 53.555 -113.725 53.885 -113.395 ;
        RECT 53.555 -115.085 53.885 -114.755 ;
        RECT 53.555 -116.445 53.885 -116.115 ;
        RECT 53.555 -117.805 53.885 -117.475 ;
        RECT 53.555 -119.165 53.885 -118.835 ;
        RECT 53.555 -120.525 53.885 -120.195 ;
        RECT 53.555 -121.885 53.885 -121.555 ;
        RECT 53.555 -123.245 53.885 -122.915 ;
        RECT 53.555 -124.605 53.885 -124.275 ;
        RECT 53.555 -125.965 53.885 -125.635 ;
        RECT 53.555 -127.325 53.885 -126.995 ;
        RECT 53.555 -128.685 53.885 -128.355 ;
        RECT 53.555 -130.045 53.885 -129.715 ;
        RECT 53.555 -131.405 53.885 -131.075 ;
        RECT 53.555 -132.765 53.885 -132.435 ;
        RECT 53.555 -134.125 53.885 -133.795 ;
        RECT 53.555 -135.485 53.885 -135.155 ;
        RECT 53.555 -136.845 53.885 -136.515 ;
        RECT 53.555 -138.205 53.885 -137.875 ;
        RECT 53.555 -139.565 53.885 -139.235 ;
        RECT 53.555 -140.925 53.885 -140.595 ;
        RECT 53.555 -142.285 53.885 -141.955 ;
        RECT 53.555 -143.645 53.885 -143.315 ;
        RECT 53.555 -145.005 53.885 -144.675 ;
        RECT 53.555 -146.365 53.885 -146.035 ;
        RECT 53.555 -147.725 53.885 -147.395 ;
        RECT 53.555 -149.085 53.885 -148.755 ;
        RECT 53.555 -150.445 53.885 -150.115 ;
        RECT 53.555 -151.805 53.885 -151.475 ;
        RECT 53.555 -153.165 53.885 -152.835 ;
        RECT 53.555 -154.525 53.885 -154.195 ;
        RECT 53.555 -155.885 53.885 -155.555 ;
        RECT 53.555 -157.245 53.885 -156.915 ;
        RECT 53.555 -162.89 53.885 -161.76 ;
        RECT 53.56 -163.005 53.88 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 129.945 55.245 131.075 ;
        RECT 54.915 125.635 55.245 125.965 ;
        RECT 54.915 124.275 55.245 124.605 ;
        RECT 54.92 123.6 55.24 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 -0.845 55.245 -0.515 ;
        RECT 54.915 -2.205 55.245 -1.875 ;
        RECT 54.915 -3.565 55.245 -3.235 ;
        RECT 54.92 -3.565 55.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 129.945 56.605 131.075 ;
        RECT 56.275 125.635 56.605 125.965 ;
        RECT 56.275 124.275 56.605 124.605 ;
        RECT 56.28 123.6 56.6 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -0.845 56.605 -0.515 ;
        RECT 56.275 -2.205 56.605 -1.875 ;
        RECT 56.275 -3.565 56.605 -3.235 ;
        RECT 56.28 -3.565 56.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -91.965 56.605 -91.635 ;
        RECT 56.275 -93.325 56.605 -92.995 ;
        RECT 56.275 -94.685 56.605 -94.355 ;
        RECT 56.275 -96.045 56.605 -95.715 ;
        RECT 56.275 -97.405 56.605 -97.075 ;
        RECT 56.275 -98.765 56.605 -98.435 ;
        RECT 56.275 -100.125 56.605 -99.795 ;
        RECT 56.275 -101.485 56.605 -101.155 ;
        RECT 56.275 -102.845 56.605 -102.515 ;
        RECT 56.275 -104.205 56.605 -103.875 ;
        RECT 56.275 -105.565 56.605 -105.235 ;
        RECT 56.275 -106.925 56.605 -106.595 ;
        RECT 56.275 -108.285 56.605 -107.955 ;
        RECT 56.275 -109.645 56.605 -109.315 ;
        RECT 56.275 -111.005 56.605 -110.675 ;
        RECT 56.275 -112.365 56.605 -112.035 ;
        RECT 56.275 -113.725 56.605 -113.395 ;
        RECT 56.275 -115.085 56.605 -114.755 ;
        RECT 56.275 -116.445 56.605 -116.115 ;
        RECT 56.275 -117.805 56.605 -117.475 ;
        RECT 56.275 -119.165 56.605 -118.835 ;
        RECT 56.275 -120.525 56.605 -120.195 ;
        RECT 56.275 -121.885 56.605 -121.555 ;
        RECT 56.275 -123.245 56.605 -122.915 ;
        RECT 56.275 -124.605 56.605 -124.275 ;
        RECT 56.275 -125.965 56.605 -125.635 ;
        RECT 56.275 -127.325 56.605 -126.995 ;
        RECT 56.275 -128.685 56.605 -128.355 ;
        RECT 56.275 -130.045 56.605 -129.715 ;
        RECT 56.275 -131.405 56.605 -131.075 ;
        RECT 56.275 -132.765 56.605 -132.435 ;
        RECT 56.275 -134.125 56.605 -133.795 ;
        RECT 56.275 -135.485 56.605 -135.155 ;
        RECT 56.275 -136.845 56.605 -136.515 ;
        RECT 56.275 -138.205 56.605 -137.875 ;
        RECT 56.275 -139.565 56.605 -139.235 ;
        RECT 56.275 -140.925 56.605 -140.595 ;
        RECT 56.275 -142.285 56.605 -141.955 ;
        RECT 56.275 -143.645 56.605 -143.315 ;
        RECT 56.275 -145.005 56.605 -144.675 ;
        RECT 56.275 -146.365 56.605 -146.035 ;
        RECT 56.275 -147.725 56.605 -147.395 ;
        RECT 56.275 -149.085 56.605 -148.755 ;
        RECT 56.275 -150.445 56.605 -150.115 ;
        RECT 56.275 -151.805 56.605 -151.475 ;
        RECT 56.275 -153.165 56.605 -152.835 ;
        RECT 56.275 -154.525 56.605 -154.195 ;
        RECT 56.275 -155.885 56.605 -155.555 ;
        RECT 56.275 -157.245 56.605 -156.915 ;
        RECT 56.275 -162.89 56.605 -161.76 ;
        RECT 56.28 -163.005 56.6 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.56 -94.075 57.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 129.945 57.965 131.075 ;
        RECT 57.635 125.635 57.965 125.965 ;
        RECT 57.635 124.275 57.965 124.605 ;
        RECT 57.64 123.6 57.96 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 -96.045 57.965 -95.715 ;
        RECT 57.635 -97.405 57.965 -97.075 ;
        RECT 57.635 -98.765 57.965 -98.435 ;
        RECT 57.635 -100.125 57.965 -99.795 ;
        RECT 57.635 -101.485 57.965 -101.155 ;
        RECT 57.635 -102.845 57.965 -102.515 ;
        RECT 57.635 -104.205 57.965 -103.875 ;
        RECT 57.635 -105.565 57.965 -105.235 ;
        RECT 57.635 -106.925 57.965 -106.595 ;
        RECT 57.635 -108.285 57.965 -107.955 ;
        RECT 57.635 -109.645 57.965 -109.315 ;
        RECT 57.635 -111.005 57.965 -110.675 ;
        RECT 57.635 -112.365 57.965 -112.035 ;
        RECT 57.635 -113.725 57.965 -113.395 ;
        RECT 57.635 -115.085 57.965 -114.755 ;
        RECT 57.635 -116.445 57.965 -116.115 ;
        RECT 57.635 -117.805 57.965 -117.475 ;
        RECT 57.635 -119.165 57.965 -118.835 ;
        RECT 57.635 -120.525 57.965 -120.195 ;
        RECT 57.635 -121.885 57.965 -121.555 ;
        RECT 57.635 -123.245 57.965 -122.915 ;
        RECT 57.635 -124.605 57.965 -124.275 ;
        RECT 57.635 -125.965 57.965 -125.635 ;
        RECT 57.635 -127.325 57.965 -126.995 ;
        RECT 57.635 -128.685 57.965 -128.355 ;
        RECT 57.635 -130.045 57.965 -129.715 ;
        RECT 57.635 -131.405 57.965 -131.075 ;
        RECT 57.635 -132.765 57.965 -132.435 ;
        RECT 57.635 -134.125 57.965 -133.795 ;
        RECT 57.635 -135.485 57.965 -135.155 ;
        RECT 57.635 -136.845 57.965 -136.515 ;
        RECT 57.635 -138.205 57.965 -137.875 ;
        RECT 57.635 -139.565 57.965 -139.235 ;
        RECT 57.635 -140.925 57.965 -140.595 ;
        RECT 57.635 -142.285 57.965 -141.955 ;
        RECT 57.635 -143.645 57.965 -143.315 ;
        RECT 57.635 -145.005 57.965 -144.675 ;
        RECT 57.635 -146.365 57.965 -146.035 ;
        RECT 57.635 -147.725 57.965 -147.395 ;
        RECT 57.635 -149.085 57.965 -148.755 ;
        RECT 57.635 -150.445 57.965 -150.115 ;
        RECT 57.635 -151.805 57.965 -151.475 ;
        RECT 57.635 -153.165 57.965 -152.835 ;
        RECT 57.635 -154.525 57.965 -154.195 ;
        RECT 57.635 -155.885 57.965 -155.555 ;
        RECT 57.635 -157.245 57.965 -156.915 ;
        RECT 57.635 -162.89 57.965 -161.76 ;
        RECT 57.64 -163.005 57.96 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 129.945 59.325 131.075 ;
        RECT 58.995 125.635 59.325 125.965 ;
        RECT 58.995 124.275 59.325 124.605 ;
        RECT 59 123.6 59.32 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 -0.845 59.325 -0.515 ;
        RECT 58.995 -2.205 59.325 -1.875 ;
        RECT 58.995 -3.565 59.325 -3.235 ;
        RECT 59 -3.565 59.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 129.945 60.685 131.075 ;
        RECT 60.355 125.635 60.685 125.965 ;
        RECT 60.355 124.275 60.685 124.605 ;
        RECT 60.36 123.6 60.68 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 -0.845 60.685 -0.515 ;
        RECT 60.355 -2.205 60.685 -1.875 ;
        RECT 60.355 -3.565 60.685 -3.235 ;
        RECT 60.36 -3.565 60.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 129.945 62.045 131.075 ;
        RECT 61.715 125.635 62.045 125.965 ;
        RECT 61.715 124.275 62.045 124.605 ;
        RECT 61.72 123.6 62.04 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -0.845 62.045 -0.515 ;
        RECT 61.715 -2.205 62.045 -1.875 ;
        RECT 61.715 -3.565 62.045 -3.235 ;
        RECT 61.72 -3.565 62.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -91.965 62.045 -91.635 ;
        RECT 61.715 -93.325 62.045 -92.995 ;
        RECT 61.715 -94.685 62.045 -94.355 ;
        RECT 61.715 -96.045 62.045 -95.715 ;
        RECT 61.715 -97.405 62.045 -97.075 ;
        RECT 61.715 -98.765 62.045 -98.435 ;
        RECT 61.715 -100.125 62.045 -99.795 ;
        RECT 61.715 -101.485 62.045 -101.155 ;
        RECT 61.715 -102.845 62.045 -102.515 ;
        RECT 61.715 -104.205 62.045 -103.875 ;
        RECT 61.715 -105.565 62.045 -105.235 ;
        RECT 61.715 -106.925 62.045 -106.595 ;
        RECT 61.715 -108.285 62.045 -107.955 ;
        RECT 61.715 -109.645 62.045 -109.315 ;
        RECT 61.715 -111.005 62.045 -110.675 ;
        RECT 61.715 -112.365 62.045 -112.035 ;
        RECT 61.715 -113.725 62.045 -113.395 ;
        RECT 61.715 -115.085 62.045 -114.755 ;
        RECT 61.715 -116.445 62.045 -116.115 ;
        RECT 61.715 -117.805 62.045 -117.475 ;
        RECT 61.715 -119.165 62.045 -118.835 ;
        RECT 61.715 -120.525 62.045 -120.195 ;
        RECT 61.715 -121.885 62.045 -121.555 ;
        RECT 61.715 -123.245 62.045 -122.915 ;
        RECT 61.715 -124.605 62.045 -124.275 ;
        RECT 61.715 -125.965 62.045 -125.635 ;
        RECT 61.715 -127.325 62.045 -126.995 ;
        RECT 61.715 -128.685 62.045 -128.355 ;
        RECT 61.715 -130.045 62.045 -129.715 ;
        RECT 61.715 -131.405 62.045 -131.075 ;
        RECT 61.715 -132.765 62.045 -132.435 ;
        RECT 61.715 -134.125 62.045 -133.795 ;
        RECT 61.715 -135.485 62.045 -135.155 ;
        RECT 61.715 -136.845 62.045 -136.515 ;
        RECT 61.715 -138.205 62.045 -137.875 ;
        RECT 61.715 -139.565 62.045 -139.235 ;
        RECT 61.715 -140.925 62.045 -140.595 ;
        RECT 61.715 -142.285 62.045 -141.955 ;
        RECT 61.715 -143.645 62.045 -143.315 ;
        RECT 61.715 -145.005 62.045 -144.675 ;
        RECT 61.715 -146.365 62.045 -146.035 ;
        RECT 61.715 -147.725 62.045 -147.395 ;
        RECT 61.715 -149.085 62.045 -148.755 ;
        RECT 61.715 -150.445 62.045 -150.115 ;
        RECT 61.715 -151.805 62.045 -151.475 ;
        RECT 61.715 -153.165 62.045 -152.835 ;
        RECT 61.715 -154.525 62.045 -154.195 ;
        RECT 61.715 -155.885 62.045 -155.555 ;
        RECT 61.715 -157.245 62.045 -156.915 ;
        RECT 61.715 -162.89 62.045 -161.76 ;
        RECT 61.72 -163.005 62.04 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 129.945 63.405 131.075 ;
        RECT 63.075 125.635 63.405 125.965 ;
        RECT 63.075 124.275 63.405 124.605 ;
        RECT 63.08 123.6 63.4 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 -96.045 63.405 -95.715 ;
        RECT 63.075 -97.405 63.405 -97.075 ;
        RECT 63.075 -98.765 63.405 -98.435 ;
        RECT 63.075 -100.125 63.405 -99.795 ;
        RECT 63.075 -101.485 63.405 -101.155 ;
        RECT 63.075 -102.845 63.405 -102.515 ;
        RECT 63.075 -104.205 63.405 -103.875 ;
        RECT 63.075 -105.565 63.405 -105.235 ;
        RECT 63.075 -106.925 63.405 -106.595 ;
        RECT 63.075 -108.285 63.405 -107.955 ;
        RECT 63.075 -109.645 63.405 -109.315 ;
        RECT 63.075 -111.005 63.405 -110.675 ;
        RECT 63.075 -112.365 63.405 -112.035 ;
        RECT 63.075 -113.725 63.405 -113.395 ;
        RECT 63.075 -115.085 63.405 -114.755 ;
        RECT 63.075 -116.445 63.405 -116.115 ;
        RECT 63.075 -117.805 63.405 -117.475 ;
        RECT 63.075 -119.165 63.405 -118.835 ;
        RECT 63.075 -120.525 63.405 -120.195 ;
        RECT 63.075 -121.885 63.405 -121.555 ;
        RECT 63.075 -123.245 63.405 -122.915 ;
        RECT 63.075 -124.605 63.405 -124.275 ;
        RECT 63.075 -125.965 63.405 -125.635 ;
        RECT 63.075 -127.325 63.405 -126.995 ;
        RECT 63.075 -128.685 63.405 -128.355 ;
        RECT 63.075 -130.045 63.405 -129.715 ;
        RECT 63.075 -131.405 63.405 -131.075 ;
        RECT 63.075 -132.765 63.405 -132.435 ;
        RECT 63.075 -134.125 63.405 -133.795 ;
        RECT 63.075 -135.485 63.405 -135.155 ;
        RECT 63.075 -136.845 63.405 -136.515 ;
        RECT 63.075 -138.205 63.405 -137.875 ;
        RECT 63.075 -139.565 63.405 -139.235 ;
        RECT 63.075 -140.925 63.405 -140.595 ;
        RECT 63.075 -142.285 63.405 -141.955 ;
        RECT 63.075 -143.645 63.405 -143.315 ;
        RECT 63.075 -145.005 63.405 -144.675 ;
        RECT 63.075 -146.365 63.405 -146.035 ;
        RECT 63.075 -147.725 63.405 -147.395 ;
        RECT 63.075 -149.085 63.405 -148.755 ;
        RECT 63.075 -150.445 63.405 -150.115 ;
        RECT 63.075 -151.805 63.405 -151.475 ;
        RECT 63.075 -153.165 63.405 -152.835 ;
        RECT 63.075 -154.525 63.405 -154.195 ;
        RECT 63.075 -155.885 63.405 -155.555 ;
        RECT 63.075 -157.245 63.405 -156.915 ;
        RECT 63.075 -162.89 63.405 -161.76 ;
        RECT 63.08 -163.005 63.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.66 -94.075 63.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 129.945 64.765 131.075 ;
        RECT 64.435 125.635 64.765 125.965 ;
        RECT 64.435 124.275 64.765 124.605 ;
        RECT 64.44 123.6 64.76 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 129.945 66.125 131.075 ;
        RECT 65.795 125.635 66.125 125.965 ;
        RECT 65.795 124.275 66.125 124.605 ;
        RECT 65.8 123.6 66.12 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -0.845 66.125 -0.515 ;
        RECT 65.795 -2.205 66.125 -1.875 ;
        RECT 65.795 -3.565 66.125 -3.235 ;
        RECT 65.8 -3.565 66.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -91.965 66.125 -91.635 ;
        RECT 65.795 -93.325 66.125 -92.995 ;
        RECT 65.795 -94.685 66.125 -94.355 ;
        RECT 65.795 -96.045 66.125 -95.715 ;
        RECT 65.795 -97.405 66.125 -97.075 ;
        RECT 65.795 -98.765 66.125 -98.435 ;
        RECT 65.795 -100.125 66.125 -99.795 ;
        RECT 65.795 -101.485 66.125 -101.155 ;
        RECT 65.795 -102.845 66.125 -102.515 ;
        RECT 65.795 -104.205 66.125 -103.875 ;
        RECT 65.795 -105.565 66.125 -105.235 ;
        RECT 65.795 -106.925 66.125 -106.595 ;
        RECT 65.795 -108.285 66.125 -107.955 ;
        RECT 65.795 -109.645 66.125 -109.315 ;
        RECT 65.795 -111.005 66.125 -110.675 ;
        RECT 65.795 -112.365 66.125 -112.035 ;
        RECT 65.795 -113.725 66.125 -113.395 ;
        RECT 65.795 -115.085 66.125 -114.755 ;
        RECT 65.795 -116.445 66.125 -116.115 ;
        RECT 65.795 -117.805 66.125 -117.475 ;
        RECT 65.795 -119.165 66.125 -118.835 ;
        RECT 65.795 -120.525 66.125 -120.195 ;
        RECT 65.795 -121.885 66.125 -121.555 ;
        RECT 65.795 -123.245 66.125 -122.915 ;
        RECT 65.795 -124.605 66.125 -124.275 ;
        RECT 65.795 -125.965 66.125 -125.635 ;
        RECT 65.795 -127.325 66.125 -126.995 ;
        RECT 65.795 -128.685 66.125 -128.355 ;
        RECT 65.795 -130.045 66.125 -129.715 ;
        RECT 65.795 -131.405 66.125 -131.075 ;
        RECT 65.795 -132.765 66.125 -132.435 ;
        RECT 65.795 -134.125 66.125 -133.795 ;
        RECT 65.795 -135.485 66.125 -135.155 ;
        RECT 65.795 -136.845 66.125 -136.515 ;
        RECT 65.795 -138.205 66.125 -137.875 ;
        RECT 65.795 -139.565 66.125 -139.235 ;
        RECT 65.795 -140.925 66.125 -140.595 ;
        RECT 65.795 -142.285 66.125 -141.955 ;
        RECT 65.795 -143.645 66.125 -143.315 ;
        RECT 65.795 -145.005 66.125 -144.675 ;
        RECT 65.795 -146.365 66.125 -146.035 ;
        RECT 65.795 -147.725 66.125 -147.395 ;
        RECT 65.795 -149.085 66.125 -148.755 ;
        RECT 65.795 -150.445 66.125 -150.115 ;
        RECT 65.795 -151.805 66.125 -151.475 ;
        RECT 65.795 -153.165 66.125 -152.835 ;
        RECT 65.795 -154.525 66.125 -154.195 ;
        RECT 65.795 -155.885 66.125 -155.555 ;
        RECT 65.795 -157.245 66.125 -156.915 ;
        RECT 65.795 -162.89 66.125 -161.76 ;
        RECT 65.8 -163.005 66.12 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 129.945 67.485 131.075 ;
        RECT 67.155 125.635 67.485 125.965 ;
        RECT 67.155 124.275 67.485 124.605 ;
        RECT 67.16 123.6 67.48 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 -0.845 67.485 -0.515 ;
        RECT 67.155 -2.205 67.485 -1.875 ;
        RECT 67.155 -3.565 67.485 -3.235 ;
        RECT 67.16 -3.565 67.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 129.945 68.845 131.075 ;
        RECT 68.515 125.635 68.845 125.965 ;
        RECT 68.515 124.275 68.845 124.605 ;
        RECT 68.52 123.6 68.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 -0.845 68.845 -0.515 ;
        RECT 68.515 -2.205 68.845 -1.875 ;
        RECT 68.515 -3.565 68.845 -3.235 ;
        RECT 68.52 -3.565 68.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 -91.965 68.845 -91.635 ;
        RECT 68.515 -93.325 68.845 -92.995 ;
        RECT 68.515 -94.685 68.845 -94.355 ;
        RECT 68.515 -96.045 68.845 -95.715 ;
        RECT 68.515 -97.405 68.845 -97.075 ;
        RECT 68.515 -98.765 68.845 -98.435 ;
        RECT 68.515 -100.125 68.845 -99.795 ;
        RECT 68.515 -101.485 68.845 -101.155 ;
        RECT 68.515 -102.845 68.845 -102.515 ;
        RECT 68.515 -104.205 68.845 -103.875 ;
        RECT 68.515 -105.565 68.845 -105.235 ;
        RECT 68.515 -106.925 68.845 -106.595 ;
        RECT 68.515 -108.285 68.845 -107.955 ;
        RECT 68.515 -109.645 68.845 -109.315 ;
        RECT 68.515 -111.005 68.845 -110.675 ;
        RECT 68.515 -112.365 68.845 -112.035 ;
        RECT 68.515 -113.725 68.845 -113.395 ;
        RECT 68.515 -115.085 68.845 -114.755 ;
        RECT 68.515 -116.445 68.845 -116.115 ;
        RECT 68.515 -117.805 68.845 -117.475 ;
        RECT 68.515 -119.165 68.845 -118.835 ;
        RECT 68.515 -120.525 68.845 -120.195 ;
        RECT 68.515 -121.885 68.845 -121.555 ;
        RECT 68.515 -123.245 68.845 -122.915 ;
        RECT 68.515 -124.605 68.845 -124.275 ;
        RECT 68.515 -125.965 68.845 -125.635 ;
        RECT 68.515 -127.325 68.845 -126.995 ;
        RECT 68.515 -128.685 68.845 -128.355 ;
        RECT 68.515 -130.045 68.845 -129.715 ;
        RECT 68.515 -131.405 68.845 -131.075 ;
        RECT 68.515 -132.765 68.845 -132.435 ;
        RECT 68.515 -134.125 68.845 -133.795 ;
        RECT 68.515 -135.485 68.845 -135.155 ;
        RECT 68.515 -136.845 68.845 -136.515 ;
        RECT 68.515 -138.205 68.845 -137.875 ;
        RECT 68.515 -139.565 68.845 -139.235 ;
        RECT 68.515 -140.925 68.845 -140.595 ;
        RECT 68.515 -142.285 68.845 -141.955 ;
        RECT 68.515 -143.645 68.845 -143.315 ;
        RECT 68.515 -145.005 68.845 -144.675 ;
        RECT 68.515 -146.365 68.845 -146.035 ;
        RECT 68.515 -147.725 68.845 -147.395 ;
        RECT 68.515 -149.085 68.845 -148.755 ;
        RECT 68.515 -150.445 68.845 -150.115 ;
        RECT 68.515 -151.805 68.845 -151.475 ;
        RECT 68.515 -153.165 68.845 -152.835 ;
        RECT 68.515 -154.525 68.845 -154.195 ;
        RECT 68.515 -155.885 68.845 -155.555 ;
        RECT 68.515 -157.245 68.845 -156.915 ;
        RECT 68.515 -162.89 68.845 -161.76 ;
        RECT 68.52 -163.005 68.84 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.76 -94.075 70.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 129.945 70.205 131.075 ;
        RECT 69.875 125.635 70.205 125.965 ;
        RECT 69.875 124.275 70.205 124.605 ;
        RECT 69.88 123.6 70.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 -96.045 70.205 -95.715 ;
        RECT 69.875 -97.405 70.205 -97.075 ;
        RECT 69.875 -98.765 70.205 -98.435 ;
        RECT 69.875 -100.125 70.205 -99.795 ;
        RECT 69.875 -101.485 70.205 -101.155 ;
        RECT 69.875 -102.845 70.205 -102.515 ;
        RECT 69.875 -104.205 70.205 -103.875 ;
        RECT 69.875 -105.565 70.205 -105.235 ;
        RECT 69.875 -106.925 70.205 -106.595 ;
        RECT 69.875 -108.285 70.205 -107.955 ;
        RECT 69.875 -109.645 70.205 -109.315 ;
        RECT 69.875 -111.005 70.205 -110.675 ;
        RECT 69.875 -112.365 70.205 -112.035 ;
        RECT 69.875 -113.725 70.205 -113.395 ;
        RECT 69.875 -115.085 70.205 -114.755 ;
        RECT 69.875 -116.445 70.205 -116.115 ;
        RECT 69.875 -117.805 70.205 -117.475 ;
        RECT 69.875 -119.165 70.205 -118.835 ;
        RECT 69.875 -120.525 70.205 -120.195 ;
        RECT 69.875 -121.885 70.205 -121.555 ;
        RECT 69.875 -123.245 70.205 -122.915 ;
        RECT 69.875 -124.605 70.205 -124.275 ;
        RECT 69.875 -125.965 70.205 -125.635 ;
        RECT 69.875 -127.325 70.205 -126.995 ;
        RECT 69.875 -128.685 70.205 -128.355 ;
        RECT 69.875 -130.045 70.205 -129.715 ;
        RECT 69.875 -131.405 70.205 -131.075 ;
        RECT 69.875 -132.765 70.205 -132.435 ;
        RECT 69.875 -134.125 70.205 -133.795 ;
        RECT 69.875 -135.485 70.205 -135.155 ;
        RECT 69.875 -136.845 70.205 -136.515 ;
        RECT 69.875 -138.205 70.205 -137.875 ;
        RECT 69.875 -139.565 70.205 -139.235 ;
        RECT 69.875 -140.925 70.205 -140.595 ;
        RECT 69.875 -142.285 70.205 -141.955 ;
        RECT 69.875 -143.645 70.205 -143.315 ;
        RECT 69.875 -145.005 70.205 -144.675 ;
        RECT 69.875 -146.365 70.205 -146.035 ;
        RECT 69.875 -147.725 70.205 -147.395 ;
        RECT 69.875 -149.085 70.205 -148.755 ;
        RECT 69.875 -150.445 70.205 -150.115 ;
        RECT 69.875 -151.805 70.205 -151.475 ;
        RECT 69.875 -153.165 70.205 -152.835 ;
        RECT 69.875 -154.525 70.205 -154.195 ;
        RECT 69.875 -155.885 70.205 -155.555 ;
        RECT 69.875 -157.245 70.205 -156.915 ;
        RECT 69.875 -162.89 70.205 -161.76 ;
        RECT 69.88 -163.005 70.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 129.945 71.565 131.075 ;
        RECT 71.235 125.635 71.565 125.965 ;
        RECT 71.235 124.275 71.565 124.605 ;
        RECT 71.24 123.6 71.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 -0.845 71.565 -0.515 ;
        RECT 71.235 -2.205 71.565 -1.875 ;
        RECT 71.235 -3.565 71.565 -3.235 ;
        RECT 71.24 -3.565 71.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 129.945 72.925 131.075 ;
        RECT 72.595 125.635 72.925 125.965 ;
        RECT 72.595 124.275 72.925 124.605 ;
        RECT 72.6 123.6 72.92 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 -0.845 72.925 -0.515 ;
        RECT 72.595 -2.205 72.925 -1.875 ;
        RECT 72.595 -3.565 72.925 -3.235 ;
        RECT 72.6 -3.565 72.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 129.945 74.285 131.075 ;
        RECT 73.955 125.635 74.285 125.965 ;
        RECT 73.955 124.275 74.285 124.605 ;
        RECT 73.96 123.6 74.28 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.96 -3.565 74.28 -0.515 ;
        RECT 73.955 -0.845 74.285 -0.515 ;
        RECT 73.955 -2.205 74.285 -1.875 ;
        RECT 73.955 -3.565 74.285 -3.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 129.945 0.845 131.075 ;
        RECT 0.515 125.635 0.845 125.965 ;
        RECT 0.515 124.275 0.845 124.605 ;
        RECT 0.52 123.6 0.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -0.845 0.845 -0.515 ;
        RECT 0.515 -2.205 0.845 -1.875 ;
        RECT 0.515 -3.565 0.845 -3.235 ;
        RECT 0.52 -3.565 0.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -91.965 0.845 -91.635 ;
        RECT 0.515 -93.325 0.845 -92.995 ;
        RECT 0.515 -94.685 0.845 -94.355 ;
        RECT 0.515 -96.045 0.845 -95.715 ;
        RECT 0.515 -97.405 0.845 -97.075 ;
        RECT 0.515 -98.765 0.845 -98.435 ;
        RECT 0.515 -100.125 0.845 -99.795 ;
        RECT 0.515 -101.485 0.845 -101.155 ;
        RECT 0.515 -102.845 0.845 -102.515 ;
        RECT 0.515 -104.205 0.845 -103.875 ;
        RECT 0.515 -105.565 0.845 -105.235 ;
        RECT 0.515 -106.925 0.845 -106.595 ;
        RECT 0.515 -108.285 0.845 -107.955 ;
        RECT 0.515 -109.645 0.845 -109.315 ;
        RECT 0.515 -111.005 0.845 -110.675 ;
        RECT 0.515 -112.365 0.845 -112.035 ;
        RECT 0.515 -113.725 0.845 -113.395 ;
        RECT 0.515 -115.085 0.845 -114.755 ;
        RECT 0.515 -116.445 0.845 -116.115 ;
        RECT 0.515 -117.805 0.845 -117.475 ;
        RECT 0.515 -119.165 0.845 -118.835 ;
        RECT 0.515 -120.525 0.845 -120.195 ;
        RECT 0.515 -121.885 0.845 -121.555 ;
        RECT 0.515 -123.245 0.845 -122.915 ;
        RECT 0.515 -124.605 0.845 -124.275 ;
        RECT 0.515 -125.965 0.845 -125.635 ;
        RECT 0.515 -127.325 0.845 -126.995 ;
        RECT 0.515 -128.685 0.845 -128.355 ;
        RECT 0.515 -130.045 0.845 -129.715 ;
        RECT 0.515 -131.405 0.845 -131.075 ;
        RECT 0.515 -132.765 0.845 -132.435 ;
        RECT 0.515 -134.125 0.845 -133.795 ;
        RECT 0.515 -135.485 0.845 -135.155 ;
        RECT 0.515 -136.845 0.845 -136.515 ;
        RECT 0.515 -138.205 0.845 -137.875 ;
        RECT 0.515 -139.565 0.845 -139.235 ;
        RECT 0.515 -140.925 0.845 -140.595 ;
        RECT 0.515 -142.285 0.845 -141.955 ;
        RECT 0.515 -143.645 0.845 -143.315 ;
        RECT 0.515 -145.005 0.845 -144.675 ;
        RECT 0.515 -146.365 0.845 -146.035 ;
        RECT 0.515 -147.725 0.845 -147.395 ;
        RECT 0.515 -149.085 0.845 -148.755 ;
        RECT 0.515 -150.445 0.845 -150.115 ;
        RECT 0.515 -151.805 0.845 -151.475 ;
        RECT 0.515 -153.165 0.845 -152.835 ;
        RECT 0.515 -154.525 0.845 -154.195 ;
        RECT 0.515 -155.885 0.845 -155.555 ;
        RECT 0.515 -157.245 0.845 -156.915 ;
        RECT 0.515 -162.89 0.845 -161.76 ;
        RECT 0.52 -163.005 0.84 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 129.945 2.205 131.075 ;
        RECT 1.875 125.635 2.205 125.965 ;
        RECT 1.875 124.275 2.205 124.605 ;
        RECT 1.88 123.6 2.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -0.845 2.205 -0.515 ;
        RECT 1.875 -2.205 2.205 -1.875 ;
        RECT 1.875 -3.565 2.205 -3.235 ;
        RECT 1.88 -3.565 2.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -91.965 2.205 -91.635 ;
        RECT 1.875 -93.325 2.205 -92.995 ;
        RECT 1.875 -94.685 2.205 -94.355 ;
        RECT 1.875 -96.045 2.205 -95.715 ;
        RECT 1.875 -97.405 2.205 -97.075 ;
        RECT 1.875 -98.765 2.205 -98.435 ;
        RECT 1.875 -100.125 2.205 -99.795 ;
        RECT 1.875 -101.485 2.205 -101.155 ;
        RECT 1.875 -102.845 2.205 -102.515 ;
        RECT 1.875 -104.205 2.205 -103.875 ;
        RECT 1.875 -105.565 2.205 -105.235 ;
        RECT 1.875 -106.925 2.205 -106.595 ;
        RECT 1.875 -108.285 2.205 -107.955 ;
        RECT 1.875 -109.645 2.205 -109.315 ;
        RECT 1.875 -111.005 2.205 -110.675 ;
        RECT 1.875 -112.365 2.205 -112.035 ;
        RECT 1.875 -113.725 2.205 -113.395 ;
        RECT 1.875 -115.085 2.205 -114.755 ;
        RECT 1.875 -116.445 2.205 -116.115 ;
        RECT 1.875 -117.805 2.205 -117.475 ;
        RECT 1.875 -119.165 2.205 -118.835 ;
        RECT 1.875 -120.525 2.205 -120.195 ;
        RECT 1.875 -121.885 2.205 -121.555 ;
        RECT 1.875 -123.245 2.205 -122.915 ;
        RECT 1.875 -124.605 2.205 -124.275 ;
        RECT 1.875 -125.965 2.205 -125.635 ;
        RECT 1.875 -127.325 2.205 -126.995 ;
        RECT 1.875 -128.685 2.205 -128.355 ;
        RECT 1.875 -130.045 2.205 -129.715 ;
        RECT 1.875 -131.405 2.205 -131.075 ;
        RECT 1.875 -132.765 2.205 -132.435 ;
        RECT 1.875 -134.125 2.205 -133.795 ;
        RECT 1.875 -135.485 2.205 -135.155 ;
        RECT 1.875 -136.845 2.205 -136.515 ;
        RECT 1.875 -138.205 2.205 -137.875 ;
        RECT 1.875 -139.565 2.205 -139.235 ;
        RECT 1.875 -140.925 2.205 -140.595 ;
        RECT 1.875 -142.285 2.205 -141.955 ;
        RECT 1.875 -143.645 2.205 -143.315 ;
        RECT 1.875 -145.005 2.205 -144.675 ;
        RECT 1.875 -146.365 2.205 -146.035 ;
        RECT 1.875 -147.725 2.205 -147.395 ;
        RECT 1.875 -149.085 2.205 -148.755 ;
        RECT 1.875 -150.445 2.205 -150.115 ;
        RECT 1.875 -151.805 2.205 -151.475 ;
        RECT 1.875 -153.165 2.205 -152.835 ;
        RECT 1.875 -154.525 2.205 -154.195 ;
        RECT 1.875 -155.885 2.205 -155.555 ;
        RECT 1.875 -157.245 2.205 -156.915 ;
        RECT 1.875 -162.89 2.205 -161.76 ;
        RECT 1.88 -163.005 2.2 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.66 -94.075 2.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 129.945 3.565 131.075 ;
        RECT 3.235 125.635 3.565 125.965 ;
        RECT 3.235 124.275 3.565 124.605 ;
        RECT 3.24 123.6 3.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 -96.045 3.565 -95.715 ;
        RECT 3.235 -97.405 3.565 -97.075 ;
        RECT 3.235 -98.765 3.565 -98.435 ;
        RECT 3.235 -100.125 3.565 -99.795 ;
        RECT 3.235 -101.485 3.565 -101.155 ;
        RECT 3.235 -102.845 3.565 -102.515 ;
        RECT 3.235 -104.205 3.565 -103.875 ;
        RECT 3.235 -105.565 3.565 -105.235 ;
        RECT 3.235 -106.925 3.565 -106.595 ;
        RECT 3.235 -108.285 3.565 -107.955 ;
        RECT 3.235 -109.645 3.565 -109.315 ;
        RECT 3.235 -111.005 3.565 -110.675 ;
        RECT 3.235 -112.365 3.565 -112.035 ;
        RECT 3.235 -113.725 3.565 -113.395 ;
        RECT 3.235 -115.085 3.565 -114.755 ;
        RECT 3.235 -116.445 3.565 -116.115 ;
        RECT 3.235 -117.805 3.565 -117.475 ;
        RECT 3.235 -119.165 3.565 -118.835 ;
        RECT 3.235 -120.525 3.565 -120.195 ;
        RECT 3.235 -121.885 3.565 -121.555 ;
        RECT 3.235 -123.245 3.565 -122.915 ;
        RECT 3.235 -124.605 3.565 -124.275 ;
        RECT 3.235 -125.965 3.565 -125.635 ;
        RECT 3.235 -127.325 3.565 -126.995 ;
        RECT 3.235 -128.685 3.565 -128.355 ;
        RECT 3.235 -130.045 3.565 -129.715 ;
        RECT 3.235 -131.405 3.565 -131.075 ;
        RECT 3.235 -132.765 3.565 -132.435 ;
        RECT 3.235 -134.125 3.565 -133.795 ;
        RECT 3.235 -135.485 3.565 -135.155 ;
        RECT 3.235 -136.845 3.565 -136.515 ;
        RECT 3.235 -138.205 3.565 -137.875 ;
        RECT 3.235 -139.565 3.565 -139.235 ;
        RECT 3.235 -140.925 3.565 -140.595 ;
        RECT 3.235 -142.285 3.565 -141.955 ;
        RECT 3.235 -143.645 3.565 -143.315 ;
        RECT 3.235 -145.005 3.565 -144.675 ;
        RECT 3.235 -146.365 3.565 -146.035 ;
        RECT 3.235 -147.725 3.565 -147.395 ;
        RECT 3.235 -149.085 3.565 -148.755 ;
        RECT 3.235 -150.445 3.565 -150.115 ;
        RECT 3.235 -151.805 3.565 -151.475 ;
        RECT 3.235 -153.165 3.565 -152.835 ;
        RECT 3.235 -154.525 3.565 -154.195 ;
        RECT 3.235 -155.885 3.565 -155.555 ;
        RECT 3.235 -157.245 3.565 -156.915 ;
        RECT 3.235 -162.89 3.565 -161.76 ;
        RECT 3.24 -163.005 3.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 129.945 4.925 131.075 ;
        RECT 4.595 125.635 4.925 125.965 ;
        RECT 4.595 124.275 4.925 124.605 ;
        RECT 4.6 123.6 4.92 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 -0.845 4.925 -0.515 ;
        RECT 4.595 -2.205 4.925 -1.875 ;
        RECT 4.595 -3.565 4.925 -3.235 ;
        RECT 4.6 -3.565 4.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 129.945 6.285 131.075 ;
        RECT 5.955 125.635 6.285 125.965 ;
        RECT 5.955 124.275 6.285 124.605 ;
        RECT 5.96 123.6 6.28 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 -0.845 6.285 -0.515 ;
        RECT 5.955 -2.205 6.285 -1.875 ;
        RECT 5.955 -3.565 6.285 -3.235 ;
        RECT 5.96 -3.565 6.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 129.945 7.645 131.075 ;
        RECT 7.315 125.635 7.645 125.965 ;
        RECT 7.315 124.275 7.645 124.605 ;
        RECT 7.32 123.6 7.64 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -0.845 7.645 -0.515 ;
        RECT 7.315 -2.205 7.645 -1.875 ;
        RECT 7.315 -3.565 7.645 -3.235 ;
        RECT 7.32 -3.565 7.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -91.965 7.645 -91.635 ;
        RECT 7.315 -93.325 7.645 -92.995 ;
        RECT 7.315 -94.685 7.645 -94.355 ;
        RECT 7.315 -96.045 7.645 -95.715 ;
        RECT 7.315 -97.405 7.645 -97.075 ;
        RECT 7.315 -98.765 7.645 -98.435 ;
        RECT 7.315 -100.125 7.645 -99.795 ;
        RECT 7.315 -101.485 7.645 -101.155 ;
        RECT 7.315 -102.845 7.645 -102.515 ;
        RECT 7.315 -104.205 7.645 -103.875 ;
        RECT 7.315 -105.565 7.645 -105.235 ;
        RECT 7.315 -106.925 7.645 -106.595 ;
        RECT 7.315 -108.285 7.645 -107.955 ;
        RECT 7.315 -109.645 7.645 -109.315 ;
        RECT 7.315 -111.005 7.645 -110.675 ;
        RECT 7.315 -112.365 7.645 -112.035 ;
        RECT 7.315 -113.725 7.645 -113.395 ;
        RECT 7.315 -115.085 7.645 -114.755 ;
        RECT 7.315 -116.445 7.645 -116.115 ;
        RECT 7.315 -117.805 7.645 -117.475 ;
        RECT 7.315 -119.165 7.645 -118.835 ;
        RECT 7.315 -120.525 7.645 -120.195 ;
        RECT 7.315 -121.885 7.645 -121.555 ;
        RECT 7.315 -123.245 7.645 -122.915 ;
        RECT 7.315 -124.605 7.645 -124.275 ;
        RECT 7.315 -125.965 7.645 -125.635 ;
        RECT 7.315 -127.325 7.645 -126.995 ;
        RECT 7.315 -128.685 7.645 -128.355 ;
        RECT 7.315 -130.045 7.645 -129.715 ;
        RECT 7.315 -131.405 7.645 -131.075 ;
        RECT 7.315 -132.765 7.645 -132.435 ;
        RECT 7.315 -134.125 7.645 -133.795 ;
        RECT 7.315 -135.485 7.645 -135.155 ;
        RECT 7.315 -136.845 7.645 -136.515 ;
        RECT 7.315 -138.205 7.645 -137.875 ;
        RECT 7.315 -139.565 7.645 -139.235 ;
        RECT 7.315 -140.925 7.645 -140.595 ;
        RECT 7.315 -142.285 7.645 -141.955 ;
        RECT 7.315 -143.645 7.645 -143.315 ;
        RECT 7.315 -145.005 7.645 -144.675 ;
        RECT 7.315 -146.365 7.645 -146.035 ;
        RECT 7.315 -147.725 7.645 -147.395 ;
        RECT 7.315 -149.085 7.645 -148.755 ;
        RECT 7.315 -150.445 7.645 -150.115 ;
        RECT 7.315 -151.805 7.645 -151.475 ;
        RECT 7.315 -153.165 7.645 -152.835 ;
        RECT 7.315 -154.525 7.645 -154.195 ;
        RECT 7.315 -155.885 7.645 -155.555 ;
        RECT 7.315 -157.245 7.645 -156.915 ;
        RECT 7.315 -162.89 7.645 -161.76 ;
        RECT 7.32 -163.005 7.64 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 129.945 9.005 131.075 ;
        RECT 8.675 125.635 9.005 125.965 ;
        RECT 8.675 124.275 9.005 124.605 ;
        RECT 8.68 123.6 9 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 -96.045 9.005 -95.715 ;
        RECT 8.675 -97.405 9.005 -97.075 ;
        RECT 8.675 -98.765 9.005 -98.435 ;
        RECT 8.675 -100.125 9.005 -99.795 ;
        RECT 8.675 -101.485 9.005 -101.155 ;
        RECT 8.675 -102.845 9.005 -102.515 ;
        RECT 8.675 -104.205 9.005 -103.875 ;
        RECT 8.675 -105.565 9.005 -105.235 ;
        RECT 8.675 -106.925 9.005 -106.595 ;
        RECT 8.675 -108.285 9.005 -107.955 ;
        RECT 8.675 -109.645 9.005 -109.315 ;
        RECT 8.675 -111.005 9.005 -110.675 ;
        RECT 8.675 -112.365 9.005 -112.035 ;
        RECT 8.675 -113.725 9.005 -113.395 ;
        RECT 8.675 -115.085 9.005 -114.755 ;
        RECT 8.675 -116.445 9.005 -116.115 ;
        RECT 8.675 -117.805 9.005 -117.475 ;
        RECT 8.675 -119.165 9.005 -118.835 ;
        RECT 8.675 -120.525 9.005 -120.195 ;
        RECT 8.675 -121.885 9.005 -121.555 ;
        RECT 8.675 -123.245 9.005 -122.915 ;
        RECT 8.675 -124.605 9.005 -124.275 ;
        RECT 8.675 -125.965 9.005 -125.635 ;
        RECT 8.675 -127.325 9.005 -126.995 ;
        RECT 8.675 -128.685 9.005 -128.355 ;
        RECT 8.675 -130.045 9.005 -129.715 ;
        RECT 8.675 -131.405 9.005 -131.075 ;
        RECT 8.675 -132.765 9.005 -132.435 ;
        RECT 8.675 -134.125 9.005 -133.795 ;
        RECT 8.675 -135.485 9.005 -135.155 ;
        RECT 8.675 -136.845 9.005 -136.515 ;
        RECT 8.675 -138.205 9.005 -137.875 ;
        RECT 8.675 -139.565 9.005 -139.235 ;
        RECT 8.675 -140.925 9.005 -140.595 ;
        RECT 8.675 -142.285 9.005 -141.955 ;
        RECT 8.675 -143.645 9.005 -143.315 ;
        RECT 8.675 -145.005 9.005 -144.675 ;
        RECT 8.675 -146.365 9.005 -146.035 ;
        RECT 8.675 -147.725 9.005 -147.395 ;
        RECT 8.675 -149.085 9.005 -148.755 ;
        RECT 8.675 -150.445 9.005 -150.115 ;
        RECT 8.675 -151.805 9.005 -151.475 ;
        RECT 8.675 -153.165 9.005 -152.835 ;
        RECT 8.675 -154.525 9.005 -154.195 ;
        RECT 8.675 -155.885 9.005 -155.555 ;
        RECT 8.675 -157.245 9.005 -156.915 ;
        RECT 8.675 -162.89 9.005 -161.76 ;
        RECT 8.68 -163.005 9 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.76 -94.075 9.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 129.945 10.365 131.075 ;
        RECT 10.035 125.635 10.365 125.965 ;
        RECT 10.035 124.275 10.365 124.605 ;
        RECT 10.04 123.6 10.36 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 129.945 11.725 131.075 ;
        RECT 11.395 125.635 11.725 125.965 ;
        RECT 11.395 124.275 11.725 124.605 ;
        RECT 11.4 123.6 11.72 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 -0.845 11.725 -0.515 ;
        RECT 11.395 -2.205 11.725 -1.875 ;
        RECT 11.395 -3.565 11.725 -3.235 ;
        RECT 11.4 -3.565 11.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 129.945 13.085 131.075 ;
        RECT 12.755 125.635 13.085 125.965 ;
        RECT 12.755 124.275 13.085 124.605 ;
        RECT 12.76 123.6 13.08 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -0.845 13.085 -0.515 ;
        RECT 12.755 -2.205 13.085 -1.875 ;
        RECT 12.755 -3.565 13.085 -3.235 ;
        RECT 12.76 -3.565 13.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -91.965 13.085 -91.635 ;
        RECT 12.755 -93.325 13.085 -92.995 ;
        RECT 12.755 -94.685 13.085 -94.355 ;
        RECT 12.755 -96.045 13.085 -95.715 ;
        RECT 12.755 -97.405 13.085 -97.075 ;
        RECT 12.755 -98.765 13.085 -98.435 ;
        RECT 12.755 -100.125 13.085 -99.795 ;
        RECT 12.755 -101.485 13.085 -101.155 ;
        RECT 12.755 -102.845 13.085 -102.515 ;
        RECT 12.755 -104.205 13.085 -103.875 ;
        RECT 12.755 -105.565 13.085 -105.235 ;
        RECT 12.755 -106.925 13.085 -106.595 ;
        RECT 12.755 -108.285 13.085 -107.955 ;
        RECT 12.755 -109.645 13.085 -109.315 ;
        RECT 12.755 -111.005 13.085 -110.675 ;
        RECT 12.755 -112.365 13.085 -112.035 ;
        RECT 12.755 -113.725 13.085 -113.395 ;
        RECT 12.755 -115.085 13.085 -114.755 ;
        RECT 12.755 -116.445 13.085 -116.115 ;
        RECT 12.755 -117.805 13.085 -117.475 ;
        RECT 12.755 -119.165 13.085 -118.835 ;
        RECT 12.755 -120.525 13.085 -120.195 ;
        RECT 12.755 -121.885 13.085 -121.555 ;
        RECT 12.755 -123.245 13.085 -122.915 ;
        RECT 12.755 -124.605 13.085 -124.275 ;
        RECT 12.755 -125.965 13.085 -125.635 ;
        RECT 12.755 -127.325 13.085 -126.995 ;
        RECT 12.755 -128.685 13.085 -128.355 ;
        RECT 12.755 -130.045 13.085 -129.715 ;
        RECT 12.755 -131.405 13.085 -131.075 ;
        RECT 12.755 -132.765 13.085 -132.435 ;
        RECT 12.755 -134.125 13.085 -133.795 ;
        RECT 12.755 -135.485 13.085 -135.155 ;
        RECT 12.755 -136.845 13.085 -136.515 ;
        RECT 12.755 -138.205 13.085 -137.875 ;
        RECT 12.755 -139.565 13.085 -139.235 ;
        RECT 12.755 -140.925 13.085 -140.595 ;
        RECT 12.755 -142.285 13.085 -141.955 ;
        RECT 12.755 -143.645 13.085 -143.315 ;
        RECT 12.755 -145.005 13.085 -144.675 ;
        RECT 12.755 -146.365 13.085 -146.035 ;
        RECT 12.755 -147.725 13.085 -147.395 ;
        RECT 12.755 -149.085 13.085 -148.755 ;
        RECT 12.755 -150.445 13.085 -150.115 ;
        RECT 12.755 -151.805 13.085 -151.475 ;
        RECT 12.755 -153.165 13.085 -152.835 ;
        RECT 12.755 -154.525 13.085 -154.195 ;
        RECT 12.755 -155.885 13.085 -155.555 ;
        RECT 12.755 -157.245 13.085 -156.915 ;
        RECT 12.755 -162.89 13.085 -161.76 ;
        RECT 12.76 -163.005 13.08 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 129.945 14.445 131.075 ;
        RECT 14.115 125.635 14.445 125.965 ;
        RECT 14.115 124.275 14.445 124.605 ;
        RECT 14.12 123.6 14.44 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -0.845 14.445 -0.515 ;
        RECT 14.115 -2.205 14.445 -1.875 ;
        RECT 14.115 -3.565 14.445 -3.235 ;
        RECT 14.12 -3.565 14.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -91.965 14.445 -91.635 ;
        RECT 14.115 -93.325 14.445 -92.995 ;
        RECT 14.115 -94.685 14.445 -94.355 ;
        RECT 14.115 -96.045 14.445 -95.715 ;
        RECT 14.115 -97.405 14.445 -97.075 ;
        RECT 14.115 -98.765 14.445 -98.435 ;
        RECT 14.115 -100.125 14.445 -99.795 ;
        RECT 14.115 -101.485 14.445 -101.155 ;
        RECT 14.115 -102.845 14.445 -102.515 ;
        RECT 14.115 -104.205 14.445 -103.875 ;
        RECT 14.115 -105.565 14.445 -105.235 ;
        RECT 14.115 -106.925 14.445 -106.595 ;
        RECT 14.115 -108.285 14.445 -107.955 ;
        RECT 14.115 -109.645 14.445 -109.315 ;
        RECT 14.115 -111.005 14.445 -110.675 ;
        RECT 14.115 -112.365 14.445 -112.035 ;
        RECT 14.115 -113.725 14.445 -113.395 ;
        RECT 14.115 -115.085 14.445 -114.755 ;
        RECT 14.115 -116.445 14.445 -116.115 ;
        RECT 14.115 -117.805 14.445 -117.475 ;
        RECT 14.115 -119.165 14.445 -118.835 ;
        RECT 14.115 -120.525 14.445 -120.195 ;
        RECT 14.115 -121.885 14.445 -121.555 ;
        RECT 14.115 -123.245 14.445 -122.915 ;
        RECT 14.115 -124.605 14.445 -124.275 ;
        RECT 14.115 -125.965 14.445 -125.635 ;
        RECT 14.115 -127.325 14.445 -126.995 ;
        RECT 14.115 -128.685 14.445 -128.355 ;
        RECT 14.115 -130.045 14.445 -129.715 ;
        RECT 14.115 -131.405 14.445 -131.075 ;
        RECT 14.115 -132.765 14.445 -132.435 ;
        RECT 14.115 -134.125 14.445 -133.795 ;
        RECT 14.115 -135.485 14.445 -135.155 ;
        RECT 14.115 -136.845 14.445 -136.515 ;
        RECT 14.115 -138.205 14.445 -137.875 ;
        RECT 14.115 -139.565 14.445 -139.235 ;
        RECT 14.115 -140.925 14.445 -140.595 ;
        RECT 14.115 -142.285 14.445 -141.955 ;
        RECT 14.115 -143.645 14.445 -143.315 ;
        RECT 14.115 -145.005 14.445 -144.675 ;
        RECT 14.115 -146.365 14.445 -146.035 ;
        RECT 14.115 -147.725 14.445 -147.395 ;
        RECT 14.115 -149.085 14.445 -148.755 ;
        RECT 14.115 -150.445 14.445 -150.115 ;
        RECT 14.115 -151.805 14.445 -151.475 ;
        RECT 14.115 -153.165 14.445 -152.835 ;
        RECT 14.115 -154.525 14.445 -154.195 ;
        RECT 14.115 -155.885 14.445 -155.555 ;
        RECT 14.115 -157.245 14.445 -156.915 ;
        RECT 14.115 -162.89 14.445 -161.76 ;
        RECT 14.12 -163.005 14.44 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.86 -94.075 15.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 129.945 15.805 131.075 ;
        RECT 15.475 125.635 15.805 125.965 ;
        RECT 15.475 124.275 15.805 124.605 ;
        RECT 15.48 123.6 15.8 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 -96.045 15.805 -95.715 ;
        RECT 15.475 -97.405 15.805 -97.075 ;
        RECT 15.475 -98.765 15.805 -98.435 ;
        RECT 15.475 -100.125 15.805 -99.795 ;
        RECT 15.475 -101.485 15.805 -101.155 ;
        RECT 15.475 -102.845 15.805 -102.515 ;
        RECT 15.475 -104.205 15.805 -103.875 ;
        RECT 15.475 -105.565 15.805 -105.235 ;
        RECT 15.475 -106.925 15.805 -106.595 ;
        RECT 15.475 -108.285 15.805 -107.955 ;
        RECT 15.475 -109.645 15.805 -109.315 ;
        RECT 15.475 -111.005 15.805 -110.675 ;
        RECT 15.475 -112.365 15.805 -112.035 ;
        RECT 15.475 -113.725 15.805 -113.395 ;
        RECT 15.475 -115.085 15.805 -114.755 ;
        RECT 15.475 -116.445 15.805 -116.115 ;
        RECT 15.475 -117.805 15.805 -117.475 ;
        RECT 15.475 -119.165 15.805 -118.835 ;
        RECT 15.475 -120.525 15.805 -120.195 ;
        RECT 15.475 -121.885 15.805 -121.555 ;
        RECT 15.475 -123.245 15.805 -122.915 ;
        RECT 15.475 -124.605 15.805 -124.275 ;
        RECT 15.475 -125.965 15.805 -125.635 ;
        RECT 15.475 -127.325 15.805 -126.995 ;
        RECT 15.475 -128.685 15.805 -128.355 ;
        RECT 15.475 -130.045 15.805 -129.715 ;
        RECT 15.475 -131.405 15.805 -131.075 ;
        RECT 15.475 -132.765 15.805 -132.435 ;
        RECT 15.475 -134.125 15.805 -133.795 ;
        RECT 15.475 -135.485 15.805 -135.155 ;
        RECT 15.475 -136.845 15.805 -136.515 ;
        RECT 15.475 -138.205 15.805 -137.875 ;
        RECT 15.475 -139.565 15.805 -139.235 ;
        RECT 15.475 -140.925 15.805 -140.595 ;
        RECT 15.475 -142.285 15.805 -141.955 ;
        RECT 15.475 -143.645 15.805 -143.315 ;
        RECT 15.475 -145.005 15.805 -144.675 ;
        RECT 15.475 -146.365 15.805 -146.035 ;
        RECT 15.475 -147.725 15.805 -147.395 ;
        RECT 15.475 -149.085 15.805 -148.755 ;
        RECT 15.475 -150.445 15.805 -150.115 ;
        RECT 15.475 -151.805 15.805 -151.475 ;
        RECT 15.475 -153.165 15.805 -152.835 ;
        RECT 15.475 -154.525 15.805 -154.195 ;
        RECT 15.475 -155.885 15.805 -155.555 ;
        RECT 15.475 -157.245 15.805 -156.915 ;
        RECT 15.475 -162.89 15.805 -161.76 ;
        RECT 15.48 -163.005 15.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 129.945 17.165 131.075 ;
        RECT 16.835 125.635 17.165 125.965 ;
        RECT 16.835 124.275 17.165 124.605 ;
        RECT 16.84 123.6 17.16 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 -0.845 17.165 -0.515 ;
        RECT 16.835 -2.205 17.165 -1.875 ;
        RECT 16.835 -3.565 17.165 -3.235 ;
        RECT 16.84 -3.565 17.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 129.945 18.525 131.075 ;
        RECT 18.195 125.635 18.525 125.965 ;
        RECT 18.195 124.275 18.525 124.605 ;
        RECT 18.2 123.6 18.52 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 -0.845 18.525 -0.515 ;
        RECT 18.195 -2.205 18.525 -1.875 ;
        RECT 18.195 -3.565 18.525 -3.235 ;
        RECT 18.2 -3.565 18.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 129.945 19.885 131.075 ;
        RECT 19.555 125.635 19.885 125.965 ;
        RECT 19.555 124.275 19.885 124.605 ;
        RECT 19.56 123.6 19.88 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -0.845 19.885 -0.515 ;
        RECT 19.555 -2.205 19.885 -1.875 ;
        RECT 19.555 -3.565 19.885 -3.235 ;
        RECT 19.56 -3.565 19.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -91.965 19.885 -91.635 ;
        RECT 19.555 -93.325 19.885 -92.995 ;
        RECT 19.555 -94.685 19.885 -94.355 ;
        RECT 19.555 -96.045 19.885 -95.715 ;
        RECT 19.555 -97.405 19.885 -97.075 ;
        RECT 19.555 -98.765 19.885 -98.435 ;
        RECT 19.555 -100.125 19.885 -99.795 ;
        RECT 19.555 -101.485 19.885 -101.155 ;
        RECT 19.555 -102.845 19.885 -102.515 ;
        RECT 19.555 -104.205 19.885 -103.875 ;
        RECT 19.555 -105.565 19.885 -105.235 ;
        RECT 19.555 -106.925 19.885 -106.595 ;
        RECT 19.555 -108.285 19.885 -107.955 ;
        RECT 19.555 -109.645 19.885 -109.315 ;
        RECT 19.555 -111.005 19.885 -110.675 ;
        RECT 19.555 -112.365 19.885 -112.035 ;
        RECT 19.555 -113.725 19.885 -113.395 ;
        RECT 19.555 -115.085 19.885 -114.755 ;
        RECT 19.555 -116.445 19.885 -116.115 ;
        RECT 19.555 -117.805 19.885 -117.475 ;
        RECT 19.555 -119.165 19.885 -118.835 ;
        RECT 19.555 -120.525 19.885 -120.195 ;
        RECT 19.555 -121.885 19.885 -121.555 ;
        RECT 19.555 -123.245 19.885 -122.915 ;
        RECT 19.555 -124.605 19.885 -124.275 ;
        RECT 19.555 -125.965 19.885 -125.635 ;
        RECT 19.555 -127.325 19.885 -126.995 ;
        RECT 19.555 -128.685 19.885 -128.355 ;
        RECT 19.555 -130.045 19.885 -129.715 ;
        RECT 19.555 -131.405 19.885 -131.075 ;
        RECT 19.555 -132.765 19.885 -132.435 ;
        RECT 19.555 -134.125 19.885 -133.795 ;
        RECT 19.555 -135.485 19.885 -135.155 ;
        RECT 19.555 -136.845 19.885 -136.515 ;
        RECT 19.555 -138.205 19.885 -137.875 ;
        RECT 19.555 -139.565 19.885 -139.235 ;
        RECT 19.555 -140.925 19.885 -140.595 ;
        RECT 19.555 -142.285 19.885 -141.955 ;
        RECT 19.555 -143.645 19.885 -143.315 ;
        RECT 19.555 -145.005 19.885 -144.675 ;
        RECT 19.555 -146.365 19.885 -146.035 ;
        RECT 19.555 -147.725 19.885 -147.395 ;
        RECT 19.555 -149.085 19.885 -148.755 ;
        RECT 19.555 -150.445 19.885 -150.115 ;
        RECT 19.555 -151.805 19.885 -151.475 ;
        RECT 19.555 -153.165 19.885 -152.835 ;
        RECT 19.555 -154.525 19.885 -154.195 ;
        RECT 19.555 -155.885 19.885 -155.555 ;
        RECT 19.555 -157.245 19.885 -156.915 ;
        RECT 19.555 -162.89 19.885 -161.76 ;
        RECT 19.56 -163.005 19.88 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 129.945 21.245 131.075 ;
        RECT 20.915 125.635 21.245 125.965 ;
        RECT 20.915 124.275 21.245 124.605 ;
        RECT 20.92 123.6 21.24 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 -96.045 21.245 -95.715 ;
        RECT 20.915 -97.405 21.245 -97.075 ;
        RECT 20.915 -98.765 21.245 -98.435 ;
        RECT 20.915 -100.125 21.245 -99.795 ;
        RECT 20.915 -101.485 21.245 -101.155 ;
        RECT 20.915 -102.845 21.245 -102.515 ;
        RECT 20.915 -104.205 21.245 -103.875 ;
        RECT 20.915 -105.565 21.245 -105.235 ;
        RECT 20.915 -106.925 21.245 -106.595 ;
        RECT 20.915 -108.285 21.245 -107.955 ;
        RECT 20.915 -109.645 21.245 -109.315 ;
        RECT 20.915 -111.005 21.245 -110.675 ;
        RECT 20.915 -112.365 21.245 -112.035 ;
        RECT 20.915 -113.725 21.245 -113.395 ;
        RECT 20.915 -115.085 21.245 -114.755 ;
        RECT 20.915 -116.445 21.245 -116.115 ;
        RECT 20.915 -117.805 21.245 -117.475 ;
        RECT 20.915 -119.165 21.245 -118.835 ;
        RECT 20.915 -120.525 21.245 -120.195 ;
        RECT 20.915 -121.885 21.245 -121.555 ;
        RECT 20.915 -123.245 21.245 -122.915 ;
        RECT 20.915 -124.605 21.245 -124.275 ;
        RECT 20.915 -125.965 21.245 -125.635 ;
        RECT 20.915 -127.325 21.245 -126.995 ;
        RECT 20.915 -128.685 21.245 -128.355 ;
        RECT 20.915 -130.045 21.245 -129.715 ;
        RECT 20.915 -131.405 21.245 -131.075 ;
        RECT 20.915 -132.765 21.245 -132.435 ;
        RECT 20.915 -134.125 21.245 -133.795 ;
        RECT 20.915 -135.485 21.245 -135.155 ;
        RECT 20.915 -136.845 21.245 -136.515 ;
        RECT 20.915 -138.205 21.245 -137.875 ;
        RECT 20.915 -139.565 21.245 -139.235 ;
        RECT 20.915 -140.925 21.245 -140.595 ;
        RECT 20.915 -142.285 21.245 -141.955 ;
        RECT 20.915 -143.645 21.245 -143.315 ;
        RECT 20.915 -145.005 21.245 -144.675 ;
        RECT 20.915 -146.365 21.245 -146.035 ;
        RECT 20.915 -147.725 21.245 -147.395 ;
        RECT 20.915 -149.085 21.245 -148.755 ;
        RECT 20.915 -150.445 21.245 -150.115 ;
        RECT 20.915 -151.805 21.245 -151.475 ;
        RECT 20.915 -153.165 21.245 -152.835 ;
        RECT 20.915 -154.525 21.245 -154.195 ;
        RECT 20.915 -155.885 21.245 -155.555 ;
        RECT 20.915 -157.245 21.245 -156.915 ;
        RECT 20.915 -162.89 21.245 -161.76 ;
        RECT 20.92 -163.005 21.24 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.96 -94.075 21.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 129.945 22.605 131.075 ;
        RECT 22.275 125.635 22.605 125.965 ;
        RECT 22.275 124.275 22.605 124.605 ;
        RECT 22.28 123.6 22.6 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 129.945 23.965 131.075 ;
        RECT 23.635 125.635 23.965 125.965 ;
        RECT 23.635 124.275 23.965 124.605 ;
        RECT 23.64 123.6 23.96 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 -0.845 23.965 -0.515 ;
        RECT 23.635 -2.205 23.965 -1.875 ;
        RECT 23.635 -3.565 23.965 -3.235 ;
        RECT 23.64 -3.565 23.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 129.945 25.325 131.075 ;
        RECT 24.995 125.635 25.325 125.965 ;
        RECT 24.995 124.275 25.325 124.605 ;
        RECT 25 123.6 25.32 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -0.845 25.325 -0.515 ;
        RECT 24.995 -2.205 25.325 -1.875 ;
        RECT 24.995 -3.565 25.325 -3.235 ;
        RECT 25 -3.565 25.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -91.965 25.325 -91.635 ;
        RECT 24.995 -93.325 25.325 -92.995 ;
        RECT 24.995 -94.685 25.325 -94.355 ;
        RECT 24.995 -96.045 25.325 -95.715 ;
        RECT 24.995 -97.405 25.325 -97.075 ;
        RECT 24.995 -98.765 25.325 -98.435 ;
        RECT 24.995 -100.125 25.325 -99.795 ;
        RECT 24.995 -101.485 25.325 -101.155 ;
        RECT 24.995 -102.845 25.325 -102.515 ;
        RECT 24.995 -104.205 25.325 -103.875 ;
        RECT 24.995 -105.565 25.325 -105.235 ;
        RECT 24.995 -106.925 25.325 -106.595 ;
        RECT 24.995 -108.285 25.325 -107.955 ;
        RECT 24.995 -109.645 25.325 -109.315 ;
        RECT 24.995 -111.005 25.325 -110.675 ;
        RECT 24.995 -112.365 25.325 -112.035 ;
        RECT 24.995 -113.725 25.325 -113.395 ;
        RECT 24.995 -115.085 25.325 -114.755 ;
        RECT 24.995 -116.445 25.325 -116.115 ;
        RECT 24.995 -117.805 25.325 -117.475 ;
        RECT 24.995 -119.165 25.325 -118.835 ;
        RECT 24.995 -120.525 25.325 -120.195 ;
        RECT 24.995 -121.885 25.325 -121.555 ;
        RECT 24.995 -123.245 25.325 -122.915 ;
        RECT 24.995 -124.605 25.325 -124.275 ;
        RECT 24.995 -125.965 25.325 -125.635 ;
        RECT 24.995 -127.325 25.325 -126.995 ;
        RECT 24.995 -128.685 25.325 -128.355 ;
        RECT 24.995 -130.045 25.325 -129.715 ;
        RECT 24.995 -131.405 25.325 -131.075 ;
        RECT 24.995 -132.765 25.325 -132.435 ;
        RECT 24.995 -134.125 25.325 -133.795 ;
        RECT 24.995 -135.485 25.325 -135.155 ;
        RECT 24.995 -136.845 25.325 -136.515 ;
        RECT 24.995 -138.205 25.325 -137.875 ;
        RECT 24.995 -139.565 25.325 -139.235 ;
        RECT 24.995 -140.925 25.325 -140.595 ;
        RECT 24.995 -142.285 25.325 -141.955 ;
        RECT 24.995 -143.645 25.325 -143.315 ;
        RECT 24.995 -145.005 25.325 -144.675 ;
        RECT 24.995 -146.365 25.325 -146.035 ;
        RECT 24.995 -147.725 25.325 -147.395 ;
        RECT 24.995 -149.085 25.325 -148.755 ;
        RECT 24.995 -150.445 25.325 -150.115 ;
        RECT 24.995 -151.805 25.325 -151.475 ;
        RECT 24.995 -153.165 25.325 -152.835 ;
        RECT 24.995 -154.525 25.325 -154.195 ;
        RECT 24.995 -155.885 25.325 -155.555 ;
        RECT 24.995 -157.245 25.325 -156.915 ;
        RECT 24.995 -162.89 25.325 -161.76 ;
        RECT 25 -163.005 25.32 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 129.945 26.685 131.075 ;
        RECT 26.355 125.635 26.685 125.965 ;
        RECT 26.355 124.275 26.685 124.605 ;
        RECT 26.36 123.6 26.68 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -0.845 26.685 -0.515 ;
        RECT 26.355 -2.205 26.685 -1.875 ;
        RECT 26.355 -3.565 26.685 -3.235 ;
        RECT 26.36 -3.565 26.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -91.965 26.685 -91.635 ;
        RECT 26.355 -93.325 26.685 -92.995 ;
        RECT 26.355 -94.685 26.685 -94.355 ;
        RECT 26.355 -96.045 26.685 -95.715 ;
        RECT 26.355 -97.405 26.685 -97.075 ;
        RECT 26.355 -98.765 26.685 -98.435 ;
        RECT 26.355 -100.125 26.685 -99.795 ;
        RECT 26.355 -101.485 26.685 -101.155 ;
        RECT 26.355 -102.845 26.685 -102.515 ;
        RECT 26.355 -104.205 26.685 -103.875 ;
        RECT 26.355 -105.565 26.685 -105.235 ;
        RECT 26.355 -106.925 26.685 -106.595 ;
        RECT 26.355 -108.285 26.685 -107.955 ;
        RECT 26.355 -109.645 26.685 -109.315 ;
        RECT 26.355 -111.005 26.685 -110.675 ;
        RECT 26.355 -112.365 26.685 -112.035 ;
        RECT 26.355 -113.725 26.685 -113.395 ;
        RECT 26.355 -115.085 26.685 -114.755 ;
        RECT 26.355 -116.445 26.685 -116.115 ;
        RECT 26.355 -117.805 26.685 -117.475 ;
        RECT 26.355 -119.165 26.685 -118.835 ;
        RECT 26.355 -120.525 26.685 -120.195 ;
        RECT 26.355 -121.885 26.685 -121.555 ;
        RECT 26.355 -123.245 26.685 -122.915 ;
        RECT 26.355 -124.605 26.685 -124.275 ;
        RECT 26.355 -125.965 26.685 -125.635 ;
        RECT 26.355 -127.325 26.685 -126.995 ;
        RECT 26.355 -128.685 26.685 -128.355 ;
        RECT 26.355 -130.045 26.685 -129.715 ;
        RECT 26.355 -131.405 26.685 -131.075 ;
        RECT 26.355 -132.765 26.685 -132.435 ;
        RECT 26.355 -134.125 26.685 -133.795 ;
        RECT 26.355 -135.485 26.685 -135.155 ;
        RECT 26.355 -136.845 26.685 -136.515 ;
        RECT 26.355 -138.205 26.685 -137.875 ;
        RECT 26.355 -139.565 26.685 -139.235 ;
        RECT 26.355 -140.925 26.685 -140.595 ;
        RECT 26.355 -142.285 26.685 -141.955 ;
        RECT 26.355 -143.645 26.685 -143.315 ;
        RECT 26.355 -145.005 26.685 -144.675 ;
        RECT 26.355 -146.365 26.685 -146.035 ;
        RECT 26.355 -147.725 26.685 -147.395 ;
        RECT 26.355 -149.085 26.685 -148.755 ;
        RECT 26.355 -150.445 26.685 -150.115 ;
        RECT 26.355 -151.805 26.685 -151.475 ;
        RECT 26.355 -153.165 26.685 -152.835 ;
        RECT 26.355 -154.525 26.685 -154.195 ;
        RECT 26.355 -155.885 26.685 -155.555 ;
        RECT 26.355 -157.245 26.685 -156.915 ;
        RECT 26.355 -162.89 26.685 -161.76 ;
        RECT 26.36 -163.005 26.68 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.06 -94.075 27.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 129.945 28.045 131.075 ;
        RECT 27.715 125.635 28.045 125.965 ;
        RECT 27.715 124.275 28.045 124.605 ;
        RECT 27.72 123.6 28.04 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 -96.045 28.045 -95.715 ;
        RECT 27.715 -97.405 28.045 -97.075 ;
        RECT 27.715 -98.765 28.045 -98.435 ;
        RECT 27.715 -100.125 28.045 -99.795 ;
        RECT 27.715 -101.485 28.045 -101.155 ;
        RECT 27.715 -102.845 28.045 -102.515 ;
        RECT 27.715 -104.205 28.045 -103.875 ;
        RECT 27.715 -105.565 28.045 -105.235 ;
        RECT 27.715 -106.925 28.045 -106.595 ;
        RECT 27.715 -108.285 28.045 -107.955 ;
        RECT 27.715 -109.645 28.045 -109.315 ;
        RECT 27.715 -111.005 28.045 -110.675 ;
        RECT 27.715 -112.365 28.045 -112.035 ;
        RECT 27.715 -113.725 28.045 -113.395 ;
        RECT 27.715 -115.085 28.045 -114.755 ;
        RECT 27.715 -116.445 28.045 -116.115 ;
        RECT 27.715 -117.805 28.045 -117.475 ;
        RECT 27.715 -119.165 28.045 -118.835 ;
        RECT 27.715 -120.525 28.045 -120.195 ;
        RECT 27.715 -121.885 28.045 -121.555 ;
        RECT 27.715 -123.245 28.045 -122.915 ;
        RECT 27.715 -124.605 28.045 -124.275 ;
        RECT 27.715 -125.965 28.045 -125.635 ;
        RECT 27.715 -127.325 28.045 -126.995 ;
        RECT 27.715 -128.685 28.045 -128.355 ;
        RECT 27.715 -130.045 28.045 -129.715 ;
        RECT 27.715 -131.405 28.045 -131.075 ;
        RECT 27.715 -132.765 28.045 -132.435 ;
        RECT 27.715 -134.125 28.045 -133.795 ;
        RECT 27.715 -135.485 28.045 -135.155 ;
        RECT 27.715 -136.845 28.045 -136.515 ;
        RECT 27.715 -138.205 28.045 -137.875 ;
        RECT 27.715 -139.565 28.045 -139.235 ;
        RECT 27.715 -140.925 28.045 -140.595 ;
        RECT 27.715 -142.285 28.045 -141.955 ;
        RECT 27.715 -143.645 28.045 -143.315 ;
        RECT 27.715 -145.005 28.045 -144.675 ;
        RECT 27.715 -146.365 28.045 -146.035 ;
        RECT 27.715 -147.725 28.045 -147.395 ;
        RECT 27.715 -149.085 28.045 -148.755 ;
        RECT 27.715 -150.445 28.045 -150.115 ;
        RECT 27.715 -151.805 28.045 -151.475 ;
        RECT 27.715 -153.165 28.045 -152.835 ;
        RECT 27.715 -154.525 28.045 -154.195 ;
        RECT 27.715 -155.885 28.045 -155.555 ;
        RECT 27.715 -157.245 28.045 -156.915 ;
        RECT 27.715 -162.89 28.045 -161.76 ;
        RECT 27.72 -163.005 28.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 129.945 29.405 131.075 ;
        RECT 29.075 125.635 29.405 125.965 ;
        RECT 29.075 124.275 29.405 124.605 ;
        RECT 29.08 123.6 29.4 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -0.845 29.405 -0.515 ;
        RECT 29.075 -2.205 29.405 -1.875 ;
        RECT 29.075 -3.565 29.405 -3.235 ;
        RECT 29.08 -3.565 29.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 129.945 30.765 131.075 ;
        RECT 30.435 125.635 30.765 125.965 ;
        RECT 30.435 124.275 30.765 124.605 ;
        RECT 30.44 123.6 30.76 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -0.845 30.765 -0.515 ;
        RECT 30.435 -2.205 30.765 -1.875 ;
        RECT 30.435 -3.565 30.765 -3.235 ;
        RECT 30.44 -3.565 30.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 129.945 32.125 131.075 ;
        RECT 31.795 125.635 32.125 125.965 ;
        RECT 31.795 124.275 32.125 124.605 ;
        RECT 31.8 123.6 32.12 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -0.845 32.125 -0.515 ;
        RECT 31.795 -2.205 32.125 -1.875 ;
        RECT 31.795 -3.565 32.125 -3.235 ;
        RECT 31.8 -3.565 32.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -151.805 32.125 -151.475 ;
        RECT 31.795 -153.165 32.125 -152.835 ;
        RECT 31.795 -154.525 32.125 -154.195 ;
        RECT 31.795 -155.885 32.125 -155.555 ;
        RECT 31.795 -157.245 32.125 -156.915 ;
        RECT 31.795 -162.89 32.125 -161.76 ;
        RECT 31.8 -163.005 32.12 -90.96 ;
        RECT 31.795 -91.965 32.125 -91.635 ;
        RECT 31.795 -93.325 32.125 -92.995 ;
        RECT 31.795 -94.685 32.125 -94.355 ;
        RECT 31.795 -96.045 32.125 -95.715 ;
        RECT 31.795 -97.405 32.125 -97.075 ;
        RECT 31.795 -98.765 32.125 -98.435 ;
        RECT 31.795 -100.125 32.125 -99.795 ;
        RECT 31.795 -101.485 32.125 -101.155 ;
        RECT 31.795 -102.845 32.125 -102.515 ;
        RECT 31.795 -104.205 32.125 -103.875 ;
        RECT 31.795 -105.565 32.125 -105.235 ;
        RECT 31.795 -106.925 32.125 -106.595 ;
        RECT 31.795 -108.285 32.125 -107.955 ;
        RECT 31.795 -109.645 32.125 -109.315 ;
        RECT 31.795 -111.005 32.125 -110.675 ;
        RECT 31.795 -112.365 32.125 -112.035 ;
        RECT 31.795 -113.725 32.125 -113.395 ;
        RECT 31.795 -115.085 32.125 -114.755 ;
        RECT 31.795 -116.445 32.125 -116.115 ;
        RECT 31.795 -117.805 32.125 -117.475 ;
        RECT 31.795 -119.165 32.125 -118.835 ;
        RECT 31.795 -120.525 32.125 -120.195 ;
        RECT 31.795 -121.885 32.125 -121.555 ;
        RECT 31.795 -123.245 32.125 -122.915 ;
        RECT 31.795 -124.605 32.125 -124.275 ;
        RECT 31.795 -125.965 32.125 -125.635 ;
        RECT 31.795 -127.325 32.125 -126.995 ;
        RECT 31.795 -128.685 32.125 -128.355 ;
        RECT 31.795 -130.045 32.125 -129.715 ;
        RECT 31.795 -131.405 32.125 -131.075 ;
        RECT 31.795 -132.765 32.125 -132.435 ;
        RECT 31.795 -134.125 32.125 -133.795 ;
        RECT 31.795 -135.485 32.125 -135.155 ;
        RECT 31.795 -136.845 32.125 -136.515 ;
        RECT 31.795 -138.205 32.125 -137.875 ;
        RECT 31.795 -139.565 32.125 -139.235 ;
        RECT 31.795 -140.925 32.125 -140.595 ;
        RECT 31.795 -142.285 32.125 -141.955 ;
        RECT 31.795 -143.645 32.125 -143.315 ;
        RECT 31.795 -145.005 32.125 -144.675 ;
        RECT 31.795 -146.365 32.125 -146.035 ;
        RECT 31.795 -147.725 32.125 -147.395 ;
        RECT 31.795 -149.085 32.125 -148.755 ;
        RECT 31.795 -150.445 32.125 -150.115 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 -154.525 -10.035 -154.195 ;
        RECT -10.365 -157.245 -10.035 -156.915 ;
        RECT -10.365 -162.89 -10.035 -161.76 ;
        RECT -10.36 -163.005 -10.04 -152.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 129.945 -8.675 131.075 ;
        RECT -9.005 125.635 -8.675 125.965 ;
        RECT -9.005 124.275 -8.675 124.605 ;
        RECT -9.005 122.915 -8.675 123.245 ;
        RECT -9.005 121.555 -8.675 121.885 ;
        RECT -9.005 120.195 -8.675 120.525 ;
        RECT -9.005 118.835 -8.675 119.165 ;
        RECT -9.005 117.475 -8.675 117.805 ;
        RECT -9.005 110.675 -8.675 111.005 ;
        RECT -9.005 107.955 -8.675 108.285 ;
        RECT -9.005 103.875 -8.675 104.205 ;
        RECT -9.005 99.795 -8.675 100.125 ;
        RECT -9.005 97.075 -8.675 97.405 ;
        RECT -9.005 90.275 -8.675 90.605 ;
        RECT -9.005 88.915 -8.675 89.245 ;
        RECT -9.005 82.115 -8.675 82.445 ;
        RECT -9.005 79.395 -8.675 79.725 ;
        RECT -9.005 75.315 -8.675 75.645 ;
        RECT -9.005 71.235 -8.675 71.565 ;
        RECT -9.005 68.515 -8.675 68.845 ;
        RECT -9.005 61.715 -8.675 62.045 ;
        RECT -9.005 60.355 -8.675 60.685 ;
        RECT -9.005 50.835 -8.675 51.165 ;
        RECT -9.005 46.755 -8.675 47.085 ;
        RECT -9.005 42.675 -8.675 43.005 ;
        RECT -9.005 39.955 -8.675 40.285 ;
        RECT -9.005 33.155 -8.675 33.485 ;
        RECT -9.005 31.795 -8.675 32.125 ;
        RECT -9.005 29.075 -8.675 29.405 ;
        RECT -9.005 22.275 -8.675 22.605 ;
        RECT -9.005 19.555 -8.675 19.885 ;
        RECT -9.005 18.195 -8.675 18.525 ;
        RECT -9.005 11.395 -8.675 11.725 ;
        RECT -9.005 4.595 -8.675 4.925 ;
        RECT -9.005 3.235 -8.675 3.565 ;
        RECT -9.005 1.875 -8.675 2.205 ;
        RECT -9.005 0.515 -8.675 0.845 ;
        RECT -9.005 -0.845 -8.675 -0.515 ;
        RECT -9.005 -2.205 -8.675 -1.875 ;
        RECT -9.005 -3.565 -8.675 -3.235 ;
        RECT -9.005 -4.925 -8.675 -4.595 ;
        RECT -9.005 -6.285 -8.675 -5.955 ;
        RECT -9.005 -7.645 -8.675 -7.315 ;
        RECT -9.005 -9.005 -8.675 -8.675 ;
        RECT -9.005 -10.365 -8.675 -10.035 ;
        RECT -9.005 -11.725 -8.675 -11.395 ;
        RECT -9.005 -13.085 -8.675 -12.755 ;
        RECT -9.005 -14.445 -8.675 -14.115 ;
        RECT -9.005 -15.805 -8.675 -15.475 ;
        RECT -9.005 -17.165 -8.675 -16.835 ;
        RECT -9 -19.88 -8.68 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 -82.445 -8.675 -82.115 ;
        RECT -9.005 -83.805 -8.675 -83.475 ;
        RECT -9.005 -85.165 -8.675 -84.835 ;
        RECT -9 -85.84 -8.68 -81.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 -138.205 -8.675 -137.875 ;
        RECT -9.005 -139.565 -8.675 -139.235 ;
        RECT -9.005 -140.925 -8.675 -140.595 ;
        RECT -9.005 -142.285 -8.675 -141.955 ;
        RECT -9.005 -143.645 -8.675 -143.315 ;
        RECT -9.005 -145.005 -8.675 -144.675 ;
        RECT -9.005 -146.365 -8.675 -146.035 ;
        RECT -9.005 -147.725 -8.675 -147.395 ;
        RECT -9.005 -149.085 -8.675 -148.755 ;
        RECT -9.005 -150.445 -8.675 -150.115 ;
        RECT -9.005 -151.805 -8.675 -151.475 ;
        RECT -9.005 -153.165 -8.675 -152.835 ;
        RECT -9.005 -154.525 -8.675 -154.195 ;
        RECT -9.005 -155.885 -8.675 -155.555 ;
        RECT -9.005 -157.245 -8.675 -156.915 ;
        RECT -9.005 -162.89 -8.675 -161.76 ;
        RECT -9 -163.005 -8.68 -137.875 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.645 129.945 -7.315 131.075 ;
        RECT -7.645 125.635 -7.315 125.965 ;
        RECT -7.645 124.275 -7.315 124.605 ;
        RECT -7.645 122.915 -7.315 123.245 ;
        RECT -7.645 121.555 -7.315 121.885 ;
        RECT -7.645 120.195 -7.315 120.525 ;
        RECT -7.645 118.835 -7.315 119.165 ;
        RECT -7.645 117.475 -7.315 117.805 ;
        RECT -7.645 110.675 -7.315 111.005 ;
        RECT -7.645 107.955 -7.315 108.285 ;
        RECT -7.645 103.875 -7.315 104.205 ;
        RECT -7.645 99.795 -7.315 100.125 ;
        RECT -7.645 97.075 -7.315 97.405 ;
        RECT -7.645 90.275 -7.315 90.605 ;
        RECT -7.645 88.915 -7.315 89.245 ;
        RECT -7.645 82.115 -7.315 82.445 ;
        RECT -7.645 79.395 -7.315 79.725 ;
        RECT -7.645 75.315 -7.315 75.645 ;
        RECT -7.645 71.235 -7.315 71.565 ;
        RECT -7.645 68.515 -7.315 68.845 ;
        RECT -7.645 61.715 -7.315 62.045 ;
        RECT -7.645 60.355 -7.315 60.685 ;
        RECT -7.645 50.835 -7.315 51.165 ;
        RECT -7.645 46.755 -7.315 47.085 ;
        RECT -7.645 42.675 -7.315 43.005 ;
        RECT -7.645 39.955 -7.315 40.285 ;
        RECT -7.645 33.155 -7.315 33.485 ;
        RECT -7.645 31.795 -7.315 32.125 ;
        RECT -7.645 29.075 -7.315 29.405 ;
        RECT -7.645 22.275 -7.315 22.605 ;
        RECT -7.645 19.555 -7.315 19.885 ;
        RECT -7.645 18.195 -7.315 18.525 ;
        RECT -7.645 11.395 -7.315 11.725 ;
        RECT -7.645 4.595 -7.315 4.925 ;
        RECT -7.645 3.235 -7.315 3.565 ;
        RECT -7.645 1.875 -7.315 2.205 ;
        RECT -7.645 0.515 -7.315 0.845 ;
        RECT -7.645 -0.845 -7.315 -0.515 ;
        RECT -7.645 -2.205 -7.315 -1.875 ;
        RECT -7.645 -3.565 -7.315 -3.235 ;
        RECT -7.645 -4.925 -7.315 -4.595 ;
        RECT -7.645 -6.285 -7.315 -5.955 ;
        RECT -7.645 -7.645 -7.315 -7.315 ;
        RECT -7.645 -9.005 -7.315 -8.675 ;
        RECT -7.645 -10.365 -7.315 -10.035 ;
        RECT -7.645 -11.725 -7.315 -11.395 ;
        RECT -7.645 -13.085 -7.315 -12.755 ;
        RECT -7.645 -14.445 -7.315 -14.115 ;
        RECT -7.645 -15.805 -7.315 -15.475 ;
        RECT -7.645 -17.165 -7.315 -16.835 ;
        RECT -7.645 -21.245 -7.315 -20.915 ;
        RECT -7.645 -22.605 -7.315 -22.275 ;
        RECT -7.645 -23.965 -7.315 -23.635 ;
        RECT -7.645 -25.325 -7.315 -24.995 ;
        RECT -7.645 -26.685 -7.315 -26.355 ;
        RECT -7.645 -28.045 -7.315 -27.715 ;
        RECT -7.645 -29.405 -7.315 -29.075 ;
        RECT -7.645 -30.765 -7.315 -30.435 ;
        RECT -7.645 -32.125 -7.315 -31.795 ;
        RECT -7.645 -33.485 -7.315 -33.155 ;
        RECT -7.645 -34.845 -7.315 -34.515 ;
        RECT -7.645 -36.205 -7.315 -35.875 ;
        RECT -7.645 -37.565 -7.315 -37.235 ;
        RECT -7.645 -38.925 -7.315 -38.595 ;
        RECT -7.645 -40.285 -7.315 -39.955 ;
        RECT -7.645 -41.645 -7.315 -41.315 ;
        RECT -7.645 -43.005 -7.315 -42.675 ;
        RECT -7.645 -44.365 -7.315 -44.035 ;
        RECT -7.645 -45.725 -7.315 -45.395 ;
        RECT -7.645 -49.805 -7.315 -49.475 ;
        RECT -7.645 -51.165 -7.315 -50.835 ;
        RECT -7.645 -52.525 -7.315 -52.195 ;
        RECT -7.645 -53.885 -7.315 -53.555 ;
        RECT -7.645 -55.245 -7.315 -54.915 ;
        RECT -7.645 -56.605 -7.315 -56.275 ;
        RECT -7.645 -57.965 -7.315 -57.635 ;
        RECT -7.645 -59.325 -7.315 -58.995 ;
        RECT -7.645 -60.685 -7.315 -60.355 ;
        RECT -7.645 -62.045 -7.315 -61.715 ;
        RECT -7.645 -63.405 -7.315 -63.075 ;
        RECT -7.645 -64.765 -7.315 -64.435 ;
        RECT -7.645 -66.125 -7.315 -65.795 ;
        RECT -7.645 -67.485 -7.315 -67.155 ;
        RECT -7.645 -68.845 -7.315 -68.515 ;
        RECT -7.645 -70.205 -7.315 -69.875 ;
        RECT -7.645 -71.565 -7.315 -71.235 ;
        RECT -7.645 -72.925 -7.315 -72.595 ;
        RECT -7.645 -74.285 -7.315 -73.955 ;
        RECT -7.645 -75.645 -7.315 -75.315 ;
        RECT -7.645 -77.005 -7.315 -76.675 ;
        RECT -7.645 -78.365 -7.315 -78.035 ;
        RECT -7.645 -79.725 -7.315 -79.395 ;
        RECT -7.645 -81.085 -7.315 -80.755 ;
        RECT -7.645 -82.445 -7.315 -82.115 ;
        RECT -7.645 -83.805 -7.315 -83.475 ;
        RECT -7.645 -85.165 -7.315 -84.835 ;
        RECT -7.645 -87.885 -7.315 -87.555 ;
        RECT -7.645 -89.245 -7.315 -88.915 ;
        RECT -7.645 -90.605 -7.315 -90.275 ;
        RECT -7.645 -91.965 -7.315 -91.635 ;
        RECT -7.645 -93.325 -7.315 -92.995 ;
        RECT -7.645 -94.685 -7.315 -94.355 ;
        RECT -7.645 -96.045 -7.315 -95.715 ;
        RECT -7.645 -97.405 -7.315 -97.075 ;
        RECT -7.645 -98.765 -7.315 -98.435 ;
        RECT -7.645 -100.125 -7.315 -99.795 ;
        RECT -7.645 -101.485 -7.315 -101.155 ;
        RECT -7.645 -102.845 -7.315 -102.515 ;
        RECT -7.645 -104.205 -7.315 -103.875 ;
        RECT -7.645 -105.565 -7.315 -105.235 ;
        RECT -7.645 -106.925 -7.315 -106.595 ;
        RECT -7.645 -108.285 -7.315 -107.955 ;
        RECT -7.645 -109.645 -7.315 -109.315 ;
        RECT -7.645 -111.005 -7.315 -110.675 ;
        RECT -7.645 -112.365 -7.315 -112.035 ;
        RECT -7.645 -113.725 -7.315 -113.395 ;
        RECT -7.645 -115.085 -7.315 -114.755 ;
        RECT -7.645 -116.445 -7.315 -116.115 ;
        RECT -7.645 -117.805 -7.315 -117.475 ;
        RECT -7.645 -119.165 -7.315 -118.835 ;
        RECT -7.645 -120.525 -7.315 -120.195 ;
        RECT -7.645 -121.885 -7.315 -121.555 ;
        RECT -7.645 -123.245 -7.315 -122.915 ;
        RECT -7.645 -124.605 -7.315 -124.275 ;
        RECT -7.645 -125.965 -7.315 -125.635 ;
        RECT -7.645 -127.325 -7.315 -126.995 ;
        RECT -7.645 -128.685 -7.315 -128.355 ;
        RECT -7.645 -130.045 -7.315 -129.715 ;
        RECT -7.645 -131.405 -7.315 -131.075 ;
        RECT -7.645 -132.765 -7.315 -132.435 ;
        RECT -7.645 -134.125 -7.315 -133.795 ;
        RECT -7.645 -135.485 -7.315 -135.155 ;
        RECT -7.645 -136.845 -7.315 -136.515 ;
        RECT -7.645 -138.205 -7.315 -137.875 ;
        RECT -7.645 -139.565 -7.315 -139.235 ;
        RECT -7.645 -140.925 -7.315 -140.595 ;
        RECT -7.645 -142.285 -7.315 -141.955 ;
        RECT -7.645 -143.645 -7.315 -143.315 ;
        RECT -7.645 -145.005 -7.315 -144.675 ;
        RECT -7.645 -146.365 -7.315 -146.035 ;
        RECT -7.645 -147.725 -7.315 -147.395 ;
        RECT -7.645 -149.085 -7.315 -148.755 ;
        RECT -7.645 -150.445 -7.315 -150.115 ;
        RECT -7.645 -151.805 -7.315 -151.475 ;
        RECT -7.645 -153.165 -7.315 -152.835 ;
        RECT -7.645 -154.525 -7.315 -154.195 ;
        RECT -7.645 -155.885 -7.315 -155.555 ;
        RECT -7.645 -157.245 -7.315 -156.915 ;
        RECT -7.645 -162.89 -7.315 -161.76 ;
        RECT -7.64 -163.005 -7.32 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.285 129.945 -5.955 131.075 ;
        RECT -6.285 125.635 -5.955 125.965 ;
        RECT -6.285 124.275 -5.955 124.605 ;
        RECT -6.285 -0.845 -5.955 -0.515 ;
        RECT -6.285 -2.205 -5.955 -1.875 ;
        RECT -6.285 -3.565 -5.955 -3.235 ;
        RECT -6.285 -4.925 -5.955 -4.595 ;
        RECT -6.285 -6.285 -5.955 -5.955 ;
        RECT -6.285 -7.645 -5.955 -7.315 ;
        RECT -6.285 -9.005 -5.955 -8.675 ;
        RECT -6.285 -10.365 -5.955 -10.035 ;
        RECT -6.285 -11.725 -5.955 -11.395 ;
        RECT -6.285 -13.085 -5.955 -12.755 ;
        RECT -6.285 -14.445 -5.955 -14.115 ;
        RECT -6.285 -15.805 -5.955 -15.475 ;
        RECT -6.285 -17.165 -5.955 -16.835 ;
        RECT -6.285 -21.245 -5.955 -20.915 ;
        RECT -6.285 -22.605 -5.955 -22.275 ;
        RECT -6.285 -23.965 -5.955 -23.635 ;
        RECT -6.285 -25.325 -5.955 -24.995 ;
        RECT -6.285 -26.685 -5.955 -26.355 ;
        RECT -6.285 -28.045 -5.955 -27.715 ;
        RECT -6.285 -29.405 -5.955 -29.075 ;
        RECT -6.285 -30.765 -5.955 -30.435 ;
        RECT -6.285 -32.125 -5.955 -31.795 ;
        RECT -6.285 -33.485 -5.955 -33.155 ;
        RECT -6.285 -34.845 -5.955 -34.515 ;
        RECT -6.285 -36.205 -5.955 -35.875 ;
        RECT -6.285 -37.565 -5.955 -37.235 ;
        RECT -6.285 -38.925 -5.955 -38.595 ;
        RECT -6.285 -40.285 -5.955 -39.955 ;
        RECT -6.285 -41.645 -5.955 -41.315 ;
        RECT -6.285 -43.005 -5.955 -42.675 ;
        RECT -6.285 -44.365 -5.955 -44.035 ;
        RECT -6.285 -45.725 -5.955 -45.395 ;
        RECT -6.285 -49.805 -5.955 -49.475 ;
        RECT -6.285 -51.165 -5.955 -50.835 ;
        RECT -6.285 -52.525 -5.955 -52.195 ;
        RECT -6.285 -53.885 -5.955 -53.555 ;
        RECT -6.285 -55.245 -5.955 -54.915 ;
        RECT -6.285 -56.605 -5.955 -56.275 ;
        RECT -6.285 -57.965 -5.955 -57.635 ;
        RECT -6.285 -59.325 -5.955 -58.995 ;
        RECT -6.285 -60.685 -5.955 -60.355 ;
        RECT -6.285 -62.045 -5.955 -61.715 ;
        RECT -6.285 -63.405 -5.955 -63.075 ;
        RECT -6.285 -64.765 -5.955 -64.435 ;
        RECT -6.285 -66.125 -5.955 -65.795 ;
        RECT -6.285 -67.485 -5.955 -67.155 ;
        RECT -6.285 -68.845 -5.955 -68.515 ;
        RECT -6.285 -70.205 -5.955 -69.875 ;
        RECT -6.285 -71.565 -5.955 -71.235 ;
        RECT -6.285 -72.925 -5.955 -72.595 ;
        RECT -6.285 -74.285 -5.955 -73.955 ;
        RECT -6.285 -75.645 -5.955 -75.315 ;
        RECT -6.285 -77.005 -5.955 -76.675 ;
        RECT -6.285 -78.365 -5.955 -78.035 ;
        RECT -6.285 -79.725 -5.955 -79.395 ;
        RECT -6.285 -81.085 -5.955 -80.755 ;
        RECT -6.285 -82.445 -5.955 -82.115 ;
        RECT -6.285 -83.805 -5.955 -83.475 ;
        RECT -6.285 -85.165 -5.955 -84.835 ;
        RECT -6.285 -87.885 -5.955 -87.555 ;
        RECT -6.285 -89.245 -5.955 -88.915 ;
        RECT -6.285 -90.605 -5.955 -90.275 ;
        RECT -6.285 -91.965 -5.955 -91.635 ;
        RECT -6.285 -93.325 -5.955 -92.995 ;
        RECT -6.285 -94.685 -5.955 -94.355 ;
        RECT -6.285 -96.045 -5.955 -95.715 ;
        RECT -6.285 -97.405 -5.955 -97.075 ;
        RECT -6.285 -98.765 -5.955 -98.435 ;
        RECT -6.285 -100.125 -5.955 -99.795 ;
        RECT -6.285 -101.485 -5.955 -101.155 ;
        RECT -6.285 -102.845 -5.955 -102.515 ;
        RECT -6.285 -104.205 -5.955 -103.875 ;
        RECT -6.285 -105.565 -5.955 -105.235 ;
        RECT -6.285 -106.925 -5.955 -106.595 ;
        RECT -6.285 -108.285 -5.955 -107.955 ;
        RECT -6.285 -109.645 -5.955 -109.315 ;
        RECT -6.285 -111.005 -5.955 -110.675 ;
        RECT -6.285 -112.365 -5.955 -112.035 ;
        RECT -6.285 -113.725 -5.955 -113.395 ;
        RECT -6.285 -115.085 -5.955 -114.755 ;
        RECT -6.285 -116.445 -5.955 -116.115 ;
        RECT -6.285 -117.805 -5.955 -117.475 ;
        RECT -6.285 -119.165 -5.955 -118.835 ;
        RECT -6.285 -120.525 -5.955 -120.195 ;
        RECT -6.285 -121.885 -5.955 -121.555 ;
        RECT -6.285 -123.245 -5.955 -122.915 ;
        RECT -6.285 -124.605 -5.955 -124.275 ;
        RECT -6.285 -125.965 -5.955 -125.635 ;
        RECT -6.285 -127.325 -5.955 -126.995 ;
        RECT -6.285 -128.685 -5.955 -128.355 ;
        RECT -6.285 -130.045 -5.955 -129.715 ;
        RECT -6.285 -131.405 -5.955 -131.075 ;
        RECT -6.285 -132.765 -5.955 -132.435 ;
        RECT -6.285 -134.125 -5.955 -133.795 ;
        RECT -6.285 -135.485 -5.955 -135.155 ;
        RECT -6.285 -136.845 -5.955 -136.515 ;
        RECT -6.285 -138.205 -5.955 -137.875 ;
        RECT -6.285 -139.565 -5.955 -139.235 ;
        RECT -6.285 -140.925 -5.955 -140.595 ;
        RECT -6.285 -142.285 -5.955 -141.955 ;
        RECT -6.285 -143.645 -5.955 -143.315 ;
        RECT -6.285 -145.005 -5.955 -144.675 ;
        RECT -6.285 -146.365 -5.955 -146.035 ;
        RECT -6.285 -147.725 -5.955 -147.395 ;
        RECT -6.285 -149.085 -5.955 -148.755 ;
        RECT -6.285 -150.445 -5.955 -150.115 ;
        RECT -6.285 -151.805 -5.955 -151.475 ;
        RECT -6.285 -153.165 -5.955 -152.835 ;
        RECT -6.285 -154.525 -5.955 -154.195 ;
        RECT -6.285 -155.885 -5.955 -155.555 ;
        RECT -6.285 -157.245 -5.955 -156.915 ;
        RECT -6.285 -162.89 -5.955 -161.76 ;
        RECT -6.28 -163.005 -5.96 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.925 129.945 -4.595 131.075 ;
        RECT -4.925 125.635 -4.595 125.965 ;
        RECT -4.925 124.275 -4.595 124.605 ;
        RECT -4.925 121.41 -4.595 121.74 ;
        RECT -4.925 119.235 -4.595 119.565 ;
        RECT -4.925 117.655 -4.595 117.985 ;
        RECT -4.925 116.805 -4.595 117.135 ;
        RECT -4.925 114.495 -4.595 114.825 ;
        RECT -4.925 113.645 -4.595 113.975 ;
        RECT -4.925 111.335 -4.595 111.665 ;
        RECT -4.925 110.485 -4.595 110.815 ;
        RECT -4.925 108.175 -4.595 108.505 ;
        RECT -4.925 107.325 -4.595 107.655 ;
        RECT -4.925 105.015 -4.595 105.345 ;
        RECT -4.925 103.435 -4.595 103.765 ;
        RECT -4.925 102.585 -4.595 102.915 ;
        RECT -4.925 100.275 -4.595 100.605 ;
        RECT -4.925 99.425 -4.595 99.755 ;
        RECT -4.925 97.115 -4.595 97.445 ;
        RECT -4.925 96.265 -4.595 96.595 ;
        RECT -4.925 93.955 -4.595 94.285 ;
        RECT -4.925 93.105 -4.595 93.435 ;
        RECT -4.925 90.795 -4.595 91.125 ;
        RECT -4.925 89.215 -4.595 89.545 ;
        RECT -4.925 88.365 -4.595 88.695 ;
        RECT -4.925 86.055 -4.595 86.385 ;
        RECT -4.925 85.205 -4.595 85.535 ;
        RECT -4.925 82.895 -4.595 83.225 ;
        RECT -4.925 82.045 -4.595 82.375 ;
        RECT -4.925 79.735 -4.595 80.065 ;
        RECT -4.925 78.885 -4.595 79.215 ;
        RECT -4.925 76.575 -4.595 76.905 ;
        RECT -4.925 74.995 -4.595 75.325 ;
        RECT -4.925 74.145 -4.595 74.475 ;
        RECT -4.925 71.835 -4.595 72.165 ;
        RECT -4.925 70.985 -4.595 71.315 ;
        RECT -4.925 68.675 -4.595 69.005 ;
        RECT -4.925 67.825 -4.595 68.155 ;
        RECT -4.925 65.515 -4.595 65.845 ;
        RECT -4.925 64.665 -4.595 64.995 ;
        RECT -4.925 62.355 -4.595 62.685 ;
        RECT -4.925 60.775 -4.595 61.105 ;
        RECT -4.925 59.925 -4.595 60.255 ;
        RECT -4.925 57.615 -4.595 57.945 ;
        RECT -4.925 56.765 -4.595 57.095 ;
        RECT -4.925 54.455 -4.595 54.785 ;
        RECT -4.925 53.605 -4.595 53.935 ;
        RECT -4.925 51.295 -4.595 51.625 ;
        RECT -4.925 50.445 -4.595 50.775 ;
        RECT -4.925 48.135 -4.595 48.465 ;
        RECT -4.925 46.555 -4.595 46.885 ;
        RECT -4.925 45.705 -4.595 46.035 ;
        RECT -4.925 43.395 -4.595 43.725 ;
        RECT -4.925 42.545 -4.595 42.875 ;
        RECT -4.925 40.235 -4.595 40.565 ;
        RECT -4.925 39.385 -4.595 39.715 ;
        RECT -4.925 37.075 -4.595 37.405 ;
        RECT -4.925 36.225 -4.595 36.555 ;
        RECT -4.925 33.915 -4.595 34.245 ;
        RECT -4.925 32.335 -4.595 32.665 ;
        RECT -4.925 31.485 -4.595 31.815 ;
        RECT -4.925 29.175 -4.595 29.505 ;
        RECT -4.925 28.325 -4.595 28.655 ;
        RECT -4.925 26.015 -4.595 26.345 ;
        RECT -4.925 25.165 -4.595 25.495 ;
        RECT -4.925 22.855 -4.595 23.185 ;
        RECT -4.925 22.005 -4.595 22.335 ;
        RECT -4.925 19.695 -4.595 20.025 ;
        RECT -4.925 18.115 -4.595 18.445 ;
        RECT -4.925 17.265 -4.595 17.595 ;
        RECT -4.925 14.955 -4.595 15.285 ;
        RECT -4.925 14.105 -4.595 14.435 ;
        RECT -4.925 11.795 -4.595 12.125 ;
        RECT -4.925 10.945 -4.595 11.275 ;
        RECT -4.925 8.635 -4.595 8.965 ;
        RECT -4.925 7.785 -4.595 8.115 ;
        RECT -4.925 5.475 -4.595 5.805 ;
        RECT -4.925 3.895 -4.595 4.225 ;
        RECT -4.925 3.045 -4.595 3.375 ;
        RECT -4.925 0.87 -4.595 1.2 ;
        RECT -4.925 -0.845 -4.595 -0.515 ;
        RECT -4.925 -2.205 -4.595 -1.875 ;
        RECT -4.925 -3.565 -4.595 -3.235 ;
        RECT -4.925 -4.925 -4.595 -4.595 ;
        RECT -4.925 -6.285 -4.595 -5.955 ;
        RECT -4.925 -7.645 -4.595 -7.315 ;
        RECT -4.925 -9.005 -4.595 -8.675 ;
        RECT -4.925 -10.365 -4.595 -10.035 ;
        RECT -4.925 -11.725 -4.595 -11.395 ;
        RECT -4.925 -13.085 -4.595 -12.755 ;
        RECT -4.925 -14.445 -4.595 -14.115 ;
        RECT -4.925 -15.805 -4.595 -15.475 ;
        RECT -4.925 -17.165 -4.595 -16.835 ;
        RECT -4.925 -21.245 -4.595 -20.915 ;
        RECT -4.925 -22.605 -4.595 -22.275 ;
        RECT -4.925 -23.965 -4.595 -23.635 ;
        RECT -4.925 -25.325 -4.595 -24.995 ;
        RECT -4.925 -26.685 -4.595 -26.355 ;
        RECT -4.925 -28.045 -4.595 -27.715 ;
        RECT -4.925 -29.405 -4.595 -29.075 ;
        RECT -4.925 -30.765 -4.595 -30.435 ;
        RECT -4.925 -32.125 -4.595 -31.795 ;
        RECT -4.925 -33.485 -4.595 -33.155 ;
        RECT -4.925 -34.845 -4.595 -34.515 ;
        RECT -4.925 -36.205 -4.595 -35.875 ;
        RECT -4.925 -37.565 -4.595 -37.235 ;
        RECT -4.925 -38.925 -4.595 -38.595 ;
        RECT -4.925 -40.285 -4.595 -39.955 ;
        RECT -4.925 -41.645 -4.595 -41.315 ;
        RECT -4.925 -43.005 -4.595 -42.675 ;
        RECT -4.925 -44.365 -4.595 -44.035 ;
        RECT -4.925 -45.725 -4.595 -45.395 ;
        RECT -4.925 -49.805 -4.595 -49.475 ;
        RECT -4.925 -51.165 -4.595 -50.835 ;
        RECT -4.925 -52.525 -4.595 -52.195 ;
        RECT -4.925 -53.885 -4.595 -53.555 ;
        RECT -4.925 -55.245 -4.595 -54.915 ;
        RECT -4.925 -56.605 -4.595 -56.275 ;
        RECT -4.925 -57.965 -4.595 -57.635 ;
        RECT -4.925 -59.325 -4.595 -58.995 ;
        RECT -4.925 -60.685 -4.595 -60.355 ;
        RECT -4.925 -62.045 -4.595 -61.715 ;
        RECT -4.925 -63.405 -4.595 -63.075 ;
        RECT -4.925 -64.765 -4.595 -64.435 ;
        RECT -4.925 -66.125 -4.595 -65.795 ;
        RECT -4.925 -67.485 -4.595 -67.155 ;
        RECT -4.925 -68.845 -4.595 -68.515 ;
        RECT -4.925 -70.205 -4.595 -69.875 ;
        RECT -4.925 -71.565 -4.595 -71.235 ;
        RECT -4.925 -72.925 -4.595 -72.595 ;
        RECT -4.925 -74.285 -4.595 -73.955 ;
        RECT -4.925 -75.645 -4.595 -75.315 ;
        RECT -4.925 -77.005 -4.595 -76.675 ;
        RECT -4.925 -78.365 -4.595 -78.035 ;
        RECT -4.925 -79.725 -4.595 -79.395 ;
        RECT -4.925 -81.085 -4.595 -80.755 ;
        RECT -4.925 -82.445 -4.595 -82.115 ;
        RECT -4.925 -83.805 -4.595 -83.475 ;
        RECT -4.925 -85.165 -4.595 -84.835 ;
        RECT -4.925 -87.885 -4.595 -87.555 ;
        RECT -4.925 -89.245 -4.595 -88.915 ;
        RECT -4.925 -90.605 -4.595 -90.275 ;
        RECT -4.925 -91.965 -4.595 -91.635 ;
        RECT -4.925 -93.325 -4.595 -92.995 ;
        RECT -4.925 -94.685 -4.595 -94.355 ;
        RECT -4.925 -96.045 -4.595 -95.715 ;
        RECT -4.925 -97.405 -4.595 -97.075 ;
        RECT -4.925 -98.765 -4.595 -98.435 ;
        RECT -4.925 -100.125 -4.595 -99.795 ;
        RECT -4.925 -101.485 -4.595 -101.155 ;
        RECT -4.925 -102.845 -4.595 -102.515 ;
        RECT -4.925 -104.205 -4.595 -103.875 ;
        RECT -4.925 -105.565 -4.595 -105.235 ;
        RECT -4.925 -106.925 -4.595 -106.595 ;
        RECT -4.925 -108.285 -4.595 -107.955 ;
        RECT -4.925 -109.645 -4.595 -109.315 ;
        RECT -4.925 -111.005 -4.595 -110.675 ;
        RECT -4.925 -112.365 -4.595 -112.035 ;
        RECT -4.925 -113.725 -4.595 -113.395 ;
        RECT -4.925 -115.085 -4.595 -114.755 ;
        RECT -4.925 -116.445 -4.595 -116.115 ;
        RECT -4.925 -117.805 -4.595 -117.475 ;
        RECT -4.925 -119.165 -4.595 -118.835 ;
        RECT -4.925 -120.525 -4.595 -120.195 ;
        RECT -4.925 -121.885 -4.595 -121.555 ;
        RECT -4.925 -123.245 -4.595 -122.915 ;
        RECT -4.925 -124.605 -4.595 -124.275 ;
        RECT -4.925 -125.965 -4.595 -125.635 ;
        RECT -4.925 -127.325 -4.595 -126.995 ;
        RECT -4.925 -128.685 -4.595 -128.355 ;
        RECT -4.925 -130.045 -4.595 -129.715 ;
        RECT -4.925 -131.405 -4.595 -131.075 ;
        RECT -4.925 -132.765 -4.595 -132.435 ;
        RECT -4.925 -134.125 -4.595 -133.795 ;
        RECT -4.925 -135.485 -4.595 -135.155 ;
        RECT -4.925 -136.845 -4.595 -136.515 ;
        RECT -4.925 -138.205 -4.595 -137.875 ;
        RECT -4.925 -139.565 -4.595 -139.235 ;
        RECT -4.925 -140.925 -4.595 -140.595 ;
        RECT -4.925 -142.285 -4.595 -141.955 ;
        RECT -4.925 -143.645 -4.595 -143.315 ;
        RECT -4.925 -145.005 -4.595 -144.675 ;
        RECT -4.925 -146.365 -4.595 -146.035 ;
        RECT -4.925 -147.725 -4.595 -147.395 ;
        RECT -4.925 -149.085 -4.595 -148.755 ;
        RECT -4.925 -150.445 -4.595 -150.115 ;
        RECT -4.925 -151.805 -4.595 -151.475 ;
        RECT -4.925 -153.165 -4.595 -152.835 ;
        RECT -4.925 -154.525 -4.595 -154.195 ;
        RECT -4.925 -155.885 -4.595 -155.555 ;
        RECT -4.925 -157.245 -4.595 -156.915 ;
        RECT -4.925 -162.89 -4.595 -161.76 ;
        RECT -4.92 -163.005 -4.6 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.565 129.945 -3.235 131.075 ;
        RECT -3.565 125.635 -3.235 125.965 ;
        RECT -3.565 124.275 -3.235 124.605 ;
        RECT -3.565 121.41 -3.235 121.74 ;
        RECT -3.565 119.235 -3.235 119.565 ;
        RECT -3.565 117.655 -3.235 117.985 ;
        RECT -3.565 116.805 -3.235 117.135 ;
        RECT -3.565 114.495 -3.235 114.825 ;
        RECT -3.565 113.645 -3.235 113.975 ;
        RECT -3.565 111.335 -3.235 111.665 ;
        RECT -3.565 110.485 -3.235 110.815 ;
        RECT -3.565 108.175 -3.235 108.505 ;
        RECT -3.565 107.325 -3.235 107.655 ;
        RECT -3.565 105.015 -3.235 105.345 ;
        RECT -3.565 103.435 -3.235 103.765 ;
        RECT -3.565 102.585 -3.235 102.915 ;
        RECT -3.565 100.275 -3.235 100.605 ;
        RECT -3.565 99.425 -3.235 99.755 ;
        RECT -3.565 97.115 -3.235 97.445 ;
        RECT -3.565 96.265 -3.235 96.595 ;
        RECT -3.565 93.955 -3.235 94.285 ;
        RECT -3.565 93.105 -3.235 93.435 ;
        RECT -3.565 90.795 -3.235 91.125 ;
        RECT -3.565 89.215 -3.235 89.545 ;
        RECT -3.565 88.365 -3.235 88.695 ;
        RECT -3.565 86.055 -3.235 86.385 ;
        RECT -3.565 85.205 -3.235 85.535 ;
        RECT -3.565 82.895 -3.235 83.225 ;
        RECT -3.565 82.045 -3.235 82.375 ;
        RECT -3.565 79.735 -3.235 80.065 ;
        RECT -3.565 78.885 -3.235 79.215 ;
        RECT -3.565 76.575 -3.235 76.905 ;
        RECT -3.565 74.995 -3.235 75.325 ;
        RECT -3.565 74.145 -3.235 74.475 ;
        RECT -3.565 71.835 -3.235 72.165 ;
        RECT -3.565 70.985 -3.235 71.315 ;
        RECT -3.565 68.675 -3.235 69.005 ;
        RECT -3.565 67.825 -3.235 68.155 ;
        RECT -3.565 65.515 -3.235 65.845 ;
        RECT -3.565 64.665 -3.235 64.995 ;
        RECT -3.565 62.355 -3.235 62.685 ;
        RECT -3.565 60.775 -3.235 61.105 ;
        RECT -3.565 59.925 -3.235 60.255 ;
        RECT -3.565 57.615 -3.235 57.945 ;
        RECT -3.565 56.765 -3.235 57.095 ;
        RECT -3.565 54.455 -3.235 54.785 ;
        RECT -3.565 53.605 -3.235 53.935 ;
        RECT -3.565 51.295 -3.235 51.625 ;
        RECT -3.565 50.445 -3.235 50.775 ;
        RECT -3.565 48.135 -3.235 48.465 ;
        RECT -3.565 46.555 -3.235 46.885 ;
        RECT -3.565 45.705 -3.235 46.035 ;
        RECT -3.565 43.395 -3.235 43.725 ;
        RECT -3.565 42.545 -3.235 42.875 ;
        RECT -3.565 40.235 -3.235 40.565 ;
        RECT -3.565 39.385 -3.235 39.715 ;
        RECT -3.565 37.075 -3.235 37.405 ;
        RECT -3.565 36.225 -3.235 36.555 ;
        RECT -3.565 33.915 -3.235 34.245 ;
        RECT -3.565 32.335 -3.235 32.665 ;
        RECT -3.565 31.485 -3.235 31.815 ;
        RECT -3.565 29.175 -3.235 29.505 ;
        RECT -3.565 28.325 -3.235 28.655 ;
        RECT -3.565 26.015 -3.235 26.345 ;
        RECT -3.565 25.165 -3.235 25.495 ;
        RECT -3.565 22.855 -3.235 23.185 ;
        RECT -3.565 22.005 -3.235 22.335 ;
        RECT -3.565 19.695 -3.235 20.025 ;
        RECT -3.565 18.115 -3.235 18.445 ;
        RECT -3.565 17.265 -3.235 17.595 ;
        RECT -3.565 14.955 -3.235 15.285 ;
        RECT -3.565 14.105 -3.235 14.435 ;
        RECT -3.565 11.795 -3.235 12.125 ;
        RECT -3.565 10.945 -3.235 11.275 ;
        RECT -3.565 8.635 -3.235 8.965 ;
        RECT -3.565 7.785 -3.235 8.115 ;
        RECT -3.565 5.475 -3.235 5.805 ;
        RECT -3.565 3.895 -3.235 4.225 ;
        RECT -3.565 3.045 -3.235 3.375 ;
        RECT -3.565 0.87 -3.235 1.2 ;
        RECT -3.565 -0.845 -3.235 -0.515 ;
        RECT -3.565 -2.205 -3.235 -1.875 ;
        RECT -3.565 -3.565 -3.235 -3.235 ;
        RECT -3.565 -4.925 -3.235 -4.595 ;
        RECT -3.565 -6.285 -3.235 -5.955 ;
        RECT -3.565 -7.645 -3.235 -7.315 ;
        RECT -3.565 -9.005 -3.235 -8.675 ;
        RECT -3.565 -10.365 -3.235 -10.035 ;
        RECT -3.565 -11.725 -3.235 -11.395 ;
        RECT -3.565 -13.085 -3.235 -12.755 ;
        RECT -3.565 -14.445 -3.235 -14.115 ;
        RECT -3.565 -15.805 -3.235 -15.475 ;
        RECT -3.565 -17.165 -3.235 -16.835 ;
        RECT -3.565 -21.245 -3.235 -20.915 ;
        RECT -3.565 -22.605 -3.235 -22.275 ;
        RECT -3.565 -23.965 -3.235 -23.635 ;
        RECT -3.565 -25.325 -3.235 -24.995 ;
        RECT -3.565 -26.685 -3.235 -26.355 ;
        RECT -3.565 -28.045 -3.235 -27.715 ;
        RECT -3.565 -29.405 -3.235 -29.075 ;
        RECT -3.565 -30.765 -3.235 -30.435 ;
        RECT -3.565 -32.125 -3.235 -31.795 ;
        RECT -3.565 -33.485 -3.235 -33.155 ;
        RECT -3.565 -34.845 -3.235 -34.515 ;
        RECT -3.565 -36.205 -3.235 -35.875 ;
        RECT -3.565 -37.565 -3.235 -37.235 ;
        RECT -3.565 -38.925 -3.235 -38.595 ;
        RECT -3.565 -40.285 -3.235 -39.955 ;
        RECT -3.565 -41.645 -3.235 -41.315 ;
        RECT -3.565 -43.005 -3.235 -42.675 ;
        RECT -3.565 -44.365 -3.235 -44.035 ;
        RECT -3.565 -45.725 -3.235 -45.395 ;
        RECT -3.565 -49.805 -3.235 -49.475 ;
        RECT -3.565 -51.165 -3.235 -50.835 ;
        RECT -3.565 -52.525 -3.235 -52.195 ;
        RECT -3.565 -53.885 -3.235 -53.555 ;
        RECT -3.565 -55.245 -3.235 -54.915 ;
        RECT -3.565 -56.605 -3.235 -56.275 ;
        RECT -3.565 -57.965 -3.235 -57.635 ;
        RECT -3.565 -59.325 -3.235 -58.995 ;
        RECT -3.565 -60.685 -3.235 -60.355 ;
        RECT -3.565 -62.045 -3.235 -61.715 ;
        RECT -3.565 -63.405 -3.235 -63.075 ;
        RECT -3.565 -64.765 -3.235 -64.435 ;
        RECT -3.565 -66.125 -3.235 -65.795 ;
        RECT -3.565 -67.485 -3.235 -67.155 ;
        RECT -3.565 -68.845 -3.235 -68.515 ;
        RECT -3.565 -70.205 -3.235 -69.875 ;
        RECT -3.565 -71.565 -3.235 -71.235 ;
        RECT -3.565 -72.925 -3.235 -72.595 ;
        RECT -3.565 -74.285 -3.235 -73.955 ;
        RECT -3.565 -75.645 -3.235 -75.315 ;
        RECT -3.565 -77.005 -3.235 -76.675 ;
        RECT -3.565 -78.365 -3.235 -78.035 ;
        RECT -3.565 -79.725 -3.235 -79.395 ;
        RECT -3.565 -81.085 -3.235 -80.755 ;
        RECT -3.565 -82.445 -3.235 -82.115 ;
        RECT -3.565 -83.805 -3.235 -83.475 ;
        RECT -3.565 -85.165 -3.235 -84.835 ;
        RECT -3.565 -87.885 -3.235 -87.555 ;
        RECT -3.565 -89.245 -3.235 -88.915 ;
        RECT -3.565 -90.605 -3.235 -90.275 ;
        RECT -3.565 -91.965 -3.235 -91.635 ;
        RECT -3.565 -93.325 -3.235 -92.995 ;
        RECT -3.565 -94.685 -3.235 -94.355 ;
        RECT -3.565 -96.045 -3.235 -95.715 ;
        RECT -3.565 -97.405 -3.235 -97.075 ;
        RECT -3.565 -98.765 -3.235 -98.435 ;
        RECT -3.565 -100.125 -3.235 -99.795 ;
        RECT -3.565 -101.485 -3.235 -101.155 ;
        RECT -3.565 -102.845 -3.235 -102.515 ;
        RECT -3.565 -104.205 -3.235 -103.875 ;
        RECT -3.565 -105.565 -3.235 -105.235 ;
        RECT -3.565 -106.925 -3.235 -106.595 ;
        RECT -3.565 -108.285 -3.235 -107.955 ;
        RECT -3.565 -109.645 -3.235 -109.315 ;
        RECT -3.565 -111.005 -3.235 -110.675 ;
        RECT -3.565 -112.365 -3.235 -112.035 ;
        RECT -3.565 -113.725 -3.235 -113.395 ;
        RECT -3.565 -115.085 -3.235 -114.755 ;
        RECT -3.565 -116.445 -3.235 -116.115 ;
        RECT -3.565 -117.805 -3.235 -117.475 ;
        RECT -3.565 -119.165 -3.235 -118.835 ;
        RECT -3.565 -120.525 -3.235 -120.195 ;
        RECT -3.565 -121.885 -3.235 -121.555 ;
        RECT -3.565 -123.245 -3.235 -122.915 ;
        RECT -3.565 -124.605 -3.235 -124.275 ;
        RECT -3.565 -125.965 -3.235 -125.635 ;
        RECT -3.565 -127.325 -3.235 -126.995 ;
        RECT -3.565 -128.685 -3.235 -128.355 ;
        RECT -3.565 -130.045 -3.235 -129.715 ;
        RECT -3.565 -131.405 -3.235 -131.075 ;
        RECT -3.565 -132.765 -3.235 -132.435 ;
        RECT -3.565 -134.125 -3.235 -133.795 ;
        RECT -3.565 -135.485 -3.235 -135.155 ;
        RECT -3.565 -136.845 -3.235 -136.515 ;
        RECT -3.565 -138.205 -3.235 -137.875 ;
        RECT -3.565 -139.565 -3.235 -139.235 ;
        RECT -3.565 -140.925 -3.235 -140.595 ;
        RECT -3.565 -142.285 -3.235 -141.955 ;
        RECT -3.565 -143.645 -3.235 -143.315 ;
        RECT -3.565 -145.005 -3.235 -144.675 ;
        RECT -3.565 -146.365 -3.235 -146.035 ;
        RECT -3.565 -147.725 -3.235 -147.395 ;
        RECT -3.565 -149.085 -3.235 -148.755 ;
        RECT -3.565 -150.445 -3.235 -150.115 ;
        RECT -3.565 -151.805 -3.235 -151.475 ;
        RECT -3.565 -153.165 -3.235 -152.835 ;
        RECT -3.565 -154.525 -3.235 -154.195 ;
        RECT -3.565 -155.885 -3.235 -155.555 ;
        RECT -3.565 -157.245 -3.235 -156.915 ;
        RECT -3.565 -162.89 -3.235 -161.76 ;
        RECT -3.56 -163.005 -3.24 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 129.945 -1.875 131.075 ;
        RECT -2.205 125.635 -1.875 125.965 ;
        RECT -2.205 124.275 -1.875 124.605 ;
        RECT -2.205 121.41 -1.875 121.74 ;
        RECT -2.205 119.235 -1.875 119.565 ;
        RECT -2.205 117.655 -1.875 117.985 ;
        RECT -2.205 116.805 -1.875 117.135 ;
        RECT -2.205 114.495 -1.875 114.825 ;
        RECT -2.205 113.645 -1.875 113.975 ;
        RECT -2.205 111.335 -1.875 111.665 ;
        RECT -2.205 110.485 -1.875 110.815 ;
        RECT -2.205 108.175 -1.875 108.505 ;
        RECT -2.205 107.325 -1.875 107.655 ;
        RECT -2.205 105.015 -1.875 105.345 ;
        RECT -2.205 103.435 -1.875 103.765 ;
        RECT -2.205 102.585 -1.875 102.915 ;
        RECT -2.205 100.275 -1.875 100.605 ;
        RECT -2.205 99.425 -1.875 99.755 ;
        RECT -2.205 97.115 -1.875 97.445 ;
        RECT -2.205 96.265 -1.875 96.595 ;
        RECT -2.205 93.955 -1.875 94.285 ;
        RECT -2.205 93.105 -1.875 93.435 ;
        RECT -2.205 90.795 -1.875 91.125 ;
        RECT -2.205 89.215 -1.875 89.545 ;
        RECT -2.205 88.365 -1.875 88.695 ;
        RECT -2.205 86.055 -1.875 86.385 ;
        RECT -2.205 85.205 -1.875 85.535 ;
        RECT -2.205 82.895 -1.875 83.225 ;
        RECT -2.205 82.045 -1.875 82.375 ;
        RECT -2.205 79.735 -1.875 80.065 ;
        RECT -2.205 78.885 -1.875 79.215 ;
        RECT -2.205 76.575 -1.875 76.905 ;
        RECT -2.205 74.995 -1.875 75.325 ;
        RECT -2.205 74.145 -1.875 74.475 ;
        RECT -2.205 71.835 -1.875 72.165 ;
        RECT -2.205 70.985 -1.875 71.315 ;
        RECT -2.205 68.675 -1.875 69.005 ;
        RECT -2.205 67.825 -1.875 68.155 ;
        RECT -2.205 65.515 -1.875 65.845 ;
        RECT -2.205 64.665 -1.875 64.995 ;
        RECT -2.205 62.355 -1.875 62.685 ;
        RECT -2.205 60.775 -1.875 61.105 ;
        RECT -2.205 59.925 -1.875 60.255 ;
        RECT -2.205 57.615 -1.875 57.945 ;
        RECT -2.205 56.765 -1.875 57.095 ;
        RECT -2.205 54.455 -1.875 54.785 ;
        RECT -2.205 53.605 -1.875 53.935 ;
        RECT -2.205 51.295 -1.875 51.625 ;
        RECT -2.205 50.445 -1.875 50.775 ;
        RECT -2.205 48.135 -1.875 48.465 ;
        RECT -2.205 46.555 -1.875 46.885 ;
        RECT -2.205 45.705 -1.875 46.035 ;
        RECT -2.205 43.395 -1.875 43.725 ;
        RECT -2.205 42.545 -1.875 42.875 ;
        RECT -2.205 40.235 -1.875 40.565 ;
        RECT -2.205 39.385 -1.875 39.715 ;
        RECT -2.205 37.075 -1.875 37.405 ;
        RECT -2.205 36.225 -1.875 36.555 ;
        RECT -2.205 33.915 -1.875 34.245 ;
        RECT -2.205 32.335 -1.875 32.665 ;
        RECT -2.205 31.485 -1.875 31.815 ;
        RECT -2.205 29.175 -1.875 29.505 ;
        RECT -2.205 28.325 -1.875 28.655 ;
        RECT -2.205 26.015 -1.875 26.345 ;
        RECT -2.205 25.165 -1.875 25.495 ;
        RECT -2.205 22.855 -1.875 23.185 ;
        RECT -2.205 22.005 -1.875 22.335 ;
        RECT -2.205 19.695 -1.875 20.025 ;
        RECT -2.205 18.115 -1.875 18.445 ;
        RECT -2.205 17.265 -1.875 17.595 ;
        RECT -2.205 14.955 -1.875 15.285 ;
        RECT -2.205 14.105 -1.875 14.435 ;
        RECT -2.205 11.795 -1.875 12.125 ;
        RECT -2.205 10.945 -1.875 11.275 ;
        RECT -2.205 8.635 -1.875 8.965 ;
        RECT -2.205 7.785 -1.875 8.115 ;
        RECT -2.205 5.475 -1.875 5.805 ;
        RECT -2.205 3.895 -1.875 4.225 ;
        RECT -2.205 3.045 -1.875 3.375 ;
        RECT -2.205 0.87 -1.875 1.2 ;
        RECT -2.205 -0.845 -1.875 -0.515 ;
        RECT -2.205 -2.205 -1.875 -1.875 ;
        RECT -2.205 -3.565 -1.875 -3.235 ;
        RECT -2.205 -4.925 -1.875 -4.595 ;
        RECT -2.205 -6.285 -1.875 -5.955 ;
        RECT -2.205 -7.645 -1.875 -7.315 ;
        RECT -2.205 -9.005 -1.875 -8.675 ;
        RECT -2.205 -10.365 -1.875 -10.035 ;
        RECT -2.205 -11.725 -1.875 -11.395 ;
        RECT -2.205 -13.085 -1.875 -12.755 ;
        RECT -2.205 -14.445 -1.875 -14.115 ;
        RECT -2.205 -15.805 -1.875 -15.475 ;
        RECT -2.205 -17.165 -1.875 -16.835 ;
        RECT -2.205 -21.245 -1.875 -20.915 ;
        RECT -2.205 -22.605 -1.875 -22.275 ;
        RECT -2.205 -23.965 -1.875 -23.635 ;
        RECT -2.205 -25.325 -1.875 -24.995 ;
        RECT -2.205 -26.685 -1.875 -26.355 ;
        RECT -2.205 -28.045 -1.875 -27.715 ;
        RECT -2.205 -29.405 -1.875 -29.075 ;
        RECT -2.205 -30.765 -1.875 -30.435 ;
        RECT -2.205 -32.125 -1.875 -31.795 ;
        RECT -2.205 -33.485 -1.875 -33.155 ;
        RECT -2.205 -34.845 -1.875 -34.515 ;
        RECT -2.205 -36.205 -1.875 -35.875 ;
        RECT -2.205 -37.565 -1.875 -37.235 ;
        RECT -2.205 -38.925 -1.875 -38.595 ;
        RECT -2.205 -40.285 -1.875 -39.955 ;
        RECT -2.205 -41.645 -1.875 -41.315 ;
        RECT -2.205 -43.005 -1.875 -42.675 ;
        RECT -2.205 -44.365 -1.875 -44.035 ;
        RECT -2.205 -45.725 -1.875 -45.395 ;
        RECT -2.205 -49.805 -1.875 -49.475 ;
        RECT -2.205 -51.165 -1.875 -50.835 ;
        RECT -2.205 -52.525 -1.875 -52.195 ;
        RECT -2.205 -53.885 -1.875 -53.555 ;
        RECT -2.205 -55.245 -1.875 -54.915 ;
        RECT -2.205 -56.605 -1.875 -56.275 ;
        RECT -2.205 -57.965 -1.875 -57.635 ;
        RECT -2.205 -59.325 -1.875 -58.995 ;
        RECT -2.205 -60.685 -1.875 -60.355 ;
        RECT -2.205 -62.045 -1.875 -61.715 ;
        RECT -2.205 -63.405 -1.875 -63.075 ;
        RECT -2.205 -64.765 -1.875 -64.435 ;
        RECT -2.205 -66.125 -1.875 -65.795 ;
        RECT -2.205 -67.485 -1.875 -67.155 ;
        RECT -2.205 -68.845 -1.875 -68.515 ;
        RECT -2.205 -70.205 -1.875 -69.875 ;
        RECT -2.205 -71.565 -1.875 -71.235 ;
        RECT -2.205 -72.925 -1.875 -72.595 ;
        RECT -2.205 -74.285 -1.875 -73.955 ;
        RECT -2.205 -75.645 -1.875 -75.315 ;
        RECT -2.205 -77.005 -1.875 -76.675 ;
        RECT -2.205 -78.365 -1.875 -78.035 ;
        RECT -2.205 -79.725 -1.875 -79.395 ;
        RECT -2.205 -81.085 -1.875 -80.755 ;
        RECT -2.205 -82.445 -1.875 -82.115 ;
        RECT -2.205 -83.805 -1.875 -83.475 ;
        RECT -2.205 -85.165 -1.875 -84.835 ;
        RECT -2.205 -87.885 -1.875 -87.555 ;
        RECT -2.205 -89.245 -1.875 -88.915 ;
        RECT -2.205 -90.605 -1.875 -90.275 ;
        RECT -2.205 -91.965 -1.875 -91.635 ;
        RECT -2.205 -93.325 -1.875 -92.995 ;
        RECT -2.205 -94.685 -1.875 -94.355 ;
        RECT -2.205 -96.045 -1.875 -95.715 ;
        RECT -2.205 -97.405 -1.875 -97.075 ;
        RECT -2.205 -98.765 -1.875 -98.435 ;
        RECT -2.205 -100.125 -1.875 -99.795 ;
        RECT -2.205 -101.485 -1.875 -101.155 ;
        RECT -2.205 -102.845 -1.875 -102.515 ;
        RECT -2.205 -104.205 -1.875 -103.875 ;
        RECT -2.205 -105.565 -1.875 -105.235 ;
        RECT -2.205 -106.925 -1.875 -106.595 ;
        RECT -2.205 -108.285 -1.875 -107.955 ;
        RECT -2.205 -109.645 -1.875 -109.315 ;
        RECT -2.205 -111.005 -1.875 -110.675 ;
        RECT -2.205 -112.365 -1.875 -112.035 ;
        RECT -2.205 -113.725 -1.875 -113.395 ;
        RECT -2.205 -115.085 -1.875 -114.755 ;
        RECT -2.205 -116.445 -1.875 -116.115 ;
        RECT -2.205 -117.805 -1.875 -117.475 ;
        RECT -2.205 -119.165 -1.875 -118.835 ;
        RECT -2.205 -120.525 -1.875 -120.195 ;
        RECT -2.205 -121.885 -1.875 -121.555 ;
        RECT -2.205 -123.245 -1.875 -122.915 ;
        RECT -2.205 -124.605 -1.875 -124.275 ;
        RECT -2.205 -125.965 -1.875 -125.635 ;
        RECT -2.205 -127.325 -1.875 -126.995 ;
        RECT -2.205 -128.685 -1.875 -128.355 ;
        RECT -2.205 -130.045 -1.875 -129.715 ;
        RECT -2.205 -131.405 -1.875 -131.075 ;
        RECT -2.205 -132.765 -1.875 -132.435 ;
        RECT -2.205 -134.125 -1.875 -133.795 ;
        RECT -2.205 -135.485 -1.875 -135.155 ;
        RECT -2.205 -136.845 -1.875 -136.515 ;
        RECT -2.205 -138.205 -1.875 -137.875 ;
        RECT -2.205 -139.565 -1.875 -139.235 ;
        RECT -2.205 -140.925 -1.875 -140.595 ;
        RECT -2.205 -142.285 -1.875 -141.955 ;
        RECT -2.205 -143.645 -1.875 -143.315 ;
        RECT -2.205 -145.005 -1.875 -144.675 ;
        RECT -2.205 -146.365 -1.875 -146.035 ;
        RECT -2.205 -147.725 -1.875 -147.395 ;
        RECT -2.205 -149.085 -1.875 -148.755 ;
        RECT -2.205 -150.445 -1.875 -150.115 ;
        RECT -2.205 -151.805 -1.875 -151.475 ;
        RECT -2.205 -153.165 -1.875 -152.835 ;
        RECT -2.205 -154.525 -1.875 -154.195 ;
        RECT -2.205 -155.885 -1.875 -155.555 ;
        RECT -2.205 -157.245 -1.875 -156.915 ;
        RECT -2.205 -162.89 -1.875 -161.76 ;
        RECT -2.2 -163.005 -1.88 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 -139.565 -0.515 -139.235 ;
        RECT -0.845 -140.925 -0.515 -140.595 ;
        RECT -0.845 -142.285 -0.515 -141.955 ;
        RECT -0.845 -143.645 -0.515 -143.315 ;
        RECT -0.845 -145.005 -0.515 -144.675 ;
        RECT -0.845 -146.365 -0.515 -146.035 ;
        RECT -0.845 -147.725 -0.515 -147.395 ;
        RECT -0.845 -149.085 -0.515 -148.755 ;
        RECT -0.845 -150.445 -0.515 -150.115 ;
        RECT -0.845 -151.805 -0.515 -151.475 ;
        RECT -0.845 -153.165 -0.515 -152.835 ;
        RECT -0.845 -154.525 -0.515 -154.195 ;
        RECT -0.845 -155.885 -0.515 -155.555 ;
        RECT -0.845 -157.245 -0.515 -156.915 ;
        RECT -0.845 -162.89 -0.515 -161.76 ;
        RECT -0.84 -163.005 -0.52 131.19 ;
        RECT -0.845 129.945 -0.515 131.075 ;
        RECT -0.845 125.635 -0.515 125.965 ;
        RECT -0.845 124.275 -0.515 124.605 ;
        RECT -0.845 121.41 -0.515 121.74 ;
        RECT -0.845 119.235 -0.515 119.565 ;
        RECT -0.845 117.655 -0.515 117.985 ;
        RECT -0.845 116.805 -0.515 117.135 ;
        RECT -0.845 114.495 -0.515 114.825 ;
        RECT -0.845 113.645 -0.515 113.975 ;
        RECT -0.845 111.335 -0.515 111.665 ;
        RECT -0.845 110.485 -0.515 110.815 ;
        RECT -0.845 108.175 -0.515 108.505 ;
        RECT -0.845 107.325 -0.515 107.655 ;
        RECT -0.845 105.015 -0.515 105.345 ;
        RECT -0.845 103.435 -0.515 103.765 ;
        RECT -0.845 102.585 -0.515 102.915 ;
        RECT -0.845 100.275 -0.515 100.605 ;
        RECT -0.845 99.425 -0.515 99.755 ;
        RECT -0.845 97.115 -0.515 97.445 ;
        RECT -0.845 96.265 -0.515 96.595 ;
        RECT -0.845 93.955 -0.515 94.285 ;
        RECT -0.845 93.105 -0.515 93.435 ;
        RECT -0.845 90.795 -0.515 91.125 ;
        RECT -0.845 89.215 -0.515 89.545 ;
        RECT -0.845 88.365 -0.515 88.695 ;
        RECT -0.845 86.055 -0.515 86.385 ;
        RECT -0.845 85.205 -0.515 85.535 ;
        RECT -0.845 82.895 -0.515 83.225 ;
        RECT -0.845 82.045 -0.515 82.375 ;
        RECT -0.845 79.735 -0.515 80.065 ;
        RECT -0.845 78.885 -0.515 79.215 ;
        RECT -0.845 76.575 -0.515 76.905 ;
        RECT -0.845 74.995 -0.515 75.325 ;
        RECT -0.845 74.145 -0.515 74.475 ;
        RECT -0.845 71.835 -0.515 72.165 ;
        RECT -0.845 70.985 -0.515 71.315 ;
        RECT -0.845 68.675 -0.515 69.005 ;
        RECT -0.845 67.825 -0.515 68.155 ;
        RECT -0.845 65.515 -0.515 65.845 ;
        RECT -0.845 64.665 -0.515 64.995 ;
        RECT -0.845 62.355 -0.515 62.685 ;
        RECT -0.845 60.775 -0.515 61.105 ;
        RECT -0.845 59.925 -0.515 60.255 ;
        RECT -0.845 57.615 -0.515 57.945 ;
        RECT -0.845 56.765 -0.515 57.095 ;
        RECT -0.845 54.455 -0.515 54.785 ;
        RECT -0.845 53.605 -0.515 53.935 ;
        RECT -0.845 51.295 -0.515 51.625 ;
        RECT -0.845 50.445 -0.515 50.775 ;
        RECT -0.845 48.135 -0.515 48.465 ;
        RECT -0.845 46.555 -0.515 46.885 ;
        RECT -0.845 45.705 -0.515 46.035 ;
        RECT -0.845 43.395 -0.515 43.725 ;
        RECT -0.845 42.545 -0.515 42.875 ;
        RECT -0.845 40.235 -0.515 40.565 ;
        RECT -0.845 39.385 -0.515 39.715 ;
        RECT -0.845 37.075 -0.515 37.405 ;
        RECT -0.845 36.225 -0.515 36.555 ;
        RECT -0.845 33.915 -0.515 34.245 ;
        RECT -0.845 32.335 -0.515 32.665 ;
        RECT -0.845 31.485 -0.515 31.815 ;
        RECT -0.845 29.175 -0.515 29.505 ;
        RECT -0.845 28.325 -0.515 28.655 ;
        RECT -0.845 26.015 -0.515 26.345 ;
        RECT -0.845 25.165 -0.515 25.495 ;
        RECT -0.845 22.855 -0.515 23.185 ;
        RECT -0.845 22.005 -0.515 22.335 ;
        RECT -0.845 19.695 -0.515 20.025 ;
        RECT -0.845 18.115 -0.515 18.445 ;
        RECT -0.845 17.265 -0.515 17.595 ;
        RECT -0.845 14.955 -0.515 15.285 ;
        RECT -0.845 14.105 -0.515 14.435 ;
        RECT -0.845 11.795 -0.515 12.125 ;
        RECT -0.845 10.945 -0.515 11.275 ;
        RECT -0.845 8.635 -0.515 8.965 ;
        RECT -0.845 7.785 -0.515 8.115 ;
        RECT -0.845 5.475 -0.515 5.805 ;
        RECT -0.845 3.895 -0.515 4.225 ;
        RECT -0.845 3.045 -0.515 3.375 ;
        RECT -0.845 0.87 -0.515 1.2 ;
        RECT -0.845 -0.845 -0.515 -0.515 ;
        RECT -0.845 -2.205 -0.515 -1.875 ;
        RECT -0.845 -3.565 -0.515 -3.235 ;
        RECT -0.845 -4.925 -0.515 -4.595 ;
        RECT -0.845 -6.285 -0.515 -5.955 ;
        RECT -0.845 -7.645 -0.515 -7.315 ;
        RECT -0.845 -9.005 -0.515 -8.675 ;
        RECT -0.845 -10.365 -0.515 -10.035 ;
        RECT -0.845 -13.085 -0.515 -12.755 ;
        RECT -0.845 -14.445 -0.515 -14.115 ;
        RECT -0.845 -15.805 -0.515 -15.475 ;
        RECT -0.845 -17.165 -0.515 -16.835 ;
        RECT -0.845 -21.245 -0.515 -20.915 ;
        RECT -0.845 -22.605 -0.515 -22.275 ;
        RECT -0.845 -23.965 -0.515 -23.635 ;
        RECT -0.845 -25.325 -0.515 -24.995 ;
        RECT -0.845 -26.685 -0.515 -26.355 ;
        RECT -0.845 -28.045 -0.515 -27.715 ;
        RECT -0.845 -29.405 -0.515 -29.075 ;
        RECT -0.845 -30.765 -0.515 -30.435 ;
        RECT -0.845 -32.125 -0.515 -31.795 ;
        RECT -0.845 -33.485 -0.515 -33.155 ;
        RECT -0.845 -34.845 -0.515 -34.515 ;
        RECT -0.845 -36.205 -0.515 -35.875 ;
        RECT -0.845 -37.565 -0.515 -37.235 ;
        RECT -0.845 -38.925 -0.515 -38.595 ;
        RECT -0.845 -40.285 -0.515 -39.955 ;
        RECT -0.845 -41.645 -0.515 -41.315 ;
        RECT -0.845 -43.005 -0.515 -42.675 ;
        RECT -0.845 -44.365 -0.515 -44.035 ;
        RECT -0.845 -45.725 -0.515 -45.395 ;
        RECT -0.845 -49.805 -0.515 -49.475 ;
        RECT -0.845 -51.165 -0.515 -50.835 ;
        RECT -0.845 -52.525 -0.515 -52.195 ;
        RECT -0.845 -53.885 -0.515 -53.555 ;
        RECT -0.845 -55.245 -0.515 -54.915 ;
        RECT -0.845 -56.605 -0.515 -56.275 ;
        RECT -0.845 -57.965 -0.515 -57.635 ;
        RECT -0.845 -59.325 -0.515 -58.995 ;
        RECT -0.845 -60.685 -0.515 -60.355 ;
        RECT -0.845 -62.045 -0.515 -61.715 ;
        RECT -0.845 -63.405 -0.515 -63.075 ;
        RECT -0.845 -64.765 -0.515 -64.435 ;
        RECT -0.845 -66.125 -0.515 -65.795 ;
        RECT -0.845 -67.485 -0.515 -67.155 ;
        RECT -0.845 -68.845 -0.515 -68.515 ;
        RECT -0.845 -70.205 -0.515 -69.875 ;
        RECT -0.845 -71.565 -0.515 -71.235 ;
        RECT -0.845 -72.925 -0.515 -72.595 ;
        RECT -0.845 -74.285 -0.515 -73.955 ;
        RECT -0.845 -75.645 -0.515 -75.315 ;
        RECT -0.845 -77.005 -0.515 -76.675 ;
        RECT -0.845 -78.365 -0.515 -78.035 ;
        RECT -0.845 -79.725 -0.515 -79.395 ;
        RECT -0.845 -81.085 -0.515 -80.755 ;
        RECT -0.845 -82.445 -0.515 -82.115 ;
        RECT -0.845 -83.805 -0.515 -83.475 ;
        RECT -0.845 -85.165 -0.515 -84.835 ;
        RECT -0.845 -87.885 -0.515 -87.555 ;
        RECT -0.845 -89.245 -0.515 -88.915 ;
        RECT -0.845 -90.605 -0.515 -90.275 ;
        RECT -0.845 -91.965 -0.515 -91.635 ;
        RECT -0.845 -93.325 -0.515 -92.995 ;
        RECT -0.845 -94.685 -0.515 -94.355 ;
        RECT -0.845 -96.045 -0.515 -95.715 ;
        RECT -0.845 -97.405 -0.515 -97.075 ;
        RECT -0.845 -98.765 -0.515 -98.435 ;
        RECT -0.845 -100.125 -0.515 -99.795 ;
        RECT -0.845 -101.485 -0.515 -101.155 ;
        RECT -0.845 -102.845 -0.515 -102.515 ;
        RECT -0.845 -104.205 -0.515 -103.875 ;
        RECT -0.845 -105.565 -0.515 -105.235 ;
        RECT -0.845 -106.925 -0.515 -106.595 ;
        RECT -0.845 -108.285 -0.515 -107.955 ;
        RECT -0.845 -109.645 -0.515 -109.315 ;
        RECT -0.845 -111.005 -0.515 -110.675 ;
        RECT -0.845 -112.365 -0.515 -112.035 ;
        RECT -0.845 -113.725 -0.515 -113.395 ;
        RECT -0.845 -115.085 -0.515 -114.755 ;
        RECT -0.845 -116.445 -0.515 -116.115 ;
        RECT -0.845 -117.805 -0.515 -117.475 ;
        RECT -0.845 -119.165 -0.515 -118.835 ;
        RECT -0.845 -120.525 -0.515 -120.195 ;
        RECT -0.845 -121.885 -0.515 -121.555 ;
        RECT -0.845 -123.245 -0.515 -122.915 ;
        RECT -0.845 -124.605 -0.515 -124.275 ;
        RECT -0.845 -125.965 -0.515 -125.635 ;
        RECT -0.845 -127.325 -0.515 -126.995 ;
        RECT -0.845 -128.685 -0.515 -128.355 ;
        RECT -0.845 -130.045 -0.515 -129.715 ;
        RECT -0.845 -131.405 -0.515 -131.075 ;
        RECT -0.845 -132.765 -0.515 -132.435 ;
        RECT -0.845 -134.125 -0.515 -133.795 ;
        RECT -0.845 -135.485 -0.515 -135.155 ;
        RECT -0.845 -136.845 -0.515 -136.515 ;
        RECT -0.845 -138.205 -0.515 -137.875 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 129.945 -18.195 131.075 ;
        RECT -18.525 125.635 -18.195 125.965 ;
        RECT -18.525 124.275 -18.195 124.605 ;
        RECT -18.525 122.915 -18.195 123.245 ;
        RECT -18.525 121.555 -18.195 121.885 ;
        RECT -18.525 120.195 -18.195 120.525 ;
        RECT -18.525 118.835 -18.195 119.165 ;
        RECT -18.525 117.475 -18.195 117.805 ;
        RECT -18.525 116.115 -18.195 116.445 ;
        RECT -18.525 114.755 -18.195 115.085 ;
        RECT -18.525 113.395 -18.195 113.725 ;
        RECT -18.525 112.035 -18.195 112.365 ;
        RECT -18.525 110.675 -18.195 111.005 ;
        RECT -18.525 109.315 -18.195 109.645 ;
        RECT -18.525 107.955 -18.195 108.285 ;
        RECT -18.525 106.595 -18.195 106.925 ;
        RECT -18.525 105.235 -18.195 105.565 ;
        RECT -18.525 103.875 -18.195 104.205 ;
        RECT -18.525 102.515 -18.195 102.845 ;
        RECT -18.525 101.155 -18.195 101.485 ;
        RECT -18.525 99.795 -18.195 100.125 ;
        RECT -18.525 98.435 -18.195 98.765 ;
        RECT -18.525 97.075 -18.195 97.405 ;
        RECT -18.525 95.715 -18.195 96.045 ;
        RECT -18.525 94.355 -18.195 94.685 ;
        RECT -18.525 92.995 -18.195 93.325 ;
        RECT -18.525 91.635 -18.195 91.965 ;
        RECT -18.525 90.275 -18.195 90.605 ;
        RECT -18.525 88.915 -18.195 89.245 ;
        RECT -18.525 87.555 -18.195 87.885 ;
        RECT -18.525 86.195 -18.195 86.525 ;
        RECT -18.525 84.835 -18.195 85.165 ;
        RECT -18.525 83.475 -18.195 83.805 ;
        RECT -18.525 82.115 -18.195 82.445 ;
        RECT -18.525 80.755 -18.195 81.085 ;
        RECT -18.525 79.395 -18.195 79.725 ;
        RECT -18.525 78.035 -18.195 78.365 ;
        RECT -18.525 76.675 -18.195 77.005 ;
        RECT -18.525 75.315 -18.195 75.645 ;
        RECT -18.525 73.955 -18.195 74.285 ;
        RECT -18.525 72.595 -18.195 72.925 ;
        RECT -18.525 71.235 -18.195 71.565 ;
        RECT -18.525 69.875 -18.195 70.205 ;
        RECT -18.525 68.515 -18.195 68.845 ;
        RECT -18.525 67.155 -18.195 67.485 ;
        RECT -18.525 65.795 -18.195 66.125 ;
        RECT -18.525 64.435 -18.195 64.765 ;
        RECT -18.525 63.075 -18.195 63.405 ;
        RECT -18.525 61.715 -18.195 62.045 ;
        RECT -18.525 60.355 -18.195 60.685 ;
        RECT -18.525 58.995 -18.195 59.325 ;
        RECT -18.525 57.635 -18.195 57.965 ;
        RECT -18.525 56.275 -18.195 56.605 ;
        RECT -18.525 54.915 -18.195 55.245 ;
        RECT -18.525 53.555 -18.195 53.885 ;
        RECT -18.525 52.195 -18.195 52.525 ;
        RECT -18.525 50.835 -18.195 51.165 ;
        RECT -18.525 49.475 -18.195 49.805 ;
        RECT -18.525 48.115 -18.195 48.445 ;
        RECT -18.525 46.755 -18.195 47.085 ;
        RECT -18.525 45.395 -18.195 45.725 ;
        RECT -18.525 44.035 -18.195 44.365 ;
        RECT -18.525 42.675 -18.195 43.005 ;
        RECT -18.525 41.315 -18.195 41.645 ;
        RECT -18.525 39.955 -18.195 40.285 ;
        RECT -18.525 38.595 -18.195 38.925 ;
        RECT -18.525 37.235 -18.195 37.565 ;
        RECT -18.525 35.875 -18.195 36.205 ;
        RECT -18.525 34.515 -18.195 34.845 ;
        RECT -18.525 33.155 -18.195 33.485 ;
        RECT -18.525 31.795 -18.195 32.125 ;
        RECT -18.525 30.435 -18.195 30.765 ;
        RECT -18.525 29.075 -18.195 29.405 ;
        RECT -18.525 27.715 -18.195 28.045 ;
        RECT -18.525 26.355 -18.195 26.685 ;
        RECT -18.525 24.995 -18.195 25.325 ;
        RECT -18.525 23.635 -18.195 23.965 ;
        RECT -18.525 22.275 -18.195 22.605 ;
        RECT -18.525 20.915 -18.195 21.245 ;
        RECT -18.525 19.555 -18.195 19.885 ;
        RECT -18.525 18.195 -18.195 18.525 ;
        RECT -18.525 16.835 -18.195 17.165 ;
        RECT -18.525 15.475 -18.195 15.805 ;
        RECT -18.525 14.115 -18.195 14.445 ;
        RECT -18.525 12.755 -18.195 13.085 ;
        RECT -18.525 11.395 -18.195 11.725 ;
        RECT -18.525 10.035 -18.195 10.365 ;
        RECT -18.525 8.675 -18.195 9.005 ;
        RECT -18.525 7.315 -18.195 7.645 ;
        RECT -18.525 5.955 -18.195 6.285 ;
        RECT -18.525 4.595 -18.195 4.925 ;
        RECT -18.525 3.235 -18.195 3.565 ;
        RECT -18.525 1.875 -18.195 2.205 ;
        RECT -18.525 0.515 -18.195 0.845 ;
        RECT -18.525 -0.845 -18.195 -0.515 ;
        RECT -18.525 -2.205 -18.195 -1.875 ;
        RECT -18.525 -6.285 -18.195 -5.955 ;
        RECT -18.525 -8.19 -18.195 -7.86 ;
        RECT -18.525 -11.725 -18.195 -11.395 ;
        RECT -18.525 -14.23 -18.195 -13.9 ;
        RECT -18.525 -15.805 -18.195 -15.475 ;
        RECT -18.525 -18.525 -18.195 -18.195 ;
        RECT -18.52 -19.2 -18.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -25.325 -18.195 -24.995 ;
        RECT -18.525 -26.685 -18.195 -26.355 ;
        RECT -18.525 -28.045 -18.195 -27.715 ;
        RECT -18.525 -29.405 -18.195 -29.075 ;
        RECT -18.525 -31.17 -18.195 -30.84 ;
        RECT -18.525 -32.125 -18.195 -31.795 ;
        RECT -18.525 -33.485 -18.195 -33.155 ;
        RECT -18.525 -36.205 -18.195 -35.875 ;
        RECT -18.525 -37.21 -18.195 -36.88 ;
        RECT -18.525 -38.925 -18.195 -38.595 ;
        RECT -18.525 -41.645 -18.195 -41.315 ;
        RECT -18.52 -42.32 -18.2 -24.32 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -48.445 -18.195 -48.115 ;
        RECT -18.525 -49.805 -18.195 -49.475 ;
        RECT -18.525 -51.165 -18.195 -50.835 ;
        RECT -18.525 -52.75 -18.195 -52.42 ;
        RECT -18.525 -53.885 -18.195 -53.555 ;
        RECT -18.525 -55.245 -18.195 -54.915 ;
        RECT -18.525 -57.965 -18.195 -57.635 ;
        RECT -18.525 -59.325 -18.195 -58.995 ;
        RECT -18.525 -60.29 -18.195 -59.96 ;
        RECT -18.525 -62.045 -18.195 -61.715 ;
        RECT -18.525 -63.405 -18.195 -63.075 ;
        RECT -18.525 -66.125 -18.195 -65.795 ;
        RECT -18.525 -68.845 -18.195 -68.515 ;
        RECT -18.525 -70.205 -18.195 -69.875 ;
        RECT -18.525 -71.565 -18.195 -71.235 ;
        RECT -18.525 -72.925 -18.195 -72.595 ;
        RECT -18.525 -74.93 -18.195 -74.6 ;
        RECT -18.525 -75.645 -18.195 -75.315 ;
        RECT -18.525 -77.005 -18.195 -76.675 ;
        RECT -18.525 -79.725 -18.195 -79.395 ;
        RECT -18.525 -81.085 -18.195 -80.755 ;
        RECT -18.525 -82.47 -18.195 -82.14 ;
        RECT -18.525 -83.805 -18.195 -83.475 ;
        RECT -18.525 -85.165 -18.195 -84.835 ;
        RECT -18.525 -87.885 -18.195 -87.555 ;
        RECT -18.525 -93.325 -18.195 -92.995 ;
        RECT -18.525 -94.685 -18.195 -94.355 ;
        RECT -18.525 -96.045 -18.195 -95.715 ;
        RECT -18.525 -100.125 -18.195 -99.795 ;
        RECT -18.525 -104.205 -18.195 -103.875 ;
        RECT -18.525 -105.565 -18.195 -105.235 ;
        RECT -18.525 -106.925 -18.195 -106.595 ;
        RECT -18.525 -117.805 -18.195 -117.475 ;
        RECT -18.525 -120.525 -18.195 -120.195 ;
        RECT -18.525 -124.605 -18.195 -124.275 ;
        RECT -18.525 -127.325 -18.195 -126.995 ;
        RECT -18.525 -131.405 -18.195 -131.075 ;
        RECT -18.525 -136.845 -18.195 -136.515 ;
        RECT -18.525 -138.205 -18.195 -137.875 ;
        RECT -18.525 -139.565 -18.195 -139.235 ;
        RECT -18.525 -140.925 -18.195 -140.595 ;
        RECT -18.525 -142.285 -18.195 -141.955 ;
        RECT -18.525 -143.645 -18.195 -143.315 ;
        RECT -18.525 -145.005 -18.195 -144.675 ;
        RECT -18.525 -146.365 -18.195 -146.035 ;
        RECT -18.525 -148.215 -18.195 -147.885 ;
        RECT -18.525 -149.085 -18.195 -148.755 ;
        RECT -18.525 -150.445 -18.195 -150.115 ;
        RECT -18.525 -151.805 -18.195 -151.475 ;
        RECT -18.525 -153.165 -18.195 -152.835 ;
        RECT -18.525 -154.525 -18.195 -154.195 ;
        RECT -18.525 -157.245 -18.195 -156.915 ;
        RECT -18.525 -162.89 -18.195 -161.76 ;
        RECT -18.52 -163.005 -18.2 -47.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 129.945 -16.835 131.075 ;
        RECT -17.165 125.635 -16.835 125.965 ;
        RECT -17.165 124.275 -16.835 124.605 ;
        RECT -17.165 122.915 -16.835 123.245 ;
        RECT -17.165 121.555 -16.835 121.885 ;
        RECT -17.165 120.195 -16.835 120.525 ;
        RECT -17.165 118.835 -16.835 119.165 ;
        RECT -17.165 117.475 -16.835 117.805 ;
        RECT -17.165 116.115 -16.835 116.445 ;
        RECT -17.165 114.755 -16.835 115.085 ;
        RECT -17.165 113.395 -16.835 113.725 ;
        RECT -17.165 112.035 -16.835 112.365 ;
        RECT -17.165 110.675 -16.835 111.005 ;
        RECT -17.165 109.315 -16.835 109.645 ;
        RECT -17.165 107.955 -16.835 108.285 ;
        RECT -17.165 106.595 -16.835 106.925 ;
        RECT -17.165 105.235 -16.835 105.565 ;
        RECT -17.165 103.875 -16.835 104.205 ;
        RECT -17.165 102.515 -16.835 102.845 ;
        RECT -17.165 101.155 -16.835 101.485 ;
        RECT -17.165 99.795 -16.835 100.125 ;
        RECT -17.165 98.435 -16.835 98.765 ;
        RECT -17.165 97.075 -16.835 97.405 ;
        RECT -17.165 95.715 -16.835 96.045 ;
        RECT -17.165 94.355 -16.835 94.685 ;
        RECT -17.165 92.995 -16.835 93.325 ;
        RECT -17.165 91.635 -16.835 91.965 ;
        RECT -17.165 90.275 -16.835 90.605 ;
        RECT -17.165 88.915 -16.835 89.245 ;
        RECT -17.165 87.555 -16.835 87.885 ;
        RECT -17.165 86.195 -16.835 86.525 ;
        RECT -17.165 84.835 -16.835 85.165 ;
        RECT -17.165 83.475 -16.835 83.805 ;
        RECT -17.165 82.115 -16.835 82.445 ;
        RECT -17.165 80.755 -16.835 81.085 ;
        RECT -17.165 79.395 -16.835 79.725 ;
        RECT -17.165 78.035 -16.835 78.365 ;
        RECT -17.165 76.675 -16.835 77.005 ;
        RECT -17.165 75.315 -16.835 75.645 ;
        RECT -17.165 73.955 -16.835 74.285 ;
        RECT -17.165 72.595 -16.835 72.925 ;
        RECT -17.165 71.235 -16.835 71.565 ;
        RECT -17.165 69.875 -16.835 70.205 ;
        RECT -17.165 68.515 -16.835 68.845 ;
        RECT -17.165 67.155 -16.835 67.485 ;
        RECT -17.165 65.795 -16.835 66.125 ;
        RECT -17.165 64.435 -16.835 64.765 ;
        RECT -17.165 63.075 -16.835 63.405 ;
        RECT -17.165 61.715 -16.835 62.045 ;
        RECT -17.165 60.355 -16.835 60.685 ;
        RECT -17.165 58.995 -16.835 59.325 ;
        RECT -17.165 57.635 -16.835 57.965 ;
        RECT -17.165 56.275 -16.835 56.605 ;
        RECT -17.165 54.915 -16.835 55.245 ;
        RECT -17.165 53.555 -16.835 53.885 ;
        RECT -17.165 52.195 -16.835 52.525 ;
        RECT -17.165 50.835 -16.835 51.165 ;
        RECT -17.165 49.475 -16.835 49.805 ;
        RECT -17.165 48.115 -16.835 48.445 ;
        RECT -17.165 46.755 -16.835 47.085 ;
        RECT -17.165 45.395 -16.835 45.725 ;
        RECT -17.165 44.035 -16.835 44.365 ;
        RECT -17.165 42.675 -16.835 43.005 ;
        RECT -17.165 41.315 -16.835 41.645 ;
        RECT -17.165 39.955 -16.835 40.285 ;
        RECT -17.165 38.595 -16.835 38.925 ;
        RECT -17.165 37.235 -16.835 37.565 ;
        RECT -17.165 35.875 -16.835 36.205 ;
        RECT -17.165 34.515 -16.835 34.845 ;
        RECT -17.165 33.155 -16.835 33.485 ;
        RECT -17.165 31.795 -16.835 32.125 ;
        RECT -17.165 30.435 -16.835 30.765 ;
        RECT -17.165 29.075 -16.835 29.405 ;
        RECT -17.165 27.715 -16.835 28.045 ;
        RECT -17.165 26.355 -16.835 26.685 ;
        RECT -17.165 24.995 -16.835 25.325 ;
        RECT -17.165 23.635 -16.835 23.965 ;
        RECT -17.165 22.275 -16.835 22.605 ;
        RECT -17.165 20.915 -16.835 21.245 ;
        RECT -17.165 19.555 -16.835 19.885 ;
        RECT -17.165 18.195 -16.835 18.525 ;
        RECT -17.165 16.835 -16.835 17.165 ;
        RECT -17.165 15.475 -16.835 15.805 ;
        RECT -17.165 14.115 -16.835 14.445 ;
        RECT -17.165 12.755 -16.835 13.085 ;
        RECT -17.165 11.395 -16.835 11.725 ;
        RECT -17.165 10.035 -16.835 10.365 ;
        RECT -17.165 8.675 -16.835 9.005 ;
        RECT -17.165 7.315 -16.835 7.645 ;
        RECT -17.165 5.955 -16.835 6.285 ;
        RECT -17.165 4.595 -16.835 4.925 ;
        RECT -17.165 3.235 -16.835 3.565 ;
        RECT -17.165 1.875 -16.835 2.205 ;
        RECT -17.165 0.515 -16.835 0.845 ;
        RECT -17.165 -0.845 -16.835 -0.515 ;
        RECT -17.165 -2.205 -16.835 -1.875 ;
        RECT -17.165 -3.565 -16.835 -3.235 ;
        RECT -17.165 -6.285 -16.835 -5.955 ;
        RECT -17.165 -8.19 -16.835 -7.86 ;
        RECT -17.16 -8.32 -16.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -23.965 -16.835 -23.635 ;
        RECT -17.165 -25.325 -16.835 -24.995 ;
        RECT -17.165 -26.685 -16.835 -26.355 ;
        RECT -17.165 -28.045 -16.835 -27.715 ;
        RECT -17.165 -29.405 -16.835 -29.075 ;
        RECT -17.165 -31.17 -16.835 -30.84 ;
        RECT -17.165 -32.125 -16.835 -31.795 ;
        RECT -17.165 -33.485 -16.835 -33.155 ;
        RECT -17.165 -36.205 -16.835 -35.875 ;
        RECT -17.165 -37.21 -16.835 -36.88 ;
        RECT -17.165 -38.925 -16.835 -38.595 ;
        RECT -17.165 -41.645 -16.835 -41.315 ;
        RECT -17.165 -48.445 -16.835 -48.115 ;
        RECT -17.165 -49.805 -16.835 -49.475 ;
        RECT -17.165 -51.165 -16.835 -50.835 ;
        RECT -17.165 -52.75 -16.835 -52.42 ;
        RECT -17.165 -53.885 -16.835 -53.555 ;
        RECT -17.165 -55.245 -16.835 -54.915 ;
        RECT -17.165 -57.965 -16.835 -57.635 ;
        RECT -17.165 -59.325 -16.835 -58.995 ;
        RECT -17.165 -60.29 -16.835 -59.96 ;
        RECT -17.165 -62.045 -16.835 -61.715 ;
        RECT -17.165 -63.405 -16.835 -63.075 ;
        RECT -17.165 -66.125 -16.835 -65.795 ;
        RECT -17.165 -68.845 -16.835 -68.515 ;
        RECT -17.165 -70.205 -16.835 -69.875 ;
        RECT -17.165 -71.565 -16.835 -71.235 ;
        RECT -17.165 -72.925 -16.835 -72.595 ;
        RECT -17.165 -74.93 -16.835 -74.6 ;
        RECT -17.165 -75.645 -16.835 -75.315 ;
        RECT -17.165 -77.005 -16.835 -76.675 ;
        RECT -17.165 -79.725 -16.835 -79.395 ;
        RECT -17.165 -82.47 -16.835 -82.14 ;
        RECT -17.165 -83.805 -16.835 -83.475 ;
        RECT -17.165 -85.165 -16.835 -84.835 ;
        RECT -17.165 -87.885 -16.835 -87.555 ;
        RECT -17.16 -92.64 -16.84 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -154.525 -16.835 -154.195 ;
        RECT -17.165 -157.245 -16.835 -156.915 ;
        RECT -17.165 -162.89 -16.835 -161.76 ;
        RECT -17.16 -163.005 -16.84 -153.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 129.945 -15.475 131.075 ;
        RECT -15.805 125.635 -15.475 125.965 ;
        RECT -15.805 124.275 -15.475 124.605 ;
        RECT -15.805 122.915 -15.475 123.245 ;
        RECT -15.805 121.555 -15.475 121.885 ;
        RECT -15.805 120.195 -15.475 120.525 ;
        RECT -15.805 118.835 -15.475 119.165 ;
        RECT -15.805 117.475 -15.475 117.805 ;
        RECT -15.805 116.115 -15.475 116.445 ;
        RECT -15.805 114.755 -15.475 115.085 ;
        RECT -15.805 113.395 -15.475 113.725 ;
        RECT -15.805 112.035 -15.475 112.365 ;
        RECT -15.805 110.675 -15.475 111.005 ;
        RECT -15.805 109.315 -15.475 109.645 ;
        RECT -15.805 107.955 -15.475 108.285 ;
        RECT -15.805 106.595 -15.475 106.925 ;
        RECT -15.805 105.235 -15.475 105.565 ;
        RECT -15.805 103.875 -15.475 104.205 ;
        RECT -15.805 102.515 -15.475 102.845 ;
        RECT -15.805 101.155 -15.475 101.485 ;
        RECT -15.805 99.795 -15.475 100.125 ;
        RECT -15.805 98.435 -15.475 98.765 ;
        RECT -15.805 97.075 -15.475 97.405 ;
        RECT -15.805 95.715 -15.475 96.045 ;
        RECT -15.805 94.355 -15.475 94.685 ;
        RECT -15.805 92.995 -15.475 93.325 ;
        RECT -15.805 91.635 -15.475 91.965 ;
        RECT -15.805 90.275 -15.475 90.605 ;
        RECT -15.805 88.915 -15.475 89.245 ;
        RECT -15.805 87.555 -15.475 87.885 ;
        RECT -15.805 86.195 -15.475 86.525 ;
        RECT -15.805 84.835 -15.475 85.165 ;
        RECT -15.805 83.475 -15.475 83.805 ;
        RECT -15.805 82.115 -15.475 82.445 ;
        RECT -15.805 80.755 -15.475 81.085 ;
        RECT -15.805 79.395 -15.475 79.725 ;
        RECT -15.805 78.035 -15.475 78.365 ;
        RECT -15.805 76.675 -15.475 77.005 ;
        RECT -15.805 75.315 -15.475 75.645 ;
        RECT -15.805 73.955 -15.475 74.285 ;
        RECT -15.805 72.595 -15.475 72.925 ;
        RECT -15.805 71.235 -15.475 71.565 ;
        RECT -15.805 69.875 -15.475 70.205 ;
        RECT -15.805 68.515 -15.475 68.845 ;
        RECT -15.805 67.155 -15.475 67.485 ;
        RECT -15.805 65.795 -15.475 66.125 ;
        RECT -15.805 64.435 -15.475 64.765 ;
        RECT -15.805 63.075 -15.475 63.405 ;
        RECT -15.805 61.715 -15.475 62.045 ;
        RECT -15.805 60.355 -15.475 60.685 ;
        RECT -15.805 58.995 -15.475 59.325 ;
        RECT -15.805 57.635 -15.475 57.965 ;
        RECT -15.805 56.275 -15.475 56.605 ;
        RECT -15.805 54.915 -15.475 55.245 ;
        RECT -15.805 53.555 -15.475 53.885 ;
        RECT -15.805 52.195 -15.475 52.525 ;
        RECT -15.805 50.835 -15.475 51.165 ;
        RECT -15.805 49.475 -15.475 49.805 ;
        RECT -15.805 48.115 -15.475 48.445 ;
        RECT -15.805 46.755 -15.475 47.085 ;
        RECT -15.805 45.395 -15.475 45.725 ;
        RECT -15.805 44.035 -15.475 44.365 ;
        RECT -15.805 42.675 -15.475 43.005 ;
        RECT -15.805 41.315 -15.475 41.645 ;
        RECT -15.805 39.955 -15.475 40.285 ;
        RECT -15.805 38.595 -15.475 38.925 ;
        RECT -15.805 37.235 -15.475 37.565 ;
        RECT -15.805 35.875 -15.475 36.205 ;
        RECT -15.805 34.515 -15.475 34.845 ;
        RECT -15.805 33.155 -15.475 33.485 ;
        RECT -15.805 31.795 -15.475 32.125 ;
        RECT -15.805 30.435 -15.475 30.765 ;
        RECT -15.805 29.075 -15.475 29.405 ;
        RECT -15.805 27.715 -15.475 28.045 ;
        RECT -15.805 26.355 -15.475 26.685 ;
        RECT -15.805 24.995 -15.475 25.325 ;
        RECT -15.805 23.635 -15.475 23.965 ;
        RECT -15.805 22.275 -15.475 22.605 ;
        RECT -15.805 20.915 -15.475 21.245 ;
        RECT -15.805 19.555 -15.475 19.885 ;
        RECT -15.805 18.195 -15.475 18.525 ;
        RECT -15.805 16.835 -15.475 17.165 ;
        RECT -15.805 15.475 -15.475 15.805 ;
        RECT -15.805 14.115 -15.475 14.445 ;
        RECT -15.805 12.755 -15.475 13.085 ;
        RECT -15.805 11.395 -15.475 11.725 ;
        RECT -15.805 10.035 -15.475 10.365 ;
        RECT -15.805 8.675 -15.475 9.005 ;
        RECT -15.805 7.315 -15.475 7.645 ;
        RECT -15.805 5.955 -15.475 6.285 ;
        RECT -15.805 4.595 -15.475 4.925 ;
        RECT -15.805 3.235 -15.475 3.565 ;
        RECT -15.805 1.875 -15.475 2.205 ;
        RECT -15.805 0.515 -15.475 0.845 ;
        RECT -15.805 -0.845 -15.475 -0.515 ;
        RECT -15.805 -2.205 -15.475 -1.875 ;
        RECT -15.805 -3.565 -15.475 -3.235 ;
        RECT -15.805 -6.285 -15.475 -5.955 ;
        RECT -15.805 -8.19 -15.475 -7.86 ;
        RECT -15.805 -9.005 -15.475 -8.675 ;
        RECT -15.805 -11.725 -15.475 -11.395 ;
        RECT -15.805 -14.23 -15.475 -13.9 ;
        RECT -15.805 -15.805 -15.475 -15.475 ;
        RECT -15.805 -18.525 -15.475 -18.195 ;
        RECT -15.805 -23.965 -15.475 -23.635 ;
        RECT -15.805 -25.325 -15.475 -24.995 ;
        RECT -15.805 -26.685 -15.475 -26.355 ;
        RECT -15.805 -28.045 -15.475 -27.715 ;
        RECT -15.805 -29.405 -15.475 -29.075 ;
        RECT -15.805 -31.17 -15.475 -30.84 ;
        RECT -15.805 -32.125 -15.475 -31.795 ;
        RECT -15.805 -33.485 -15.475 -33.155 ;
        RECT -15.805 -36.205 -15.475 -35.875 ;
        RECT -15.805 -37.21 -15.475 -36.88 ;
        RECT -15.805 -38.925 -15.475 -38.595 ;
        RECT -15.805 -41.645 -15.475 -41.315 ;
        RECT -15.805 -48.445 -15.475 -48.115 ;
        RECT -15.805 -49.805 -15.475 -49.475 ;
        RECT -15.805 -51.165 -15.475 -50.835 ;
        RECT -15.805 -52.75 -15.475 -52.42 ;
        RECT -15.805 -53.885 -15.475 -53.555 ;
        RECT -15.805 -55.245 -15.475 -54.915 ;
        RECT -15.805 -57.965 -15.475 -57.635 ;
        RECT -15.805 -59.325 -15.475 -58.995 ;
        RECT -15.805 -60.29 -15.475 -59.96 ;
        RECT -15.805 -62.045 -15.475 -61.715 ;
        RECT -15.805 -63.405 -15.475 -63.075 ;
        RECT -15.805 -66.125 -15.475 -65.795 ;
        RECT -15.805 -68.845 -15.475 -68.515 ;
        RECT -15.805 -70.205 -15.475 -69.875 ;
        RECT -15.805 -71.565 -15.475 -71.235 ;
        RECT -15.805 -72.925 -15.475 -72.595 ;
        RECT -15.805 -74.93 -15.475 -74.6 ;
        RECT -15.805 -75.645 -15.475 -75.315 ;
        RECT -15.805 -77.005 -15.475 -76.675 ;
        RECT -15.805 -79.725 -15.475 -79.395 ;
        RECT -15.805 -82.47 -15.475 -82.14 ;
        RECT -15.805 -83.805 -15.475 -83.475 ;
        RECT -15.805 -85.165 -15.475 -84.835 ;
        RECT -15.805 -87.885 -15.475 -87.555 ;
        RECT -15.8 -89.92 -15.48 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 -94.685 -15.475 -94.355 ;
        RECT -15.805 -96.045 -15.475 -95.715 ;
        RECT -15.805 -105.565 -15.475 -105.235 ;
        RECT -15.805 -106.925 -15.475 -106.595 ;
        RECT -15.805 -117.805 -15.475 -117.475 ;
        RECT -15.805 -120.525 -15.475 -120.195 ;
        RECT -15.805 -131.405 -15.475 -131.075 ;
        RECT -15.805 -136.845 -15.475 -136.515 ;
        RECT -15.805 -138.205 -15.475 -137.875 ;
        RECT -15.805 -139.565 -15.475 -139.235 ;
        RECT -15.805 -140.925 -15.475 -140.595 ;
        RECT -15.805 -142.285 -15.475 -141.955 ;
        RECT -15.805 -143.645 -15.475 -143.315 ;
        RECT -15.805 -145.005 -15.475 -144.675 ;
        RECT -15.805 -146.365 -15.475 -146.035 ;
        RECT -15.805 -148.215 -15.475 -147.885 ;
        RECT -15.805 -149.085 -15.475 -148.755 ;
        RECT -15.805 -150.445 -15.475 -150.115 ;
        RECT -15.805 -153.165 -15.475 -152.835 ;
        RECT -15.805 -154.525 -15.475 -154.195 ;
        RECT -15.805 -157.245 -15.475 -156.915 ;
        RECT -15.805 -162.89 -15.475 -161.76 ;
        RECT -15.8 -163.005 -15.48 -93.68 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 129.945 -14.115 131.075 ;
        RECT -14.445 125.635 -14.115 125.965 ;
        RECT -14.445 124.275 -14.115 124.605 ;
        RECT -14.445 122.915 -14.115 123.245 ;
        RECT -14.445 121.555 -14.115 121.885 ;
        RECT -14.445 120.195 -14.115 120.525 ;
        RECT -14.445 118.835 -14.115 119.165 ;
        RECT -14.445 117.475 -14.115 117.805 ;
        RECT -14.445 116.115 -14.115 116.445 ;
        RECT -14.445 114.755 -14.115 115.085 ;
        RECT -14.445 113.395 -14.115 113.725 ;
        RECT -14.445 112.035 -14.115 112.365 ;
        RECT -14.445 110.675 -14.115 111.005 ;
        RECT -14.445 109.315 -14.115 109.645 ;
        RECT -14.445 107.955 -14.115 108.285 ;
        RECT -14.445 106.595 -14.115 106.925 ;
        RECT -14.445 105.235 -14.115 105.565 ;
        RECT -14.445 103.875 -14.115 104.205 ;
        RECT -14.445 102.515 -14.115 102.845 ;
        RECT -14.445 101.155 -14.115 101.485 ;
        RECT -14.445 99.795 -14.115 100.125 ;
        RECT -14.445 98.435 -14.115 98.765 ;
        RECT -14.445 97.075 -14.115 97.405 ;
        RECT -14.445 95.715 -14.115 96.045 ;
        RECT -14.445 94.355 -14.115 94.685 ;
        RECT -14.445 92.995 -14.115 93.325 ;
        RECT -14.445 91.635 -14.115 91.965 ;
        RECT -14.445 90.275 -14.115 90.605 ;
        RECT -14.445 88.915 -14.115 89.245 ;
        RECT -14.445 87.555 -14.115 87.885 ;
        RECT -14.445 86.195 -14.115 86.525 ;
        RECT -14.445 84.835 -14.115 85.165 ;
        RECT -14.445 83.475 -14.115 83.805 ;
        RECT -14.445 82.115 -14.115 82.445 ;
        RECT -14.445 80.755 -14.115 81.085 ;
        RECT -14.445 79.395 -14.115 79.725 ;
        RECT -14.445 78.035 -14.115 78.365 ;
        RECT -14.445 76.675 -14.115 77.005 ;
        RECT -14.445 75.315 -14.115 75.645 ;
        RECT -14.445 73.955 -14.115 74.285 ;
        RECT -14.445 72.595 -14.115 72.925 ;
        RECT -14.445 71.235 -14.115 71.565 ;
        RECT -14.445 69.875 -14.115 70.205 ;
        RECT -14.445 68.515 -14.115 68.845 ;
        RECT -14.445 67.155 -14.115 67.485 ;
        RECT -14.445 65.795 -14.115 66.125 ;
        RECT -14.445 64.435 -14.115 64.765 ;
        RECT -14.445 63.075 -14.115 63.405 ;
        RECT -14.445 61.715 -14.115 62.045 ;
        RECT -14.445 60.355 -14.115 60.685 ;
        RECT -14.445 58.995 -14.115 59.325 ;
        RECT -14.445 57.635 -14.115 57.965 ;
        RECT -14.445 56.275 -14.115 56.605 ;
        RECT -14.445 54.915 -14.115 55.245 ;
        RECT -14.445 53.555 -14.115 53.885 ;
        RECT -14.445 52.195 -14.115 52.525 ;
        RECT -14.445 50.835 -14.115 51.165 ;
        RECT -14.445 49.475 -14.115 49.805 ;
        RECT -14.445 48.115 -14.115 48.445 ;
        RECT -14.445 46.755 -14.115 47.085 ;
        RECT -14.445 45.395 -14.115 45.725 ;
        RECT -14.445 44.035 -14.115 44.365 ;
        RECT -14.445 42.675 -14.115 43.005 ;
        RECT -14.445 41.315 -14.115 41.645 ;
        RECT -14.445 39.955 -14.115 40.285 ;
        RECT -14.445 38.595 -14.115 38.925 ;
        RECT -14.445 37.235 -14.115 37.565 ;
        RECT -14.445 35.875 -14.115 36.205 ;
        RECT -14.445 34.515 -14.115 34.845 ;
        RECT -14.445 33.155 -14.115 33.485 ;
        RECT -14.445 31.795 -14.115 32.125 ;
        RECT -14.445 30.435 -14.115 30.765 ;
        RECT -14.445 29.075 -14.115 29.405 ;
        RECT -14.445 27.715 -14.115 28.045 ;
        RECT -14.445 26.355 -14.115 26.685 ;
        RECT -14.445 24.995 -14.115 25.325 ;
        RECT -14.445 23.635 -14.115 23.965 ;
        RECT -14.445 22.275 -14.115 22.605 ;
        RECT -14.445 20.915 -14.115 21.245 ;
        RECT -14.445 19.555 -14.115 19.885 ;
        RECT -14.445 18.195 -14.115 18.525 ;
        RECT -14.445 16.835 -14.115 17.165 ;
        RECT -14.445 15.475 -14.115 15.805 ;
        RECT -14.445 14.115 -14.115 14.445 ;
        RECT -14.445 12.755 -14.115 13.085 ;
        RECT -14.445 11.395 -14.115 11.725 ;
        RECT -14.445 10.035 -14.115 10.365 ;
        RECT -14.445 8.675 -14.115 9.005 ;
        RECT -14.445 7.315 -14.115 7.645 ;
        RECT -14.445 5.955 -14.115 6.285 ;
        RECT -14.445 4.595 -14.115 4.925 ;
        RECT -14.445 3.235 -14.115 3.565 ;
        RECT -14.445 1.875 -14.115 2.205 ;
        RECT -14.445 0.515 -14.115 0.845 ;
        RECT -14.445 -0.845 -14.115 -0.515 ;
        RECT -14.445 -2.205 -14.115 -1.875 ;
        RECT -14.445 -3.565 -14.115 -3.235 ;
        RECT -14.445 -6.285 -14.115 -5.955 ;
        RECT -14.445 -8.19 -14.115 -7.86 ;
        RECT -14.445 -9.005 -14.115 -8.675 ;
        RECT -14.445 -11.725 -14.115 -11.395 ;
        RECT -14.445 -14.23 -14.115 -13.9 ;
        RECT -14.445 -15.805 -14.115 -15.475 ;
        RECT -14.445 -18.525 -14.115 -18.195 ;
        RECT -14.445 -23.965 -14.115 -23.635 ;
        RECT -14.445 -25.325 -14.115 -24.995 ;
        RECT -14.445 -26.685 -14.115 -26.355 ;
        RECT -14.445 -28.045 -14.115 -27.715 ;
        RECT -14.445 -29.405 -14.115 -29.075 ;
        RECT -14.445 -31.17 -14.115 -30.84 ;
        RECT -14.445 -32.125 -14.115 -31.795 ;
        RECT -14.445 -33.485 -14.115 -33.155 ;
        RECT -14.445 -36.205 -14.115 -35.875 ;
        RECT -14.445 -37.21 -14.115 -36.88 ;
        RECT -14.445 -38.925 -14.115 -38.595 ;
        RECT -14.445 -41.645 -14.115 -41.315 ;
        RECT -14.445 -48.445 -14.115 -48.115 ;
        RECT -14.445 -49.805 -14.115 -49.475 ;
        RECT -14.445 -51.165 -14.115 -50.835 ;
        RECT -14.445 -52.75 -14.115 -52.42 ;
        RECT -14.445 -53.885 -14.115 -53.555 ;
        RECT -14.445 -55.245 -14.115 -54.915 ;
        RECT -14.445 -57.965 -14.115 -57.635 ;
        RECT -14.445 -59.325 -14.115 -58.995 ;
        RECT -14.445 -60.29 -14.115 -59.96 ;
        RECT -14.445 -62.045 -14.115 -61.715 ;
        RECT -14.445 -63.405 -14.115 -63.075 ;
        RECT -14.445 -66.125 -14.115 -65.795 ;
        RECT -14.445 -68.845 -14.115 -68.515 ;
        RECT -14.445 -70.205 -14.115 -69.875 ;
        RECT -14.445 -71.565 -14.115 -71.235 ;
        RECT -14.445 -72.925 -14.115 -72.595 ;
        RECT -14.445 -74.93 -14.115 -74.6 ;
        RECT -14.445 -75.645 -14.115 -75.315 ;
        RECT -14.445 -77.005 -14.115 -76.675 ;
        RECT -14.445 -79.725 -14.115 -79.395 ;
        RECT -14.445 -82.47 -14.115 -82.14 ;
        RECT -14.445 -83.805 -14.115 -83.475 ;
        RECT -14.445 -85.165 -14.115 -84.835 ;
        RECT -14.445 -87.885 -14.115 -87.555 ;
        RECT -14.44 -89.24 -14.12 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -93.325 -14.115 -92.995 ;
        RECT -14.445 -94.685 -14.115 -94.355 ;
        RECT -14.445 -96.045 -14.115 -95.715 ;
        RECT -14.445 -98.765 -14.115 -98.435 ;
        RECT -14.445 -106.925 -14.115 -106.595 ;
        RECT -14.445 -112.365 -14.115 -112.035 ;
        RECT -14.445 -113.725 -14.115 -113.395 ;
        RECT -14.445 -120.525 -14.115 -120.195 ;
        RECT -14.445 -121.885 -14.115 -121.555 ;
        RECT -14.445 -125.965 -14.115 -125.635 ;
        RECT -14.445 -127.325 -14.115 -126.995 ;
        RECT -14.445 -131.405 -14.115 -131.075 ;
        RECT -14.445 -134.125 -14.115 -133.795 ;
        RECT -14.445 -136.845 -14.115 -136.515 ;
        RECT -14.445 -138.205 -14.115 -137.875 ;
        RECT -14.445 -139.565 -14.115 -139.235 ;
        RECT -14.445 -140.925 -14.115 -140.595 ;
        RECT -14.445 -142.285 -14.115 -141.955 ;
        RECT -14.445 -143.645 -14.115 -143.315 ;
        RECT -14.445 -145.005 -14.115 -144.675 ;
        RECT -14.445 -146.365 -14.115 -146.035 ;
        RECT -14.445 -148.215 -14.115 -147.885 ;
        RECT -14.445 -149.085 -14.115 -148.755 ;
        RECT -14.445 -150.445 -14.115 -150.115 ;
        RECT -14.445 -153.165 -14.115 -152.835 ;
        RECT -14.445 -154.525 -14.115 -154.195 ;
        RECT -14.445 -157.245 -14.115 -156.915 ;
        RECT -14.445 -162.89 -14.115 -161.76 ;
        RECT -14.44 -163.005 -14.12 -92.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 129.945 -12.755 131.075 ;
        RECT -13.085 125.635 -12.755 125.965 ;
        RECT -13.085 124.275 -12.755 124.605 ;
        RECT -13.085 122.915 -12.755 123.245 ;
        RECT -13.085 121.555 -12.755 121.885 ;
        RECT -13.085 120.195 -12.755 120.525 ;
        RECT -13.085 118.835 -12.755 119.165 ;
        RECT -13.085 117.475 -12.755 117.805 ;
        RECT -13.085 116.115 -12.755 116.445 ;
        RECT -13.085 114.755 -12.755 115.085 ;
        RECT -13.085 113.395 -12.755 113.725 ;
        RECT -13.085 112.035 -12.755 112.365 ;
        RECT -13.085 110.675 -12.755 111.005 ;
        RECT -13.085 109.315 -12.755 109.645 ;
        RECT -13.085 107.955 -12.755 108.285 ;
        RECT -13.085 106.595 -12.755 106.925 ;
        RECT -13.085 105.235 -12.755 105.565 ;
        RECT -13.085 103.875 -12.755 104.205 ;
        RECT -13.085 102.515 -12.755 102.845 ;
        RECT -13.085 101.155 -12.755 101.485 ;
        RECT -13.085 99.795 -12.755 100.125 ;
        RECT -13.085 98.435 -12.755 98.765 ;
        RECT -13.085 97.075 -12.755 97.405 ;
        RECT -13.085 95.715 -12.755 96.045 ;
        RECT -13.085 94.355 -12.755 94.685 ;
        RECT -13.085 92.995 -12.755 93.325 ;
        RECT -13.085 91.635 -12.755 91.965 ;
        RECT -13.085 90.275 -12.755 90.605 ;
        RECT -13.085 88.915 -12.755 89.245 ;
        RECT -13.085 87.555 -12.755 87.885 ;
        RECT -13.085 86.195 -12.755 86.525 ;
        RECT -13.085 84.835 -12.755 85.165 ;
        RECT -13.085 83.475 -12.755 83.805 ;
        RECT -13.085 82.115 -12.755 82.445 ;
        RECT -13.085 80.755 -12.755 81.085 ;
        RECT -13.085 79.395 -12.755 79.725 ;
        RECT -13.085 78.035 -12.755 78.365 ;
        RECT -13.085 76.675 -12.755 77.005 ;
        RECT -13.085 75.315 -12.755 75.645 ;
        RECT -13.085 73.955 -12.755 74.285 ;
        RECT -13.085 72.595 -12.755 72.925 ;
        RECT -13.085 71.235 -12.755 71.565 ;
        RECT -13.085 69.875 -12.755 70.205 ;
        RECT -13.085 68.515 -12.755 68.845 ;
        RECT -13.085 67.155 -12.755 67.485 ;
        RECT -13.085 65.795 -12.755 66.125 ;
        RECT -13.085 64.435 -12.755 64.765 ;
        RECT -13.085 63.075 -12.755 63.405 ;
        RECT -13.085 61.715 -12.755 62.045 ;
        RECT -13.085 60.355 -12.755 60.685 ;
        RECT -13.085 58.995 -12.755 59.325 ;
        RECT -13.085 57.635 -12.755 57.965 ;
        RECT -13.085 56.275 -12.755 56.605 ;
        RECT -13.085 54.915 -12.755 55.245 ;
        RECT -13.085 53.555 -12.755 53.885 ;
        RECT -13.085 52.195 -12.755 52.525 ;
        RECT -13.085 50.835 -12.755 51.165 ;
        RECT -13.085 49.475 -12.755 49.805 ;
        RECT -13.085 48.115 -12.755 48.445 ;
        RECT -13.085 46.755 -12.755 47.085 ;
        RECT -13.085 45.395 -12.755 45.725 ;
        RECT -13.085 44.035 -12.755 44.365 ;
        RECT -13.085 42.675 -12.755 43.005 ;
        RECT -13.085 41.315 -12.755 41.645 ;
        RECT -13.085 39.955 -12.755 40.285 ;
        RECT -13.085 38.595 -12.755 38.925 ;
        RECT -13.085 37.235 -12.755 37.565 ;
        RECT -13.085 35.875 -12.755 36.205 ;
        RECT -13.085 34.515 -12.755 34.845 ;
        RECT -13.085 33.155 -12.755 33.485 ;
        RECT -13.085 31.795 -12.755 32.125 ;
        RECT -13.085 30.435 -12.755 30.765 ;
        RECT -13.085 29.075 -12.755 29.405 ;
        RECT -13.085 27.715 -12.755 28.045 ;
        RECT -13.085 26.355 -12.755 26.685 ;
        RECT -13.085 24.995 -12.755 25.325 ;
        RECT -13.085 23.635 -12.755 23.965 ;
        RECT -13.085 22.275 -12.755 22.605 ;
        RECT -13.085 20.915 -12.755 21.245 ;
        RECT -13.085 19.555 -12.755 19.885 ;
        RECT -13.085 18.195 -12.755 18.525 ;
        RECT -13.085 16.835 -12.755 17.165 ;
        RECT -13.085 15.475 -12.755 15.805 ;
        RECT -13.085 14.115 -12.755 14.445 ;
        RECT -13.085 12.755 -12.755 13.085 ;
        RECT -13.085 11.395 -12.755 11.725 ;
        RECT -13.085 10.035 -12.755 10.365 ;
        RECT -13.085 8.675 -12.755 9.005 ;
        RECT -13.085 7.315 -12.755 7.645 ;
        RECT -13.085 5.955 -12.755 6.285 ;
        RECT -13.085 4.595 -12.755 4.925 ;
        RECT -13.085 3.235 -12.755 3.565 ;
        RECT -13.085 1.875 -12.755 2.205 ;
        RECT -13.085 0.515 -12.755 0.845 ;
        RECT -13.085 -0.845 -12.755 -0.515 ;
        RECT -13.085 -2.205 -12.755 -1.875 ;
        RECT -13.085 -3.565 -12.755 -3.235 ;
        RECT -13.085 -6.285 -12.755 -5.955 ;
        RECT -13.085 -8.19 -12.755 -7.86 ;
        RECT -13.085 -9.005 -12.755 -8.675 ;
        RECT -13.085 -11.725 -12.755 -11.395 ;
        RECT -13.085 -14.23 -12.755 -13.9 ;
        RECT -13.085 -15.805 -12.755 -15.475 ;
        RECT -13.085 -18.525 -12.755 -18.195 ;
        RECT -13.08 -18.525 -12.76 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 -82.47 -12.755 -82.14 ;
        RECT -13.085 -83.805 -12.755 -83.475 ;
        RECT -13.085 -85.165 -12.755 -84.835 ;
        RECT -13.085 -87.885 -12.755 -87.555 ;
        RECT -13.085 -91.965 -12.755 -91.635 ;
        RECT -13.085 -93.325 -12.755 -92.995 ;
        RECT -13.085 -94.685 -12.755 -94.355 ;
        RECT -13.085 -96.045 -12.755 -95.715 ;
        RECT -13.085 -97.405 -12.755 -97.075 ;
        RECT -13.085 -98.765 -12.755 -98.435 ;
        RECT -13.085 -113.725 -12.755 -113.395 ;
        RECT -13.085 -116.445 -12.755 -116.115 ;
        RECT -13.085 -120.525 -12.755 -120.195 ;
        RECT -13.085 -121.885 -12.755 -121.555 ;
        RECT -13.085 -125.965 -12.755 -125.635 ;
        RECT -13.085 -127.325 -12.755 -126.995 ;
        RECT -13.085 -128.685 -12.755 -128.355 ;
        RECT -13.085 -131.405 -12.755 -131.075 ;
        RECT -13.085 -132.765 -12.755 -132.435 ;
        RECT -13.085 -134.125 -12.755 -133.795 ;
        RECT -13.085 -135.485 -12.755 -135.155 ;
        RECT -13.085 -136.845 -12.755 -136.515 ;
        RECT -13.085 -138.205 -12.755 -137.875 ;
        RECT -13.085 -139.565 -12.755 -139.235 ;
        RECT -13.085 -140.925 -12.755 -140.595 ;
        RECT -13.085 -142.285 -12.755 -141.955 ;
        RECT -13.085 -143.645 -12.755 -143.315 ;
        RECT -13.085 -145.005 -12.755 -144.675 ;
        RECT -13.085 -146.365 -12.755 -146.035 ;
        RECT -13.085 -148.215 -12.755 -147.885 ;
        RECT -13.085 -149.085 -12.755 -148.755 ;
        RECT -13.085 -150.445 -12.755 -150.115 ;
        RECT -13.085 -151.805 -12.755 -151.475 ;
        RECT -13.085 -153.165 -12.755 -152.835 ;
        RECT -13.085 -154.525 -12.755 -154.195 ;
        RECT -13.085 -157.245 -12.755 -156.915 ;
        RECT -13.085 -162.89 -12.755 -161.76 ;
        RECT -13.08 -163.005 -12.76 -80.76 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.725 129.945 -11.395 131.075 ;
        RECT -11.725 125.635 -11.395 125.965 ;
        RECT -11.725 124.275 -11.395 124.605 ;
        RECT -11.725 122.915 -11.395 123.245 ;
        RECT -11.725 121.555 -11.395 121.885 ;
        RECT -11.725 120.195 -11.395 120.525 ;
        RECT -11.725 118.835 -11.395 119.165 ;
        RECT -11.725 117.475 -11.395 117.805 ;
        RECT -11.725 116.115 -11.395 116.445 ;
        RECT -11.725 114.755 -11.395 115.085 ;
        RECT -11.725 113.395 -11.395 113.725 ;
        RECT -11.725 112.035 -11.395 112.365 ;
        RECT -11.725 110.675 -11.395 111.005 ;
        RECT -11.725 109.315 -11.395 109.645 ;
        RECT -11.725 107.955 -11.395 108.285 ;
        RECT -11.725 106.595 -11.395 106.925 ;
        RECT -11.725 105.235 -11.395 105.565 ;
        RECT -11.725 103.875 -11.395 104.205 ;
        RECT -11.725 102.515 -11.395 102.845 ;
        RECT -11.725 101.155 -11.395 101.485 ;
        RECT -11.725 99.795 -11.395 100.125 ;
        RECT -11.725 98.435 -11.395 98.765 ;
        RECT -11.725 97.075 -11.395 97.405 ;
        RECT -11.725 95.715 -11.395 96.045 ;
        RECT -11.725 94.355 -11.395 94.685 ;
        RECT -11.725 92.995 -11.395 93.325 ;
        RECT -11.725 91.635 -11.395 91.965 ;
        RECT -11.725 90.275 -11.395 90.605 ;
        RECT -11.725 88.915 -11.395 89.245 ;
        RECT -11.725 87.555 -11.395 87.885 ;
        RECT -11.725 86.195 -11.395 86.525 ;
        RECT -11.725 84.835 -11.395 85.165 ;
        RECT -11.725 83.475 -11.395 83.805 ;
        RECT -11.725 82.115 -11.395 82.445 ;
        RECT -11.725 80.755 -11.395 81.085 ;
        RECT -11.725 79.395 -11.395 79.725 ;
        RECT -11.725 78.035 -11.395 78.365 ;
        RECT -11.725 76.675 -11.395 77.005 ;
        RECT -11.725 75.315 -11.395 75.645 ;
        RECT -11.725 73.955 -11.395 74.285 ;
        RECT -11.725 72.595 -11.395 72.925 ;
        RECT -11.725 71.235 -11.395 71.565 ;
        RECT -11.725 69.875 -11.395 70.205 ;
        RECT -11.725 68.515 -11.395 68.845 ;
        RECT -11.725 67.155 -11.395 67.485 ;
        RECT -11.725 65.795 -11.395 66.125 ;
        RECT -11.725 64.435 -11.395 64.765 ;
        RECT -11.725 63.075 -11.395 63.405 ;
        RECT -11.725 61.715 -11.395 62.045 ;
        RECT -11.725 60.355 -11.395 60.685 ;
        RECT -11.725 58.995 -11.395 59.325 ;
        RECT -11.725 57.635 -11.395 57.965 ;
        RECT -11.725 56.275 -11.395 56.605 ;
        RECT -11.725 54.915 -11.395 55.245 ;
        RECT -11.725 53.555 -11.395 53.885 ;
        RECT -11.725 52.195 -11.395 52.525 ;
        RECT -11.725 50.835 -11.395 51.165 ;
        RECT -11.725 49.475 -11.395 49.805 ;
        RECT -11.725 48.115 -11.395 48.445 ;
        RECT -11.725 46.755 -11.395 47.085 ;
        RECT -11.725 45.395 -11.395 45.725 ;
        RECT -11.725 44.035 -11.395 44.365 ;
        RECT -11.725 42.675 -11.395 43.005 ;
        RECT -11.725 41.315 -11.395 41.645 ;
        RECT -11.725 39.955 -11.395 40.285 ;
        RECT -11.725 38.595 -11.395 38.925 ;
        RECT -11.725 37.235 -11.395 37.565 ;
        RECT -11.725 35.875 -11.395 36.205 ;
        RECT -11.725 34.515 -11.395 34.845 ;
        RECT -11.725 33.155 -11.395 33.485 ;
        RECT -11.725 31.795 -11.395 32.125 ;
        RECT -11.725 30.435 -11.395 30.765 ;
        RECT -11.725 29.075 -11.395 29.405 ;
        RECT -11.725 27.715 -11.395 28.045 ;
        RECT -11.725 26.355 -11.395 26.685 ;
        RECT -11.725 24.995 -11.395 25.325 ;
        RECT -11.725 23.635 -11.395 23.965 ;
        RECT -11.725 22.275 -11.395 22.605 ;
        RECT -11.725 20.915 -11.395 21.245 ;
        RECT -11.725 19.555 -11.395 19.885 ;
        RECT -11.725 18.195 -11.395 18.525 ;
        RECT -11.725 16.835 -11.395 17.165 ;
        RECT -11.725 15.475 -11.395 15.805 ;
        RECT -11.725 14.115 -11.395 14.445 ;
        RECT -11.725 12.755 -11.395 13.085 ;
        RECT -11.725 11.395 -11.395 11.725 ;
        RECT -11.725 10.035 -11.395 10.365 ;
        RECT -11.725 8.675 -11.395 9.005 ;
        RECT -11.725 7.315 -11.395 7.645 ;
        RECT -11.725 5.955 -11.395 6.285 ;
        RECT -11.725 4.595 -11.395 4.925 ;
        RECT -11.725 3.235 -11.395 3.565 ;
        RECT -11.725 1.875 -11.395 2.205 ;
        RECT -11.725 0.515 -11.395 0.845 ;
        RECT -11.725 -0.845 -11.395 -0.515 ;
        RECT -11.725 -2.205 -11.395 -1.875 ;
        RECT -11.725 -3.565 -11.395 -3.235 ;
        RECT -11.725 -4.925 -11.395 -4.595 ;
        RECT -11.725 -6.285 -11.395 -5.955 ;
        RECT -11.725 -8.19 -11.395 -7.86 ;
        RECT -11.725 -9.005 -11.395 -8.675 ;
        RECT -11.725 -10.365 -11.395 -10.035 ;
        RECT -11.725 -11.725 -11.395 -11.395 ;
        RECT -11.725 -14.23 -11.395 -13.9 ;
        RECT -11.725 -15.805 -11.395 -15.475 ;
        RECT -11.72 -17.84 -11.4 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.725 -91.965 -11.395 -91.635 ;
        RECT -11.725 -93.325 -11.395 -92.995 ;
        RECT -11.725 -94.685 -11.395 -94.355 ;
        RECT -11.725 -96.045 -11.395 -95.715 ;
        RECT -11.725 -97.405 -11.395 -97.075 ;
        RECT -11.725 -98.765 -11.395 -98.435 ;
        RECT -11.725 -101.485 -11.395 -101.155 ;
        RECT -11.725 -105.565 -11.395 -105.235 ;
        RECT -11.725 -106.925 -11.395 -106.595 ;
        RECT -11.725 -109.645 -11.395 -109.315 ;
        RECT -11.725 -111.005 -11.395 -110.675 ;
        RECT -11.725 -113.725 -11.395 -113.395 ;
        RECT -11.725 -115.085 -11.395 -114.755 ;
        RECT -11.725 -116.445 -11.395 -116.115 ;
        RECT -11.725 -117.805 -11.395 -117.475 ;
        RECT -11.725 -119.165 -11.395 -118.835 ;
        RECT -11.725 -120.525 -11.395 -120.195 ;
        RECT -11.725 -121.885 -11.395 -121.555 ;
        RECT -11.725 -125.965 -11.395 -125.635 ;
        RECT -11.725 -127.325 -11.395 -126.995 ;
        RECT -11.725 -128.685 -11.395 -128.355 ;
        RECT -11.725 -130.045 -11.395 -129.715 ;
        RECT -11.725 -131.405 -11.395 -131.075 ;
        RECT -11.725 -132.765 -11.395 -132.435 ;
        RECT -11.725 -134.125 -11.395 -133.795 ;
        RECT -11.725 -135.485 -11.395 -135.155 ;
        RECT -11.725 -136.845 -11.395 -136.515 ;
        RECT -11.725 -138.205 -11.395 -137.875 ;
        RECT -11.725 -139.565 -11.395 -139.235 ;
        RECT -11.725 -140.925 -11.395 -140.595 ;
        RECT -11.725 -142.285 -11.395 -141.955 ;
        RECT -11.725 -143.645 -11.395 -143.315 ;
        RECT -11.725 -145.005 -11.395 -144.675 ;
        RECT -11.725 -146.365 -11.395 -146.035 ;
        RECT -11.725 -148.215 -11.395 -147.885 ;
        RECT -11.725 -149.085 -11.395 -148.755 ;
        RECT -11.725 -150.445 -11.395 -150.115 ;
        RECT -11.725 -151.805 -11.395 -151.475 ;
        RECT -11.725 -153.165 -11.395 -152.835 ;
        RECT -11.725 -154.525 -11.395 -154.195 ;
        RECT -11.725 -157.245 -11.395 -156.915 ;
        RECT -11.725 -162.89 -11.395 -161.76 ;
        RECT -11.72 -163.005 -11.4 -88.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 -53.885 -10.035 -53.555 ;
        RECT -10.365 -55.245 -10.035 -54.915 ;
        RECT -10.365 -57.965 -10.035 -57.635 ;
        RECT -10.365 -59.325 -10.035 -58.995 ;
        RECT -10.365 -60.29 -10.035 -59.96 ;
        RECT -10.365 -62.045 -10.035 -61.715 ;
        RECT -10.365 -63.405 -10.035 -63.075 ;
        RECT -10.365 -66.125 -10.035 -65.795 ;
        RECT -10.365 -68.845 -10.035 -68.515 ;
        RECT -10.365 -70.205 -10.035 -69.875 ;
        RECT -10.365 -71.565 -10.035 -71.235 ;
        RECT -10.365 -72.925 -10.035 -72.595 ;
        RECT -10.365 -74.93 -10.035 -74.6 ;
        RECT -10.365 -75.645 -10.035 -75.315 ;
        RECT -10.365 -77.005 -10.035 -76.675 ;
        RECT -10.365 -79.725 -10.035 -79.395 ;
        RECT -10.365 -82.47 -10.035 -82.14 ;
        RECT -10.365 -83.805 -10.035 -83.475 ;
        RECT -10.365 -85.165 -10.035 -84.835 ;
        RECT -10.365 -87.885 -10.035 -87.555 ;
        RECT -10.365 -91.965 -10.035 -91.635 ;
        RECT -10.365 -93.325 -10.035 -92.995 ;
        RECT -10.365 -94.685 -10.035 -94.355 ;
        RECT -10.365 -96.045 -10.035 -95.715 ;
        RECT -10.365 -97.405 -10.035 -97.075 ;
        RECT -10.365 -98.765 -10.035 -98.435 ;
        RECT -10.365 -101.485 -10.035 -101.155 ;
        RECT -10.365 -105.565 -10.035 -105.235 ;
        RECT -10.365 -106.925 -10.035 -106.595 ;
        RECT -10.365 -109.645 -10.035 -109.315 ;
        RECT -10.365 -111.005 -10.035 -110.675 ;
        RECT -10.365 -113.725 -10.035 -113.395 ;
        RECT -10.365 -115.085 -10.035 -114.755 ;
        RECT -10.365 -116.445 -10.035 -116.115 ;
        RECT -10.365 -117.805 -10.035 -117.475 ;
        RECT -10.365 -119.165 -10.035 -118.835 ;
        RECT -10.365 -120.525 -10.035 -120.195 ;
        RECT -10.365 -121.885 -10.035 -121.555 ;
        RECT -10.365 -125.965 -10.035 -125.635 ;
        RECT -10.365 -127.325 -10.035 -126.995 ;
        RECT -10.365 -128.685 -10.035 -128.355 ;
        RECT -10.365 -130.045 -10.035 -129.715 ;
        RECT -10.365 -131.405 -10.035 -131.075 ;
        RECT -10.365 -132.765 -10.035 -132.435 ;
        RECT -10.365 -134.125 -10.035 -133.795 ;
        RECT -10.365 -135.485 -10.035 -135.155 ;
        RECT -10.365 -136.845 -10.035 -136.515 ;
        RECT -10.365 -138.205 -10.035 -137.875 ;
        RECT -10.365 -139.565 -10.035 -139.235 ;
        RECT -10.365 -140.925 -10.035 -140.595 ;
        RECT -10.365 -142.285 -10.035 -141.955 ;
        RECT -10.365 -143.645 -10.035 -143.315 ;
        RECT -10.365 -145.005 -10.035 -144.675 ;
        RECT -10.365 -146.365 -10.035 -146.035 ;
        RECT -10.36 -146.365 -10.04 131.19 ;
        RECT -10.365 129.945 -10.035 131.075 ;
        RECT -10.365 125.635 -10.035 125.965 ;
        RECT -10.365 124.275 -10.035 124.605 ;
        RECT -10.365 122.915 -10.035 123.245 ;
        RECT -10.365 121.555 -10.035 121.885 ;
        RECT -10.365 120.195 -10.035 120.525 ;
        RECT -10.365 118.835 -10.035 119.165 ;
        RECT -10.365 117.475 -10.035 117.805 ;
        RECT -10.365 110.675 -10.035 111.005 ;
        RECT -10.365 107.955 -10.035 108.285 ;
        RECT -10.365 103.875 -10.035 104.205 ;
        RECT -10.365 99.795 -10.035 100.125 ;
        RECT -10.365 97.075 -10.035 97.405 ;
        RECT -10.365 90.275 -10.035 90.605 ;
        RECT -10.365 88.915 -10.035 89.245 ;
        RECT -10.365 82.115 -10.035 82.445 ;
        RECT -10.365 79.395 -10.035 79.725 ;
        RECT -10.365 75.315 -10.035 75.645 ;
        RECT -10.365 71.235 -10.035 71.565 ;
        RECT -10.365 68.515 -10.035 68.845 ;
        RECT -10.365 61.715 -10.035 62.045 ;
        RECT -10.365 60.355 -10.035 60.685 ;
        RECT -10.365 50.835 -10.035 51.165 ;
        RECT -10.365 46.755 -10.035 47.085 ;
        RECT -10.365 42.675 -10.035 43.005 ;
        RECT -10.365 39.955 -10.035 40.285 ;
        RECT -10.365 33.155 -10.035 33.485 ;
        RECT -10.365 31.795 -10.035 32.125 ;
        RECT -10.365 29.075 -10.035 29.405 ;
        RECT -10.365 22.275 -10.035 22.605 ;
        RECT -10.365 19.555 -10.035 19.885 ;
        RECT -10.365 18.195 -10.035 18.525 ;
        RECT -10.365 11.395 -10.035 11.725 ;
        RECT -10.365 4.595 -10.035 4.925 ;
        RECT -10.365 3.235 -10.035 3.565 ;
        RECT -10.365 1.875 -10.035 2.205 ;
        RECT -10.365 0.515 -10.035 0.845 ;
        RECT -10.365 -0.845 -10.035 -0.515 ;
        RECT -10.365 -2.205 -10.035 -1.875 ;
        RECT -10.365 -3.565 -10.035 -3.235 ;
        RECT -10.365 -4.925 -10.035 -4.595 ;
        RECT -10.365 -6.285 -10.035 -5.955 ;
        RECT -10.365 -8.19 -10.035 -7.86 ;
        RECT -10.365 -9.005 -10.035 -8.675 ;
        RECT -10.365 -10.365 -10.035 -10.035 ;
        RECT -10.365 -11.725 -10.035 -11.395 ;
        RECT -10.365 -14.23 -10.035 -13.9 ;
        RECT -10.365 -15.805 -10.035 -15.475 ;
        RECT -10.365 -23.965 -10.035 -23.635 ;
        RECT -10.365 -25.325 -10.035 -24.995 ;
        RECT -10.365 -26.685 -10.035 -26.355 ;
        RECT -10.365 -28.045 -10.035 -27.715 ;
        RECT -10.365 -29.405 -10.035 -29.075 ;
        RECT -10.365 -31.17 -10.035 -30.84 ;
        RECT -10.365 -32.125 -10.035 -31.795 ;
        RECT -10.365 -33.485 -10.035 -33.155 ;
        RECT -10.365 -36.205 -10.035 -35.875 ;
        RECT -10.365 -37.21 -10.035 -36.88 ;
        RECT -10.365 -38.925 -10.035 -38.595 ;
        RECT -10.365 -41.645 -10.035 -41.315 ;
        RECT -10.365 -49.805 -10.035 -49.475 ;
        RECT -10.365 -51.165 -10.035 -50.835 ;
        RECT -10.365 -52.75 -10.035 -52.42 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 129.945 -26.355 131.075 ;
        RECT -26.685 125.635 -26.355 125.965 ;
        RECT -26.685 124.275 -26.355 124.605 ;
        RECT -26.685 122.915 -26.355 123.245 ;
        RECT -26.685 121.555 -26.355 121.885 ;
        RECT -26.685 120.195 -26.355 120.525 ;
        RECT -26.685 118.835 -26.355 119.165 ;
        RECT -26.685 117.475 -26.355 117.805 ;
        RECT -26.685 116.115 -26.355 116.445 ;
        RECT -26.685 114.755 -26.355 115.085 ;
        RECT -26.685 113.395 -26.355 113.725 ;
        RECT -26.685 112.035 -26.355 112.365 ;
        RECT -26.685 110.675 -26.355 111.005 ;
        RECT -26.685 109.315 -26.355 109.645 ;
        RECT -26.685 107.955 -26.355 108.285 ;
        RECT -26.685 106.595 -26.355 106.925 ;
        RECT -26.685 105.235 -26.355 105.565 ;
        RECT -26.685 103.875 -26.355 104.205 ;
        RECT -26.685 102.515 -26.355 102.845 ;
        RECT -26.685 101.155 -26.355 101.485 ;
        RECT -26.685 99.795 -26.355 100.125 ;
        RECT -26.685 98.435 -26.355 98.765 ;
        RECT -26.685 97.075 -26.355 97.405 ;
        RECT -26.685 95.715 -26.355 96.045 ;
        RECT -26.685 94.355 -26.355 94.685 ;
        RECT -26.685 92.995 -26.355 93.325 ;
        RECT -26.685 91.635 -26.355 91.965 ;
        RECT -26.685 90.275 -26.355 90.605 ;
        RECT -26.685 88.915 -26.355 89.245 ;
        RECT -26.685 87.555 -26.355 87.885 ;
        RECT -26.685 86.195 -26.355 86.525 ;
        RECT -26.685 84.835 -26.355 85.165 ;
        RECT -26.685 83.475 -26.355 83.805 ;
        RECT -26.685 82.115 -26.355 82.445 ;
        RECT -26.685 80.755 -26.355 81.085 ;
        RECT -26.685 79.395 -26.355 79.725 ;
        RECT -26.685 78.035 -26.355 78.365 ;
        RECT -26.685 76.675 -26.355 77.005 ;
        RECT -26.685 75.315 -26.355 75.645 ;
        RECT -26.685 73.955 -26.355 74.285 ;
        RECT -26.685 72.595 -26.355 72.925 ;
        RECT -26.685 71.235 -26.355 71.565 ;
        RECT -26.685 69.875 -26.355 70.205 ;
        RECT -26.685 68.515 -26.355 68.845 ;
        RECT -26.685 67.155 -26.355 67.485 ;
        RECT -26.685 65.795 -26.355 66.125 ;
        RECT -26.685 64.435 -26.355 64.765 ;
        RECT -26.685 63.075 -26.355 63.405 ;
        RECT -26.685 61.715 -26.355 62.045 ;
        RECT -26.685 60.355 -26.355 60.685 ;
        RECT -26.685 58.995 -26.355 59.325 ;
        RECT -26.685 57.635 -26.355 57.965 ;
        RECT -26.685 56.275 -26.355 56.605 ;
        RECT -26.685 54.915 -26.355 55.245 ;
        RECT -26.685 53.555 -26.355 53.885 ;
        RECT -26.685 52.195 -26.355 52.525 ;
        RECT -26.685 50.835 -26.355 51.165 ;
        RECT -26.685 49.475 -26.355 49.805 ;
        RECT -26.685 48.115 -26.355 48.445 ;
        RECT -26.685 46.755 -26.355 47.085 ;
        RECT -26.685 45.395 -26.355 45.725 ;
        RECT -26.685 44.035 -26.355 44.365 ;
        RECT -26.685 42.675 -26.355 43.005 ;
        RECT -26.685 41.315 -26.355 41.645 ;
        RECT -26.685 39.955 -26.355 40.285 ;
        RECT -26.685 38.595 -26.355 38.925 ;
        RECT -26.685 37.235 -26.355 37.565 ;
        RECT -26.685 35.875 -26.355 36.205 ;
        RECT -26.685 34.515 -26.355 34.845 ;
        RECT -26.685 33.155 -26.355 33.485 ;
        RECT -26.685 31.795 -26.355 32.125 ;
        RECT -26.685 30.435 -26.355 30.765 ;
        RECT -26.685 29.075 -26.355 29.405 ;
        RECT -26.685 27.715 -26.355 28.045 ;
        RECT -26.685 26.355 -26.355 26.685 ;
        RECT -26.685 24.995 -26.355 25.325 ;
        RECT -26.685 23.635 -26.355 23.965 ;
        RECT -26.685 22.275 -26.355 22.605 ;
        RECT -26.685 20.915 -26.355 21.245 ;
        RECT -26.685 19.555 -26.355 19.885 ;
        RECT -26.685 18.195 -26.355 18.525 ;
        RECT -26.685 16.835 -26.355 17.165 ;
        RECT -26.685 15.475 -26.355 15.805 ;
        RECT -26.685 14.115 -26.355 14.445 ;
        RECT -26.685 12.755 -26.355 13.085 ;
        RECT -26.685 11.395 -26.355 11.725 ;
        RECT -26.685 10.035 -26.355 10.365 ;
        RECT -26.685 8.675 -26.355 9.005 ;
        RECT -26.685 7.315 -26.355 7.645 ;
        RECT -26.685 5.955 -26.355 6.285 ;
        RECT -26.685 4.595 -26.355 4.925 ;
        RECT -26.685 3.235 -26.355 3.565 ;
        RECT -26.685 1.875 -26.355 2.205 ;
        RECT -26.685 0.515 -26.355 0.845 ;
        RECT -26.685 -0.845 -26.355 -0.515 ;
        RECT -26.68 -5.6 -26.36 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 -29.405 -26.355 -29.075 ;
        RECT -26.685 -31.17 -26.355 -30.84 ;
        RECT -26.685 -32.125 -26.355 -31.795 ;
        RECT -26.685 -33.485 -26.355 -33.155 ;
        RECT -26.685 -36.205 -26.355 -35.875 ;
        RECT -26.685 -37.21 -26.355 -36.88 ;
        RECT -26.685 -38.925 -26.355 -38.595 ;
        RECT -26.685 -41.645 -26.355 -41.315 ;
        RECT -26.685 -51.165 -26.355 -50.835 ;
        RECT -26.685 -52.525 -26.355 -52.195 ;
        RECT -26.685 -53.885 -26.355 -53.555 ;
        RECT -26.685 -55.245 -26.355 -54.915 ;
        RECT -26.685 -56.605 -26.355 -56.275 ;
        RECT -26.685 -57.965 -26.355 -57.635 ;
        RECT -26.685 -59.325 -26.355 -58.995 ;
        RECT -26.685 -60.685 -26.355 -60.355 ;
        RECT -26.685 -62.045 -26.355 -61.715 ;
        RECT -26.685 -63.405 -26.355 -63.075 ;
        RECT -26.685 -64.765 -26.355 -64.435 ;
        RECT -26.685 -66.125 -26.355 -65.795 ;
        RECT -26.685 -67.485 -26.355 -67.155 ;
        RECT -26.685 -68.845 -26.355 -68.515 ;
        RECT -26.685 -71.565 -26.355 -71.235 ;
        RECT -26.685 -72.925 -26.355 -72.595 ;
        RECT -26.685 -74.285 -26.355 -73.955 ;
        RECT -26.685 -75.645 -26.355 -75.315 ;
        RECT -26.685 -77.005 -26.355 -76.675 ;
        RECT -26.685 -79.725 -26.355 -79.395 ;
        RECT -26.685 -82.445 -26.355 -82.115 ;
        RECT -26.685 -83.805 -26.355 -83.475 ;
        RECT -26.685 -85.165 -26.355 -84.835 ;
        RECT -26.685 -87.885 -26.355 -87.555 ;
        RECT -26.685 -89.245 -26.355 -88.915 ;
        RECT -26.685 -91.965 -26.355 -91.635 ;
        RECT -26.685 -93.325 -26.355 -92.995 ;
        RECT -26.685 -94.685 -26.355 -94.355 ;
        RECT -26.685 -96.045 -26.355 -95.715 ;
        RECT -26.685 -98.765 -26.355 -98.435 ;
        RECT -26.685 -100.125 -26.355 -99.795 ;
        RECT -26.685 -101.485 -26.355 -101.155 ;
        RECT -26.685 -102.845 -26.355 -102.515 ;
        RECT -26.685 -105.565 -26.355 -105.235 ;
        RECT -26.685 -106.925 -26.355 -106.595 ;
        RECT -26.685 -108.285 -26.355 -107.955 ;
        RECT -26.685 -113.725 -26.355 -113.395 ;
        RECT -26.685 -115.085 -26.355 -114.755 ;
        RECT -26.685 -117.805 -26.355 -117.475 ;
        RECT -26.685 -120.525 -26.355 -120.195 ;
        RECT -26.685 -121.885 -26.355 -121.555 ;
        RECT -26.685 -123.245 -26.355 -122.915 ;
        RECT -26.685 -125.965 -26.355 -125.635 ;
        RECT -26.685 -127.325 -26.355 -126.995 ;
        RECT -26.685 -131.405 -26.355 -131.075 ;
        RECT -26.685 -135.485 -26.355 -135.155 ;
        RECT -26.685 -136.845 -26.355 -136.515 ;
        RECT -26.685 -138.205 -26.355 -137.875 ;
        RECT -26.685 -139.565 -26.355 -139.235 ;
        RECT -26.685 -140.925 -26.355 -140.595 ;
        RECT -26.685 -142.285 -26.355 -141.955 ;
        RECT -26.685 -143.645 -26.355 -143.315 ;
        RECT -26.685 -145.005 -26.355 -144.675 ;
        RECT -26.685 -146.365 -26.355 -146.035 ;
        RECT -26.685 -148.215 -26.355 -147.885 ;
        RECT -26.685 -149.085 -26.355 -148.755 ;
        RECT -26.685 -150.445 -26.355 -150.115 ;
        RECT -26.685 -153.165 -26.355 -152.835 ;
        RECT -26.685 -154.525 -26.355 -154.195 ;
        RECT -26.685 -157.245 -26.355 -156.915 ;
        RECT -26.685 -162.89 -26.355 -161.76 ;
        RECT -26.68 -163.005 -26.36 -27.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.325 129.945 -24.995 131.075 ;
        RECT -25.325 125.635 -24.995 125.965 ;
        RECT -25.325 124.275 -24.995 124.605 ;
        RECT -25.325 122.915 -24.995 123.245 ;
        RECT -25.325 121.555 -24.995 121.885 ;
        RECT -25.325 120.195 -24.995 120.525 ;
        RECT -25.325 118.835 -24.995 119.165 ;
        RECT -25.325 117.475 -24.995 117.805 ;
        RECT -25.325 116.115 -24.995 116.445 ;
        RECT -25.325 114.755 -24.995 115.085 ;
        RECT -25.325 113.395 -24.995 113.725 ;
        RECT -25.325 112.035 -24.995 112.365 ;
        RECT -25.325 110.675 -24.995 111.005 ;
        RECT -25.325 109.315 -24.995 109.645 ;
        RECT -25.325 107.955 -24.995 108.285 ;
        RECT -25.325 106.595 -24.995 106.925 ;
        RECT -25.325 105.235 -24.995 105.565 ;
        RECT -25.325 103.875 -24.995 104.205 ;
        RECT -25.325 102.515 -24.995 102.845 ;
        RECT -25.325 101.155 -24.995 101.485 ;
        RECT -25.325 99.795 -24.995 100.125 ;
        RECT -25.325 98.435 -24.995 98.765 ;
        RECT -25.325 97.075 -24.995 97.405 ;
        RECT -25.325 95.715 -24.995 96.045 ;
        RECT -25.325 94.355 -24.995 94.685 ;
        RECT -25.325 92.995 -24.995 93.325 ;
        RECT -25.325 91.635 -24.995 91.965 ;
        RECT -25.325 90.275 -24.995 90.605 ;
        RECT -25.325 88.915 -24.995 89.245 ;
        RECT -25.325 87.555 -24.995 87.885 ;
        RECT -25.325 86.195 -24.995 86.525 ;
        RECT -25.325 84.835 -24.995 85.165 ;
        RECT -25.325 83.475 -24.995 83.805 ;
        RECT -25.325 82.115 -24.995 82.445 ;
        RECT -25.325 80.755 -24.995 81.085 ;
        RECT -25.325 79.395 -24.995 79.725 ;
        RECT -25.325 78.035 -24.995 78.365 ;
        RECT -25.325 76.675 -24.995 77.005 ;
        RECT -25.325 75.315 -24.995 75.645 ;
        RECT -25.325 73.955 -24.995 74.285 ;
        RECT -25.325 72.595 -24.995 72.925 ;
        RECT -25.325 71.235 -24.995 71.565 ;
        RECT -25.325 69.875 -24.995 70.205 ;
        RECT -25.325 68.515 -24.995 68.845 ;
        RECT -25.325 67.155 -24.995 67.485 ;
        RECT -25.325 65.795 -24.995 66.125 ;
        RECT -25.325 64.435 -24.995 64.765 ;
        RECT -25.325 63.075 -24.995 63.405 ;
        RECT -25.325 61.715 -24.995 62.045 ;
        RECT -25.325 60.355 -24.995 60.685 ;
        RECT -25.325 58.995 -24.995 59.325 ;
        RECT -25.325 57.635 -24.995 57.965 ;
        RECT -25.325 56.275 -24.995 56.605 ;
        RECT -25.325 54.915 -24.995 55.245 ;
        RECT -25.325 53.555 -24.995 53.885 ;
        RECT -25.325 52.195 -24.995 52.525 ;
        RECT -25.325 50.835 -24.995 51.165 ;
        RECT -25.325 49.475 -24.995 49.805 ;
        RECT -25.325 48.115 -24.995 48.445 ;
        RECT -25.325 46.755 -24.995 47.085 ;
        RECT -25.325 45.395 -24.995 45.725 ;
        RECT -25.325 44.035 -24.995 44.365 ;
        RECT -25.325 42.675 -24.995 43.005 ;
        RECT -25.325 41.315 -24.995 41.645 ;
        RECT -25.325 39.955 -24.995 40.285 ;
        RECT -25.325 38.595 -24.995 38.925 ;
        RECT -25.325 37.235 -24.995 37.565 ;
        RECT -25.325 35.875 -24.995 36.205 ;
        RECT -25.325 34.515 -24.995 34.845 ;
        RECT -25.325 33.155 -24.995 33.485 ;
        RECT -25.325 31.795 -24.995 32.125 ;
        RECT -25.325 30.435 -24.995 30.765 ;
        RECT -25.325 29.075 -24.995 29.405 ;
        RECT -25.325 27.715 -24.995 28.045 ;
        RECT -25.325 26.355 -24.995 26.685 ;
        RECT -25.325 24.995 -24.995 25.325 ;
        RECT -25.325 23.635 -24.995 23.965 ;
        RECT -25.325 22.275 -24.995 22.605 ;
        RECT -25.325 20.915 -24.995 21.245 ;
        RECT -25.325 19.555 -24.995 19.885 ;
        RECT -25.325 18.195 -24.995 18.525 ;
        RECT -25.325 16.835 -24.995 17.165 ;
        RECT -25.325 15.475 -24.995 15.805 ;
        RECT -25.325 14.115 -24.995 14.445 ;
        RECT -25.325 12.755 -24.995 13.085 ;
        RECT -25.325 11.395 -24.995 11.725 ;
        RECT -25.325 10.035 -24.995 10.365 ;
        RECT -25.325 8.675 -24.995 9.005 ;
        RECT -25.325 7.315 -24.995 7.645 ;
        RECT -25.325 5.955 -24.995 6.285 ;
        RECT -25.325 4.595 -24.995 4.925 ;
        RECT -25.325 3.235 -24.995 3.565 ;
        RECT -25.325 1.875 -24.995 2.205 ;
        RECT -25.325 0.515 -24.995 0.845 ;
        RECT -25.325 -0.845 -24.995 -0.515 ;
        RECT -25.325 -6.285 -24.995 -5.955 ;
        RECT -25.325 -8.19 -24.995 -7.86 ;
        RECT -25.325 -11.725 -24.995 -11.395 ;
        RECT -25.325 -14.23 -24.995 -13.9 ;
        RECT -25.325 -15.805 -24.995 -15.475 ;
        RECT -25.325 -28.045 -24.995 -27.715 ;
        RECT -25.325 -29.405 -24.995 -29.075 ;
        RECT -25.325 -31.17 -24.995 -30.84 ;
        RECT -25.325 -32.125 -24.995 -31.795 ;
        RECT -25.325 -33.485 -24.995 -33.155 ;
        RECT -25.325 -36.205 -24.995 -35.875 ;
        RECT -25.325 -37.21 -24.995 -36.88 ;
        RECT -25.325 -38.925 -24.995 -38.595 ;
        RECT -25.325 -41.645 -24.995 -41.315 ;
        RECT -25.325 -51.165 -24.995 -50.835 ;
        RECT -25.325 -52.525 -24.995 -52.195 ;
        RECT -25.325 -53.885 -24.995 -53.555 ;
        RECT -25.325 -55.245 -24.995 -54.915 ;
        RECT -25.325 -56.605 -24.995 -56.275 ;
        RECT -25.325 -57.965 -24.995 -57.635 ;
        RECT -25.325 -59.325 -24.995 -58.995 ;
        RECT -25.325 -60.685 -24.995 -60.355 ;
        RECT -25.325 -62.045 -24.995 -61.715 ;
        RECT -25.325 -63.405 -24.995 -63.075 ;
        RECT -25.325 -64.765 -24.995 -64.435 ;
        RECT -25.325 -66.125 -24.995 -65.795 ;
        RECT -25.325 -67.485 -24.995 -67.155 ;
        RECT -25.325 -68.845 -24.995 -68.515 ;
        RECT -25.325 -70.205 -24.995 -69.875 ;
        RECT -25.325 -71.565 -24.995 -71.235 ;
        RECT -25.325 -72.925 -24.995 -72.595 ;
        RECT -25.325 -74.285 -24.995 -73.955 ;
        RECT -25.325 -75.645 -24.995 -75.315 ;
        RECT -25.325 -77.005 -24.995 -76.675 ;
        RECT -25.325 -78.365 -24.995 -78.035 ;
        RECT -25.325 -79.725 -24.995 -79.395 ;
        RECT -25.325 -81.085 -24.995 -80.755 ;
        RECT -25.325 -82.445 -24.995 -82.115 ;
        RECT -25.325 -83.805 -24.995 -83.475 ;
        RECT -25.325 -85.165 -24.995 -84.835 ;
        RECT -25.325 -86.525 -24.995 -86.195 ;
        RECT -25.325 -87.885 -24.995 -87.555 ;
        RECT -25.325 -89.245 -24.995 -88.915 ;
        RECT -25.325 -90.605 -24.995 -90.275 ;
        RECT -25.325 -91.965 -24.995 -91.635 ;
        RECT -25.325 -93.325 -24.995 -92.995 ;
        RECT -25.325 -94.685 -24.995 -94.355 ;
        RECT -25.325 -96.045 -24.995 -95.715 ;
        RECT -25.325 -98.765 -24.995 -98.435 ;
        RECT -25.325 -100.125 -24.995 -99.795 ;
        RECT -25.325 -101.485 -24.995 -101.155 ;
        RECT -25.325 -102.845 -24.995 -102.515 ;
        RECT -25.325 -104.205 -24.995 -103.875 ;
        RECT -25.325 -105.565 -24.995 -105.235 ;
        RECT -25.325 -106.925 -24.995 -106.595 ;
        RECT -25.325 -108.285 -24.995 -107.955 ;
        RECT -25.325 -113.725 -24.995 -113.395 ;
        RECT -25.325 -115.085 -24.995 -114.755 ;
        RECT -25.325 -117.805 -24.995 -117.475 ;
        RECT -25.325 -120.525 -24.995 -120.195 ;
        RECT -25.325 -121.885 -24.995 -121.555 ;
        RECT -25.325 -123.245 -24.995 -122.915 ;
        RECT -25.325 -125.965 -24.995 -125.635 ;
        RECT -25.325 -127.325 -24.995 -126.995 ;
        RECT -25.325 -131.405 -24.995 -131.075 ;
        RECT -25.325 -135.485 -24.995 -135.155 ;
        RECT -25.325 -136.845 -24.995 -136.515 ;
        RECT -25.325 -138.205 -24.995 -137.875 ;
        RECT -25.325 -139.565 -24.995 -139.235 ;
        RECT -25.325 -140.925 -24.995 -140.595 ;
        RECT -25.325 -142.285 -24.995 -141.955 ;
        RECT -25.325 -143.645 -24.995 -143.315 ;
        RECT -25.325 -145.005 -24.995 -144.675 ;
        RECT -25.325 -146.365 -24.995 -146.035 ;
        RECT -25.325 -148.215 -24.995 -147.885 ;
        RECT -25.325 -149.085 -24.995 -148.755 ;
        RECT -25.325 -150.445 -24.995 -150.115 ;
        RECT -25.325 -151.805 -24.995 -151.475 ;
        RECT -25.325 -153.165 -24.995 -152.835 ;
        RECT -25.325 -154.525 -24.995 -154.195 ;
        RECT -25.325 -157.245 -24.995 -156.915 ;
        RECT -25.325 -162.89 -24.995 -161.76 ;
        RECT -25.32 -163.005 -25 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.965 129.945 -23.635 131.075 ;
        RECT -23.965 125.635 -23.635 125.965 ;
        RECT -23.965 124.275 -23.635 124.605 ;
        RECT -23.965 122.915 -23.635 123.245 ;
        RECT -23.965 121.555 -23.635 121.885 ;
        RECT -23.965 120.195 -23.635 120.525 ;
        RECT -23.965 118.835 -23.635 119.165 ;
        RECT -23.965 117.475 -23.635 117.805 ;
        RECT -23.965 116.115 -23.635 116.445 ;
        RECT -23.965 114.755 -23.635 115.085 ;
        RECT -23.965 113.395 -23.635 113.725 ;
        RECT -23.965 112.035 -23.635 112.365 ;
        RECT -23.965 110.675 -23.635 111.005 ;
        RECT -23.965 109.315 -23.635 109.645 ;
        RECT -23.965 107.955 -23.635 108.285 ;
        RECT -23.965 106.595 -23.635 106.925 ;
        RECT -23.965 105.235 -23.635 105.565 ;
        RECT -23.965 103.875 -23.635 104.205 ;
        RECT -23.965 102.515 -23.635 102.845 ;
        RECT -23.965 101.155 -23.635 101.485 ;
        RECT -23.965 99.795 -23.635 100.125 ;
        RECT -23.965 98.435 -23.635 98.765 ;
        RECT -23.965 97.075 -23.635 97.405 ;
        RECT -23.965 95.715 -23.635 96.045 ;
        RECT -23.965 94.355 -23.635 94.685 ;
        RECT -23.965 92.995 -23.635 93.325 ;
        RECT -23.965 91.635 -23.635 91.965 ;
        RECT -23.965 90.275 -23.635 90.605 ;
        RECT -23.965 88.915 -23.635 89.245 ;
        RECT -23.965 87.555 -23.635 87.885 ;
        RECT -23.965 86.195 -23.635 86.525 ;
        RECT -23.965 84.835 -23.635 85.165 ;
        RECT -23.965 83.475 -23.635 83.805 ;
        RECT -23.965 82.115 -23.635 82.445 ;
        RECT -23.965 80.755 -23.635 81.085 ;
        RECT -23.965 79.395 -23.635 79.725 ;
        RECT -23.965 78.035 -23.635 78.365 ;
        RECT -23.965 76.675 -23.635 77.005 ;
        RECT -23.965 75.315 -23.635 75.645 ;
        RECT -23.965 73.955 -23.635 74.285 ;
        RECT -23.965 72.595 -23.635 72.925 ;
        RECT -23.965 71.235 -23.635 71.565 ;
        RECT -23.965 69.875 -23.635 70.205 ;
        RECT -23.965 68.515 -23.635 68.845 ;
        RECT -23.965 67.155 -23.635 67.485 ;
        RECT -23.965 65.795 -23.635 66.125 ;
        RECT -23.965 64.435 -23.635 64.765 ;
        RECT -23.965 63.075 -23.635 63.405 ;
        RECT -23.965 61.715 -23.635 62.045 ;
        RECT -23.965 60.355 -23.635 60.685 ;
        RECT -23.965 58.995 -23.635 59.325 ;
        RECT -23.965 57.635 -23.635 57.965 ;
        RECT -23.965 56.275 -23.635 56.605 ;
        RECT -23.965 54.915 -23.635 55.245 ;
        RECT -23.965 53.555 -23.635 53.885 ;
        RECT -23.965 52.195 -23.635 52.525 ;
        RECT -23.965 50.835 -23.635 51.165 ;
        RECT -23.965 49.475 -23.635 49.805 ;
        RECT -23.965 48.115 -23.635 48.445 ;
        RECT -23.965 46.755 -23.635 47.085 ;
        RECT -23.965 45.395 -23.635 45.725 ;
        RECT -23.965 44.035 -23.635 44.365 ;
        RECT -23.965 42.675 -23.635 43.005 ;
        RECT -23.965 41.315 -23.635 41.645 ;
        RECT -23.965 39.955 -23.635 40.285 ;
        RECT -23.965 38.595 -23.635 38.925 ;
        RECT -23.965 37.235 -23.635 37.565 ;
        RECT -23.965 35.875 -23.635 36.205 ;
        RECT -23.965 34.515 -23.635 34.845 ;
        RECT -23.965 33.155 -23.635 33.485 ;
        RECT -23.965 31.795 -23.635 32.125 ;
        RECT -23.965 30.435 -23.635 30.765 ;
        RECT -23.965 29.075 -23.635 29.405 ;
        RECT -23.965 27.715 -23.635 28.045 ;
        RECT -23.965 26.355 -23.635 26.685 ;
        RECT -23.965 24.995 -23.635 25.325 ;
        RECT -23.965 23.635 -23.635 23.965 ;
        RECT -23.965 22.275 -23.635 22.605 ;
        RECT -23.965 20.915 -23.635 21.245 ;
        RECT -23.965 19.555 -23.635 19.885 ;
        RECT -23.965 18.195 -23.635 18.525 ;
        RECT -23.965 16.835 -23.635 17.165 ;
        RECT -23.965 15.475 -23.635 15.805 ;
        RECT -23.965 14.115 -23.635 14.445 ;
        RECT -23.965 12.755 -23.635 13.085 ;
        RECT -23.965 11.395 -23.635 11.725 ;
        RECT -23.965 10.035 -23.635 10.365 ;
        RECT -23.965 8.675 -23.635 9.005 ;
        RECT -23.965 7.315 -23.635 7.645 ;
        RECT -23.965 5.955 -23.635 6.285 ;
        RECT -23.965 4.595 -23.635 4.925 ;
        RECT -23.965 3.235 -23.635 3.565 ;
        RECT -23.965 1.875 -23.635 2.205 ;
        RECT -23.965 0.515 -23.635 0.845 ;
        RECT -23.965 -0.845 -23.635 -0.515 ;
        RECT -23.965 -6.285 -23.635 -5.955 ;
        RECT -23.965 -8.19 -23.635 -7.86 ;
        RECT -23.965 -11.725 -23.635 -11.395 ;
        RECT -23.965 -14.23 -23.635 -13.9 ;
        RECT -23.965 -15.805 -23.635 -15.475 ;
        RECT -23.965 -28.045 -23.635 -27.715 ;
        RECT -23.965 -29.405 -23.635 -29.075 ;
        RECT -23.965 -31.17 -23.635 -30.84 ;
        RECT -23.965 -32.125 -23.635 -31.795 ;
        RECT -23.965 -33.485 -23.635 -33.155 ;
        RECT -23.965 -36.205 -23.635 -35.875 ;
        RECT -23.965 -37.21 -23.635 -36.88 ;
        RECT -23.965 -38.925 -23.635 -38.595 ;
        RECT -23.965 -41.645 -23.635 -41.315 ;
        RECT -23.965 -51.165 -23.635 -50.835 ;
        RECT -23.965 -52.525 -23.635 -52.195 ;
        RECT -23.965 -53.885 -23.635 -53.555 ;
        RECT -23.965 -55.245 -23.635 -54.915 ;
        RECT -23.965 -56.605 -23.635 -56.275 ;
        RECT -23.965 -57.965 -23.635 -57.635 ;
        RECT -23.965 -59.325 -23.635 -58.995 ;
        RECT -23.965 -60.685 -23.635 -60.355 ;
        RECT -23.965 -62.045 -23.635 -61.715 ;
        RECT -23.965 -63.405 -23.635 -63.075 ;
        RECT -23.965 -64.765 -23.635 -64.435 ;
        RECT -23.965 -66.125 -23.635 -65.795 ;
        RECT -23.965 -67.485 -23.635 -67.155 ;
        RECT -23.965 -68.845 -23.635 -68.515 ;
        RECT -23.965 -70.205 -23.635 -69.875 ;
        RECT -23.965 -71.565 -23.635 -71.235 ;
        RECT -23.965 -72.925 -23.635 -72.595 ;
        RECT -23.965 -74.285 -23.635 -73.955 ;
        RECT -23.965 -75.645 -23.635 -75.315 ;
        RECT -23.965 -77.005 -23.635 -76.675 ;
        RECT -23.965 -78.365 -23.635 -78.035 ;
        RECT -23.965 -79.725 -23.635 -79.395 ;
        RECT -23.965 -81.085 -23.635 -80.755 ;
        RECT -23.965 -82.445 -23.635 -82.115 ;
        RECT -23.965 -83.805 -23.635 -83.475 ;
        RECT -23.965 -85.165 -23.635 -84.835 ;
        RECT -23.965 -86.525 -23.635 -86.195 ;
        RECT -23.965 -87.885 -23.635 -87.555 ;
        RECT -23.965 -89.245 -23.635 -88.915 ;
        RECT -23.965 -90.605 -23.635 -90.275 ;
        RECT -23.965 -91.965 -23.635 -91.635 ;
        RECT -23.965 -93.325 -23.635 -92.995 ;
        RECT -23.965 -94.685 -23.635 -94.355 ;
        RECT -23.965 -96.045 -23.635 -95.715 ;
        RECT -23.965 -98.765 -23.635 -98.435 ;
        RECT -23.965 -100.125 -23.635 -99.795 ;
        RECT -23.965 -101.485 -23.635 -101.155 ;
        RECT -23.965 -102.845 -23.635 -102.515 ;
        RECT -23.965 -104.205 -23.635 -103.875 ;
        RECT -23.965 -105.565 -23.635 -105.235 ;
        RECT -23.965 -106.925 -23.635 -106.595 ;
        RECT -23.965 -113.725 -23.635 -113.395 ;
        RECT -23.965 -115.085 -23.635 -114.755 ;
        RECT -23.965 -117.805 -23.635 -117.475 ;
        RECT -23.965 -120.525 -23.635 -120.195 ;
        RECT -23.965 -121.885 -23.635 -121.555 ;
        RECT -23.965 -125.965 -23.635 -125.635 ;
        RECT -23.965 -127.325 -23.635 -126.995 ;
        RECT -23.965 -131.405 -23.635 -131.075 ;
        RECT -23.965 -136.845 -23.635 -136.515 ;
        RECT -23.965 -138.205 -23.635 -137.875 ;
        RECT -23.965 -139.565 -23.635 -139.235 ;
        RECT -23.965 -140.925 -23.635 -140.595 ;
        RECT -23.965 -142.285 -23.635 -141.955 ;
        RECT -23.965 -143.645 -23.635 -143.315 ;
        RECT -23.965 -145.005 -23.635 -144.675 ;
        RECT -23.965 -146.365 -23.635 -146.035 ;
        RECT -23.965 -148.215 -23.635 -147.885 ;
        RECT -23.965 -149.085 -23.635 -148.755 ;
        RECT -23.965 -150.445 -23.635 -150.115 ;
        RECT -23.965 -151.805 -23.635 -151.475 ;
        RECT -23.965 -153.165 -23.635 -152.835 ;
        RECT -23.965 -154.525 -23.635 -154.195 ;
        RECT -23.965 -157.245 -23.635 -156.915 ;
        RECT -23.965 -162.89 -23.635 -161.76 ;
        RECT -23.96 -163.005 -23.64 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.605 129.945 -22.275 131.075 ;
        RECT -22.605 125.635 -22.275 125.965 ;
        RECT -22.605 124.275 -22.275 124.605 ;
        RECT -22.605 122.915 -22.275 123.245 ;
        RECT -22.605 121.555 -22.275 121.885 ;
        RECT -22.605 120.195 -22.275 120.525 ;
        RECT -22.605 118.835 -22.275 119.165 ;
        RECT -22.605 117.475 -22.275 117.805 ;
        RECT -22.605 116.115 -22.275 116.445 ;
        RECT -22.605 114.755 -22.275 115.085 ;
        RECT -22.605 113.395 -22.275 113.725 ;
        RECT -22.605 112.035 -22.275 112.365 ;
        RECT -22.605 110.675 -22.275 111.005 ;
        RECT -22.605 109.315 -22.275 109.645 ;
        RECT -22.605 107.955 -22.275 108.285 ;
        RECT -22.605 106.595 -22.275 106.925 ;
        RECT -22.605 105.235 -22.275 105.565 ;
        RECT -22.605 103.875 -22.275 104.205 ;
        RECT -22.605 102.515 -22.275 102.845 ;
        RECT -22.605 101.155 -22.275 101.485 ;
        RECT -22.605 99.795 -22.275 100.125 ;
        RECT -22.605 98.435 -22.275 98.765 ;
        RECT -22.605 97.075 -22.275 97.405 ;
        RECT -22.605 95.715 -22.275 96.045 ;
        RECT -22.605 94.355 -22.275 94.685 ;
        RECT -22.605 92.995 -22.275 93.325 ;
        RECT -22.605 91.635 -22.275 91.965 ;
        RECT -22.605 90.275 -22.275 90.605 ;
        RECT -22.605 88.915 -22.275 89.245 ;
        RECT -22.605 87.555 -22.275 87.885 ;
        RECT -22.605 86.195 -22.275 86.525 ;
        RECT -22.605 84.835 -22.275 85.165 ;
        RECT -22.605 83.475 -22.275 83.805 ;
        RECT -22.605 82.115 -22.275 82.445 ;
        RECT -22.605 80.755 -22.275 81.085 ;
        RECT -22.605 79.395 -22.275 79.725 ;
        RECT -22.605 78.035 -22.275 78.365 ;
        RECT -22.605 76.675 -22.275 77.005 ;
        RECT -22.605 75.315 -22.275 75.645 ;
        RECT -22.605 73.955 -22.275 74.285 ;
        RECT -22.605 72.595 -22.275 72.925 ;
        RECT -22.605 71.235 -22.275 71.565 ;
        RECT -22.605 69.875 -22.275 70.205 ;
        RECT -22.605 68.515 -22.275 68.845 ;
        RECT -22.605 67.155 -22.275 67.485 ;
        RECT -22.605 65.795 -22.275 66.125 ;
        RECT -22.605 64.435 -22.275 64.765 ;
        RECT -22.605 63.075 -22.275 63.405 ;
        RECT -22.605 61.715 -22.275 62.045 ;
        RECT -22.605 60.355 -22.275 60.685 ;
        RECT -22.605 58.995 -22.275 59.325 ;
        RECT -22.605 57.635 -22.275 57.965 ;
        RECT -22.605 56.275 -22.275 56.605 ;
        RECT -22.605 54.915 -22.275 55.245 ;
        RECT -22.605 53.555 -22.275 53.885 ;
        RECT -22.605 52.195 -22.275 52.525 ;
        RECT -22.605 50.835 -22.275 51.165 ;
        RECT -22.605 49.475 -22.275 49.805 ;
        RECT -22.605 48.115 -22.275 48.445 ;
        RECT -22.605 46.755 -22.275 47.085 ;
        RECT -22.605 45.395 -22.275 45.725 ;
        RECT -22.605 44.035 -22.275 44.365 ;
        RECT -22.605 42.675 -22.275 43.005 ;
        RECT -22.605 41.315 -22.275 41.645 ;
        RECT -22.605 39.955 -22.275 40.285 ;
        RECT -22.605 38.595 -22.275 38.925 ;
        RECT -22.605 37.235 -22.275 37.565 ;
        RECT -22.605 35.875 -22.275 36.205 ;
        RECT -22.605 34.515 -22.275 34.845 ;
        RECT -22.605 33.155 -22.275 33.485 ;
        RECT -22.605 31.795 -22.275 32.125 ;
        RECT -22.605 30.435 -22.275 30.765 ;
        RECT -22.605 29.075 -22.275 29.405 ;
        RECT -22.605 27.715 -22.275 28.045 ;
        RECT -22.605 26.355 -22.275 26.685 ;
        RECT -22.605 24.995 -22.275 25.325 ;
        RECT -22.605 23.635 -22.275 23.965 ;
        RECT -22.605 22.275 -22.275 22.605 ;
        RECT -22.605 20.915 -22.275 21.245 ;
        RECT -22.605 19.555 -22.275 19.885 ;
        RECT -22.605 18.195 -22.275 18.525 ;
        RECT -22.605 16.835 -22.275 17.165 ;
        RECT -22.605 15.475 -22.275 15.805 ;
        RECT -22.605 14.115 -22.275 14.445 ;
        RECT -22.605 12.755 -22.275 13.085 ;
        RECT -22.605 11.395 -22.275 11.725 ;
        RECT -22.605 10.035 -22.275 10.365 ;
        RECT -22.605 8.675 -22.275 9.005 ;
        RECT -22.605 7.315 -22.275 7.645 ;
        RECT -22.605 5.955 -22.275 6.285 ;
        RECT -22.605 4.595 -22.275 4.925 ;
        RECT -22.605 3.235 -22.275 3.565 ;
        RECT -22.605 1.875 -22.275 2.205 ;
        RECT -22.605 0.515 -22.275 0.845 ;
        RECT -22.605 -0.845 -22.275 -0.515 ;
        RECT -22.605 -6.285 -22.275 -5.955 ;
        RECT -22.605 -8.19 -22.275 -7.86 ;
        RECT -22.605 -11.725 -22.275 -11.395 ;
        RECT -22.605 -14.23 -22.275 -13.9 ;
        RECT -22.605 -15.805 -22.275 -15.475 ;
        RECT -22.605 -28.045 -22.275 -27.715 ;
        RECT -22.605 -29.405 -22.275 -29.075 ;
        RECT -22.605 -31.17 -22.275 -30.84 ;
        RECT -22.605 -32.125 -22.275 -31.795 ;
        RECT -22.605 -33.485 -22.275 -33.155 ;
        RECT -22.605 -36.205 -22.275 -35.875 ;
        RECT -22.605 -37.21 -22.275 -36.88 ;
        RECT -22.605 -38.925 -22.275 -38.595 ;
        RECT -22.605 -41.645 -22.275 -41.315 ;
        RECT -22.605 -51.165 -22.275 -50.835 ;
        RECT -22.605 -52.525 -22.275 -52.195 ;
        RECT -22.605 -53.885 -22.275 -53.555 ;
        RECT -22.605 -55.245 -22.275 -54.915 ;
        RECT -22.605 -56.605 -22.275 -56.275 ;
        RECT -22.605 -57.965 -22.275 -57.635 ;
        RECT -22.605 -59.325 -22.275 -58.995 ;
        RECT -22.605 -60.685 -22.275 -60.355 ;
        RECT -22.605 -62.045 -22.275 -61.715 ;
        RECT -22.605 -63.405 -22.275 -63.075 ;
        RECT -22.605 -64.765 -22.275 -64.435 ;
        RECT -22.605 -66.125 -22.275 -65.795 ;
        RECT -22.605 -67.485 -22.275 -67.155 ;
        RECT -22.605 -68.845 -22.275 -68.515 ;
        RECT -22.605 -70.205 -22.275 -69.875 ;
        RECT -22.605 -71.565 -22.275 -71.235 ;
        RECT -22.605 -72.925 -22.275 -72.595 ;
        RECT -22.605 -74.285 -22.275 -73.955 ;
        RECT -22.605 -75.645 -22.275 -75.315 ;
        RECT -22.605 -77.005 -22.275 -76.675 ;
        RECT -22.605 -78.365 -22.275 -78.035 ;
        RECT -22.605 -79.725 -22.275 -79.395 ;
        RECT -22.605 -81.085 -22.275 -80.755 ;
        RECT -22.605 -82.445 -22.275 -82.115 ;
        RECT -22.605 -83.805 -22.275 -83.475 ;
        RECT -22.605 -85.165 -22.275 -84.835 ;
        RECT -22.605 -86.525 -22.275 -86.195 ;
        RECT -22.605 -87.885 -22.275 -87.555 ;
        RECT -22.605 -89.245 -22.275 -88.915 ;
        RECT -22.605 -90.605 -22.275 -90.275 ;
        RECT -22.605 -91.965 -22.275 -91.635 ;
        RECT -22.605 -93.325 -22.275 -92.995 ;
        RECT -22.605 -94.685 -22.275 -94.355 ;
        RECT -22.605 -96.045 -22.275 -95.715 ;
        RECT -22.605 -98.765 -22.275 -98.435 ;
        RECT -22.605 -100.125 -22.275 -99.795 ;
        RECT -22.605 -101.485 -22.275 -101.155 ;
        RECT -22.605 -102.845 -22.275 -102.515 ;
        RECT -22.605 -104.205 -22.275 -103.875 ;
        RECT -22.605 -105.565 -22.275 -105.235 ;
        RECT -22.605 -106.925 -22.275 -106.595 ;
        RECT -22.605 -113.725 -22.275 -113.395 ;
        RECT -22.605 -115.085 -22.275 -114.755 ;
        RECT -22.605 -117.805 -22.275 -117.475 ;
        RECT -22.605 -120.525 -22.275 -120.195 ;
        RECT -22.605 -121.885 -22.275 -121.555 ;
        RECT -22.605 -123.245 -22.275 -122.915 ;
        RECT -22.605 -125.965 -22.275 -125.635 ;
        RECT -22.605 -127.325 -22.275 -126.995 ;
        RECT -22.605 -131.405 -22.275 -131.075 ;
        RECT -22.605 -135.485 -22.275 -135.155 ;
        RECT -22.605 -136.845 -22.275 -136.515 ;
        RECT -22.605 -138.205 -22.275 -137.875 ;
        RECT -22.605 -139.565 -22.275 -139.235 ;
        RECT -22.605 -140.925 -22.275 -140.595 ;
        RECT -22.605 -142.285 -22.275 -141.955 ;
        RECT -22.605 -143.645 -22.275 -143.315 ;
        RECT -22.605 -145.005 -22.275 -144.675 ;
        RECT -22.605 -146.365 -22.275 -146.035 ;
        RECT -22.605 -149.085 -22.275 -148.755 ;
        RECT -22.605 -150.445 -22.275 -150.115 ;
        RECT -22.605 -154.525 -22.275 -154.195 ;
        RECT -22.605 -157.245 -22.275 -156.915 ;
        RECT -22.605 -162.89 -22.275 -161.76 ;
        RECT -22.6 -163.005 -22.28 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 129.945 -20.915 131.075 ;
        RECT -21.245 125.635 -20.915 125.965 ;
        RECT -21.245 124.275 -20.915 124.605 ;
        RECT -21.245 122.915 -20.915 123.245 ;
        RECT -21.245 121.555 -20.915 121.885 ;
        RECT -21.245 120.195 -20.915 120.525 ;
        RECT -21.245 118.835 -20.915 119.165 ;
        RECT -21.245 117.475 -20.915 117.805 ;
        RECT -21.245 116.115 -20.915 116.445 ;
        RECT -21.245 114.755 -20.915 115.085 ;
        RECT -21.245 113.395 -20.915 113.725 ;
        RECT -21.245 112.035 -20.915 112.365 ;
        RECT -21.245 110.675 -20.915 111.005 ;
        RECT -21.245 109.315 -20.915 109.645 ;
        RECT -21.245 107.955 -20.915 108.285 ;
        RECT -21.245 106.595 -20.915 106.925 ;
        RECT -21.245 105.235 -20.915 105.565 ;
        RECT -21.245 103.875 -20.915 104.205 ;
        RECT -21.245 102.515 -20.915 102.845 ;
        RECT -21.245 101.155 -20.915 101.485 ;
        RECT -21.245 99.795 -20.915 100.125 ;
        RECT -21.245 98.435 -20.915 98.765 ;
        RECT -21.245 97.075 -20.915 97.405 ;
        RECT -21.245 95.715 -20.915 96.045 ;
        RECT -21.245 94.355 -20.915 94.685 ;
        RECT -21.245 92.995 -20.915 93.325 ;
        RECT -21.245 91.635 -20.915 91.965 ;
        RECT -21.245 90.275 -20.915 90.605 ;
        RECT -21.245 88.915 -20.915 89.245 ;
        RECT -21.245 87.555 -20.915 87.885 ;
        RECT -21.245 86.195 -20.915 86.525 ;
        RECT -21.245 84.835 -20.915 85.165 ;
        RECT -21.245 83.475 -20.915 83.805 ;
        RECT -21.245 82.115 -20.915 82.445 ;
        RECT -21.245 80.755 -20.915 81.085 ;
        RECT -21.245 79.395 -20.915 79.725 ;
        RECT -21.245 78.035 -20.915 78.365 ;
        RECT -21.245 76.675 -20.915 77.005 ;
        RECT -21.245 75.315 -20.915 75.645 ;
        RECT -21.245 73.955 -20.915 74.285 ;
        RECT -21.245 72.595 -20.915 72.925 ;
        RECT -21.245 71.235 -20.915 71.565 ;
        RECT -21.245 69.875 -20.915 70.205 ;
        RECT -21.245 68.515 -20.915 68.845 ;
        RECT -21.245 67.155 -20.915 67.485 ;
        RECT -21.245 65.795 -20.915 66.125 ;
        RECT -21.245 64.435 -20.915 64.765 ;
        RECT -21.245 63.075 -20.915 63.405 ;
        RECT -21.245 61.715 -20.915 62.045 ;
        RECT -21.245 60.355 -20.915 60.685 ;
        RECT -21.245 58.995 -20.915 59.325 ;
        RECT -21.245 57.635 -20.915 57.965 ;
        RECT -21.245 56.275 -20.915 56.605 ;
        RECT -21.245 54.915 -20.915 55.245 ;
        RECT -21.245 53.555 -20.915 53.885 ;
        RECT -21.245 52.195 -20.915 52.525 ;
        RECT -21.245 50.835 -20.915 51.165 ;
        RECT -21.245 49.475 -20.915 49.805 ;
        RECT -21.245 48.115 -20.915 48.445 ;
        RECT -21.245 46.755 -20.915 47.085 ;
        RECT -21.245 45.395 -20.915 45.725 ;
        RECT -21.245 44.035 -20.915 44.365 ;
        RECT -21.245 42.675 -20.915 43.005 ;
        RECT -21.245 41.315 -20.915 41.645 ;
        RECT -21.245 39.955 -20.915 40.285 ;
        RECT -21.245 38.595 -20.915 38.925 ;
        RECT -21.245 37.235 -20.915 37.565 ;
        RECT -21.245 35.875 -20.915 36.205 ;
        RECT -21.245 34.515 -20.915 34.845 ;
        RECT -21.245 33.155 -20.915 33.485 ;
        RECT -21.245 31.795 -20.915 32.125 ;
        RECT -21.245 30.435 -20.915 30.765 ;
        RECT -21.245 29.075 -20.915 29.405 ;
        RECT -21.245 27.715 -20.915 28.045 ;
        RECT -21.245 26.355 -20.915 26.685 ;
        RECT -21.245 24.995 -20.915 25.325 ;
        RECT -21.245 23.635 -20.915 23.965 ;
        RECT -21.245 22.275 -20.915 22.605 ;
        RECT -21.245 20.915 -20.915 21.245 ;
        RECT -21.245 19.555 -20.915 19.885 ;
        RECT -21.245 18.195 -20.915 18.525 ;
        RECT -21.245 16.835 -20.915 17.165 ;
        RECT -21.245 15.475 -20.915 15.805 ;
        RECT -21.245 14.115 -20.915 14.445 ;
        RECT -21.245 12.755 -20.915 13.085 ;
        RECT -21.245 11.395 -20.915 11.725 ;
        RECT -21.245 10.035 -20.915 10.365 ;
        RECT -21.245 8.675 -20.915 9.005 ;
        RECT -21.245 7.315 -20.915 7.645 ;
        RECT -21.245 5.955 -20.915 6.285 ;
        RECT -21.245 4.595 -20.915 4.925 ;
        RECT -21.245 3.235 -20.915 3.565 ;
        RECT -21.245 1.875 -20.915 2.205 ;
        RECT -21.245 0.515 -20.915 0.845 ;
        RECT -21.245 -0.845 -20.915 -0.515 ;
        RECT -21.245 -2.205 -20.915 -1.875 ;
        RECT -21.245 -6.285 -20.915 -5.955 ;
        RECT -21.245 -8.19 -20.915 -7.86 ;
        RECT -21.245 -11.725 -20.915 -11.395 ;
        RECT -21.245 -14.23 -20.915 -13.9 ;
        RECT -21.245 -15.805 -20.915 -15.475 ;
        RECT -21.24 -21.24 -20.92 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -28.045 -20.915 -27.715 ;
        RECT -21.245 -29.405 -20.915 -29.075 ;
        RECT -21.245 -31.17 -20.915 -30.84 ;
        RECT -21.245 -32.125 -20.915 -31.795 ;
        RECT -21.245 -33.485 -20.915 -33.155 ;
        RECT -21.245 -36.205 -20.915 -35.875 ;
        RECT -21.245 -37.21 -20.915 -36.88 ;
        RECT -21.245 -38.925 -20.915 -38.595 ;
        RECT -21.245 -41.645 -20.915 -41.315 ;
        RECT -21.24 -44.36 -20.92 -27.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -51.165 -20.915 -50.835 ;
        RECT -21.245 -52.525 -20.915 -52.195 ;
        RECT -21.245 -53.885 -20.915 -53.555 ;
        RECT -21.245 -55.245 -20.915 -54.915 ;
        RECT -21.245 -56.605 -20.915 -56.275 ;
        RECT -21.245 -57.965 -20.915 -57.635 ;
        RECT -21.245 -59.325 -20.915 -58.995 ;
        RECT -21.245 -60.685 -20.915 -60.355 ;
        RECT -21.245 -62.045 -20.915 -61.715 ;
        RECT -21.245 -63.405 -20.915 -63.075 ;
        RECT -21.245 -64.765 -20.915 -64.435 ;
        RECT -21.245 -66.125 -20.915 -65.795 ;
        RECT -21.245 -67.485 -20.915 -67.155 ;
        RECT -21.245 -68.845 -20.915 -68.515 ;
        RECT -21.245 -70.205 -20.915 -69.875 ;
        RECT -21.245 -71.565 -20.915 -71.235 ;
        RECT -21.245 -72.925 -20.915 -72.595 ;
        RECT -21.245 -74.285 -20.915 -73.955 ;
        RECT -21.245 -75.645 -20.915 -75.315 ;
        RECT -21.245 -77.005 -20.915 -76.675 ;
        RECT -21.245 -78.365 -20.915 -78.035 ;
        RECT -21.245 -79.725 -20.915 -79.395 ;
        RECT -21.245 -81.085 -20.915 -80.755 ;
        RECT -21.245 -82.445 -20.915 -82.115 ;
        RECT -21.245 -83.805 -20.915 -83.475 ;
        RECT -21.245 -85.165 -20.915 -84.835 ;
        RECT -21.245 -86.525 -20.915 -86.195 ;
        RECT -21.245 -87.885 -20.915 -87.555 ;
        RECT -21.245 -89.245 -20.915 -88.915 ;
        RECT -21.245 -90.605 -20.915 -90.275 ;
        RECT -21.24 -91.28 -20.92 -50.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 129.945 -19.555 131.075 ;
        RECT -19.885 125.635 -19.555 125.965 ;
        RECT -19.885 124.275 -19.555 124.605 ;
        RECT -19.885 122.915 -19.555 123.245 ;
        RECT -19.885 121.555 -19.555 121.885 ;
        RECT -19.885 120.195 -19.555 120.525 ;
        RECT -19.885 118.835 -19.555 119.165 ;
        RECT -19.885 117.475 -19.555 117.805 ;
        RECT -19.885 116.115 -19.555 116.445 ;
        RECT -19.885 114.755 -19.555 115.085 ;
        RECT -19.885 113.395 -19.555 113.725 ;
        RECT -19.885 112.035 -19.555 112.365 ;
        RECT -19.885 110.675 -19.555 111.005 ;
        RECT -19.885 109.315 -19.555 109.645 ;
        RECT -19.885 107.955 -19.555 108.285 ;
        RECT -19.885 106.595 -19.555 106.925 ;
        RECT -19.885 105.235 -19.555 105.565 ;
        RECT -19.885 103.875 -19.555 104.205 ;
        RECT -19.885 102.515 -19.555 102.845 ;
        RECT -19.885 101.155 -19.555 101.485 ;
        RECT -19.885 99.795 -19.555 100.125 ;
        RECT -19.885 98.435 -19.555 98.765 ;
        RECT -19.885 97.075 -19.555 97.405 ;
        RECT -19.885 95.715 -19.555 96.045 ;
        RECT -19.885 94.355 -19.555 94.685 ;
        RECT -19.885 92.995 -19.555 93.325 ;
        RECT -19.885 91.635 -19.555 91.965 ;
        RECT -19.885 90.275 -19.555 90.605 ;
        RECT -19.885 88.915 -19.555 89.245 ;
        RECT -19.885 87.555 -19.555 87.885 ;
        RECT -19.885 86.195 -19.555 86.525 ;
        RECT -19.885 84.835 -19.555 85.165 ;
        RECT -19.885 83.475 -19.555 83.805 ;
        RECT -19.885 82.115 -19.555 82.445 ;
        RECT -19.885 80.755 -19.555 81.085 ;
        RECT -19.885 79.395 -19.555 79.725 ;
        RECT -19.885 78.035 -19.555 78.365 ;
        RECT -19.885 76.675 -19.555 77.005 ;
        RECT -19.885 75.315 -19.555 75.645 ;
        RECT -19.885 73.955 -19.555 74.285 ;
        RECT -19.885 72.595 -19.555 72.925 ;
        RECT -19.885 71.235 -19.555 71.565 ;
        RECT -19.885 69.875 -19.555 70.205 ;
        RECT -19.885 68.515 -19.555 68.845 ;
        RECT -19.885 67.155 -19.555 67.485 ;
        RECT -19.885 65.795 -19.555 66.125 ;
        RECT -19.885 64.435 -19.555 64.765 ;
        RECT -19.885 63.075 -19.555 63.405 ;
        RECT -19.885 61.715 -19.555 62.045 ;
        RECT -19.885 60.355 -19.555 60.685 ;
        RECT -19.885 58.995 -19.555 59.325 ;
        RECT -19.885 57.635 -19.555 57.965 ;
        RECT -19.885 56.275 -19.555 56.605 ;
        RECT -19.885 54.915 -19.555 55.245 ;
        RECT -19.885 53.555 -19.555 53.885 ;
        RECT -19.885 52.195 -19.555 52.525 ;
        RECT -19.885 50.835 -19.555 51.165 ;
        RECT -19.885 49.475 -19.555 49.805 ;
        RECT -19.885 48.115 -19.555 48.445 ;
        RECT -19.885 46.755 -19.555 47.085 ;
        RECT -19.885 45.395 -19.555 45.725 ;
        RECT -19.885 44.035 -19.555 44.365 ;
        RECT -19.885 42.675 -19.555 43.005 ;
        RECT -19.885 41.315 -19.555 41.645 ;
        RECT -19.885 39.955 -19.555 40.285 ;
        RECT -19.885 38.595 -19.555 38.925 ;
        RECT -19.885 37.235 -19.555 37.565 ;
        RECT -19.885 35.875 -19.555 36.205 ;
        RECT -19.885 34.515 -19.555 34.845 ;
        RECT -19.885 33.155 -19.555 33.485 ;
        RECT -19.885 31.795 -19.555 32.125 ;
        RECT -19.885 30.435 -19.555 30.765 ;
        RECT -19.885 29.075 -19.555 29.405 ;
        RECT -19.885 27.715 -19.555 28.045 ;
        RECT -19.885 26.355 -19.555 26.685 ;
        RECT -19.885 24.995 -19.555 25.325 ;
        RECT -19.885 23.635 -19.555 23.965 ;
        RECT -19.885 22.275 -19.555 22.605 ;
        RECT -19.885 20.915 -19.555 21.245 ;
        RECT -19.885 19.555 -19.555 19.885 ;
        RECT -19.885 18.195 -19.555 18.525 ;
        RECT -19.885 16.835 -19.555 17.165 ;
        RECT -19.885 15.475 -19.555 15.805 ;
        RECT -19.885 14.115 -19.555 14.445 ;
        RECT -19.885 12.755 -19.555 13.085 ;
        RECT -19.885 11.395 -19.555 11.725 ;
        RECT -19.885 10.035 -19.555 10.365 ;
        RECT -19.885 8.675 -19.555 9.005 ;
        RECT -19.885 7.315 -19.555 7.645 ;
        RECT -19.885 5.955 -19.555 6.285 ;
        RECT -19.885 4.595 -19.555 4.925 ;
        RECT -19.885 3.235 -19.555 3.565 ;
        RECT -19.885 1.875 -19.555 2.205 ;
        RECT -19.885 0.515 -19.555 0.845 ;
        RECT -19.885 -0.845 -19.555 -0.515 ;
        RECT -19.885 -2.205 -19.555 -1.875 ;
        RECT -19.885 -6.285 -19.555 -5.955 ;
        RECT -19.885 -8.19 -19.555 -7.86 ;
        RECT -19.885 -11.725 -19.555 -11.395 ;
        RECT -19.885 -14.23 -19.555 -13.9 ;
        RECT -19.885 -15.805 -19.555 -15.475 ;
        RECT -19.88 -20.56 -19.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -26.685 -19.555 -26.355 ;
        RECT -19.885 -28.045 -19.555 -27.715 ;
        RECT -19.885 -29.405 -19.555 -29.075 ;
        RECT -19.885 -31.17 -19.555 -30.84 ;
        RECT -19.885 -32.125 -19.555 -31.795 ;
        RECT -19.885 -33.485 -19.555 -33.155 ;
        RECT -19.885 -36.205 -19.555 -35.875 ;
        RECT -19.885 -37.21 -19.555 -36.88 ;
        RECT -19.885 -38.925 -19.555 -38.595 ;
        RECT -19.885 -41.645 -19.555 -41.315 ;
        RECT -19.88 -43.68 -19.56 -25.68 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -63.405 -19.555 -63.075 ;
        RECT -19.885 -66.125 -19.555 -65.795 ;
        RECT -19.885 -68.845 -19.555 -68.515 ;
        RECT -19.885 -70.205 -19.555 -69.875 ;
        RECT -19.885 -71.565 -19.555 -71.235 ;
        RECT -19.885 -72.925 -19.555 -72.595 ;
        RECT -19.885 -74.93 -19.555 -74.6 ;
        RECT -19.885 -75.645 -19.555 -75.315 ;
        RECT -19.885 -77.005 -19.555 -76.675 ;
        RECT -19.885 -79.725 -19.555 -79.395 ;
        RECT -19.885 -81.085 -19.555 -80.755 ;
        RECT -19.885 -82.47 -19.555 -82.14 ;
        RECT -19.885 -83.805 -19.555 -83.475 ;
        RECT -19.885 -85.165 -19.555 -84.835 ;
        RECT -19.885 -87.885 -19.555 -87.555 ;
        RECT -19.885 -93.325 -19.555 -92.995 ;
        RECT -19.885 -94.685 -19.555 -94.355 ;
        RECT -19.885 -96.045 -19.555 -95.715 ;
        RECT -19.885 -100.125 -19.555 -99.795 ;
        RECT -19.885 -104.205 -19.555 -103.875 ;
        RECT -19.885 -105.565 -19.555 -105.235 ;
        RECT -19.885 -106.925 -19.555 -106.595 ;
        RECT -19.885 -117.805 -19.555 -117.475 ;
        RECT -19.885 -120.525 -19.555 -120.195 ;
        RECT -19.885 -123.245 -19.555 -122.915 ;
        RECT -19.885 -124.605 -19.555 -124.275 ;
        RECT -19.885 -125.965 -19.555 -125.635 ;
        RECT -19.885 -127.325 -19.555 -126.995 ;
        RECT -19.885 -131.405 -19.555 -131.075 ;
        RECT -19.885 -136.845 -19.555 -136.515 ;
        RECT -19.885 -138.205 -19.555 -137.875 ;
        RECT -19.885 -139.565 -19.555 -139.235 ;
        RECT -19.885 -140.925 -19.555 -140.595 ;
        RECT -19.885 -142.285 -19.555 -141.955 ;
        RECT -19.885 -143.645 -19.555 -143.315 ;
        RECT -19.885 -145.005 -19.555 -144.675 ;
        RECT -19.885 -146.365 -19.555 -146.035 ;
        RECT -19.885 -148.215 -19.555 -147.885 ;
        RECT -19.885 -149.085 -19.555 -148.755 ;
        RECT -19.885 -150.445 -19.555 -150.115 ;
        RECT -19.885 -153.165 -19.555 -152.835 ;
        RECT -19.885 -154.525 -19.555 -154.195 ;
        RECT -19.885 -157.245 -19.555 -156.915 ;
        RECT -19.885 -162.89 -19.555 -161.76 ;
        RECT -19.88 -163.005 -19.56 -48.8 ;
        RECT -19.885 -49.805 -19.555 -49.475 ;
        RECT -19.885 -51.165 -19.555 -50.835 ;
        RECT -19.885 -52.75 -19.555 -52.42 ;
        RECT -19.885 -53.885 -19.555 -53.555 ;
        RECT -19.885 -55.245 -19.555 -54.915 ;
        RECT -19.885 -57.965 -19.555 -57.635 ;
        RECT -19.885 -59.325 -19.555 -58.995 ;
        RECT -19.885 -60.29 -19.555 -59.96 ;
        RECT -19.885 -62.045 -19.555 -61.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.485 129.945 -33.155 131.075 ;
        RECT -33.485 125.635 -33.155 125.965 ;
        RECT -33.485 124.275 -33.155 124.605 ;
        RECT -33.485 122.915 -33.155 123.245 ;
        RECT -33.485 121.555 -33.155 121.885 ;
        RECT -33.485 120.195 -33.155 120.525 ;
        RECT -33.485 118.835 -33.155 119.165 ;
        RECT -33.485 117.475 -33.155 117.805 ;
        RECT -33.485 116.115 -33.155 116.445 ;
        RECT -33.485 114.755 -33.155 115.085 ;
        RECT -33.485 113.395 -33.155 113.725 ;
        RECT -33.485 112.035 -33.155 112.365 ;
        RECT -33.485 110.675 -33.155 111.005 ;
        RECT -33.485 109.315 -33.155 109.645 ;
        RECT -33.485 107.955 -33.155 108.285 ;
        RECT -33.485 106.595 -33.155 106.925 ;
        RECT -33.485 105.235 -33.155 105.565 ;
        RECT -33.485 103.875 -33.155 104.205 ;
        RECT -33.485 102.515 -33.155 102.845 ;
        RECT -33.485 101.155 -33.155 101.485 ;
        RECT -33.485 99.795 -33.155 100.125 ;
        RECT -33.485 98.435 -33.155 98.765 ;
        RECT -33.485 97.075 -33.155 97.405 ;
        RECT -33.485 95.715 -33.155 96.045 ;
        RECT -33.485 94.355 -33.155 94.685 ;
        RECT -33.485 92.995 -33.155 93.325 ;
        RECT -33.485 91.635 -33.155 91.965 ;
        RECT -33.485 90.275 -33.155 90.605 ;
        RECT -33.485 88.915 -33.155 89.245 ;
        RECT -33.485 87.555 -33.155 87.885 ;
        RECT -33.485 86.195 -33.155 86.525 ;
        RECT -33.485 84.835 -33.155 85.165 ;
        RECT -33.485 83.475 -33.155 83.805 ;
        RECT -33.485 82.115 -33.155 82.445 ;
        RECT -33.485 80.755 -33.155 81.085 ;
        RECT -33.485 79.395 -33.155 79.725 ;
        RECT -33.485 78.035 -33.155 78.365 ;
        RECT -33.485 76.675 -33.155 77.005 ;
        RECT -33.485 75.315 -33.155 75.645 ;
        RECT -33.485 73.955 -33.155 74.285 ;
        RECT -33.485 72.595 -33.155 72.925 ;
        RECT -33.485 71.235 -33.155 71.565 ;
        RECT -33.485 69.875 -33.155 70.205 ;
        RECT -33.485 68.515 -33.155 68.845 ;
        RECT -33.485 67.155 -33.155 67.485 ;
        RECT -33.485 65.795 -33.155 66.125 ;
        RECT -33.485 64.435 -33.155 64.765 ;
        RECT -33.485 63.075 -33.155 63.405 ;
        RECT -33.485 61.715 -33.155 62.045 ;
        RECT -33.485 60.355 -33.155 60.685 ;
        RECT -33.485 58.995 -33.155 59.325 ;
        RECT -33.485 57.635 -33.155 57.965 ;
        RECT -33.485 56.275 -33.155 56.605 ;
        RECT -33.485 54.915 -33.155 55.245 ;
        RECT -33.485 53.555 -33.155 53.885 ;
        RECT -33.485 52.195 -33.155 52.525 ;
        RECT -33.485 50.835 -33.155 51.165 ;
        RECT -33.485 49.475 -33.155 49.805 ;
        RECT -33.485 48.115 -33.155 48.445 ;
        RECT -33.485 46.755 -33.155 47.085 ;
        RECT -33.485 45.395 -33.155 45.725 ;
        RECT -33.485 44.035 -33.155 44.365 ;
        RECT -33.485 42.675 -33.155 43.005 ;
        RECT -33.485 41.315 -33.155 41.645 ;
        RECT -33.485 39.955 -33.155 40.285 ;
        RECT -33.485 38.595 -33.155 38.925 ;
        RECT -33.485 37.235 -33.155 37.565 ;
        RECT -33.485 35.875 -33.155 36.205 ;
        RECT -33.485 34.515 -33.155 34.845 ;
        RECT -33.485 33.155 -33.155 33.485 ;
        RECT -33.485 31.795 -33.155 32.125 ;
        RECT -33.485 30.435 -33.155 30.765 ;
        RECT -33.485 29.075 -33.155 29.405 ;
        RECT -33.485 27.715 -33.155 28.045 ;
        RECT -33.485 26.355 -33.155 26.685 ;
        RECT -33.485 24.995 -33.155 25.325 ;
        RECT -33.485 23.635 -33.155 23.965 ;
        RECT -33.485 22.275 -33.155 22.605 ;
        RECT -33.485 20.915 -33.155 21.245 ;
        RECT -33.485 19.555 -33.155 19.885 ;
        RECT -33.485 18.195 -33.155 18.525 ;
        RECT -33.485 16.835 -33.155 17.165 ;
        RECT -33.485 15.475 -33.155 15.805 ;
        RECT -33.485 14.115 -33.155 14.445 ;
        RECT -33.485 12.755 -33.155 13.085 ;
        RECT -33.485 11.395 -33.155 11.725 ;
        RECT -33.485 10.035 -33.155 10.365 ;
        RECT -33.485 8.675 -33.155 9.005 ;
        RECT -33.485 7.315 -33.155 7.645 ;
        RECT -33.485 5.955 -33.155 6.285 ;
        RECT -33.485 4.595 -33.155 4.925 ;
        RECT -33.485 3.235 -33.155 3.565 ;
        RECT -33.485 1.875 -33.155 2.205 ;
        RECT -33.485 0.515 -33.155 0.845 ;
        RECT -33.485 -7.645 -33.155 -7.315 ;
        RECT -33.485 -11.725 -33.155 -11.395 ;
        RECT -33.485 -13.085 -33.155 -12.755 ;
        RECT -33.485 -14.445 -33.155 -14.115 ;
        RECT -33.485 -15.805 -33.155 -15.475 ;
        RECT -33.485 -17.165 -33.155 -16.835 ;
        RECT -33.485 -19.885 -33.155 -19.555 ;
        RECT -33.485 -21.245 -33.155 -20.915 ;
        RECT -33.485 -22.605 -33.155 -22.275 ;
        RECT -33.485 -29.405 -33.155 -29.075 ;
        RECT -33.485 -30.765 -33.155 -30.435 ;
        RECT -33.485 -32.125 -33.155 -31.795 ;
        RECT -33.485 -33.485 -33.155 -33.155 ;
        RECT -33.485 -34.845 -33.155 -34.515 ;
        RECT -33.485 -36.205 -33.155 -35.875 ;
        RECT -33.485 -37.565 -33.155 -37.235 ;
        RECT -33.485 -38.925 -33.155 -38.595 ;
        RECT -33.485 -40.285 -33.155 -39.955 ;
        RECT -33.485 -41.645 -33.155 -41.315 ;
        RECT -33.485 -43.005 -33.155 -42.675 ;
        RECT -33.485 -44.365 -33.155 -44.035 ;
        RECT -33.485 -45.725 -33.155 -45.395 ;
        RECT -33.485 -49.805 -33.155 -49.475 ;
        RECT -33.485 -51.165 -33.155 -50.835 ;
        RECT -33.485 -52.525 -33.155 -52.195 ;
        RECT -33.485 -53.885 -33.155 -53.555 ;
        RECT -33.485 -55.245 -33.155 -54.915 ;
        RECT -33.485 -56.605 -33.155 -56.275 ;
        RECT -33.485 -57.965 -33.155 -57.635 ;
        RECT -33.485 -59.325 -33.155 -58.995 ;
        RECT -33.485 -60.685 -33.155 -60.355 ;
        RECT -33.485 -62.045 -33.155 -61.715 ;
        RECT -33.485 -63.405 -33.155 -63.075 ;
        RECT -33.485 -64.765 -33.155 -64.435 ;
        RECT -33.485 -66.125 -33.155 -65.795 ;
        RECT -33.485 -67.485 -33.155 -67.155 ;
        RECT -33.485 -68.845 -33.155 -68.515 ;
        RECT -33.485 -70.37 -33.155 -70.04 ;
        RECT -33.485 -71.565 -33.155 -71.235 ;
        RECT -33.485 -72.925 -33.155 -72.595 ;
        RECT -33.485 -74.285 -33.155 -73.955 ;
        RECT -33.485 -75.645 -33.155 -75.315 ;
        RECT -33.485 -77.005 -33.155 -76.675 ;
        RECT -33.485 -79.725 -33.155 -79.395 ;
        RECT -33.485 -80.91 -33.155 -80.58 ;
        RECT -33.485 -82.445 -33.155 -82.115 ;
        RECT -33.485 -83.805 -33.155 -83.475 ;
        RECT -33.485 -85.165 -33.155 -84.835 ;
        RECT -33.485 -87.885 -33.155 -87.555 ;
        RECT -33.485 -89.245 -33.155 -88.915 ;
        RECT -33.485 -91.965 -33.155 -91.635 ;
        RECT -33.485 -93.325 -33.155 -92.995 ;
        RECT -33.485 -94.685 -33.155 -94.355 ;
        RECT -33.485 -96.045 -33.155 -95.715 ;
        RECT -33.485 -98.765 -33.155 -98.435 ;
        RECT -33.485 -100.125 -33.155 -99.795 ;
        RECT -33.485 -101.485 -33.155 -101.155 ;
        RECT -33.485 -102.845 -33.155 -102.515 ;
        RECT -33.485 -105.565 -33.155 -105.235 ;
        RECT -33.485 -106.925 -33.155 -106.595 ;
        RECT -33.485 -108.285 -33.155 -107.955 ;
        RECT -33.485 -112.365 -33.155 -112.035 ;
        RECT -33.485 -113.725 -33.155 -113.395 ;
        RECT -33.485 -115.085 -33.155 -114.755 ;
        RECT -33.485 -116.445 -33.155 -116.115 ;
        RECT -33.485 -117.805 -33.155 -117.475 ;
        RECT -33.485 -120.525 -33.155 -120.195 ;
        RECT -33.485 -121.885 -33.155 -121.555 ;
        RECT -33.485 -123.245 -33.155 -122.915 ;
        RECT -33.485 -124.605 -33.155 -124.275 ;
        RECT -33.485 -125.965 -33.155 -125.635 ;
        RECT -33.485 -127.325 -33.155 -126.995 ;
        RECT -33.485 -130.045 -33.155 -129.715 ;
        RECT -33.485 -131.405 -33.155 -131.075 ;
        RECT -33.485 -135.485 -33.155 -135.155 ;
        RECT -33.485 -136.845 -33.155 -136.515 ;
        RECT -33.485 -138.205 -33.155 -137.875 ;
        RECT -33.485 -139.565 -33.155 -139.235 ;
        RECT -33.485 -140.925 -33.155 -140.595 ;
        RECT -33.485 -142.285 -33.155 -141.955 ;
        RECT -33.485 -143.645 -33.155 -143.315 ;
        RECT -33.485 -145.005 -33.155 -144.675 ;
        RECT -33.485 -146.365 -33.155 -146.035 ;
        RECT -33.485 -148.215 -33.155 -147.885 ;
        RECT -33.485 -149.085 -33.155 -148.755 ;
        RECT -33.485 -150.445 -33.155 -150.115 ;
        RECT -33.485 -151.805 -33.155 -151.475 ;
        RECT -33.48 -151.805 -33.16 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.125 129.945 -31.795 131.075 ;
        RECT -32.125 125.635 -31.795 125.965 ;
        RECT -32.125 124.275 -31.795 124.605 ;
        RECT -32.125 122.915 -31.795 123.245 ;
        RECT -32.125 121.555 -31.795 121.885 ;
        RECT -32.125 120.195 -31.795 120.525 ;
        RECT -32.125 118.835 -31.795 119.165 ;
        RECT -32.125 117.475 -31.795 117.805 ;
        RECT -32.125 116.115 -31.795 116.445 ;
        RECT -32.125 114.755 -31.795 115.085 ;
        RECT -32.125 113.395 -31.795 113.725 ;
        RECT -32.125 112.035 -31.795 112.365 ;
        RECT -32.125 110.675 -31.795 111.005 ;
        RECT -32.125 109.315 -31.795 109.645 ;
        RECT -32.125 107.955 -31.795 108.285 ;
        RECT -32.125 106.595 -31.795 106.925 ;
        RECT -32.125 105.235 -31.795 105.565 ;
        RECT -32.125 103.875 -31.795 104.205 ;
        RECT -32.125 102.515 -31.795 102.845 ;
        RECT -32.125 101.155 -31.795 101.485 ;
        RECT -32.125 99.795 -31.795 100.125 ;
        RECT -32.125 98.435 -31.795 98.765 ;
        RECT -32.125 97.075 -31.795 97.405 ;
        RECT -32.125 95.715 -31.795 96.045 ;
        RECT -32.125 94.355 -31.795 94.685 ;
        RECT -32.125 92.995 -31.795 93.325 ;
        RECT -32.125 91.635 -31.795 91.965 ;
        RECT -32.125 90.275 -31.795 90.605 ;
        RECT -32.125 88.915 -31.795 89.245 ;
        RECT -32.125 87.555 -31.795 87.885 ;
        RECT -32.125 86.195 -31.795 86.525 ;
        RECT -32.125 84.835 -31.795 85.165 ;
        RECT -32.125 83.475 -31.795 83.805 ;
        RECT -32.125 82.115 -31.795 82.445 ;
        RECT -32.125 80.755 -31.795 81.085 ;
        RECT -32.125 79.395 -31.795 79.725 ;
        RECT -32.125 78.035 -31.795 78.365 ;
        RECT -32.125 76.675 -31.795 77.005 ;
        RECT -32.125 75.315 -31.795 75.645 ;
        RECT -32.125 73.955 -31.795 74.285 ;
        RECT -32.125 72.595 -31.795 72.925 ;
        RECT -32.125 71.235 -31.795 71.565 ;
        RECT -32.125 69.875 -31.795 70.205 ;
        RECT -32.125 68.515 -31.795 68.845 ;
        RECT -32.125 67.155 -31.795 67.485 ;
        RECT -32.125 65.795 -31.795 66.125 ;
        RECT -32.125 64.435 -31.795 64.765 ;
        RECT -32.125 63.075 -31.795 63.405 ;
        RECT -32.125 61.715 -31.795 62.045 ;
        RECT -32.125 60.355 -31.795 60.685 ;
        RECT -32.125 58.995 -31.795 59.325 ;
        RECT -32.125 57.635 -31.795 57.965 ;
        RECT -32.125 56.275 -31.795 56.605 ;
        RECT -32.125 54.915 -31.795 55.245 ;
        RECT -32.125 53.555 -31.795 53.885 ;
        RECT -32.125 52.195 -31.795 52.525 ;
        RECT -32.125 50.835 -31.795 51.165 ;
        RECT -32.125 49.475 -31.795 49.805 ;
        RECT -32.125 48.115 -31.795 48.445 ;
        RECT -32.125 46.755 -31.795 47.085 ;
        RECT -32.125 45.395 -31.795 45.725 ;
        RECT -32.125 44.035 -31.795 44.365 ;
        RECT -32.125 42.675 -31.795 43.005 ;
        RECT -32.125 41.315 -31.795 41.645 ;
        RECT -32.125 39.955 -31.795 40.285 ;
        RECT -32.125 38.595 -31.795 38.925 ;
        RECT -32.125 37.235 -31.795 37.565 ;
        RECT -32.125 35.875 -31.795 36.205 ;
        RECT -32.125 34.515 -31.795 34.845 ;
        RECT -32.125 33.155 -31.795 33.485 ;
        RECT -32.125 31.795 -31.795 32.125 ;
        RECT -32.125 30.435 -31.795 30.765 ;
        RECT -32.125 29.075 -31.795 29.405 ;
        RECT -32.125 27.715 -31.795 28.045 ;
        RECT -32.125 26.355 -31.795 26.685 ;
        RECT -32.125 24.995 -31.795 25.325 ;
        RECT -32.125 23.635 -31.795 23.965 ;
        RECT -32.125 22.275 -31.795 22.605 ;
        RECT -32.125 20.915 -31.795 21.245 ;
        RECT -32.125 19.555 -31.795 19.885 ;
        RECT -32.125 18.195 -31.795 18.525 ;
        RECT -32.125 16.835 -31.795 17.165 ;
        RECT -32.125 15.475 -31.795 15.805 ;
        RECT -32.125 14.115 -31.795 14.445 ;
        RECT -32.125 12.755 -31.795 13.085 ;
        RECT -32.125 11.395 -31.795 11.725 ;
        RECT -32.125 10.035 -31.795 10.365 ;
        RECT -32.125 8.675 -31.795 9.005 ;
        RECT -32.125 7.315 -31.795 7.645 ;
        RECT -32.125 5.955 -31.795 6.285 ;
        RECT -32.125 4.595 -31.795 4.925 ;
        RECT -32.125 3.235 -31.795 3.565 ;
        RECT -32.125 1.875 -31.795 2.205 ;
        RECT -32.125 0.515 -31.795 0.845 ;
        RECT -32.125 -7.645 -31.795 -7.315 ;
        RECT -32.125 -11.725 -31.795 -11.395 ;
        RECT -32.125 -13.085 -31.795 -12.755 ;
        RECT -32.125 -14.445 -31.795 -14.115 ;
        RECT -32.125 -15.805 -31.795 -15.475 ;
        RECT -32.125 -17.165 -31.795 -16.835 ;
        RECT -32.125 -19.885 -31.795 -19.555 ;
        RECT -32.125 -21.245 -31.795 -20.915 ;
        RECT -32.125 -22.605 -31.795 -22.275 ;
        RECT -32.125 -29.405 -31.795 -29.075 ;
        RECT -32.125 -30.765 -31.795 -30.435 ;
        RECT -32.125 -32.125 -31.795 -31.795 ;
        RECT -32.125 -33.485 -31.795 -33.155 ;
        RECT -32.125 -34.845 -31.795 -34.515 ;
        RECT -32.125 -36.205 -31.795 -35.875 ;
        RECT -32.125 -37.565 -31.795 -37.235 ;
        RECT -32.125 -38.925 -31.795 -38.595 ;
        RECT -32.125 -40.285 -31.795 -39.955 ;
        RECT -32.125 -41.645 -31.795 -41.315 ;
        RECT -32.125 -43.005 -31.795 -42.675 ;
        RECT -32.125 -44.365 -31.795 -44.035 ;
        RECT -32.125 -45.725 -31.795 -45.395 ;
        RECT -32.125 -49.805 -31.795 -49.475 ;
        RECT -32.125 -51.165 -31.795 -50.835 ;
        RECT -32.125 -52.525 -31.795 -52.195 ;
        RECT -32.125 -53.885 -31.795 -53.555 ;
        RECT -32.125 -55.245 -31.795 -54.915 ;
        RECT -32.125 -56.605 -31.795 -56.275 ;
        RECT -32.125 -57.965 -31.795 -57.635 ;
        RECT -32.125 -59.325 -31.795 -58.995 ;
        RECT -32.125 -60.685 -31.795 -60.355 ;
        RECT -32.125 -62.045 -31.795 -61.715 ;
        RECT -32.125 -63.405 -31.795 -63.075 ;
        RECT -32.125 -64.765 -31.795 -64.435 ;
        RECT -32.125 -66.125 -31.795 -65.795 ;
        RECT -32.125 -67.485 -31.795 -67.155 ;
        RECT -32.125 -68.845 -31.795 -68.515 ;
        RECT -32.125 -70.37 -31.795 -70.04 ;
        RECT -32.125 -71.565 -31.795 -71.235 ;
        RECT -32.125 -72.925 -31.795 -72.595 ;
        RECT -32.125 -74.285 -31.795 -73.955 ;
        RECT -32.125 -75.645 -31.795 -75.315 ;
        RECT -32.125 -77.005 -31.795 -76.675 ;
        RECT -32.125 -79.725 -31.795 -79.395 ;
        RECT -32.125 -80.91 -31.795 -80.58 ;
        RECT -32.125 -82.445 -31.795 -82.115 ;
        RECT -32.125 -83.805 -31.795 -83.475 ;
        RECT -32.125 -85.165 -31.795 -84.835 ;
        RECT -32.125 -87.885 -31.795 -87.555 ;
        RECT -32.125 -89.245 -31.795 -88.915 ;
        RECT -32.125 -91.965 -31.795 -91.635 ;
        RECT -32.125 -93.325 -31.795 -92.995 ;
        RECT -32.125 -94.685 -31.795 -94.355 ;
        RECT -32.125 -96.045 -31.795 -95.715 ;
        RECT -32.125 -98.765 -31.795 -98.435 ;
        RECT -32.125 -100.125 -31.795 -99.795 ;
        RECT -32.125 -101.485 -31.795 -101.155 ;
        RECT -32.125 -102.845 -31.795 -102.515 ;
        RECT -32.125 -105.565 -31.795 -105.235 ;
        RECT -32.125 -106.925 -31.795 -106.595 ;
        RECT -32.125 -108.285 -31.795 -107.955 ;
        RECT -32.125 -112.365 -31.795 -112.035 ;
        RECT -32.125 -113.725 -31.795 -113.395 ;
        RECT -32.125 -115.085 -31.795 -114.755 ;
        RECT -32.125 -117.805 -31.795 -117.475 ;
        RECT -32.125 -120.525 -31.795 -120.195 ;
        RECT -32.125 -121.885 -31.795 -121.555 ;
        RECT -32.125 -123.245 -31.795 -122.915 ;
        RECT -32.125 -124.605 -31.795 -124.275 ;
        RECT -32.125 -125.965 -31.795 -125.635 ;
        RECT -32.125 -127.325 -31.795 -126.995 ;
        RECT -32.125 -130.045 -31.795 -129.715 ;
        RECT -32.125 -131.405 -31.795 -131.075 ;
        RECT -32.125 -135.485 -31.795 -135.155 ;
        RECT -32.125 -136.845 -31.795 -136.515 ;
        RECT -32.125 -138.205 -31.795 -137.875 ;
        RECT -32.125 -139.565 -31.795 -139.235 ;
        RECT -32.125 -140.925 -31.795 -140.595 ;
        RECT -32.125 -142.285 -31.795 -141.955 ;
        RECT -32.125 -143.645 -31.795 -143.315 ;
        RECT -32.125 -145.005 -31.795 -144.675 ;
        RECT -32.125 -146.365 -31.795 -146.035 ;
        RECT -32.125 -148.215 -31.795 -147.885 ;
        RECT -32.125 -149.085 -31.795 -148.755 ;
        RECT -32.125 -150.445 -31.795 -150.115 ;
        RECT -32.125 -153.165 -31.795 -152.835 ;
        RECT -32.125 -154.525 -31.795 -154.195 ;
        RECT -32.125 -157.245 -31.795 -156.915 ;
        RECT -32.125 -162.89 -31.795 -161.76 ;
        RECT -32.12 -163.005 -31.8 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 129.945 -30.435 131.075 ;
        RECT -30.765 125.635 -30.435 125.965 ;
        RECT -30.765 124.275 -30.435 124.605 ;
        RECT -30.765 122.915 -30.435 123.245 ;
        RECT -30.765 121.555 -30.435 121.885 ;
        RECT -30.765 120.195 -30.435 120.525 ;
        RECT -30.765 118.835 -30.435 119.165 ;
        RECT -30.765 117.475 -30.435 117.805 ;
        RECT -30.765 116.115 -30.435 116.445 ;
        RECT -30.765 114.755 -30.435 115.085 ;
        RECT -30.765 113.395 -30.435 113.725 ;
        RECT -30.765 112.035 -30.435 112.365 ;
        RECT -30.765 110.675 -30.435 111.005 ;
        RECT -30.765 109.315 -30.435 109.645 ;
        RECT -30.765 107.955 -30.435 108.285 ;
        RECT -30.765 106.595 -30.435 106.925 ;
        RECT -30.765 105.235 -30.435 105.565 ;
        RECT -30.765 103.875 -30.435 104.205 ;
        RECT -30.765 102.515 -30.435 102.845 ;
        RECT -30.765 101.155 -30.435 101.485 ;
        RECT -30.765 99.795 -30.435 100.125 ;
        RECT -30.765 98.435 -30.435 98.765 ;
        RECT -30.765 97.075 -30.435 97.405 ;
        RECT -30.765 95.715 -30.435 96.045 ;
        RECT -30.765 94.355 -30.435 94.685 ;
        RECT -30.765 92.995 -30.435 93.325 ;
        RECT -30.765 91.635 -30.435 91.965 ;
        RECT -30.765 90.275 -30.435 90.605 ;
        RECT -30.765 88.915 -30.435 89.245 ;
        RECT -30.765 87.555 -30.435 87.885 ;
        RECT -30.765 86.195 -30.435 86.525 ;
        RECT -30.765 84.835 -30.435 85.165 ;
        RECT -30.765 83.475 -30.435 83.805 ;
        RECT -30.765 82.115 -30.435 82.445 ;
        RECT -30.765 80.755 -30.435 81.085 ;
        RECT -30.765 79.395 -30.435 79.725 ;
        RECT -30.765 78.035 -30.435 78.365 ;
        RECT -30.765 76.675 -30.435 77.005 ;
        RECT -30.765 75.315 -30.435 75.645 ;
        RECT -30.765 73.955 -30.435 74.285 ;
        RECT -30.765 72.595 -30.435 72.925 ;
        RECT -30.765 71.235 -30.435 71.565 ;
        RECT -30.765 69.875 -30.435 70.205 ;
        RECT -30.765 68.515 -30.435 68.845 ;
        RECT -30.765 67.155 -30.435 67.485 ;
        RECT -30.765 65.795 -30.435 66.125 ;
        RECT -30.765 64.435 -30.435 64.765 ;
        RECT -30.765 63.075 -30.435 63.405 ;
        RECT -30.765 61.715 -30.435 62.045 ;
        RECT -30.765 60.355 -30.435 60.685 ;
        RECT -30.765 58.995 -30.435 59.325 ;
        RECT -30.765 57.635 -30.435 57.965 ;
        RECT -30.765 56.275 -30.435 56.605 ;
        RECT -30.765 54.915 -30.435 55.245 ;
        RECT -30.765 53.555 -30.435 53.885 ;
        RECT -30.765 52.195 -30.435 52.525 ;
        RECT -30.765 50.835 -30.435 51.165 ;
        RECT -30.765 49.475 -30.435 49.805 ;
        RECT -30.765 48.115 -30.435 48.445 ;
        RECT -30.765 46.755 -30.435 47.085 ;
        RECT -30.765 45.395 -30.435 45.725 ;
        RECT -30.765 44.035 -30.435 44.365 ;
        RECT -30.765 42.675 -30.435 43.005 ;
        RECT -30.765 41.315 -30.435 41.645 ;
        RECT -30.765 39.955 -30.435 40.285 ;
        RECT -30.765 38.595 -30.435 38.925 ;
        RECT -30.765 37.235 -30.435 37.565 ;
        RECT -30.765 35.875 -30.435 36.205 ;
        RECT -30.765 34.515 -30.435 34.845 ;
        RECT -30.765 33.155 -30.435 33.485 ;
        RECT -30.765 31.795 -30.435 32.125 ;
        RECT -30.765 30.435 -30.435 30.765 ;
        RECT -30.765 29.075 -30.435 29.405 ;
        RECT -30.765 27.715 -30.435 28.045 ;
        RECT -30.765 26.355 -30.435 26.685 ;
        RECT -30.765 24.995 -30.435 25.325 ;
        RECT -30.765 23.635 -30.435 23.965 ;
        RECT -30.765 22.275 -30.435 22.605 ;
        RECT -30.765 20.915 -30.435 21.245 ;
        RECT -30.765 19.555 -30.435 19.885 ;
        RECT -30.765 18.195 -30.435 18.525 ;
        RECT -30.765 16.835 -30.435 17.165 ;
        RECT -30.765 15.475 -30.435 15.805 ;
        RECT -30.765 14.115 -30.435 14.445 ;
        RECT -30.765 12.755 -30.435 13.085 ;
        RECT -30.765 11.395 -30.435 11.725 ;
        RECT -30.765 10.035 -30.435 10.365 ;
        RECT -30.765 8.675 -30.435 9.005 ;
        RECT -30.765 7.315 -30.435 7.645 ;
        RECT -30.765 5.955 -30.435 6.285 ;
        RECT -30.765 4.595 -30.435 4.925 ;
        RECT -30.765 3.235 -30.435 3.565 ;
        RECT -30.765 1.875 -30.435 2.205 ;
        RECT -30.765 0.515 -30.435 0.845 ;
        RECT -30.765 -7.645 -30.435 -7.315 ;
        RECT -30.765 -11.725 -30.435 -11.395 ;
        RECT -30.765 -13.085 -30.435 -12.755 ;
        RECT -30.765 -14.445 -30.435 -14.115 ;
        RECT -30.765 -15.805 -30.435 -15.475 ;
        RECT -30.765 -17.165 -30.435 -16.835 ;
        RECT -30.765 -19.885 -30.435 -19.555 ;
        RECT -30.765 -21.245 -30.435 -20.915 ;
        RECT -30.765 -22.605 -30.435 -22.275 ;
        RECT -30.765 -29.405 -30.435 -29.075 ;
        RECT -30.765 -30.765 -30.435 -30.435 ;
        RECT -30.765 -32.125 -30.435 -31.795 ;
        RECT -30.765 -33.485 -30.435 -33.155 ;
        RECT -30.765 -34.845 -30.435 -34.515 ;
        RECT -30.765 -36.205 -30.435 -35.875 ;
        RECT -30.765 -37.565 -30.435 -37.235 ;
        RECT -30.765 -38.925 -30.435 -38.595 ;
        RECT -30.765 -40.285 -30.435 -39.955 ;
        RECT -30.765 -41.645 -30.435 -41.315 ;
        RECT -30.765 -43.005 -30.435 -42.675 ;
        RECT -30.765 -44.365 -30.435 -44.035 ;
        RECT -30.765 -45.725 -30.435 -45.395 ;
        RECT -30.765 -49.805 -30.435 -49.475 ;
        RECT -30.765 -51.165 -30.435 -50.835 ;
        RECT -30.765 -52.525 -30.435 -52.195 ;
        RECT -30.765 -53.885 -30.435 -53.555 ;
        RECT -30.765 -55.245 -30.435 -54.915 ;
        RECT -30.765 -56.605 -30.435 -56.275 ;
        RECT -30.765 -57.965 -30.435 -57.635 ;
        RECT -30.765 -59.325 -30.435 -58.995 ;
        RECT -30.765 -60.685 -30.435 -60.355 ;
        RECT -30.765 -62.045 -30.435 -61.715 ;
        RECT -30.765 -63.405 -30.435 -63.075 ;
        RECT -30.765 -64.765 -30.435 -64.435 ;
        RECT -30.765 -66.125 -30.435 -65.795 ;
        RECT -30.765 -67.485 -30.435 -67.155 ;
        RECT -30.765 -68.845 -30.435 -68.515 ;
        RECT -30.765 -70.37 -30.435 -70.04 ;
        RECT -30.765 -71.565 -30.435 -71.235 ;
        RECT -30.765 -72.925 -30.435 -72.595 ;
        RECT -30.765 -74.285 -30.435 -73.955 ;
        RECT -30.765 -75.645 -30.435 -75.315 ;
        RECT -30.765 -77.005 -30.435 -76.675 ;
        RECT -30.765 -79.725 -30.435 -79.395 ;
        RECT -30.765 -80.91 -30.435 -80.58 ;
        RECT -30.765 -82.445 -30.435 -82.115 ;
        RECT -30.765 -83.805 -30.435 -83.475 ;
        RECT -30.765 -85.165 -30.435 -84.835 ;
        RECT -30.765 -87.885 -30.435 -87.555 ;
        RECT -30.765 -89.245 -30.435 -88.915 ;
        RECT -30.765 -91.965 -30.435 -91.635 ;
        RECT -30.765 -93.325 -30.435 -92.995 ;
        RECT -30.765 -94.685 -30.435 -94.355 ;
        RECT -30.765 -96.045 -30.435 -95.715 ;
        RECT -30.765 -98.765 -30.435 -98.435 ;
        RECT -30.765 -100.125 -30.435 -99.795 ;
        RECT -30.765 -101.485 -30.435 -101.155 ;
        RECT -30.765 -102.845 -30.435 -102.515 ;
        RECT -30.765 -105.565 -30.435 -105.235 ;
        RECT -30.765 -106.925 -30.435 -106.595 ;
        RECT -30.765 -108.285 -30.435 -107.955 ;
        RECT -30.765 -112.365 -30.435 -112.035 ;
        RECT -30.765 -113.725 -30.435 -113.395 ;
        RECT -30.765 -115.085 -30.435 -114.755 ;
        RECT -30.765 -117.805 -30.435 -117.475 ;
        RECT -30.765 -120.525 -30.435 -120.195 ;
        RECT -30.765 -121.885 -30.435 -121.555 ;
        RECT -30.765 -123.245 -30.435 -122.915 ;
        RECT -30.765 -124.605 -30.435 -124.275 ;
        RECT -30.765 -125.965 -30.435 -125.635 ;
        RECT -30.765 -127.325 -30.435 -126.995 ;
        RECT -30.765 -130.045 -30.435 -129.715 ;
        RECT -30.765 -131.405 -30.435 -131.075 ;
        RECT -30.765 -135.485 -30.435 -135.155 ;
        RECT -30.765 -136.845 -30.435 -136.515 ;
        RECT -30.765 -138.205 -30.435 -137.875 ;
        RECT -30.765 -139.565 -30.435 -139.235 ;
        RECT -30.765 -140.925 -30.435 -140.595 ;
        RECT -30.765 -142.285 -30.435 -141.955 ;
        RECT -30.765 -143.645 -30.435 -143.315 ;
        RECT -30.765 -145.005 -30.435 -144.675 ;
        RECT -30.765 -146.365 -30.435 -146.035 ;
        RECT -30.765 -148.215 -30.435 -147.885 ;
        RECT -30.765 -149.085 -30.435 -148.755 ;
        RECT -30.765 -150.445 -30.435 -150.115 ;
        RECT -30.765 -151.805 -30.435 -151.475 ;
        RECT -30.765 -153.165 -30.435 -152.835 ;
        RECT -30.765 -154.525 -30.435 -154.195 ;
        RECT -30.765 -157.245 -30.435 -156.915 ;
        RECT -30.765 -162.89 -30.435 -161.76 ;
        RECT -30.76 -163.005 -30.44 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 129.945 -29.075 131.075 ;
        RECT -29.405 125.635 -29.075 125.965 ;
        RECT -29.405 124.275 -29.075 124.605 ;
        RECT -29.405 122.915 -29.075 123.245 ;
        RECT -29.405 121.555 -29.075 121.885 ;
        RECT -29.405 120.195 -29.075 120.525 ;
        RECT -29.405 118.835 -29.075 119.165 ;
        RECT -29.405 117.475 -29.075 117.805 ;
        RECT -29.405 116.115 -29.075 116.445 ;
        RECT -29.405 114.755 -29.075 115.085 ;
        RECT -29.405 113.395 -29.075 113.725 ;
        RECT -29.405 112.035 -29.075 112.365 ;
        RECT -29.405 110.675 -29.075 111.005 ;
        RECT -29.405 109.315 -29.075 109.645 ;
        RECT -29.405 107.955 -29.075 108.285 ;
        RECT -29.405 106.595 -29.075 106.925 ;
        RECT -29.405 105.235 -29.075 105.565 ;
        RECT -29.405 103.875 -29.075 104.205 ;
        RECT -29.405 102.515 -29.075 102.845 ;
        RECT -29.405 101.155 -29.075 101.485 ;
        RECT -29.405 99.795 -29.075 100.125 ;
        RECT -29.405 98.435 -29.075 98.765 ;
        RECT -29.405 97.075 -29.075 97.405 ;
        RECT -29.405 95.715 -29.075 96.045 ;
        RECT -29.405 94.355 -29.075 94.685 ;
        RECT -29.405 92.995 -29.075 93.325 ;
        RECT -29.405 91.635 -29.075 91.965 ;
        RECT -29.405 90.275 -29.075 90.605 ;
        RECT -29.405 88.915 -29.075 89.245 ;
        RECT -29.405 87.555 -29.075 87.885 ;
        RECT -29.405 86.195 -29.075 86.525 ;
        RECT -29.405 84.835 -29.075 85.165 ;
        RECT -29.405 83.475 -29.075 83.805 ;
        RECT -29.405 82.115 -29.075 82.445 ;
        RECT -29.405 80.755 -29.075 81.085 ;
        RECT -29.405 79.395 -29.075 79.725 ;
        RECT -29.405 78.035 -29.075 78.365 ;
        RECT -29.405 76.675 -29.075 77.005 ;
        RECT -29.405 75.315 -29.075 75.645 ;
        RECT -29.405 73.955 -29.075 74.285 ;
        RECT -29.405 72.595 -29.075 72.925 ;
        RECT -29.405 71.235 -29.075 71.565 ;
        RECT -29.405 69.875 -29.075 70.205 ;
        RECT -29.405 68.515 -29.075 68.845 ;
        RECT -29.405 67.155 -29.075 67.485 ;
        RECT -29.405 65.795 -29.075 66.125 ;
        RECT -29.405 64.435 -29.075 64.765 ;
        RECT -29.405 63.075 -29.075 63.405 ;
        RECT -29.405 61.715 -29.075 62.045 ;
        RECT -29.405 60.355 -29.075 60.685 ;
        RECT -29.405 58.995 -29.075 59.325 ;
        RECT -29.405 57.635 -29.075 57.965 ;
        RECT -29.405 56.275 -29.075 56.605 ;
        RECT -29.405 54.915 -29.075 55.245 ;
        RECT -29.405 53.555 -29.075 53.885 ;
        RECT -29.405 52.195 -29.075 52.525 ;
        RECT -29.405 50.835 -29.075 51.165 ;
        RECT -29.405 49.475 -29.075 49.805 ;
        RECT -29.405 48.115 -29.075 48.445 ;
        RECT -29.405 46.755 -29.075 47.085 ;
        RECT -29.405 45.395 -29.075 45.725 ;
        RECT -29.405 44.035 -29.075 44.365 ;
        RECT -29.405 42.675 -29.075 43.005 ;
        RECT -29.405 41.315 -29.075 41.645 ;
        RECT -29.405 39.955 -29.075 40.285 ;
        RECT -29.405 38.595 -29.075 38.925 ;
        RECT -29.405 37.235 -29.075 37.565 ;
        RECT -29.405 35.875 -29.075 36.205 ;
        RECT -29.405 34.515 -29.075 34.845 ;
        RECT -29.405 33.155 -29.075 33.485 ;
        RECT -29.405 31.795 -29.075 32.125 ;
        RECT -29.405 30.435 -29.075 30.765 ;
        RECT -29.405 29.075 -29.075 29.405 ;
        RECT -29.405 27.715 -29.075 28.045 ;
        RECT -29.405 26.355 -29.075 26.685 ;
        RECT -29.405 24.995 -29.075 25.325 ;
        RECT -29.405 23.635 -29.075 23.965 ;
        RECT -29.405 22.275 -29.075 22.605 ;
        RECT -29.405 20.915 -29.075 21.245 ;
        RECT -29.405 19.555 -29.075 19.885 ;
        RECT -29.405 18.195 -29.075 18.525 ;
        RECT -29.405 16.835 -29.075 17.165 ;
        RECT -29.405 15.475 -29.075 15.805 ;
        RECT -29.405 14.115 -29.075 14.445 ;
        RECT -29.405 12.755 -29.075 13.085 ;
        RECT -29.405 11.395 -29.075 11.725 ;
        RECT -29.405 10.035 -29.075 10.365 ;
        RECT -29.405 8.675 -29.075 9.005 ;
        RECT -29.405 7.315 -29.075 7.645 ;
        RECT -29.405 5.955 -29.075 6.285 ;
        RECT -29.405 4.595 -29.075 4.925 ;
        RECT -29.405 3.235 -29.075 3.565 ;
        RECT -29.405 1.875 -29.075 2.205 ;
        RECT -29.405 0.515 -29.075 0.845 ;
        RECT -29.405 -8.19 -29.075 -7.86 ;
        RECT -29.405 -11.725 -29.075 -11.395 ;
        RECT -29.405 -14.23 -29.075 -13.9 ;
        RECT -29.405 -15.805 -29.075 -15.475 ;
        RECT -29.405 -29.405 -29.075 -29.075 ;
        RECT -29.405 -31.17 -29.075 -30.84 ;
        RECT -29.405 -32.125 -29.075 -31.795 ;
        RECT -29.405 -33.485 -29.075 -33.155 ;
        RECT -29.405 -36.205 -29.075 -35.875 ;
        RECT -29.405 -37.21 -29.075 -36.88 ;
        RECT -29.405 -38.925 -29.075 -38.595 ;
        RECT -29.405 -41.645 -29.075 -41.315 ;
        RECT -29.405 -51.165 -29.075 -50.835 ;
        RECT -29.405 -52.525 -29.075 -52.195 ;
        RECT -29.405 -53.885 -29.075 -53.555 ;
        RECT -29.405 -55.245 -29.075 -54.915 ;
        RECT -29.405 -56.605 -29.075 -56.275 ;
        RECT -29.405 -57.965 -29.075 -57.635 ;
        RECT -29.405 -59.325 -29.075 -58.995 ;
        RECT -29.405 -60.685 -29.075 -60.355 ;
        RECT -29.405 -62.045 -29.075 -61.715 ;
        RECT -29.405 -63.405 -29.075 -63.075 ;
        RECT -29.405 -64.765 -29.075 -64.435 ;
        RECT -29.405 -66.125 -29.075 -65.795 ;
        RECT -29.405 -67.485 -29.075 -67.155 ;
        RECT -29.405 -68.845 -29.075 -68.515 ;
        RECT -29.405 -70.37 -29.075 -70.04 ;
        RECT -29.405 -71.565 -29.075 -71.235 ;
        RECT -29.405 -72.925 -29.075 -72.595 ;
        RECT -29.405 -74.285 -29.075 -73.955 ;
        RECT -29.405 -75.645 -29.075 -75.315 ;
        RECT -29.405 -77.005 -29.075 -76.675 ;
        RECT -29.405 -79.725 -29.075 -79.395 ;
        RECT -29.405 -80.91 -29.075 -80.58 ;
        RECT -29.405 -82.445 -29.075 -82.115 ;
        RECT -29.405 -83.805 -29.075 -83.475 ;
        RECT -29.405 -85.165 -29.075 -84.835 ;
        RECT -29.405 -87.885 -29.075 -87.555 ;
        RECT -29.405 -89.245 -29.075 -88.915 ;
        RECT -29.4 -91.96 -29.08 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -154.525 -29.075 -154.195 ;
        RECT -29.405 -157.245 -29.075 -156.915 ;
        RECT -29.405 -162.89 -29.075 -161.76 ;
        RECT -29.4 -163.005 -29.08 -153.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.045 118.835 -27.715 119.165 ;
        RECT -28.045 117.475 -27.715 117.805 ;
        RECT -28.045 116.115 -27.715 116.445 ;
        RECT -28.045 114.755 -27.715 115.085 ;
        RECT -28.045 113.395 -27.715 113.725 ;
        RECT -28.045 112.035 -27.715 112.365 ;
        RECT -28.045 110.675 -27.715 111.005 ;
        RECT -28.045 109.315 -27.715 109.645 ;
        RECT -28.045 107.955 -27.715 108.285 ;
        RECT -28.045 106.595 -27.715 106.925 ;
        RECT -28.045 105.235 -27.715 105.565 ;
        RECT -28.045 103.875 -27.715 104.205 ;
        RECT -28.045 102.515 -27.715 102.845 ;
        RECT -28.045 101.155 -27.715 101.485 ;
        RECT -28.045 99.795 -27.715 100.125 ;
        RECT -28.045 98.435 -27.715 98.765 ;
        RECT -28.045 97.075 -27.715 97.405 ;
        RECT -28.045 95.715 -27.715 96.045 ;
        RECT -28.045 94.355 -27.715 94.685 ;
        RECT -28.045 92.995 -27.715 93.325 ;
        RECT -28.045 91.635 -27.715 91.965 ;
        RECT -28.045 90.275 -27.715 90.605 ;
        RECT -28.045 88.915 -27.715 89.245 ;
        RECT -28.045 87.555 -27.715 87.885 ;
        RECT -28.045 86.195 -27.715 86.525 ;
        RECT -28.045 84.835 -27.715 85.165 ;
        RECT -28.045 83.475 -27.715 83.805 ;
        RECT -28.045 82.115 -27.715 82.445 ;
        RECT -28.045 80.755 -27.715 81.085 ;
        RECT -28.045 79.395 -27.715 79.725 ;
        RECT -28.045 78.035 -27.715 78.365 ;
        RECT -28.045 76.675 -27.715 77.005 ;
        RECT -28.045 75.315 -27.715 75.645 ;
        RECT -28.045 73.955 -27.715 74.285 ;
        RECT -28.045 72.595 -27.715 72.925 ;
        RECT -28.045 71.235 -27.715 71.565 ;
        RECT -28.045 69.875 -27.715 70.205 ;
        RECT -28.045 68.515 -27.715 68.845 ;
        RECT -28.045 67.155 -27.715 67.485 ;
        RECT -28.045 65.795 -27.715 66.125 ;
        RECT -28.045 64.435 -27.715 64.765 ;
        RECT -28.045 63.075 -27.715 63.405 ;
        RECT -28.045 61.715 -27.715 62.045 ;
        RECT -28.045 60.355 -27.715 60.685 ;
        RECT -28.045 58.995 -27.715 59.325 ;
        RECT -28.045 57.635 -27.715 57.965 ;
        RECT -28.045 56.275 -27.715 56.605 ;
        RECT -28.045 54.915 -27.715 55.245 ;
        RECT -28.045 53.555 -27.715 53.885 ;
        RECT -28.045 52.195 -27.715 52.525 ;
        RECT -28.045 50.835 -27.715 51.165 ;
        RECT -28.045 49.475 -27.715 49.805 ;
        RECT -28.045 48.115 -27.715 48.445 ;
        RECT -28.045 46.755 -27.715 47.085 ;
        RECT -28.045 45.395 -27.715 45.725 ;
        RECT -28.045 44.035 -27.715 44.365 ;
        RECT -28.045 42.675 -27.715 43.005 ;
        RECT -28.045 41.315 -27.715 41.645 ;
        RECT -28.045 39.955 -27.715 40.285 ;
        RECT -28.045 38.595 -27.715 38.925 ;
        RECT -28.045 37.235 -27.715 37.565 ;
        RECT -28.045 35.875 -27.715 36.205 ;
        RECT -28.045 34.515 -27.715 34.845 ;
        RECT -28.045 33.155 -27.715 33.485 ;
        RECT -28.045 31.795 -27.715 32.125 ;
        RECT -28.045 30.435 -27.715 30.765 ;
        RECT -28.045 29.075 -27.715 29.405 ;
        RECT -28.045 27.715 -27.715 28.045 ;
        RECT -28.045 26.355 -27.715 26.685 ;
        RECT -28.045 24.995 -27.715 25.325 ;
        RECT -28.045 23.635 -27.715 23.965 ;
        RECT -28.045 22.275 -27.715 22.605 ;
        RECT -28.045 20.915 -27.715 21.245 ;
        RECT -28.045 19.555 -27.715 19.885 ;
        RECT -28.045 18.195 -27.715 18.525 ;
        RECT -28.045 16.835 -27.715 17.165 ;
        RECT -28.045 15.475 -27.715 15.805 ;
        RECT -28.045 14.115 -27.715 14.445 ;
        RECT -28.045 12.755 -27.715 13.085 ;
        RECT -28.045 11.395 -27.715 11.725 ;
        RECT -28.045 10.035 -27.715 10.365 ;
        RECT -28.045 8.675 -27.715 9.005 ;
        RECT -28.045 7.315 -27.715 7.645 ;
        RECT -28.045 5.955 -27.715 6.285 ;
        RECT -28.045 4.595 -27.715 4.925 ;
        RECT -28.045 3.235 -27.715 3.565 ;
        RECT -28.045 1.875 -27.715 2.205 ;
        RECT -28.045 0.515 -27.715 0.845 ;
        RECT -28.045 -8.19 -27.715 -7.86 ;
        RECT -28.045 -11.725 -27.715 -11.395 ;
        RECT -28.045 -14.23 -27.715 -13.9 ;
        RECT -28.045 -15.805 -27.715 -15.475 ;
        RECT -28.045 -29.405 -27.715 -29.075 ;
        RECT -28.045 -31.17 -27.715 -30.84 ;
        RECT -28.045 -32.125 -27.715 -31.795 ;
        RECT -28.045 -33.485 -27.715 -33.155 ;
        RECT -28.045 -36.205 -27.715 -35.875 ;
        RECT -28.045 -37.21 -27.715 -36.88 ;
        RECT -28.045 -38.925 -27.715 -38.595 ;
        RECT -28.045 -41.645 -27.715 -41.315 ;
        RECT -28.045 -51.165 -27.715 -50.835 ;
        RECT -28.045 -52.525 -27.715 -52.195 ;
        RECT -28.045 -53.885 -27.715 -53.555 ;
        RECT -28.045 -55.245 -27.715 -54.915 ;
        RECT -28.045 -56.605 -27.715 -56.275 ;
        RECT -28.045 -57.965 -27.715 -57.635 ;
        RECT -28.045 -59.325 -27.715 -58.995 ;
        RECT -28.045 -60.685 -27.715 -60.355 ;
        RECT -28.045 -62.045 -27.715 -61.715 ;
        RECT -28.045 -63.405 -27.715 -63.075 ;
        RECT -28.045 -64.765 -27.715 -64.435 ;
        RECT -28.045 -66.125 -27.715 -65.795 ;
        RECT -28.045 -67.485 -27.715 -67.155 ;
        RECT -28.045 -68.845 -27.715 -68.515 ;
        RECT -28.045 -70.37 -27.715 -70.04 ;
        RECT -28.045 -71.565 -27.715 -71.235 ;
        RECT -28.045 -72.925 -27.715 -72.595 ;
        RECT -28.045 -74.285 -27.715 -73.955 ;
        RECT -28.045 -75.645 -27.715 -75.315 ;
        RECT -28.045 -77.005 -27.715 -76.675 ;
        RECT -28.045 -79.725 -27.715 -79.395 ;
        RECT -28.045 -80.91 -27.715 -80.58 ;
        RECT -28.045 -82.445 -27.715 -82.115 ;
        RECT -28.045 -83.805 -27.715 -83.475 ;
        RECT -28.045 -85.165 -27.715 -84.835 ;
        RECT -28.045 -87.885 -27.715 -87.555 ;
        RECT -28.045 -89.245 -27.715 -88.915 ;
        RECT -28.045 -91.965 -27.715 -91.635 ;
        RECT -28.045 -93.325 -27.715 -92.995 ;
        RECT -28.045 -94.685 -27.715 -94.355 ;
        RECT -28.045 -96.045 -27.715 -95.715 ;
        RECT -28.045 -98.765 -27.715 -98.435 ;
        RECT -28.045 -100.125 -27.715 -99.795 ;
        RECT -28.045 -101.485 -27.715 -101.155 ;
        RECT -28.045 -102.845 -27.715 -102.515 ;
        RECT -28.045 -105.565 -27.715 -105.235 ;
        RECT -28.045 -106.925 -27.715 -106.595 ;
        RECT -28.045 -108.285 -27.715 -107.955 ;
        RECT -28.045 -112.365 -27.715 -112.035 ;
        RECT -28.045 -113.725 -27.715 -113.395 ;
        RECT -28.045 -115.085 -27.715 -114.755 ;
        RECT -28.045 -117.805 -27.715 -117.475 ;
        RECT -28.045 -120.525 -27.715 -120.195 ;
        RECT -28.045 -121.885 -27.715 -121.555 ;
        RECT -28.045 -123.245 -27.715 -122.915 ;
        RECT -28.045 -124.605 -27.715 -124.275 ;
        RECT -28.045 -125.965 -27.715 -125.635 ;
        RECT -28.045 -127.325 -27.715 -126.995 ;
        RECT -28.045 -131.405 -27.715 -131.075 ;
        RECT -28.045 -135.485 -27.715 -135.155 ;
        RECT -28.045 -136.845 -27.715 -136.515 ;
        RECT -28.045 -138.205 -27.715 -137.875 ;
        RECT -28.045 -139.565 -27.715 -139.235 ;
        RECT -28.045 -140.925 -27.715 -140.595 ;
        RECT -28.045 -142.285 -27.715 -141.955 ;
        RECT -28.045 -143.645 -27.715 -143.315 ;
        RECT -28.045 -145.005 -27.715 -144.675 ;
        RECT -28.045 -146.365 -27.715 -146.035 ;
        RECT -28.045 -148.215 -27.715 -147.885 ;
        RECT -28.045 -149.085 -27.715 -148.755 ;
        RECT -28.045 -150.445 -27.715 -150.115 ;
        RECT -28.045 -151.805 -27.715 -151.475 ;
        RECT -28.045 -153.165 -27.715 -152.835 ;
        RECT -28.045 -154.525 -27.715 -154.195 ;
        RECT -28.045 -157.245 -27.715 -156.915 ;
        RECT -28.045 -162.89 -27.715 -161.76 ;
        RECT -28.04 -163.005 -27.72 131.19 ;
        RECT -28.045 129.945 -27.715 131.075 ;
        RECT -28.045 125.635 -27.715 125.965 ;
        RECT -28.045 124.275 -27.715 124.605 ;
        RECT -28.045 122.915 -27.715 123.245 ;
        RECT -28.045 121.555 -27.715 121.885 ;
        RECT -28.045 120.195 -27.715 120.525 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 129.945 -41.315 131.075 ;
        RECT -41.645 125.635 -41.315 125.965 ;
        RECT -41.645 124.275 -41.315 124.605 ;
        RECT -41.645 122.915 -41.315 123.245 ;
        RECT -41.645 121.555 -41.315 121.885 ;
        RECT -41.645 120.195 -41.315 120.525 ;
        RECT -41.645 118.835 -41.315 119.165 ;
        RECT -41.645 117.475 -41.315 117.805 ;
        RECT -41.645 116.115 -41.315 116.445 ;
        RECT -41.645 114.755 -41.315 115.085 ;
        RECT -41.645 113.395 -41.315 113.725 ;
        RECT -41.645 112.035 -41.315 112.365 ;
        RECT -41.645 110.675 -41.315 111.005 ;
        RECT -41.645 109.315 -41.315 109.645 ;
        RECT -41.645 107.955 -41.315 108.285 ;
        RECT -41.645 106.595 -41.315 106.925 ;
        RECT -41.645 105.235 -41.315 105.565 ;
        RECT -41.645 103.875 -41.315 104.205 ;
        RECT -41.645 102.515 -41.315 102.845 ;
        RECT -41.645 101.155 -41.315 101.485 ;
        RECT -41.645 99.795 -41.315 100.125 ;
        RECT -41.645 98.435 -41.315 98.765 ;
        RECT -41.645 97.075 -41.315 97.405 ;
        RECT -41.645 95.715 -41.315 96.045 ;
        RECT -41.645 94.355 -41.315 94.685 ;
        RECT -41.645 92.995 -41.315 93.325 ;
        RECT -41.645 91.635 -41.315 91.965 ;
        RECT -41.645 90.275 -41.315 90.605 ;
        RECT -41.645 88.915 -41.315 89.245 ;
        RECT -41.645 87.555 -41.315 87.885 ;
        RECT -41.645 86.195 -41.315 86.525 ;
        RECT -41.645 84.835 -41.315 85.165 ;
        RECT -41.645 83.475 -41.315 83.805 ;
        RECT -41.645 82.115 -41.315 82.445 ;
        RECT -41.645 80.755 -41.315 81.085 ;
        RECT -41.645 79.395 -41.315 79.725 ;
        RECT -41.645 78.035 -41.315 78.365 ;
        RECT -41.645 76.675 -41.315 77.005 ;
        RECT -41.645 75.315 -41.315 75.645 ;
        RECT -41.645 73.955 -41.315 74.285 ;
        RECT -41.645 72.595 -41.315 72.925 ;
        RECT -41.645 71.235 -41.315 71.565 ;
        RECT -41.645 69.875 -41.315 70.205 ;
        RECT -41.645 68.515 -41.315 68.845 ;
        RECT -41.645 67.155 -41.315 67.485 ;
        RECT -41.645 65.795 -41.315 66.125 ;
        RECT -41.645 64.435 -41.315 64.765 ;
        RECT -41.645 63.075 -41.315 63.405 ;
        RECT -41.645 61.715 -41.315 62.045 ;
        RECT -41.645 60.355 -41.315 60.685 ;
        RECT -41.645 58.995 -41.315 59.325 ;
        RECT -41.645 57.635 -41.315 57.965 ;
        RECT -41.645 56.275 -41.315 56.605 ;
        RECT -41.645 54.915 -41.315 55.245 ;
        RECT -41.645 53.555 -41.315 53.885 ;
        RECT -41.645 52.195 -41.315 52.525 ;
        RECT -41.645 50.835 -41.315 51.165 ;
        RECT -41.645 49.475 -41.315 49.805 ;
        RECT -41.645 48.115 -41.315 48.445 ;
        RECT -41.645 46.755 -41.315 47.085 ;
        RECT -41.645 45.395 -41.315 45.725 ;
        RECT -41.645 44.035 -41.315 44.365 ;
        RECT -41.645 42.675 -41.315 43.005 ;
        RECT -41.645 41.315 -41.315 41.645 ;
        RECT -41.645 39.955 -41.315 40.285 ;
        RECT -41.645 38.595 -41.315 38.925 ;
        RECT -41.645 37.235 -41.315 37.565 ;
        RECT -41.645 35.875 -41.315 36.205 ;
        RECT -41.645 34.515 -41.315 34.845 ;
        RECT -41.645 33.155 -41.315 33.485 ;
        RECT -41.645 31.795 -41.315 32.125 ;
        RECT -41.645 30.435 -41.315 30.765 ;
        RECT -41.645 29.075 -41.315 29.405 ;
        RECT -41.645 27.715 -41.315 28.045 ;
        RECT -41.645 26.355 -41.315 26.685 ;
        RECT -41.645 24.995 -41.315 25.325 ;
        RECT -41.645 23.635 -41.315 23.965 ;
        RECT -41.645 22.275 -41.315 22.605 ;
        RECT -41.645 20.915 -41.315 21.245 ;
        RECT -41.645 19.555 -41.315 19.885 ;
        RECT -41.645 18.195 -41.315 18.525 ;
        RECT -41.645 16.835 -41.315 17.165 ;
        RECT -41.645 15.475 -41.315 15.805 ;
        RECT -41.645 14.115 -41.315 14.445 ;
        RECT -41.645 12.755 -41.315 13.085 ;
        RECT -41.645 11.395 -41.315 11.725 ;
        RECT -41.645 10.035 -41.315 10.365 ;
        RECT -41.645 8.675 -41.315 9.005 ;
        RECT -41.645 7.315 -41.315 7.645 ;
        RECT -41.645 5.955 -41.315 6.285 ;
        RECT -41.645 4.595 -41.315 4.925 ;
        RECT -41.645 3.235 -41.315 3.565 ;
        RECT -41.645 1.875 -41.315 2.205 ;
        RECT -41.645 0.515 -41.315 0.845 ;
        RECT -41.645 -0.845 -41.315 -0.515 ;
        RECT -41.645 -2.205 -41.315 -1.875 ;
        RECT -41.645 -3.565 -41.315 -3.235 ;
        RECT -41.645 -4.925 -41.315 -4.595 ;
        RECT -41.645 -7.645 -41.315 -7.315 ;
        RECT -41.645 -11.725 -41.315 -11.395 ;
        RECT -41.645 -13.085 -41.315 -12.755 ;
        RECT -41.645 -14.445 -41.315 -14.115 ;
        RECT -41.645 -15.805 -41.315 -15.475 ;
        RECT -41.645 -17.165 -41.315 -16.835 ;
        RECT -41.645 -19.885 -41.315 -19.555 ;
        RECT -41.645 -21.245 -41.315 -20.915 ;
        RECT -41.645 -22.605 -41.315 -22.275 ;
        RECT -41.645 -29.405 -41.315 -29.075 ;
        RECT -41.645 -30.765 -41.315 -30.435 ;
        RECT -41.645 -32.125 -41.315 -31.795 ;
        RECT -41.645 -33.485 -41.315 -33.155 ;
        RECT -41.645 -34.845 -41.315 -34.515 ;
        RECT -41.645 -36.205 -41.315 -35.875 ;
        RECT -41.645 -37.565 -41.315 -37.235 ;
        RECT -41.645 -38.925 -41.315 -38.595 ;
        RECT -41.645 -40.285 -41.315 -39.955 ;
        RECT -41.645 -41.645 -41.315 -41.315 ;
        RECT -41.645 -43.005 -41.315 -42.675 ;
        RECT -41.645 -44.365 -41.315 -44.035 ;
        RECT -41.645 -45.725 -41.315 -45.395 ;
        RECT -41.645 -47.085 -41.315 -46.755 ;
        RECT -41.645 -48.445 -41.315 -48.115 ;
        RECT -41.645 -49.805 -41.315 -49.475 ;
        RECT -41.645 -51.165 -41.315 -50.835 ;
        RECT -41.645 -52.525 -41.315 -52.195 ;
        RECT -41.645 -53.885 -41.315 -53.555 ;
        RECT -41.645 -55.245 -41.315 -54.915 ;
        RECT -41.645 -56.605 -41.315 -56.275 ;
        RECT -41.645 -57.965 -41.315 -57.635 ;
        RECT -41.645 -59.325 -41.315 -58.995 ;
        RECT -41.645 -60.685 -41.315 -60.355 ;
        RECT -41.645 -62.045 -41.315 -61.715 ;
        RECT -41.645 -63.405 -41.315 -63.075 ;
        RECT -41.645 -64.765 -41.315 -64.435 ;
        RECT -41.645 -66.125 -41.315 -65.795 ;
        RECT -41.645 -67.485 -41.315 -67.155 ;
        RECT -41.645 -68.845 -41.315 -68.515 ;
        RECT -41.645 -70.37 -41.315 -70.04 ;
        RECT -41.645 -71.565 -41.315 -71.235 ;
        RECT -41.645 -72.925 -41.315 -72.595 ;
        RECT -41.645 -74.285 -41.315 -73.955 ;
        RECT -41.645 -75.645 -41.315 -75.315 ;
        RECT -41.645 -77.005 -41.315 -76.675 ;
        RECT -41.645 -79.725 -41.315 -79.395 ;
        RECT -41.645 -80.91 -41.315 -80.58 ;
        RECT -41.645 -82.445 -41.315 -82.115 ;
        RECT -41.645 -83.805 -41.315 -83.475 ;
        RECT -41.645 -85.165 -41.315 -84.835 ;
        RECT -41.645 -87.885 -41.315 -87.555 ;
        RECT -41.645 -89.245 -41.315 -88.915 ;
        RECT -41.64 -91.28 -41.32 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 -154.525 -41.315 -154.195 ;
        RECT -41.645 -157.245 -41.315 -156.915 ;
        RECT -41.645 -162.89 -41.315 -161.76 ;
        RECT -41.64 -163.005 -41.32 -152.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.285 129.945 -39.955 131.075 ;
        RECT -40.285 125.635 -39.955 125.965 ;
        RECT -40.285 124.275 -39.955 124.605 ;
        RECT -40.285 122.915 -39.955 123.245 ;
        RECT -40.285 121.555 -39.955 121.885 ;
        RECT -40.285 120.195 -39.955 120.525 ;
        RECT -40.285 118.835 -39.955 119.165 ;
        RECT -40.285 117.475 -39.955 117.805 ;
        RECT -40.285 116.115 -39.955 116.445 ;
        RECT -40.285 114.755 -39.955 115.085 ;
        RECT -40.285 113.395 -39.955 113.725 ;
        RECT -40.285 112.035 -39.955 112.365 ;
        RECT -40.285 110.675 -39.955 111.005 ;
        RECT -40.285 109.315 -39.955 109.645 ;
        RECT -40.285 107.955 -39.955 108.285 ;
        RECT -40.285 106.595 -39.955 106.925 ;
        RECT -40.285 105.235 -39.955 105.565 ;
        RECT -40.285 103.875 -39.955 104.205 ;
        RECT -40.285 102.515 -39.955 102.845 ;
        RECT -40.285 101.155 -39.955 101.485 ;
        RECT -40.285 99.795 -39.955 100.125 ;
        RECT -40.285 98.435 -39.955 98.765 ;
        RECT -40.285 97.075 -39.955 97.405 ;
        RECT -40.285 95.715 -39.955 96.045 ;
        RECT -40.285 94.355 -39.955 94.685 ;
        RECT -40.285 92.995 -39.955 93.325 ;
        RECT -40.285 91.635 -39.955 91.965 ;
        RECT -40.285 90.275 -39.955 90.605 ;
        RECT -40.285 88.915 -39.955 89.245 ;
        RECT -40.285 87.555 -39.955 87.885 ;
        RECT -40.285 86.195 -39.955 86.525 ;
        RECT -40.285 84.835 -39.955 85.165 ;
        RECT -40.285 83.475 -39.955 83.805 ;
        RECT -40.285 82.115 -39.955 82.445 ;
        RECT -40.285 80.755 -39.955 81.085 ;
        RECT -40.285 79.395 -39.955 79.725 ;
        RECT -40.285 78.035 -39.955 78.365 ;
        RECT -40.285 76.675 -39.955 77.005 ;
        RECT -40.285 75.315 -39.955 75.645 ;
        RECT -40.285 73.955 -39.955 74.285 ;
        RECT -40.285 72.595 -39.955 72.925 ;
        RECT -40.285 71.235 -39.955 71.565 ;
        RECT -40.285 69.875 -39.955 70.205 ;
        RECT -40.285 68.515 -39.955 68.845 ;
        RECT -40.285 67.155 -39.955 67.485 ;
        RECT -40.285 65.795 -39.955 66.125 ;
        RECT -40.285 64.435 -39.955 64.765 ;
        RECT -40.285 63.075 -39.955 63.405 ;
        RECT -40.285 61.715 -39.955 62.045 ;
        RECT -40.285 60.355 -39.955 60.685 ;
        RECT -40.285 58.995 -39.955 59.325 ;
        RECT -40.285 57.635 -39.955 57.965 ;
        RECT -40.285 56.275 -39.955 56.605 ;
        RECT -40.285 54.915 -39.955 55.245 ;
        RECT -40.285 53.555 -39.955 53.885 ;
        RECT -40.285 52.195 -39.955 52.525 ;
        RECT -40.285 50.835 -39.955 51.165 ;
        RECT -40.285 49.475 -39.955 49.805 ;
        RECT -40.285 48.115 -39.955 48.445 ;
        RECT -40.285 46.755 -39.955 47.085 ;
        RECT -40.285 45.395 -39.955 45.725 ;
        RECT -40.285 44.035 -39.955 44.365 ;
        RECT -40.285 42.675 -39.955 43.005 ;
        RECT -40.285 41.315 -39.955 41.645 ;
        RECT -40.285 39.955 -39.955 40.285 ;
        RECT -40.285 38.595 -39.955 38.925 ;
        RECT -40.285 37.235 -39.955 37.565 ;
        RECT -40.285 35.875 -39.955 36.205 ;
        RECT -40.285 34.515 -39.955 34.845 ;
        RECT -40.285 33.155 -39.955 33.485 ;
        RECT -40.285 31.795 -39.955 32.125 ;
        RECT -40.285 30.435 -39.955 30.765 ;
        RECT -40.285 29.075 -39.955 29.405 ;
        RECT -40.285 27.715 -39.955 28.045 ;
        RECT -40.285 26.355 -39.955 26.685 ;
        RECT -40.285 24.995 -39.955 25.325 ;
        RECT -40.285 23.635 -39.955 23.965 ;
        RECT -40.285 22.275 -39.955 22.605 ;
        RECT -40.285 20.915 -39.955 21.245 ;
        RECT -40.285 19.555 -39.955 19.885 ;
        RECT -40.285 18.195 -39.955 18.525 ;
        RECT -40.285 16.835 -39.955 17.165 ;
        RECT -40.285 15.475 -39.955 15.805 ;
        RECT -40.285 14.115 -39.955 14.445 ;
        RECT -40.285 12.755 -39.955 13.085 ;
        RECT -40.285 11.395 -39.955 11.725 ;
        RECT -40.285 10.035 -39.955 10.365 ;
        RECT -40.285 8.675 -39.955 9.005 ;
        RECT -40.285 7.315 -39.955 7.645 ;
        RECT -40.285 5.955 -39.955 6.285 ;
        RECT -40.285 4.595 -39.955 4.925 ;
        RECT -40.285 3.235 -39.955 3.565 ;
        RECT -40.285 1.875 -39.955 2.205 ;
        RECT -40.285 0.515 -39.955 0.845 ;
        RECT -40.285 -0.845 -39.955 -0.515 ;
        RECT -40.285 -2.205 -39.955 -1.875 ;
        RECT -40.285 -3.565 -39.955 -3.235 ;
        RECT -40.285 -7.645 -39.955 -7.315 ;
        RECT -40.285 -11.725 -39.955 -11.395 ;
        RECT -40.285 -13.085 -39.955 -12.755 ;
        RECT -40.285 -14.445 -39.955 -14.115 ;
        RECT -40.285 -15.805 -39.955 -15.475 ;
        RECT -40.285 -17.165 -39.955 -16.835 ;
        RECT -40.285 -19.885 -39.955 -19.555 ;
        RECT -40.285 -21.245 -39.955 -20.915 ;
        RECT -40.285 -22.605 -39.955 -22.275 ;
        RECT -40.285 -29.405 -39.955 -29.075 ;
        RECT -40.285 -30.765 -39.955 -30.435 ;
        RECT -40.285 -32.125 -39.955 -31.795 ;
        RECT -40.285 -33.485 -39.955 -33.155 ;
        RECT -40.285 -34.845 -39.955 -34.515 ;
        RECT -40.285 -36.205 -39.955 -35.875 ;
        RECT -40.285 -37.565 -39.955 -37.235 ;
        RECT -40.285 -38.925 -39.955 -38.595 ;
        RECT -40.285 -40.285 -39.955 -39.955 ;
        RECT -40.285 -41.645 -39.955 -41.315 ;
        RECT -40.285 -43.005 -39.955 -42.675 ;
        RECT -40.285 -44.365 -39.955 -44.035 ;
        RECT -40.285 -45.725 -39.955 -45.395 ;
        RECT -40.285 -47.085 -39.955 -46.755 ;
        RECT -40.285 -48.445 -39.955 -48.115 ;
        RECT -40.285 -49.805 -39.955 -49.475 ;
        RECT -40.285 -51.165 -39.955 -50.835 ;
        RECT -40.285 -52.525 -39.955 -52.195 ;
        RECT -40.285 -53.885 -39.955 -53.555 ;
        RECT -40.285 -55.245 -39.955 -54.915 ;
        RECT -40.285 -56.605 -39.955 -56.275 ;
        RECT -40.285 -57.965 -39.955 -57.635 ;
        RECT -40.285 -59.325 -39.955 -58.995 ;
        RECT -40.285 -60.685 -39.955 -60.355 ;
        RECT -40.285 -62.045 -39.955 -61.715 ;
        RECT -40.285 -63.405 -39.955 -63.075 ;
        RECT -40.285 -64.765 -39.955 -64.435 ;
        RECT -40.285 -66.125 -39.955 -65.795 ;
        RECT -40.285 -67.485 -39.955 -67.155 ;
        RECT -40.285 -68.845 -39.955 -68.515 ;
        RECT -40.285 -70.37 -39.955 -70.04 ;
        RECT -40.285 -71.565 -39.955 -71.235 ;
        RECT -40.285 -72.925 -39.955 -72.595 ;
        RECT -40.285 -74.285 -39.955 -73.955 ;
        RECT -40.285 -75.645 -39.955 -75.315 ;
        RECT -40.285 -77.005 -39.955 -76.675 ;
        RECT -40.285 -79.725 -39.955 -79.395 ;
        RECT -40.285 -80.91 -39.955 -80.58 ;
        RECT -40.285 -82.445 -39.955 -82.115 ;
        RECT -40.285 -83.805 -39.955 -83.475 ;
        RECT -40.285 -85.165 -39.955 -84.835 ;
        RECT -40.285 -87.885 -39.955 -87.555 ;
        RECT -40.285 -89.245 -39.955 -88.915 ;
        RECT -40.285 -93.325 -39.955 -92.995 ;
        RECT -40.285 -94.685 -39.955 -94.355 ;
        RECT -40.285 -96.045 -39.955 -95.715 ;
        RECT -40.285 -98.765 -39.955 -98.435 ;
        RECT -40.285 -100.125 -39.955 -99.795 ;
        RECT -40.285 -101.485 -39.955 -101.155 ;
        RECT -40.285 -102.845 -39.955 -102.515 ;
        RECT -40.285 -104.205 -39.955 -103.875 ;
        RECT -40.285 -105.565 -39.955 -105.235 ;
        RECT -40.285 -106.925 -39.955 -106.595 ;
        RECT -40.285 -108.285 -39.955 -107.955 ;
        RECT -40.285 -109.645 -39.955 -109.315 ;
        RECT -40.285 -111.005 -39.955 -110.675 ;
        RECT -40.285 -112.365 -39.955 -112.035 ;
        RECT -40.285 -113.725 -39.955 -113.395 ;
        RECT -40.285 -115.085 -39.955 -114.755 ;
        RECT -40.285 -116.445 -39.955 -116.115 ;
        RECT -40.285 -117.805 -39.955 -117.475 ;
        RECT -40.285 -119.165 -39.955 -118.835 ;
        RECT -40.285 -120.525 -39.955 -120.195 ;
        RECT -40.285 -121.885 -39.955 -121.555 ;
        RECT -40.285 -123.245 -39.955 -122.915 ;
        RECT -40.285 -124.605 -39.955 -124.275 ;
        RECT -40.285 -125.965 -39.955 -125.635 ;
        RECT -40.285 -127.325 -39.955 -126.995 ;
        RECT -40.285 -130.045 -39.955 -129.715 ;
        RECT -40.285 -131.405 -39.955 -131.075 ;
        RECT -40.285 -132.765 -39.955 -132.435 ;
        RECT -40.285 -134.125 -39.955 -133.795 ;
        RECT -40.285 -136.845 -39.955 -136.515 ;
        RECT -40.285 -138.205 -39.955 -137.875 ;
        RECT -40.285 -139.565 -39.955 -139.235 ;
        RECT -40.285 -140.925 -39.955 -140.595 ;
        RECT -40.285 -142.285 -39.955 -141.955 ;
        RECT -40.285 -143.645 -39.955 -143.315 ;
        RECT -40.285 -145.005 -39.955 -144.675 ;
        RECT -40.285 -146.365 -39.955 -146.035 ;
        RECT -40.285 -148.215 -39.955 -147.885 ;
        RECT -40.285 -149.085 -39.955 -148.755 ;
        RECT -40.285 -150.445 -39.955 -150.115 ;
        RECT -40.285 -151.805 -39.955 -151.475 ;
        RECT -40.285 -154.525 -39.955 -154.195 ;
        RECT -40.285 -157.245 -39.955 -156.915 ;
        RECT -40.285 -162.89 -39.955 -161.76 ;
        RECT -40.28 -163.005 -39.96 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 129.945 -38.595 131.075 ;
        RECT -38.925 125.635 -38.595 125.965 ;
        RECT -38.925 124.275 -38.595 124.605 ;
        RECT -38.925 122.915 -38.595 123.245 ;
        RECT -38.925 121.555 -38.595 121.885 ;
        RECT -38.925 120.195 -38.595 120.525 ;
        RECT -38.925 118.835 -38.595 119.165 ;
        RECT -38.925 117.475 -38.595 117.805 ;
        RECT -38.925 116.115 -38.595 116.445 ;
        RECT -38.925 114.755 -38.595 115.085 ;
        RECT -38.925 113.395 -38.595 113.725 ;
        RECT -38.925 112.035 -38.595 112.365 ;
        RECT -38.925 110.675 -38.595 111.005 ;
        RECT -38.925 109.315 -38.595 109.645 ;
        RECT -38.925 107.955 -38.595 108.285 ;
        RECT -38.925 106.595 -38.595 106.925 ;
        RECT -38.925 105.235 -38.595 105.565 ;
        RECT -38.925 103.875 -38.595 104.205 ;
        RECT -38.925 102.515 -38.595 102.845 ;
        RECT -38.925 101.155 -38.595 101.485 ;
        RECT -38.925 99.795 -38.595 100.125 ;
        RECT -38.925 98.435 -38.595 98.765 ;
        RECT -38.925 97.075 -38.595 97.405 ;
        RECT -38.925 95.715 -38.595 96.045 ;
        RECT -38.925 94.355 -38.595 94.685 ;
        RECT -38.925 92.995 -38.595 93.325 ;
        RECT -38.925 91.635 -38.595 91.965 ;
        RECT -38.925 90.275 -38.595 90.605 ;
        RECT -38.925 88.915 -38.595 89.245 ;
        RECT -38.925 87.555 -38.595 87.885 ;
        RECT -38.925 86.195 -38.595 86.525 ;
        RECT -38.925 84.835 -38.595 85.165 ;
        RECT -38.925 83.475 -38.595 83.805 ;
        RECT -38.925 82.115 -38.595 82.445 ;
        RECT -38.925 80.755 -38.595 81.085 ;
        RECT -38.925 79.395 -38.595 79.725 ;
        RECT -38.925 78.035 -38.595 78.365 ;
        RECT -38.925 76.675 -38.595 77.005 ;
        RECT -38.925 75.315 -38.595 75.645 ;
        RECT -38.925 73.955 -38.595 74.285 ;
        RECT -38.925 72.595 -38.595 72.925 ;
        RECT -38.925 71.235 -38.595 71.565 ;
        RECT -38.925 69.875 -38.595 70.205 ;
        RECT -38.925 68.515 -38.595 68.845 ;
        RECT -38.925 67.155 -38.595 67.485 ;
        RECT -38.925 65.795 -38.595 66.125 ;
        RECT -38.925 64.435 -38.595 64.765 ;
        RECT -38.925 63.075 -38.595 63.405 ;
        RECT -38.925 61.715 -38.595 62.045 ;
        RECT -38.925 60.355 -38.595 60.685 ;
        RECT -38.925 58.995 -38.595 59.325 ;
        RECT -38.925 57.635 -38.595 57.965 ;
        RECT -38.925 56.275 -38.595 56.605 ;
        RECT -38.925 54.915 -38.595 55.245 ;
        RECT -38.925 53.555 -38.595 53.885 ;
        RECT -38.925 52.195 -38.595 52.525 ;
        RECT -38.925 50.835 -38.595 51.165 ;
        RECT -38.925 49.475 -38.595 49.805 ;
        RECT -38.925 48.115 -38.595 48.445 ;
        RECT -38.925 46.755 -38.595 47.085 ;
        RECT -38.925 45.395 -38.595 45.725 ;
        RECT -38.925 44.035 -38.595 44.365 ;
        RECT -38.925 42.675 -38.595 43.005 ;
        RECT -38.925 41.315 -38.595 41.645 ;
        RECT -38.925 39.955 -38.595 40.285 ;
        RECT -38.925 38.595 -38.595 38.925 ;
        RECT -38.925 37.235 -38.595 37.565 ;
        RECT -38.925 35.875 -38.595 36.205 ;
        RECT -38.925 34.515 -38.595 34.845 ;
        RECT -38.925 33.155 -38.595 33.485 ;
        RECT -38.925 31.795 -38.595 32.125 ;
        RECT -38.925 30.435 -38.595 30.765 ;
        RECT -38.925 29.075 -38.595 29.405 ;
        RECT -38.925 27.715 -38.595 28.045 ;
        RECT -38.925 26.355 -38.595 26.685 ;
        RECT -38.925 24.995 -38.595 25.325 ;
        RECT -38.925 23.635 -38.595 23.965 ;
        RECT -38.925 22.275 -38.595 22.605 ;
        RECT -38.925 20.915 -38.595 21.245 ;
        RECT -38.925 19.555 -38.595 19.885 ;
        RECT -38.925 18.195 -38.595 18.525 ;
        RECT -38.925 16.835 -38.595 17.165 ;
        RECT -38.925 15.475 -38.595 15.805 ;
        RECT -38.925 14.115 -38.595 14.445 ;
        RECT -38.925 12.755 -38.595 13.085 ;
        RECT -38.925 11.395 -38.595 11.725 ;
        RECT -38.925 10.035 -38.595 10.365 ;
        RECT -38.925 8.675 -38.595 9.005 ;
        RECT -38.925 7.315 -38.595 7.645 ;
        RECT -38.925 5.955 -38.595 6.285 ;
        RECT -38.925 4.595 -38.595 4.925 ;
        RECT -38.925 3.235 -38.595 3.565 ;
        RECT -38.925 1.875 -38.595 2.205 ;
        RECT -38.925 0.515 -38.595 0.845 ;
        RECT -38.925 -0.845 -38.595 -0.515 ;
        RECT -38.925 -2.205 -38.595 -1.875 ;
        RECT -38.925 -7.645 -38.595 -7.315 ;
        RECT -38.925 -11.725 -38.595 -11.395 ;
        RECT -38.925 -13.085 -38.595 -12.755 ;
        RECT -38.925 -14.445 -38.595 -14.115 ;
        RECT -38.925 -15.805 -38.595 -15.475 ;
        RECT -38.925 -17.165 -38.595 -16.835 ;
        RECT -38.925 -19.885 -38.595 -19.555 ;
        RECT -38.925 -21.245 -38.595 -20.915 ;
        RECT -38.925 -22.605 -38.595 -22.275 ;
        RECT -38.925 -29.405 -38.595 -29.075 ;
        RECT -38.925 -30.765 -38.595 -30.435 ;
        RECT -38.925 -32.125 -38.595 -31.795 ;
        RECT -38.925 -33.485 -38.595 -33.155 ;
        RECT -38.925 -34.845 -38.595 -34.515 ;
        RECT -38.925 -36.205 -38.595 -35.875 ;
        RECT -38.925 -37.565 -38.595 -37.235 ;
        RECT -38.925 -38.925 -38.595 -38.595 ;
        RECT -38.925 -40.285 -38.595 -39.955 ;
        RECT -38.925 -41.645 -38.595 -41.315 ;
        RECT -38.925 -43.005 -38.595 -42.675 ;
        RECT -38.925 -44.365 -38.595 -44.035 ;
        RECT -38.925 -45.725 -38.595 -45.395 ;
        RECT -38.925 -48.445 -38.595 -48.115 ;
        RECT -38.925 -49.805 -38.595 -49.475 ;
        RECT -38.925 -51.165 -38.595 -50.835 ;
        RECT -38.925 -52.525 -38.595 -52.195 ;
        RECT -38.925 -53.885 -38.595 -53.555 ;
        RECT -38.925 -55.245 -38.595 -54.915 ;
        RECT -38.925 -56.605 -38.595 -56.275 ;
        RECT -38.925 -57.965 -38.595 -57.635 ;
        RECT -38.925 -59.325 -38.595 -58.995 ;
        RECT -38.925 -60.685 -38.595 -60.355 ;
        RECT -38.925 -62.045 -38.595 -61.715 ;
        RECT -38.925 -63.405 -38.595 -63.075 ;
        RECT -38.925 -64.765 -38.595 -64.435 ;
        RECT -38.925 -66.125 -38.595 -65.795 ;
        RECT -38.925 -67.485 -38.595 -67.155 ;
        RECT -38.925 -68.845 -38.595 -68.515 ;
        RECT -38.925 -70.37 -38.595 -70.04 ;
        RECT -38.925 -71.565 -38.595 -71.235 ;
        RECT -38.925 -72.925 -38.595 -72.595 ;
        RECT -38.925 -74.285 -38.595 -73.955 ;
        RECT -38.925 -75.645 -38.595 -75.315 ;
        RECT -38.925 -77.005 -38.595 -76.675 ;
        RECT -38.925 -79.725 -38.595 -79.395 ;
        RECT -38.925 -80.91 -38.595 -80.58 ;
        RECT -38.925 -82.445 -38.595 -82.115 ;
        RECT -38.925 -83.805 -38.595 -83.475 ;
        RECT -38.925 -85.165 -38.595 -84.835 ;
        RECT -38.925 -87.885 -38.595 -87.555 ;
        RECT -38.925 -89.245 -38.595 -88.915 ;
        RECT -38.92 -91.28 -38.6 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 -154.525 -38.595 -154.195 ;
        RECT -38.925 -157.245 -38.595 -156.915 ;
        RECT -38.925 -162.89 -38.595 -161.76 ;
        RECT -38.92 -163.005 -38.6 -153.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.565 129.945 -37.235 131.075 ;
        RECT -37.565 125.635 -37.235 125.965 ;
        RECT -37.565 124.275 -37.235 124.605 ;
        RECT -37.565 122.915 -37.235 123.245 ;
        RECT -37.565 121.555 -37.235 121.885 ;
        RECT -37.565 120.195 -37.235 120.525 ;
        RECT -37.565 118.835 -37.235 119.165 ;
        RECT -37.565 117.475 -37.235 117.805 ;
        RECT -37.565 116.115 -37.235 116.445 ;
        RECT -37.565 114.755 -37.235 115.085 ;
        RECT -37.565 113.395 -37.235 113.725 ;
        RECT -37.565 112.035 -37.235 112.365 ;
        RECT -37.565 110.675 -37.235 111.005 ;
        RECT -37.565 109.315 -37.235 109.645 ;
        RECT -37.565 107.955 -37.235 108.285 ;
        RECT -37.565 106.595 -37.235 106.925 ;
        RECT -37.565 105.235 -37.235 105.565 ;
        RECT -37.565 103.875 -37.235 104.205 ;
        RECT -37.565 102.515 -37.235 102.845 ;
        RECT -37.565 101.155 -37.235 101.485 ;
        RECT -37.565 99.795 -37.235 100.125 ;
        RECT -37.565 98.435 -37.235 98.765 ;
        RECT -37.565 97.075 -37.235 97.405 ;
        RECT -37.565 95.715 -37.235 96.045 ;
        RECT -37.565 94.355 -37.235 94.685 ;
        RECT -37.565 92.995 -37.235 93.325 ;
        RECT -37.565 91.635 -37.235 91.965 ;
        RECT -37.565 90.275 -37.235 90.605 ;
        RECT -37.565 88.915 -37.235 89.245 ;
        RECT -37.565 87.555 -37.235 87.885 ;
        RECT -37.565 86.195 -37.235 86.525 ;
        RECT -37.565 84.835 -37.235 85.165 ;
        RECT -37.565 83.475 -37.235 83.805 ;
        RECT -37.565 82.115 -37.235 82.445 ;
        RECT -37.565 80.755 -37.235 81.085 ;
        RECT -37.565 79.395 -37.235 79.725 ;
        RECT -37.565 78.035 -37.235 78.365 ;
        RECT -37.565 76.675 -37.235 77.005 ;
        RECT -37.565 75.315 -37.235 75.645 ;
        RECT -37.565 73.955 -37.235 74.285 ;
        RECT -37.565 72.595 -37.235 72.925 ;
        RECT -37.565 71.235 -37.235 71.565 ;
        RECT -37.565 69.875 -37.235 70.205 ;
        RECT -37.565 68.515 -37.235 68.845 ;
        RECT -37.565 67.155 -37.235 67.485 ;
        RECT -37.565 65.795 -37.235 66.125 ;
        RECT -37.565 64.435 -37.235 64.765 ;
        RECT -37.565 63.075 -37.235 63.405 ;
        RECT -37.565 61.715 -37.235 62.045 ;
        RECT -37.565 60.355 -37.235 60.685 ;
        RECT -37.565 58.995 -37.235 59.325 ;
        RECT -37.565 57.635 -37.235 57.965 ;
        RECT -37.565 56.275 -37.235 56.605 ;
        RECT -37.565 54.915 -37.235 55.245 ;
        RECT -37.565 53.555 -37.235 53.885 ;
        RECT -37.565 52.195 -37.235 52.525 ;
        RECT -37.565 50.835 -37.235 51.165 ;
        RECT -37.565 49.475 -37.235 49.805 ;
        RECT -37.565 48.115 -37.235 48.445 ;
        RECT -37.565 46.755 -37.235 47.085 ;
        RECT -37.565 45.395 -37.235 45.725 ;
        RECT -37.565 44.035 -37.235 44.365 ;
        RECT -37.565 42.675 -37.235 43.005 ;
        RECT -37.565 41.315 -37.235 41.645 ;
        RECT -37.565 39.955 -37.235 40.285 ;
        RECT -37.565 38.595 -37.235 38.925 ;
        RECT -37.565 37.235 -37.235 37.565 ;
        RECT -37.565 35.875 -37.235 36.205 ;
        RECT -37.565 34.515 -37.235 34.845 ;
        RECT -37.565 33.155 -37.235 33.485 ;
        RECT -37.565 31.795 -37.235 32.125 ;
        RECT -37.565 30.435 -37.235 30.765 ;
        RECT -37.565 29.075 -37.235 29.405 ;
        RECT -37.565 27.715 -37.235 28.045 ;
        RECT -37.565 26.355 -37.235 26.685 ;
        RECT -37.565 24.995 -37.235 25.325 ;
        RECT -37.565 23.635 -37.235 23.965 ;
        RECT -37.565 22.275 -37.235 22.605 ;
        RECT -37.565 20.915 -37.235 21.245 ;
        RECT -37.565 19.555 -37.235 19.885 ;
        RECT -37.565 18.195 -37.235 18.525 ;
        RECT -37.565 16.835 -37.235 17.165 ;
        RECT -37.565 15.475 -37.235 15.805 ;
        RECT -37.565 14.115 -37.235 14.445 ;
        RECT -37.565 12.755 -37.235 13.085 ;
        RECT -37.565 11.395 -37.235 11.725 ;
        RECT -37.565 10.035 -37.235 10.365 ;
        RECT -37.565 8.675 -37.235 9.005 ;
        RECT -37.565 7.315 -37.235 7.645 ;
        RECT -37.565 5.955 -37.235 6.285 ;
        RECT -37.565 4.595 -37.235 4.925 ;
        RECT -37.565 3.235 -37.235 3.565 ;
        RECT -37.565 1.875 -37.235 2.205 ;
        RECT -37.565 0.515 -37.235 0.845 ;
        RECT -37.565 -0.845 -37.235 -0.515 ;
        RECT -37.565 -7.645 -37.235 -7.315 ;
        RECT -37.565 -11.725 -37.235 -11.395 ;
        RECT -37.565 -13.085 -37.235 -12.755 ;
        RECT -37.565 -14.445 -37.235 -14.115 ;
        RECT -37.565 -15.805 -37.235 -15.475 ;
        RECT -37.565 -17.165 -37.235 -16.835 ;
        RECT -37.565 -19.885 -37.235 -19.555 ;
        RECT -37.565 -21.245 -37.235 -20.915 ;
        RECT -37.565 -22.605 -37.235 -22.275 ;
        RECT -37.565 -29.405 -37.235 -29.075 ;
        RECT -37.565 -30.765 -37.235 -30.435 ;
        RECT -37.565 -32.125 -37.235 -31.795 ;
        RECT -37.565 -33.485 -37.235 -33.155 ;
        RECT -37.565 -34.845 -37.235 -34.515 ;
        RECT -37.565 -36.205 -37.235 -35.875 ;
        RECT -37.565 -37.565 -37.235 -37.235 ;
        RECT -37.565 -38.925 -37.235 -38.595 ;
        RECT -37.565 -40.285 -37.235 -39.955 ;
        RECT -37.565 -41.645 -37.235 -41.315 ;
        RECT -37.565 -43.005 -37.235 -42.675 ;
        RECT -37.565 -44.365 -37.235 -44.035 ;
        RECT -37.565 -45.725 -37.235 -45.395 ;
        RECT -37.565 -48.445 -37.235 -48.115 ;
        RECT -37.565 -49.805 -37.235 -49.475 ;
        RECT -37.565 -51.165 -37.235 -50.835 ;
        RECT -37.565 -52.525 -37.235 -52.195 ;
        RECT -37.565 -53.885 -37.235 -53.555 ;
        RECT -37.565 -55.245 -37.235 -54.915 ;
        RECT -37.565 -56.605 -37.235 -56.275 ;
        RECT -37.565 -57.965 -37.235 -57.635 ;
        RECT -37.565 -59.325 -37.235 -58.995 ;
        RECT -37.565 -60.685 -37.235 -60.355 ;
        RECT -37.565 -62.045 -37.235 -61.715 ;
        RECT -37.565 -63.405 -37.235 -63.075 ;
        RECT -37.565 -64.765 -37.235 -64.435 ;
        RECT -37.565 -66.125 -37.235 -65.795 ;
        RECT -37.565 -67.485 -37.235 -67.155 ;
        RECT -37.565 -68.845 -37.235 -68.515 ;
        RECT -37.565 -70.37 -37.235 -70.04 ;
        RECT -37.565 -71.565 -37.235 -71.235 ;
        RECT -37.565 -72.925 -37.235 -72.595 ;
        RECT -37.565 -74.285 -37.235 -73.955 ;
        RECT -37.565 -75.645 -37.235 -75.315 ;
        RECT -37.565 -77.005 -37.235 -76.675 ;
        RECT -37.565 -79.725 -37.235 -79.395 ;
        RECT -37.565 -80.91 -37.235 -80.58 ;
        RECT -37.565 -82.445 -37.235 -82.115 ;
        RECT -37.565 -83.805 -37.235 -83.475 ;
        RECT -37.565 -85.165 -37.235 -84.835 ;
        RECT -37.565 -87.885 -37.235 -87.555 ;
        RECT -37.565 -89.245 -37.235 -88.915 ;
        RECT -37.565 -91.965 -37.235 -91.635 ;
        RECT -37.565 -93.325 -37.235 -92.995 ;
        RECT -37.565 -94.685 -37.235 -94.355 ;
        RECT -37.565 -96.045 -37.235 -95.715 ;
        RECT -37.565 -98.765 -37.235 -98.435 ;
        RECT -37.565 -100.125 -37.235 -99.795 ;
        RECT -37.565 -101.485 -37.235 -101.155 ;
        RECT -37.565 -102.845 -37.235 -102.515 ;
        RECT -37.565 -104.205 -37.235 -103.875 ;
        RECT -37.565 -105.565 -37.235 -105.235 ;
        RECT -37.565 -106.925 -37.235 -106.595 ;
        RECT -37.565 -108.285 -37.235 -107.955 ;
        RECT -37.565 -112.365 -37.235 -112.035 ;
        RECT -37.565 -113.725 -37.235 -113.395 ;
        RECT -37.565 -115.085 -37.235 -114.755 ;
        RECT -37.565 -116.445 -37.235 -116.115 ;
        RECT -37.565 -117.805 -37.235 -117.475 ;
        RECT -37.565 -119.165 -37.235 -118.835 ;
        RECT -37.565 -120.525 -37.235 -120.195 ;
        RECT -37.565 -121.885 -37.235 -121.555 ;
        RECT -37.565 -123.245 -37.235 -122.915 ;
        RECT -37.565 -124.605 -37.235 -124.275 ;
        RECT -37.565 -125.965 -37.235 -125.635 ;
        RECT -37.565 -127.325 -37.235 -126.995 ;
        RECT -37.565 -130.045 -37.235 -129.715 ;
        RECT -37.565 -131.405 -37.235 -131.075 ;
        RECT -37.565 -135.485 -37.235 -135.155 ;
        RECT -37.565 -136.845 -37.235 -136.515 ;
        RECT -37.565 -138.205 -37.235 -137.875 ;
        RECT -37.565 -139.565 -37.235 -139.235 ;
        RECT -37.565 -140.925 -37.235 -140.595 ;
        RECT -37.565 -142.285 -37.235 -141.955 ;
        RECT -37.565 -143.645 -37.235 -143.315 ;
        RECT -37.565 -145.005 -37.235 -144.675 ;
        RECT -37.565 -146.365 -37.235 -146.035 ;
        RECT -37.565 -148.215 -37.235 -147.885 ;
        RECT -37.565 -149.085 -37.235 -148.755 ;
        RECT -37.565 -150.445 -37.235 -150.115 ;
        RECT -37.565 -151.805 -37.235 -151.475 ;
        RECT -37.565 -153.165 -37.235 -152.835 ;
        RECT -37.565 -154.525 -37.235 -154.195 ;
        RECT -37.565 -157.245 -37.235 -156.915 ;
        RECT -37.565 -162.89 -37.235 -161.76 ;
        RECT -37.56 -163.005 -37.24 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.205 129.945 -35.875 131.075 ;
        RECT -36.205 125.635 -35.875 125.965 ;
        RECT -36.205 124.275 -35.875 124.605 ;
        RECT -36.205 122.915 -35.875 123.245 ;
        RECT -36.205 121.555 -35.875 121.885 ;
        RECT -36.205 120.195 -35.875 120.525 ;
        RECT -36.205 118.835 -35.875 119.165 ;
        RECT -36.205 117.475 -35.875 117.805 ;
        RECT -36.205 116.115 -35.875 116.445 ;
        RECT -36.205 114.755 -35.875 115.085 ;
        RECT -36.205 113.395 -35.875 113.725 ;
        RECT -36.205 112.035 -35.875 112.365 ;
        RECT -36.205 110.675 -35.875 111.005 ;
        RECT -36.205 109.315 -35.875 109.645 ;
        RECT -36.205 107.955 -35.875 108.285 ;
        RECT -36.205 106.595 -35.875 106.925 ;
        RECT -36.205 105.235 -35.875 105.565 ;
        RECT -36.205 103.875 -35.875 104.205 ;
        RECT -36.205 102.515 -35.875 102.845 ;
        RECT -36.205 101.155 -35.875 101.485 ;
        RECT -36.205 99.795 -35.875 100.125 ;
        RECT -36.205 98.435 -35.875 98.765 ;
        RECT -36.205 97.075 -35.875 97.405 ;
        RECT -36.205 95.715 -35.875 96.045 ;
        RECT -36.205 94.355 -35.875 94.685 ;
        RECT -36.205 92.995 -35.875 93.325 ;
        RECT -36.205 91.635 -35.875 91.965 ;
        RECT -36.205 90.275 -35.875 90.605 ;
        RECT -36.205 88.915 -35.875 89.245 ;
        RECT -36.205 87.555 -35.875 87.885 ;
        RECT -36.205 86.195 -35.875 86.525 ;
        RECT -36.205 84.835 -35.875 85.165 ;
        RECT -36.205 83.475 -35.875 83.805 ;
        RECT -36.205 82.115 -35.875 82.445 ;
        RECT -36.205 80.755 -35.875 81.085 ;
        RECT -36.205 79.395 -35.875 79.725 ;
        RECT -36.205 78.035 -35.875 78.365 ;
        RECT -36.205 76.675 -35.875 77.005 ;
        RECT -36.205 75.315 -35.875 75.645 ;
        RECT -36.205 73.955 -35.875 74.285 ;
        RECT -36.205 72.595 -35.875 72.925 ;
        RECT -36.205 71.235 -35.875 71.565 ;
        RECT -36.205 69.875 -35.875 70.205 ;
        RECT -36.205 68.515 -35.875 68.845 ;
        RECT -36.205 67.155 -35.875 67.485 ;
        RECT -36.205 65.795 -35.875 66.125 ;
        RECT -36.205 64.435 -35.875 64.765 ;
        RECT -36.205 63.075 -35.875 63.405 ;
        RECT -36.205 61.715 -35.875 62.045 ;
        RECT -36.205 60.355 -35.875 60.685 ;
        RECT -36.205 58.995 -35.875 59.325 ;
        RECT -36.205 57.635 -35.875 57.965 ;
        RECT -36.205 56.275 -35.875 56.605 ;
        RECT -36.205 54.915 -35.875 55.245 ;
        RECT -36.205 53.555 -35.875 53.885 ;
        RECT -36.205 52.195 -35.875 52.525 ;
        RECT -36.205 50.835 -35.875 51.165 ;
        RECT -36.205 49.475 -35.875 49.805 ;
        RECT -36.205 48.115 -35.875 48.445 ;
        RECT -36.205 46.755 -35.875 47.085 ;
        RECT -36.205 45.395 -35.875 45.725 ;
        RECT -36.205 44.035 -35.875 44.365 ;
        RECT -36.205 42.675 -35.875 43.005 ;
        RECT -36.205 41.315 -35.875 41.645 ;
        RECT -36.205 39.955 -35.875 40.285 ;
        RECT -36.205 38.595 -35.875 38.925 ;
        RECT -36.205 37.235 -35.875 37.565 ;
        RECT -36.205 35.875 -35.875 36.205 ;
        RECT -36.205 34.515 -35.875 34.845 ;
        RECT -36.205 33.155 -35.875 33.485 ;
        RECT -36.205 31.795 -35.875 32.125 ;
        RECT -36.205 30.435 -35.875 30.765 ;
        RECT -36.205 29.075 -35.875 29.405 ;
        RECT -36.205 27.715 -35.875 28.045 ;
        RECT -36.205 26.355 -35.875 26.685 ;
        RECT -36.205 24.995 -35.875 25.325 ;
        RECT -36.205 23.635 -35.875 23.965 ;
        RECT -36.205 22.275 -35.875 22.605 ;
        RECT -36.205 20.915 -35.875 21.245 ;
        RECT -36.205 19.555 -35.875 19.885 ;
        RECT -36.205 18.195 -35.875 18.525 ;
        RECT -36.205 16.835 -35.875 17.165 ;
        RECT -36.205 15.475 -35.875 15.805 ;
        RECT -36.205 14.115 -35.875 14.445 ;
        RECT -36.205 12.755 -35.875 13.085 ;
        RECT -36.205 11.395 -35.875 11.725 ;
        RECT -36.205 10.035 -35.875 10.365 ;
        RECT -36.205 8.675 -35.875 9.005 ;
        RECT -36.205 7.315 -35.875 7.645 ;
        RECT -36.205 5.955 -35.875 6.285 ;
        RECT -36.205 4.595 -35.875 4.925 ;
        RECT -36.205 3.235 -35.875 3.565 ;
        RECT -36.205 1.875 -35.875 2.205 ;
        RECT -36.205 0.515 -35.875 0.845 ;
        RECT -36.205 -7.645 -35.875 -7.315 ;
        RECT -36.205 -11.725 -35.875 -11.395 ;
        RECT -36.205 -13.085 -35.875 -12.755 ;
        RECT -36.205 -14.445 -35.875 -14.115 ;
        RECT -36.205 -15.805 -35.875 -15.475 ;
        RECT -36.205 -17.165 -35.875 -16.835 ;
        RECT -36.205 -19.885 -35.875 -19.555 ;
        RECT -36.205 -21.245 -35.875 -20.915 ;
        RECT -36.205 -22.605 -35.875 -22.275 ;
        RECT -36.205 -29.405 -35.875 -29.075 ;
        RECT -36.205 -30.765 -35.875 -30.435 ;
        RECT -36.205 -32.125 -35.875 -31.795 ;
        RECT -36.205 -33.485 -35.875 -33.155 ;
        RECT -36.205 -34.845 -35.875 -34.515 ;
        RECT -36.205 -36.205 -35.875 -35.875 ;
        RECT -36.205 -37.565 -35.875 -37.235 ;
        RECT -36.205 -38.925 -35.875 -38.595 ;
        RECT -36.205 -40.285 -35.875 -39.955 ;
        RECT -36.205 -41.645 -35.875 -41.315 ;
        RECT -36.205 -43.005 -35.875 -42.675 ;
        RECT -36.205 -44.365 -35.875 -44.035 ;
        RECT -36.205 -45.725 -35.875 -45.395 ;
        RECT -36.205 -48.445 -35.875 -48.115 ;
        RECT -36.205 -49.805 -35.875 -49.475 ;
        RECT -36.205 -51.165 -35.875 -50.835 ;
        RECT -36.205 -52.525 -35.875 -52.195 ;
        RECT -36.205 -53.885 -35.875 -53.555 ;
        RECT -36.205 -55.245 -35.875 -54.915 ;
        RECT -36.205 -56.605 -35.875 -56.275 ;
        RECT -36.205 -57.965 -35.875 -57.635 ;
        RECT -36.205 -59.325 -35.875 -58.995 ;
        RECT -36.205 -60.685 -35.875 -60.355 ;
        RECT -36.205 -62.045 -35.875 -61.715 ;
        RECT -36.205 -63.405 -35.875 -63.075 ;
        RECT -36.205 -64.765 -35.875 -64.435 ;
        RECT -36.205 -66.125 -35.875 -65.795 ;
        RECT -36.205 -67.485 -35.875 -67.155 ;
        RECT -36.205 -68.845 -35.875 -68.515 ;
        RECT -36.205 -70.37 -35.875 -70.04 ;
        RECT -36.205 -71.565 -35.875 -71.235 ;
        RECT -36.205 -72.925 -35.875 -72.595 ;
        RECT -36.205 -74.285 -35.875 -73.955 ;
        RECT -36.205 -75.645 -35.875 -75.315 ;
        RECT -36.205 -77.005 -35.875 -76.675 ;
        RECT -36.205 -79.725 -35.875 -79.395 ;
        RECT -36.205 -80.91 -35.875 -80.58 ;
        RECT -36.205 -82.445 -35.875 -82.115 ;
        RECT -36.205 -83.805 -35.875 -83.475 ;
        RECT -36.205 -85.165 -35.875 -84.835 ;
        RECT -36.205 -87.885 -35.875 -87.555 ;
        RECT -36.205 -89.245 -35.875 -88.915 ;
        RECT -36.205 -91.965 -35.875 -91.635 ;
        RECT -36.205 -93.325 -35.875 -92.995 ;
        RECT -36.205 -94.685 -35.875 -94.355 ;
        RECT -36.205 -96.045 -35.875 -95.715 ;
        RECT -36.205 -98.765 -35.875 -98.435 ;
        RECT -36.205 -100.125 -35.875 -99.795 ;
        RECT -36.205 -101.485 -35.875 -101.155 ;
        RECT -36.205 -102.845 -35.875 -102.515 ;
        RECT -36.205 -104.205 -35.875 -103.875 ;
        RECT -36.205 -105.565 -35.875 -105.235 ;
        RECT -36.205 -106.925 -35.875 -106.595 ;
        RECT -36.205 -108.285 -35.875 -107.955 ;
        RECT -36.205 -112.365 -35.875 -112.035 ;
        RECT -36.205 -113.725 -35.875 -113.395 ;
        RECT -36.205 -115.085 -35.875 -114.755 ;
        RECT -36.205 -116.445 -35.875 -116.115 ;
        RECT -36.205 -117.805 -35.875 -117.475 ;
        RECT -36.205 -119.165 -35.875 -118.835 ;
        RECT -36.205 -120.525 -35.875 -120.195 ;
        RECT -36.205 -121.885 -35.875 -121.555 ;
        RECT -36.205 -123.245 -35.875 -122.915 ;
        RECT -36.205 -124.605 -35.875 -124.275 ;
        RECT -36.205 -125.965 -35.875 -125.635 ;
        RECT -36.205 -127.325 -35.875 -126.995 ;
        RECT -36.205 -130.045 -35.875 -129.715 ;
        RECT -36.205 -131.405 -35.875 -131.075 ;
        RECT -36.205 -135.485 -35.875 -135.155 ;
        RECT -36.205 -136.845 -35.875 -136.515 ;
        RECT -36.205 -138.205 -35.875 -137.875 ;
        RECT -36.205 -139.565 -35.875 -139.235 ;
        RECT -36.205 -140.925 -35.875 -140.595 ;
        RECT -36.205 -142.285 -35.875 -141.955 ;
        RECT -36.205 -143.645 -35.875 -143.315 ;
        RECT -36.205 -145.005 -35.875 -144.675 ;
        RECT -36.205 -146.365 -35.875 -146.035 ;
        RECT -36.205 -148.215 -35.875 -147.885 ;
        RECT -36.205 -149.085 -35.875 -148.755 ;
        RECT -36.205 -150.445 -35.875 -150.115 ;
        RECT -36.205 -151.805 -35.875 -151.475 ;
        RECT -36.205 -154.525 -35.875 -154.195 ;
        RECT -36.205 -157.245 -35.875 -156.915 ;
        RECT -36.205 -162.89 -35.875 -161.76 ;
        RECT -36.2 -163.005 -35.88 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 -89.245 -34.515 -88.915 ;
        RECT -34.845 -93.325 -34.515 -92.995 ;
        RECT -34.845 -94.685 -34.515 -94.355 ;
        RECT -34.845 -96.045 -34.515 -95.715 ;
        RECT -34.845 -98.765 -34.515 -98.435 ;
        RECT -34.845 -100.125 -34.515 -99.795 ;
        RECT -34.845 -101.485 -34.515 -101.155 ;
        RECT -34.845 -105.565 -34.515 -105.235 ;
        RECT -34.845 -106.925 -34.515 -106.595 ;
        RECT -34.845 -108.285 -34.515 -107.955 ;
        RECT -34.845 -112.365 -34.515 -112.035 ;
        RECT -34.845 -113.725 -34.515 -113.395 ;
        RECT -34.845 -115.085 -34.515 -114.755 ;
        RECT -34.845 -116.445 -34.515 -116.115 ;
        RECT -34.845 -117.805 -34.515 -117.475 ;
        RECT -34.845 -120.525 -34.515 -120.195 ;
        RECT -34.845 -121.885 -34.515 -121.555 ;
        RECT -34.845 -123.245 -34.515 -122.915 ;
        RECT -34.845 -124.605 -34.515 -124.275 ;
        RECT -34.845 -125.965 -34.515 -125.635 ;
        RECT -34.845 -127.325 -34.515 -126.995 ;
        RECT -34.845 -130.045 -34.515 -129.715 ;
        RECT -34.845 -131.405 -34.515 -131.075 ;
        RECT -34.845 -135.485 -34.515 -135.155 ;
        RECT -34.845 -136.845 -34.515 -136.515 ;
        RECT -34.845 -138.205 -34.515 -137.875 ;
        RECT -34.845 -139.565 -34.515 -139.235 ;
        RECT -34.845 -140.925 -34.515 -140.595 ;
        RECT -34.845 -142.285 -34.515 -141.955 ;
        RECT -34.845 -143.645 -34.515 -143.315 ;
        RECT -34.845 -145.005 -34.515 -144.675 ;
        RECT -34.845 -146.365 -34.515 -146.035 ;
        RECT -34.845 -149.085 -34.515 -148.755 ;
        RECT -34.845 -150.445 -34.515 -150.115 ;
        RECT -34.845 -154.525 -34.515 -154.195 ;
        RECT -34.845 -157.245 -34.515 -156.915 ;
        RECT -34.845 -162.89 -34.515 -161.76 ;
        RECT -34.84 -163.005 -34.52 131.19 ;
        RECT -34.845 129.945 -34.515 131.075 ;
        RECT -34.845 125.635 -34.515 125.965 ;
        RECT -34.845 124.275 -34.515 124.605 ;
        RECT -34.845 122.915 -34.515 123.245 ;
        RECT -34.845 121.555 -34.515 121.885 ;
        RECT -34.845 120.195 -34.515 120.525 ;
        RECT -34.845 118.835 -34.515 119.165 ;
        RECT -34.845 117.475 -34.515 117.805 ;
        RECT -34.845 116.115 -34.515 116.445 ;
        RECT -34.845 114.755 -34.515 115.085 ;
        RECT -34.845 113.395 -34.515 113.725 ;
        RECT -34.845 112.035 -34.515 112.365 ;
        RECT -34.845 110.675 -34.515 111.005 ;
        RECT -34.845 109.315 -34.515 109.645 ;
        RECT -34.845 107.955 -34.515 108.285 ;
        RECT -34.845 106.595 -34.515 106.925 ;
        RECT -34.845 105.235 -34.515 105.565 ;
        RECT -34.845 103.875 -34.515 104.205 ;
        RECT -34.845 102.515 -34.515 102.845 ;
        RECT -34.845 101.155 -34.515 101.485 ;
        RECT -34.845 99.795 -34.515 100.125 ;
        RECT -34.845 98.435 -34.515 98.765 ;
        RECT -34.845 97.075 -34.515 97.405 ;
        RECT -34.845 95.715 -34.515 96.045 ;
        RECT -34.845 94.355 -34.515 94.685 ;
        RECT -34.845 92.995 -34.515 93.325 ;
        RECT -34.845 91.635 -34.515 91.965 ;
        RECT -34.845 90.275 -34.515 90.605 ;
        RECT -34.845 88.915 -34.515 89.245 ;
        RECT -34.845 87.555 -34.515 87.885 ;
        RECT -34.845 86.195 -34.515 86.525 ;
        RECT -34.845 84.835 -34.515 85.165 ;
        RECT -34.845 83.475 -34.515 83.805 ;
        RECT -34.845 82.115 -34.515 82.445 ;
        RECT -34.845 80.755 -34.515 81.085 ;
        RECT -34.845 79.395 -34.515 79.725 ;
        RECT -34.845 78.035 -34.515 78.365 ;
        RECT -34.845 76.675 -34.515 77.005 ;
        RECT -34.845 75.315 -34.515 75.645 ;
        RECT -34.845 73.955 -34.515 74.285 ;
        RECT -34.845 72.595 -34.515 72.925 ;
        RECT -34.845 71.235 -34.515 71.565 ;
        RECT -34.845 69.875 -34.515 70.205 ;
        RECT -34.845 68.515 -34.515 68.845 ;
        RECT -34.845 67.155 -34.515 67.485 ;
        RECT -34.845 65.795 -34.515 66.125 ;
        RECT -34.845 64.435 -34.515 64.765 ;
        RECT -34.845 63.075 -34.515 63.405 ;
        RECT -34.845 61.715 -34.515 62.045 ;
        RECT -34.845 60.355 -34.515 60.685 ;
        RECT -34.845 58.995 -34.515 59.325 ;
        RECT -34.845 57.635 -34.515 57.965 ;
        RECT -34.845 56.275 -34.515 56.605 ;
        RECT -34.845 54.915 -34.515 55.245 ;
        RECT -34.845 53.555 -34.515 53.885 ;
        RECT -34.845 52.195 -34.515 52.525 ;
        RECT -34.845 50.835 -34.515 51.165 ;
        RECT -34.845 49.475 -34.515 49.805 ;
        RECT -34.845 48.115 -34.515 48.445 ;
        RECT -34.845 46.755 -34.515 47.085 ;
        RECT -34.845 45.395 -34.515 45.725 ;
        RECT -34.845 44.035 -34.515 44.365 ;
        RECT -34.845 42.675 -34.515 43.005 ;
        RECT -34.845 41.315 -34.515 41.645 ;
        RECT -34.845 39.955 -34.515 40.285 ;
        RECT -34.845 38.595 -34.515 38.925 ;
        RECT -34.845 37.235 -34.515 37.565 ;
        RECT -34.845 35.875 -34.515 36.205 ;
        RECT -34.845 34.515 -34.515 34.845 ;
        RECT -34.845 33.155 -34.515 33.485 ;
        RECT -34.845 31.795 -34.515 32.125 ;
        RECT -34.845 30.435 -34.515 30.765 ;
        RECT -34.845 29.075 -34.515 29.405 ;
        RECT -34.845 27.715 -34.515 28.045 ;
        RECT -34.845 26.355 -34.515 26.685 ;
        RECT -34.845 24.995 -34.515 25.325 ;
        RECT -34.845 23.635 -34.515 23.965 ;
        RECT -34.845 22.275 -34.515 22.605 ;
        RECT -34.845 20.915 -34.515 21.245 ;
        RECT -34.845 19.555 -34.515 19.885 ;
        RECT -34.845 18.195 -34.515 18.525 ;
        RECT -34.845 16.835 -34.515 17.165 ;
        RECT -34.845 15.475 -34.515 15.805 ;
        RECT -34.845 14.115 -34.515 14.445 ;
        RECT -34.845 12.755 -34.515 13.085 ;
        RECT -34.845 11.395 -34.515 11.725 ;
        RECT -34.845 10.035 -34.515 10.365 ;
        RECT -34.845 8.675 -34.515 9.005 ;
        RECT -34.845 7.315 -34.515 7.645 ;
        RECT -34.845 5.955 -34.515 6.285 ;
        RECT -34.845 4.595 -34.515 4.925 ;
        RECT -34.845 3.235 -34.515 3.565 ;
        RECT -34.845 1.875 -34.515 2.205 ;
        RECT -34.845 0.515 -34.515 0.845 ;
        RECT -34.845 -7.645 -34.515 -7.315 ;
        RECT -34.845 -11.725 -34.515 -11.395 ;
        RECT -34.845 -13.085 -34.515 -12.755 ;
        RECT -34.845 -14.445 -34.515 -14.115 ;
        RECT -34.845 -15.805 -34.515 -15.475 ;
        RECT -34.845 -17.165 -34.515 -16.835 ;
        RECT -34.845 -19.885 -34.515 -19.555 ;
        RECT -34.845 -21.245 -34.515 -20.915 ;
        RECT -34.845 -22.605 -34.515 -22.275 ;
        RECT -34.845 -29.405 -34.515 -29.075 ;
        RECT -34.845 -30.765 -34.515 -30.435 ;
        RECT -34.845 -32.125 -34.515 -31.795 ;
        RECT -34.845 -33.485 -34.515 -33.155 ;
        RECT -34.845 -34.845 -34.515 -34.515 ;
        RECT -34.845 -36.205 -34.515 -35.875 ;
        RECT -34.845 -37.565 -34.515 -37.235 ;
        RECT -34.845 -38.925 -34.515 -38.595 ;
        RECT -34.845 -40.285 -34.515 -39.955 ;
        RECT -34.845 -41.645 -34.515 -41.315 ;
        RECT -34.845 -43.005 -34.515 -42.675 ;
        RECT -34.845 -44.365 -34.515 -44.035 ;
        RECT -34.845 -45.725 -34.515 -45.395 ;
        RECT -34.845 -48.445 -34.515 -48.115 ;
        RECT -34.845 -49.805 -34.515 -49.475 ;
        RECT -34.845 -51.165 -34.515 -50.835 ;
        RECT -34.845 -52.525 -34.515 -52.195 ;
        RECT -34.845 -53.885 -34.515 -53.555 ;
        RECT -34.845 -55.245 -34.515 -54.915 ;
        RECT -34.845 -56.605 -34.515 -56.275 ;
        RECT -34.845 -57.965 -34.515 -57.635 ;
        RECT -34.845 -59.325 -34.515 -58.995 ;
        RECT -34.845 -60.685 -34.515 -60.355 ;
        RECT -34.845 -62.045 -34.515 -61.715 ;
        RECT -34.845 -63.405 -34.515 -63.075 ;
        RECT -34.845 -64.765 -34.515 -64.435 ;
        RECT -34.845 -66.125 -34.515 -65.795 ;
        RECT -34.845 -67.485 -34.515 -67.155 ;
        RECT -34.845 -68.845 -34.515 -68.515 ;
        RECT -34.845 -70.37 -34.515 -70.04 ;
        RECT -34.845 -71.565 -34.515 -71.235 ;
        RECT -34.845 -72.925 -34.515 -72.595 ;
        RECT -34.845 -74.285 -34.515 -73.955 ;
        RECT -34.845 -75.645 -34.515 -75.315 ;
        RECT -34.845 -77.005 -34.515 -76.675 ;
        RECT -34.845 -79.725 -34.515 -79.395 ;
        RECT -34.845 -80.91 -34.515 -80.58 ;
        RECT -34.845 -82.445 -34.515 -82.115 ;
        RECT -34.845 -83.805 -34.515 -83.475 ;
        RECT -34.845 -85.165 -34.515 -84.835 ;
        RECT -34.845 -87.885 -34.515 -87.555 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 129.945 -49.475 131.075 ;
        RECT -49.805 125.635 -49.475 125.965 ;
        RECT -49.805 124.275 -49.475 124.605 ;
        RECT -49.805 122.915 -49.475 123.245 ;
        RECT -49.805 121.555 -49.475 121.885 ;
        RECT -49.805 120.195 -49.475 120.525 ;
        RECT -49.805 118.835 -49.475 119.165 ;
        RECT -49.805 117.475 -49.475 117.805 ;
        RECT -49.805 116.115 -49.475 116.445 ;
        RECT -49.805 114.755 -49.475 115.085 ;
        RECT -49.805 113.395 -49.475 113.725 ;
        RECT -49.805 112.035 -49.475 112.365 ;
        RECT -49.805 110.675 -49.475 111.005 ;
        RECT -49.805 109.315 -49.475 109.645 ;
        RECT -49.805 107.955 -49.475 108.285 ;
        RECT -49.805 106.595 -49.475 106.925 ;
        RECT -49.805 105.235 -49.475 105.565 ;
        RECT -49.805 103.875 -49.475 104.205 ;
        RECT -49.805 102.515 -49.475 102.845 ;
        RECT -49.805 101.155 -49.475 101.485 ;
        RECT -49.805 99.795 -49.475 100.125 ;
        RECT -49.805 98.435 -49.475 98.765 ;
        RECT -49.805 97.075 -49.475 97.405 ;
        RECT -49.805 95.715 -49.475 96.045 ;
        RECT -49.805 94.355 -49.475 94.685 ;
        RECT -49.805 92.995 -49.475 93.325 ;
        RECT -49.805 91.635 -49.475 91.965 ;
        RECT -49.805 90.275 -49.475 90.605 ;
        RECT -49.805 88.915 -49.475 89.245 ;
        RECT -49.805 87.555 -49.475 87.885 ;
        RECT -49.805 86.195 -49.475 86.525 ;
        RECT -49.805 84.835 -49.475 85.165 ;
        RECT -49.805 83.475 -49.475 83.805 ;
        RECT -49.805 82.115 -49.475 82.445 ;
        RECT -49.805 80.755 -49.475 81.085 ;
        RECT -49.805 79.395 -49.475 79.725 ;
        RECT -49.805 78.035 -49.475 78.365 ;
        RECT -49.805 76.675 -49.475 77.005 ;
        RECT -49.805 75.315 -49.475 75.645 ;
        RECT -49.805 73.955 -49.475 74.285 ;
        RECT -49.8 73.28 -49.48 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 48.115 -49.475 48.445 ;
        RECT -49.805 46.755 -49.475 47.085 ;
        RECT -49.805 45.395 -49.475 45.725 ;
        RECT -49.805 44.035 -49.475 44.365 ;
        RECT -49.805 39.955 -49.475 40.285 ;
        RECT -49.805 38.595 -49.475 38.925 ;
        RECT -49.805 35.875 -49.475 36.205 ;
        RECT -49.805 34.515 -49.475 34.845 ;
        RECT -49.805 33.155 -49.475 33.485 ;
        RECT -49.805 31.795 -49.475 32.125 ;
        RECT -49.805 30.435 -49.475 30.765 ;
        RECT -49.805 29.075 -49.475 29.405 ;
        RECT -49.805 27.715 -49.475 28.045 ;
        RECT -49.805 26.355 -49.475 26.685 ;
        RECT -49.805 24.995 -49.475 25.325 ;
        RECT -49.805 23.635 -49.475 23.965 ;
        RECT -49.805 22.275 -49.475 22.605 ;
        RECT -49.805 20.915 -49.475 21.245 ;
        RECT -49.805 19.555 -49.475 19.885 ;
        RECT -49.805 18.195 -49.475 18.525 ;
        RECT -49.805 16.835 -49.475 17.165 ;
        RECT -49.805 15.475 -49.475 15.805 ;
        RECT -49.805 14.115 -49.475 14.445 ;
        RECT -49.805 12.755 -49.475 13.085 ;
        RECT -49.805 11.395 -49.475 11.725 ;
        RECT -49.805 10.035 -49.475 10.365 ;
        RECT -49.805 8.675 -49.475 9.005 ;
        RECT -49.805 7.315 -49.475 7.645 ;
        RECT -49.805 5.955 -49.475 6.285 ;
        RECT -49.805 4.595 -49.475 4.925 ;
        RECT -49.805 3.235 -49.475 3.565 ;
        RECT -49.805 1.875 -49.475 2.205 ;
        RECT -49.805 0.515 -49.475 0.845 ;
        RECT -49.805 -0.845 -49.475 -0.515 ;
        RECT -49.805 -2.205 -49.475 -1.875 ;
        RECT -49.805 -3.565 -49.475 -3.235 ;
        RECT -49.805 -4.925 -49.475 -4.595 ;
        RECT -49.805 -6.285 -49.475 -5.955 ;
        RECT -49.805 -7.645 -49.475 -7.315 ;
        RECT -49.805 -9.005 -49.475 -8.675 ;
        RECT -49.805 -10.365 -49.475 -10.035 ;
        RECT -49.805 -11.725 -49.475 -11.395 ;
        RECT -49.805 -13.085 -49.475 -12.755 ;
        RECT -49.805 -14.445 -49.475 -14.115 ;
        RECT -49.805 -15.805 -49.475 -15.475 ;
        RECT -49.805 -17.165 -49.475 -16.835 ;
        RECT -49.805 -18.525 -49.475 -18.195 ;
        RECT -49.805 -19.885 -49.475 -19.555 ;
        RECT -49.805 -21.245 -49.475 -20.915 ;
        RECT -49.805 -22.605 -49.475 -22.275 ;
        RECT -49.805 -25.325 -49.475 -24.995 ;
        RECT -49.805 -26.685 -49.475 -26.355 ;
        RECT -49.805 -28.045 -49.475 -27.715 ;
        RECT -49.805 -29.405 -49.475 -29.075 ;
        RECT -49.805 -30.765 -49.475 -30.435 ;
        RECT -49.805 -32.125 -49.475 -31.795 ;
        RECT -49.805 -33.485 -49.475 -33.155 ;
        RECT -49.805 -34.845 -49.475 -34.515 ;
        RECT -49.805 -36.205 -49.475 -35.875 ;
        RECT -49.805 -37.565 -49.475 -37.235 ;
        RECT -49.805 -38.925 -49.475 -38.595 ;
        RECT -49.805 -40.285 -49.475 -39.955 ;
        RECT -49.805 -41.645 -49.475 -41.315 ;
        RECT -49.805 -43.005 -49.475 -42.675 ;
        RECT -49.805 -44.365 -49.475 -44.035 ;
        RECT -49.805 -45.725 -49.475 -45.395 ;
        RECT -49.805 -47.085 -49.475 -46.755 ;
        RECT -49.805 -48.445 -49.475 -48.115 ;
        RECT -49.805 -49.805 -49.475 -49.475 ;
        RECT -49.805 -51.165 -49.475 -50.835 ;
        RECT -49.805 -52.525 -49.475 -52.195 ;
        RECT -49.805 -53.885 -49.475 -53.555 ;
        RECT -49.805 -55.245 -49.475 -54.915 ;
        RECT -49.805 -56.605 -49.475 -56.275 ;
        RECT -49.805 -57.965 -49.475 -57.635 ;
        RECT -49.805 -59.325 -49.475 -58.995 ;
        RECT -49.805 -60.685 -49.475 -60.355 ;
        RECT -49.805 -62.045 -49.475 -61.715 ;
        RECT -49.805 -63.405 -49.475 -63.075 ;
        RECT -49.805 -64.765 -49.475 -64.435 ;
        RECT -49.805 -66.125 -49.475 -65.795 ;
        RECT -49.805 -67.485 -49.475 -67.155 ;
        RECT -49.805 -68.845 -49.475 -68.515 ;
        RECT -49.805 -70.37 -49.475 -70.04 ;
        RECT -49.805 -71.565 -49.475 -71.235 ;
        RECT -49.805 -72.925 -49.475 -72.595 ;
        RECT -49.805 -74.285 -49.475 -73.955 ;
        RECT -49.805 -75.645 -49.475 -75.315 ;
        RECT -49.805 -77.005 -49.475 -76.675 ;
        RECT -49.805 -79.725 -49.475 -79.395 ;
        RECT -49.805 -80.91 -49.475 -80.58 ;
        RECT -49.805 -82.445 -49.475 -82.115 ;
        RECT -49.805 -83.805 -49.475 -83.475 ;
        RECT -49.805 -85.165 -49.475 -84.835 ;
        RECT -49.805 -87.885 -49.475 -87.555 ;
        RECT -49.805 -89.245 -49.475 -88.915 ;
        RECT -49.805 -91.965 -49.475 -91.635 ;
        RECT -49.805 -94.685 -49.475 -94.355 ;
        RECT -49.805 -96.045 -49.475 -95.715 ;
        RECT -49.805 -97.405 -49.475 -97.075 ;
        RECT -49.805 -98.765 -49.475 -98.435 ;
        RECT -49.805 -100.125 -49.475 -99.795 ;
        RECT -49.805 -101.485 -49.475 -101.155 ;
        RECT -49.805 -102.845 -49.475 -102.515 ;
        RECT -49.805 -104.205 -49.475 -103.875 ;
        RECT -49.805 -105.565 -49.475 -105.235 ;
        RECT -49.805 -106.925 -49.475 -106.595 ;
        RECT -49.805 -108.285 -49.475 -107.955 ;
        RECT -49.805 -109.645 -49.475 -109.315 ;
        RECT -49.805 -111.005 -49.475 -110.675 ;
        RECT -49.805 -112.365 -49.475 -112.035 ;
        RECT -49.805 -113.725 -49.475 -113.395 ;
        RECT -49.805 -115.085 -49.475 -114.755 ;
        RECT -49.805 -116.445 -49.475 -116.115 ;
        RECT -49.805 -117.805 -49.475 -117.475 ;
        RECT -49.805 -119.165 -49.475 -118.835 ;
        RECT -49.805 -120.525 -49.475 -120.195 ;
        RECT -49.805 -121.885 -49.475 -121.555 ;
        RECT -49.805 -123.245 -49.475 -122.915 ;
        RECT -49.805 -124.605 -49.475 -124.275 ;
        RECT -49.805 -125.965 -49.475 -125.635 ;
        RECT -49.805 -127.325 -49.475 -126.995 ;
        RECT -49.805 -128.685 -49.475 -128.355 ;
        RECT -49.805 -130.045 -49.475 -129.715 ;
        RECT -49.805 -131.405 -49.475 -131.075 ;
        RECT -49.805 -132.765 -49.475 -132.435 ;
        RECT -49.805 -134.125 -49.475 -133.795 ;
        RECT -49.805 -135.485 -49.475 -135.155 ;
        RECT -49.805 -136.845 -49.475 -136.515 ;
        RECT -49.805 -138.205 -49.475 -137.875 ;
        RECT -49.805 -139.565 -49.475 -139.235 ;
        RECT -49.805 -140.925 -49.475 -140.595 ;
        RECT -49.805 -142.285 -49.475 -141.955 ;
        RECT -49.805 -143.645 -49.475 -143.315 ;
        RECT -49.805 -145.005 -49.475 -144.675 ;
        RECT -49.805 -146.365 -49.475 -146.035 ;
        RECT -49.805 -148.215 -49.475 -147.885 ;
        RECT -49.805 -149.085 -49.475 -148.755 ;
        RECT -49.805 -150.445 -49.475 -150.115 ;
        RECT -49.805 -151.805 -49.475 -151.475 ;
        RECT -49.805 -154.525 -49.475 -154.195 ;
        RECT -49.805 -157.245 -49.475 -156.915 ;
        RECT -49.805 -162.89 -49.475 -161.76 ;
        RECT -49.8 -163.005 -49.48 49.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 129.945 -48.115 131.075 ;
        RECT -48.445 125.635 -48.115 125.965 ;
        RECT -48.445 124.275 -48.115 124.605 ;
        RECT -48.445 122.915 -48.115 123.245 ;
        RECT -48.445 121.555 -48.115 121.885 ;
        RECT -48.445 120.195 -48.115 120.525 ;
        RECT -48.445 118.835 -48.115 119.165 ;
        RECT -48.445 117.475 -48.115 117.805 ;
        RECT -48.445 116.115 -48.115 116.445 ;
        RECT -48.445 114.755 -48.115 115.085 ;
        RECT -48.445 113.395 -48.115 113.725 ;
        RECT -48.445 112.035 -48.115 112.365 ;
        RECT -48.445 110.675 -48.115 111.005 ;
        RECT -48.445 109.315 -48.115 109.645 ;
        RECT -48.445 107.955 -48.115 108.285 ;
        RECT -48.445 106.595 -48.115 106.925 ;
        RECT -48.445 105.235 -48.115 105.565 ;
        RECT -48.445 103.875 -48.115 104.205 ;
        RECT -48.445 102.515 -48.115 102.845 ;
        RECT -48.445 101.155 -48.115 101.485 ;
        RECT -48.445 99.795 -48.115 100.125 ;
        RECT -48.445 98.435 -48.115 98.765 ;
        RECT -48.445 97.075 -48.115 97.405 ;
        RECT -48.445 95.715 -48.115 96.045 ;
        RECT -48.445 94.355 -48.115 94.685 ;
        RECT -48.445 92.995 -48.115 93.325 ;
        RECT -48.445 91.635 -48.115 91.965 ;
        RECT -48.445 90.275 -48.115 90.605 ;
        RECT -48.445 88.915 -48.115 89.245 ;
        RECT -48.445 87.555 -48.115 87.885 ;
        RECT -48.445 86.195 -48.115 86.525 ;
        RECT -48.445 84.835 -48.115 85.165 ;
        RECT -48.445 83.475 -48.115 83.805 ;
        RECT -48.445 82.115 -48.115 82.445 ;
        RECT -48.445 80.755 -48.115 81.085 ;
        RECT -48.445 79.395 -48.115 79.725 ;
        RECT -48.445 78.035 -48.115 78.365 ;
        RECT -48.445 76.675 -48.115 77.005 ;
        RECT -48.445 75.315 -48.115 75.645 ;
        RECT -48.445 73.955 -48.115 74.285 ;
        RECT -48.445 71.64 -48.115 71.97 ;
        RECT -48.445 69.465 -48.115 69.795 ;
        RECT -48.445 68.615 -48.115 68.945 ;
        RECT -48.445 66.305 -48.115 66.635 ;
        RECT -48.445 65.455 -48.115 65.785 ;
        RECT -48.445 63.145 -48.115 63.475 ;
        RECT -48.44 62.4 -48.12 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 -98.765 -48.115 -98.435 ;
        RECT -48.445 -100.125 -48.115 -99.795 ;
        RECT -48.445 -101.485 -48.115 -101.155 ;
        RECT -48.445 -102.845 -48.115 -102.515 ;
        RECT -48.445 -104.205 -48.115 -103.875 ;
        RECT -48.445 -105.565 -48.115 -105.235 ;
        RECT -48.445 -106.925 -48.115 -106.595 ;
        RECT -48.445 -108.285 -48.115 -107.955 ;
        RECT -48.445 -109.645 -48.115 -109.315 ;
        RECT -48.445 -111.005 -48.115 -110.675 ;
        RECT -48.445 -112.365 -48.115 -112.035 ;
        RECT -48.445 -113.725 -48.115 -113.395 ;
        RECT -48.445 -115.085 -48.115 -114.755 ;
        RECT -48.445 -116.445 -48.115 -116.115 ;
        RECT -48.445 -117.805 -48.115 -117.475 ;
        RECT -48.445 -119.165 -48.115 -118.835 ;
        RECT -48.445 -120.525 -48.115 -120.195 ;
        RECT -48.445 -121.885 -48.115 -121.555 ;
        RECT -48.445 -123.245 -48.115 -122.915 ;
        RECT -48.445 -124.605 -48.115 -124.275 ;
        RECT -48.445 -125.965 -48.115 -125.635 ;
        RECT -48.445 -127.325 -48.115 -126.995 ;
        RECT -48.445 -128.685 -48.115 -128.355 ;
        RECT -48.445 -130.045 -48.115 -129.715 ;
        RECT -48.445 -131.405 -48.115 -131.075 ;
        RECT -48.445 -132.765 -48.115 -132.435 ;
        RECT -48.445 -134.125 -48.115 -133.795 ;
        RECT -48.445 -135.485 -48.115 -135.155 ;
        RECT -48.445 -136.845 -48.115 -136.515 ;
        RECT -48.445 -138.205 -48.115 -137.875 ;
        RECT -48.445 -139.565 -48.115 -139.235 ;
        RECT -48.445 -140.925 -48.115 -140.595 ;
        RECT -48.445 -142.285 -48.115 -141.955 ;
        RECT -48.445 -143.645 -48.115 -143.315 ;
        RECT -48.445 -145.005 -48.115 -144.675 ;
        RECT -48.445 -146.365 -48.115 -146.035 ;
        RECT -48.445 -148.215 -48.115 -147.885 ;
        RECT -48.445 -149.085 -48.115 -148.755 ;
        RECT -48.445 -150.445 -48.115 -150.115 ;
        RECT -48.445 -151.805 -48.115 -151.475 ;
        RECT -48.445 -154.525 -48.115 -154.195 ;
        RECT -48.445 -157.245 -48.115 -156.915 ;
        RECT -48.445 -162.89 -48.115 -161.76 ;
        RECT -48.44 -163.005 -48.12 -97.76 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 129.945 -46.755 131.075 ;
        RECT -47.085 125.635 -46.755 125.965 ;
        RECT -47.085 124.275 -46.755 124.605 ;
        RECT -47.085 122.915 -46.755 123.245 ;
        RECT -47.085 121.555 -46.755 121.885 ;
        RECT -47.085 120.195 -46.755 120.525 ;
        RECT -47.085 118.835 -46.755 119.165 ;
        RECT -47.085 117.475 -46.755 117.805 ;
        RECT -47.085 116.115 -46.755 116.445 ;
        RECT -47.085 114.755 -46.755 115.085 ;
        RECT -47.085 113.395 -46.755 113.725 ;
        RECT -47.085 112.035 -46.755 112.365 ;
        RECT -47.085 110.675 -46.755 111.005 ;
        RECT -47.085 109.315 -46.755 109.645 ;
        RECT -47.085 107.955 -46.755 108.285 ;
        RECT -47.085 106.595 -46.755 106.925 ;
        RECT -47.085 105.235 -46.755 105.565 ;
        RECT -47.085 103.875 -46.755 104.205 ;
        RECT -47.085 102.515 -46.755 102.845 ;
        RECT -47.085 101.155 -46.755 101.485 ;
        RECT -47.085 99.795 -46.755 100.125 ;
        RECT -47.085 98.435 -46.755 98.765 ;
        RECT -47.085 97.075 -46.755 97.405 ;
        RECT -47.085 95.715 -46.755 96.045 ;
        RECT -47.085 94.355 -46.755 94.685 ;
        RECT -47.085 92.995 -46.755 93.325 ;
        RECT -47.085 91.635 -46.755 91.965 ;
        RECT -47.085 90.275 -46.755 90.605 ;
        RECT -47.085 88.915 -46.755 89.245 ;
        RECT -47.085 87.555 -46.755 87.885 ;
        RECT -47.085 86.195 -46.755 86.525 ;
        RECT -47.085 84.835 -46.755 85.165 ;
        RECT -47.085 83.475 -46.755 83.805 ;
        RECT -47.085 82.115 -46.755 82.445 ;
        RECT -47.085 80.755 -46.755 81.085 ;
        RECT -47.085 79.395 -46.755 79.725 ;
        RECT -47.085 78.035 -46.755 78.365 ;
        RECT -47.085 76.675 -46.755 77.005 ;
        RECT -47.085 75.315 -46.755 75.645 ;
        RECT -47.085 73.955 -46.755 74.285 ;
        RECT -47.085 71.64 -46.755 71.97 ;
        RECT -47.085 69.465 -46.755 69.795 ;
        RECT -47.085 68.615 -46.755 68.945 ;
        RECT -47.085 66.305 -46.755 66.635 ;
        RECT -47.085 65.455 -46.755 65.785 ;
        RECT -47.085 63.145 -46.755 63.475 ;
        RECT -47.085 62.295 -46.755 62.625 ;
        RECT -47.085 59.985 -46.755 60.315 ;
        RECT -47.085 59.135 -46.755 59.465 ;
        RECT -47.085 56.825 -46.755 57.155 ;
        RECT -47.085 55.975 -46.755 56.305 ;
        RECT -47.085 53.665 -46.755 53.995 ;
        RECT -47.085 52.815 -46.755 53.145 ;
        RECT -47.085 50.64 -46.755 50.97 ;
        RECT -47.085 48.115 -46.755 48.445 ;
        RECT -47.085 46.755 -46.755 47.085 ;
        RECT -47.085 45.395 -46.755 45.725 ;
        RECT -47.085 44.035 -46.755 44.365 ;
        RECT -47.085 42.675 -46.755 43.005 ;
        RECT -47.085 41.315 -46.755 41.645 ;
        RECT -47.085 39.955 -46.755 40.285 ;
        RECT -47.085 38.595 -46.755 38.925 ;
        RECT -47.085 37.235 -46.755 37.565 ;
        RECT -47.085 35.875 -46.755 36.205 ;
        RECT -47.085 34.515 -46.755 34.845 ;
        RECT -47.085 33.155 -46.755 33.485 ;
        RECT -47.085 31.795 -46.755 32.125 ;
        RECT -47.085 30.435 -46.755 30.765 ;
        RECT -47.085 29.075 -46.755 29.405 ;
        RECT -47.085 27.715 -46.755 28.045 ;
        RECT -47.085 26.355 -46.755 26.685 ;
        RECT -47.085 24.995 -46.755 25.325 ;
        RECT -47.085 23.635 -46.755 23.965 ;
        RECT -47.085 22.275 -46.755 22.605 ;
        RECT -47.085 20.915 -46.755 21.245 ;
        RECT -47.085 19.555 -46.755 19.885 ;
        RECT -47.085 18.195 -46.755 18.525 ;
        RECT -47.085 16.835 -46.755 17.165 ;
        RECT -47.085 15.475 -46.755 15.805 ;
        RECT -47.085 14.115 -46.755 14.445 ;
        RECT -47.085 12.755 -46.755 13.085 ;
        RECT -47.085 11.395 -46.755 11.725 ;
        RECT -47.085 10.035 -46.755 10.365 ;
        RECT -47.085 8.675 -46.755 9.005 ;
        RECT -47.085 7.315 -46.755 7.645 ;
        RECT -47.085 5.955 -46.755 6.285 ;
        RECT -47.085 4.595 -46.755 4.925 ;
        RECT -47.085 3.235 -46.755 3.565 ;
        RECT -47.085 1.875 -46.755 2.205 ;
        RECT -47.085 0.515 -46.755 0.845 ;
        RECT -47.085 -0.845 -46.755 -0.515 ;
        RECT -47.085 -2.205 -46.755 -1.875 ;
        RECT -47.085 -3.565 -46.755 -3.235 ;
        RECT -47.085 -4.925 -46.755 -4.595 ;
        RECT -47.085 -6.285 -46.755 -5.955 ;
        RECT -47.085 -7.645 -46.755 -7.315 ;
        RECT -47.085 -9.005 -46.755 -8.675 ;
        RECT -47.085 -10.365 -46.755 -10.035 ;
        RECT -47.085 -11.725 -46.755 -11.395 ;
        RECT -47.085 -13.085 -46.755 -12.755 ;
        RECT -47.085 -14.445 -46.755 -14.115 ;
        RECT -47.085 -15.805 -46.755 -15.475 ;
        RECT -47.085 -17.165 -46.755 -16.835 ;
        RECT -47.085 -18.525 -46.755 -18.195 ;
        RECT -47.085 -19.885 -46.755 -19.555 ;
        RECT -47.085 -21.245 -46.755 -20.915 ;
        RECT -47.085 -22.605 -46.755 -22.275 ;
        RECT -47.085 -26.685 -46.755 -26.355 ;
        RECT -47.085 -28.045 -46.755 -27.715 ;
        RECT -47.085 -29.405 -46.755 -29.075 ;
        RECT -47.085 -30.765 -46.755 -30.435 ;
        RECT -47.085 -32.125 -46.755 -31.795 ;
        RECT -47.085 -33.485 -46.755 -33.155 ;
        RECT -47.085 -34.845 -46.755 -34.515 ;
        RECT -47.085 -36.205 -46.755 -35.875 ;
        RECT -47.085 -37.565 -46.755 -37.235 ;
        RECT -47.085 -38.925 -46.755 -38.595 ;
        RECT -47.085 -40.285 -46.755 -39.955 ;
        RECT -47.085 -41.645 -46.755 -41.315 ;
        RECT -47.085 -43.005 -46.755 -42.675 ;
        RECT -47.085 -44.365 -46.755 -44.035 ;
        RECT -47.085 -45.725 -46.755 -45.395 ;
        RECT -47.085 -47.085 -46.755 -46.755 ;
        RECT -47.085 -48.445 -46.755 -48.115 ;
        RECT -47.085 -49.805 -46.755 -49.475 ;
        RECT -47.085 -51.165 -46.755 -50.835 ;
        RECT -47.085 -52.525 -46.755 -52.195 ;
        RECT -47.085 -53.885 -46.755 -53.555 ;
        RECT -47.085 -55.245 -46.755 -54.915 ;
        RECT -47.085 -56.605 -46.755 -56.275 ;
        RECT -47.085 -57.965 -46.755 -57.635 ;
        RECT -47.085 -59.325 -46.755 -58.995 ;
        RECT -47.085 -60.685 -46.755 -60.355 ;
        RECT -47.085 -62.045 -46.755 -61.715 ;
        RECT -47.085 -63.405 -46.755 -63.075 ;
        RECT -47.085 -64.765 -46.755 -64.435 ;
        RECT -47.085 -66.125 -46.755 -65.795 ;
        RECT -47.085 -67.485 -46.755 -67.155 ;
        RECT -47.085 -68.845 -46.755 -68.515 ;
        RECT -47.085 -70.37 -46.755 -70.04 ;
        RECT -47.085 -71.565 -46.755 -71.235 ;
        RECT -47.085 -72.925 -46.755 -72.595 ;
        RECT -47.085 -74.285 -46.755 -73.955 ;
        RECT -47.085 -75.645 -46.755 -75.315 ;
        RECT -47.085 -77.005 -46.755 -76.675 ;
        RECT -47.085 -79.725 -46.755 -79.395 ;
        RECT -47.085 -80.91 -46.755 -80.58 ;
        RECT -47.085 -82.445 -46.755 -82.115 ;
        RECT -47.085 -83.805 -46.755 -83.475 ;
        RECT -47.085 -85.165 -46.755 -84.835 ;
        RECT -47.085 -87.885 -46.755 -87.555 ;
        RECT -47.085 -89.245 -46.755 -88.915 ;
        RECT -47.085 -93.325 -46.755 -92.995 ;
        RECT -47.085 -94.685 -46.755 -94.355 ;
        RECT -47.085 -96.045 -46.755 -95.715 ;
        RECT -47.085 -98.765 -46.755 -98.435 ;
        RECT -47.085 -100.125 -46.755 -99.795 ;
        RECT -47.085 -101.485 -46.755 -101.155 ;
        RECT -47.085 -102.845 -46.755 -102.515 ;
        RECT -47.085 -104.205 -46.755 -103.875 ;
        RECT -47.085 -105.565 -46.755 -105.235 ;
        RECT -47.085 -106.925 -46.755 -106.595 ;
        RECT -47.085 -108.285 -46.755 -107.955 ;
        RECT -47.085 -109.645 -46.755 -109.315 ;
        RECT -47.085 -111.005 -46.755 -110.675 ;
        RECT -47.085 -112.365 -46.755 -112.035 ;
        RECT -47.085 -113.725 -46.755 -113.395 ;
        RECT -47.085 -115.085 -46.755 -114.755 ;
        RECT -47.085 -116.445 -46.755 -116.115 ;
        RECT -47.085 -117.805 -46.755 -117.475 ;
        RECT -47.085 -119.165 -46.755 -118.835 ;
        RECT -47.085 -120.525 -46.755 -120.195 ;
        RECT -47.085 -121.885 -46.755 -121.555 ;
        RECT -47.085 -123.245 -46.755 -122.915 ;
        RECT -47.085 -124.605 -46.755 -124.275 ;
        RECT -47.085 -125.965 -46.755 -125.635 ;
        RECT -47.085 -127.325 -46.755 -126.995 ;
        RECT -47.085 -128.685 -46.755 -128.355 ;
        RECT -47.085 -130.045 -46.755 -129.715 ;
        RECT -47.085 -131.405 -46.755 -131.075 ;
        RECT -47.085 -132.765 -46.755 -132.435 ;
        RECT -47.085 -134.125 -46.755 -133.795 ;
        RECT -47.085 -135.485 -46.755 -135.155 ;
        RECT -47.085 -136.845 -46.755 -136.515 ;
        RECT -47.085 -138.205 -46.755 -137.875 ;
        RECT -47.085 -139.565 -46.755 -139.235 ;
        RECT -47.085 -140.925 -46.755 -140.595 ;
        RECT -47.085 -142.285 -46.755 -141.955 ;
        RECT -47.085 -143.645 -46.755 -143.315 ;
        RECT -47.085 -145.005 -46.755 -144.675 ;
        RECT -47.085 -146.365 -46.755 -146.035 ;
        RECT -47.085 -149.085 -46.755 -148.755 ;
        RECT -47.085 -150.445 -46.755 -150.115 ;
        RECT -47.085 -154.525 -46.755 -154.195 ;
        RECT -47.085 -157.245 -46.755 -156.915 ;
        RECT -47.085 -162.89 -46.755 -161.76 ;
        RECT -47.08 -163.005 -46.76 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 129.945 -45.395 131.075 ;
        RECT -45.725 125.635 -45.395 125.965 ;
        RECT -45.725 124.275 -45.395 124.605 ;
        RECT -45.725 122.915 -45.395 123.245 ;
        RECT -45.725 121.555 -45.395 121.885 ;
        RECT -45.725 120.195 -45.395 120.525 ;
        RECT -45.725 118.835 -45.395 119.165 ;
        RECT -45.725 117.475 -45.395 117.805 ;
        RECT -45.725 116.115 -45.395 116.445 ;
        RECT -45.725 114.755 -45.395 115.085 ;
        RECT -45.725 113.395 -45.395 113.725 ;
        RECT -45.725 112.035 -45.395 112.365 ;
        RECT -45.725 110.675 -45.395 111.005 ;
        RECT -45.725 109.315 -45.395 109.645 ;
        RECT -45.725 107.955 -45.395 108.285 ;
        RECT -45.725 106.595 -45.395 106.925 ;
        RECT -45.725 105.235 -45.395 105.565 ;
        RECT -45.725 103.875 -45.395 104.205 ;
        RECT -45.725 102.515 -45.395 102.845 ;
        RECT -45.725 101.155 -45.395 101.485 ;
        RECT -45.725 99.795 -45.395 100.125 ;
        RECT -45.725 98.435 -45.395 98.765 ;
        RECT -45.725 97.075 -45.395 97.405 ;
        RECT -45.725 95.715 -45.395 96.045 ;
        RECT -45.725 94.355 -45.395 94.685 ;
        RECT -45.725 92.995 -45.395 93.325 ;
        RECT -45.725 91.635 -45.395 91.965 ;
        RECT -45.725 90.275 -45.395 90.605 ;
        RECT -45.725 88.915 -45.395 89.245 ;
        RECT -45.725 87.555 -45.395 87.885 ;
        RECT -45.725 86.195 -45.395 86.525 ;
        RECT -45.725 84.835 -45.395 85.165 ;
        RECT -45.725 83.475 -45.395 83.805 ;
        RECT -45.725 82.115 -45.395 82.445 ;
        RECT -45.725 80.755 -45.395 81.085 ;
        RECT -45.725 79.395 -45.395 79.725 ;
        RECT -45.725 78.035 -45.395 78.365 ;
        RECT -45.725 76.675 -45.395 77.005 ;
        RECT -45.725 75.315 -45.395 75.645 ;
        RECT -45.725 73.955 -45.395 74.285 ;
        RECT -45.725 71.64 -45.395 71.97 ;
        RECT -45.725 69.465 -45.395 69.795 ;
        RECT -45.725 68.615 -45.395 68.945 ;
        RECT -45.725 66.305 -45.395 66.635 ;
        RECT -45.725 65.455 -45.395 65.785 ;
        RECT -45.725 63.145 -45.395 63.475 ;
        RECT -45.725 62.295 -45.395 62.625 ;
        RECT -45.725 59.985 -45.395 60.315 ;
        RECT -45.725 59.135 -45.395 59.465 ;
        RECT -45.725 56.825 -45.395 57.155 ;
        RECT -45.725 55.975 -45.395 56.305 ;
        RECT -45.725 53.665 -45.395 53.995 ;
        RECT -45.725 52.815 -45.395 53.145 ;
        RECT -45.725 50.64 -45.395 50.97 ;
        RECT -45.725 48.115 -45.395 48.445 ;
        RECT -45.725 46.755 -45.395 47.085 ;
        RECT -45.725 45.395 -45.395 45.725 ;
        RECT -45.725 44.035 -45.395 44.365 ;
        RECT -45.725 42.675 -45.395 43.005 ;
        RECT -45.725 41.315 -45.395 41.645 ;
        RECT -45.725 39.955 -45.395 40.285 ;
        RECT -45.725 38.595 -45.395 38.925 ;
        RECT -45.725 37.235 -45.395 37.565 ;
        RECT -45.725 35.875 -45.395 36.205 ;
        RECT -45.725 34.515 -45.395 34.845 ;
        RECT -45.725 33.155 -45.395 33.485 ;
        RECT -45.725 31.795 -45.395 32.125 ;
        RECT -45.725 30.435 -45.395 30.765 ;
        RECT -45.725 29.075 -45.395 29.405 ;
        RECT -45.725 27.715 -45.395 28.045 ;
        RECT -45.725 26.355 -45.395 26.685 ;
        RECT -45.725 24.995 -45.395 25.325 ;
        RECT -45.725 23.635 -45.395 23.965 ;
        RECT -45.725 22.275 -45.395 22.605 ;
        RECT -45.725 20.915 -45.395 21.245 ;
        RECT -45.725 19.555 -45.395 19.885 ;
        RECT -45.725 18.195 -45.395 18.525 ;
        RECT -45.725 16.835 -45.395 17.165 ;
        RECT -45.725 15.475 -45.395 15.805 ;
        RECT -45.725 14.115 -45.395 14.445 ;
        RECT -45.725 12.755 -45.395 13.085 ;
        RECT -45.725 11.395 -45.395 11.725 ;
        RECT -45.725 10.035 -45.395 10.365 ;
        RECT -45.725 8.675 -45.395 9.005 ;
        RECT -45.725 7.315 -45.395 7.645 ;
        RECT -45.725 5.955 -45.395 6.285 ;
        RECT -45.725 4.595 -45.395 4.925 ;
        RECT -45.725 3.235 -45.395 3.565 ;
        RECT -45.725 1.875 -45.395 2.205 ;
        RECT -45.725 0.515 -45.395 0.845 ;
        RECT -45.725 -0.845 -45.395 -0.515 ;
        RECT -45.725 -2.205 -45.395 -1.875 ;
        RECT -45.725 -3.565 -45.395 -3.235 ;
        RECT -45.725 -4.925 -45.395 -4.595 ;
        RECT -45.725 -6.285 -45.395 -5.955 ;
        RECT -45.725 -7.645 -45.395 -7.315 ;
        RECT -45.725 -9.005 -45.395 -8.675 ;
        RECT -45.725 -11.725 -45.395 -11.395 ;
        RECT -45.725 -13.085 -45.395 -12.755 ;
        RECT -45.725 -14.445 -45.395 -14.115 ;
        RECT -45.725 -15.805 -45.395 -15.475 ;
        RECT -45.725 -17.165 -45.395 -16.835 ;
        RECT -45.725 -18.525 -45.395 -18.195 ;
        RECT -45.725 -19.885 -45.395 -19.555 ;
        RECT -45.725 -21.245 -45.395 -20.915 ;
        RECT -45.725 -22.605 -45.395 -22.275 ;
        RECT -45.725 -26.685 -45.395 -26.355 ;
        RECT -45.725 -28.045 -45.395 -27.715 ;
        RECT -45.725 -29.405 -45.395 -29.075 ;
        RECT -45.725 -30.765 -45.395 -30.435 ;
        RECT -45.725 -32.125 -45.395 -31.795 ;
        RECT -45.725 -33.485 -45.395 -33.155 ;
        RECT -45.725 -34.845 -45.395 -34.515 ;
        RECT -45.725 -36.205 -45.395 -35.875 ;
        RECT -45.725 -37.565 -45.395 -37.235 ;
        RECT -45.725 -38.925 -45.395 -38.595 ;
        RECT -45.725 -40.285 -45.395 -39.955 ;
        RECT -45.725 -41.645 -45.395 -41.315 ;
        RECT -45.725 -43.005 -45.395 -42.675 ;
        RECT -45.725 -44.365 -45.395 -44.035 ;
        RECT -45.725 -45.725 -45.395 -45.395 ;
        RECT -45.725 -47.085 -45.395 -46.755 ;
        RECT -45.725 -48.445 -45.395 -48.115 ;
        RECT -45.725 -49.805 -45.395 -49.475 ;
        RECT -45.725 -51.165 -45.395 -50.835 ;
        RECT -45.725 -52.525 -45.395 -52.195 ;
        RECT -45.725 -53.885 -45.395 -53.555 ;
        RECT -45.725 -55.245 -45.395 -54.915 ;
        RECT -45.725 -56.605 -45.395 -56.275 ;
        RECT -45.725 -57.965 -45.395 -57.635 ;
        RECT -45.725 -59.325 -45.395 -58.995 ;
        RECT -45.725 -60.685 -45.395 -60.355 ;
        RECT -45.725 -62.045 -45.395 -61.715 ;
        RECT -45.725 -63.405 -45.395 -63.075 ;
        RECT -45.725 -64.765 -45.395 -64.435 ;
        RECT -45.725 -66.125 -45.395 -65.795 ;
        RECT -45.725 -67.485 -45.395 -67.155 ;
        RECT -45.725 -68.845 -45.395 -68.515 ;
        RECT -45.725 -70.37 -45.395 -70.04 ;
        RECT -45.725 -71.565 -45.395 -71.235 ;
        RECT -45.725 -72.925 -45.395 -72.595 ;
        RECT -45.725 -74.285 -45.395 -73.955 ;
        RECT -45.725 -75.645 -45.395 -75.315 ;
        RECT -45.725 -77.005 -45.395 -76.675 ;
        RECT -45.725 -79.725 -45.395 -79.395 ;
        RECT -45.725 -80.91 -45.395 -80.58 ;
        RECT -45.725 -82.445 -45.395 -82.115 ;
        RECT -45.725 -83.805 -45.395 -83.475 ;
        RECT -45.725 -85.165 -45.395 -84.835 ;
        RECT -45.725 -87.885 -45.395 -87.555 ;
        RECT -45.725 -89.245 -45.395 -88.915 ;
        RECT -45.725 -93.325 -45.395 -92.995 ;
        RECT -45.725 -94.685 -45.395 -94.355 ;
        RECT -45.725 -96.045 -45.395 -95.715 ;
        RECT -45.725 -98.765 -45.395 -98.435 ;
        RECT -45.725 -100.125 -45.395 -99.795 ;
        RECT -45.725 -101.485 -45.395 -101.155 ;
        RECT -45.725 -102.845 -45.395 -102.515 ;
        RECT -45.725 -104.205 -45.395 -103.875 ;
        RECT -45.725 -105.565 -45.395 -105.235 ;
        RECT -45.725 -106.925 -45.395 -106.595 ;
        RECT -45.725 -108.285 -45.395 -107.955 ;
        RECT -45.725 -109.645 -45.395 -109.315 ;
        RECT -45.725 -111.005 -45.395 -110.675 ;
        RECT -45.725 -112.365 -45.395 -112.035 ;
        RECT -45.725 -113.725 -45.395 -113.395 ;
        RECT -45.725 -115.085 -45.395 -114.755 ;
        RECT -45.725 -116.445 -45.395 -116.115 ;
        RECT -45.725 -117.805 -45.395 -117.475 ;
        RECT -45.725 -119.165 -45.395 -118.835 ;
        RECT -45.725 -120.525 -45.395 -120.195 ;
        RECT -45.725 -121.885 -45.395 -121.555 ;
        RECT -45.725 -123.245 -45.395 -122.915 ;
        RECT -45.725 -124.605 -45.395 -124.275 ;
        RECT -45.725 -125.965 -45.395 -125.635 ;
        RECT -45.725 -127.325 -45.395 -126.995 ;
        RECT -45.725 -128.685 -45.395 -128.355 ;
        RECT -45.725 -130.045 -45.395 -129.715 ;
        RECT -45.725 -131.405 -45.395 -131.075 ;
        RECT -45.725 -132.765 -45.395 -132.435 ;
        RECT -45.725 -134.125 -45.395 -133.795 ;
        RECT -45.725 -135.485 -45.395 -135.155 ;
        RECT -45.725 -136.845 -45.395 -136.515 ;
        RECT -45.725 -138.205 -45.395 -137.875 ;
        RECT -45.725 -139.565 -45.395 -139.235 ;
        RECT -45.725 -140.925 -45.395 -140.595 ;
        RECT -45.725 -142.285 -45.395 -141.955 ;
        RECT -45.725 -143.645 -45.395 -143.315 ;
        RECT -45.725 -145.005 -45.395 -144.675 ;
        RECT -45.725 -146.365 -45.395 -146.035 ;
        RECT -45.725 -148.215 -45.395 -147.885 ;
        RECT -45.725 -149.085 -45.395 -148.755 ;
        RECT -45.725 -150.445 -45.395 -150.115 ;
        RECT -45.725 -151.805 -45.395 -151.475 ;
        RECT -45.725 -154.525 -45.395 -154.195 ;
        RECT -45.725 -157.245 -45.395 -156.915 ;
        RECT -45.725 -162.89 -45.395 -161.76 ;
        RECT -45.72 -163.005 -45.4 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 129.945 -44.035 131.075 ;
        RECT -44.365 125.635 -44.035 125.965 ;
        RECT -44.365 124.275 -44.035 124.605 ;
        RECT -44.365 122.915 -44.035 123.245 ;
        RECT -44.365 121.555 -44.035 121.885 ;
        RECT -44.365 120.195 -44.035 120.525 ;
        RECT -44.365 118.835 -44.035 119.165 ;
        RECT -44.365 117.475 -44.035 117.805 ;
        RECT -44.365 116.115 -44.035 116.445 ;
        RECT -44.365 114.755 -44.035 115.085 ;
        RECT -44.365 113.395 -44.035 113.725 ;
        RECT -44.365 112.035 -44.035 112.365 ;
        RECT -44.365 110.675 -44.035 111.005 ;
        RECT -44.365 109.315 -44.035 109.645 ;
        RECT -44.365 107.955 -44.035 108.285 ;
        RECT -44.365 106.595 -44.035 106.925 ;
        RECT -44.365 105.235 -44.035 105.565 ;
        RECT -44.365 103.875 -44.035 104.205 ;
        RECT -44.365 102.515 -44.035 102.845 ;
        RECT -44.365 101.155 -44.035 101.485 ;
        RECT -44.365 99.795 -44.035 100.125 ;
        RECT -44.365 98.435 -44.035 98.765 ;
        RECT -44.365 97.075 -44.035 97.405 ;
        RECT -44.365 95.715 -44.035 96.045 ;
        RECT -44.365 94.355 -44.035 94.685 ;
        RECT -44.365 92.995 -44.035 93.325 ;
        RECT -44.365 91.635 -44.035 91.965 ;
        RECT -44.365 90.275 -44.035 90.605 ;
        RECT -44.365 88.915 -44.035 89.245 ;
        RECT -44.365 87.555 -44.035 87.885 ;
        RECT -44.365 86.195 -44.035 86.525 ;
        RECT -44.365 84.835 -44.035 85.165 ;
        RECT -44.365 83.475 -44.035 83.805 ;
        RECT -44.365 82.115 -44.035 82.445 ;
        RECT -44.365 80.755 -44.035 81.085 ;
        RECT -44.365 79.395 -44.035 79.725 ;
        RECT -44.365 78.035 -44.035 78.365 ;
        RECT -44.365 76.675 -44.035 77.005 ;
        RECT -44.365 75.315 -44.035 75.645 ;
        RECT -44.365 73.955 -44.035 74.285 ;
        RECT -44.365 71.64 -44.035 71.97 ;
        RECT -44.365 69.465 -44.035 69.795 ;
        RECT -44.365 68.615 -44.035 68.945 ;
        RECT -44.365 66.305 -44.035 66.635 ;
        RECT -44.365 65.455 -44.035 65.785 ;
        RECT -44.365 63.145 -44.035 63.475 ;
        RECT -44.365 62.295 -44.035 62.625 ;
        RECT -44.365 59.985 -44.035 60.315 ;
        RECT -44.365 59.135 -44.035 59.465 ;
        RECT -44.365 56.825 -44.035 57.155 ;
        RECT -44.365 55.975 -44.035 56.305 ;
        RECT -44.365 53.665 -44.035 53.995 ;
        RECT -44.365 52.815 -44.035 53.145 ;
        RECT -44.365 50.64 -44.035 50.97 ;
        RECT -44.365 48.115 -44.035 48.445 ;
        RECT -44.365 46.755 -44.035 47.085 ;
        RECT -44.365 45.395 -44.035 45.725 ;
        RECT -44.365 44.035 -44.035 44.365 ;
        RECT -44.365 42.675 -44.035 43.005 ;
        RECT -44.365 41.315 -44.035 41.645 ;
        RECT -44.365 39.955 -44.035 40.285 ;
        RECT -44.365 38.595 -44.035 38.925 ;
        RECT -44.365 37.235 -44.035 37.565 ;
        RECT -44.365 35.875 -44.035 36.205 ;
        RECT -44.365 34.515 -44.035 34.845 ;
        RECT -44.365 33.155 -44.035 33.485 ;
        RECT -44.365 31.795 -44.035 32.125 ;
        RECT -44.365 30.435 -44.035 30.765 ;
        RECT -44.365 29.075 -44.035 29.405 ;
        RECT -44.365 27.715 -44.035 28.045 ;
        RECT -44.365 26.355 -44.035 26.685 ;
        RECT -44.365 24.995 -44.035 25.325 ;
        RECT -44.365 23.635 -44.035 23.965 ;
        RECT -44.365 22.275 -44.035 22.605 ;
        RECT -44.365 20.915 -44.035 21.245 ;
        RECT -44.365 19.555 -44.035 19.885 ;
        RECT -44.365 18.195 -44.035 18.525 ;
        RECT -44.365 16.835 -44.035 17.165 ;
        RECT -44.365 15.475 -44.035 15.805 ;
        RECT -44.365 14.115 -44.035 14.445 ;
        RECT -44.365 12.755 -44.035 13.085 ;
        RECT -44.365 11.395 -44.035 11.725 ;
        RECT -44.365 10.035 -44.035 10.365 ;
        RECT -44.365 8.675 -44.035 9.005 ;
        RECT -44.365 7.315 -44.035 7.645 ;
        RECT -44.365 5.955 -44.035 6.285 ;
        RECT -44.365 4.595 -44.035 4.925 ;
        RECT -44.365 3.235 -44.035 3.565 ;
        RECT -44.365 1.875 -44.035 2.205 ;
        RECT -44.365 0.515 -44.035 0.845 ;
        RECT -44.365 -0.845 -44.035 -0.515 ;
        RECT -44.365 -2.205 -44.035 -1.875 ;
        RECT -44.365 -3.565 -44.035 -3.235 ;
        RECT -44.365 -4.925 -44.035 -4.595 ;
        RECT -44.365 -6.285 -44.035 -5.955 ;
        RECT -44.365 -7.645 -44.035 -7.315 ;
        RECT -44.365 -11.725 -44.035 -11.395 ;
        RECT -44.365 -13.085 -44.035 -12.755 ;
        RECT -44.365 -14.445 -44.035 -14.115 ;
        RECT -44.365 -15.805 -44.035 -15.475 ;
        RECT -44.365 -17.165 -44.035 -16.835 ;
        RECT -44.365 -19.885 -44.035 -19.555 ;
        RECT -44.365 -21.245 -44.035 -20.915 ;
        RECT -44.365 -22.605 -44.035 -22.275 ;
        RECT -44.365 -26.685 -44.035 -26.355 ;
        RECT -44.365 -28.045 -44.035 -27.715 ;
        RECT -44.365 -29.405 -44.035 -29.075 ;
        RECT -44.365 -30.765 -44.035 -30.435 ;
        RECT -44.365 -32.125 -44.035 -31.795 ;
        RECT -44.365 -33.485 -44.035 -33.155 ;
        RECT -44.365 -34.845 -44.035 -34.515 ;
        RECT -44.365 -36.205 -44.035 -35.875 ;
        RECT -44.365 -37.565 -44.035 -37.235 ;
        RECT -44.365 -38.925 -44.035 -38.595 ;
        RECT -44.365 -40.285 -44.035 -39.955 ;
        RECT -44.365 -41.645 -44.035 -41.315 ;
        RECT -44.365 -43.005 -44.035 -42.675 ;
        RECT -44.365 -44.365 -44.035 -44.035 ;
        RECT -44.365 -45.725 -44.035 -45.395 ;
        RECT -44.365 -47.085 -44.035 -46.755 ;
        RECT -44.365 -48.445 -44.035 -48.115 ;
        RECT -44.365 -49.805 -44.035 -49.475 ;
        RECT -44.365 -51.165 -44.035 -50.835 ;
        RECT -44.365 -52.525 -44.035 -52.195 ;
        RECT -44.365 -53.885 -44.035 -53.555 ;
        RECT -44.365 -55.245 -44.035 -54.915 ;
        RECT -44.365 -56.605 -44.035 -56.275 ;
        RECT -44.365 -57.965 -44.035 -57.635 ;
        RECT -44.365 -59.325 -44.035 -58.995 ;
        RECT -44.365 -60.685 -44.035 -60.355 ;
        RECT -44.365 -62.045 -44.035 -61.715 ;
        RECT -44.365 -63.405 -44.035 -63.075 ;
        RECT -44.365 -64.765 -44.035 -64.435 ;
        RECT -44.365 -66.125 -44.035 -65.795 ;
        RECT -44.365 -67.485 -44.035 -67.155 ;
        RECT -44.365 -68.845 -44.035 -68.515 ;
        RECT -44.365 -70.37 -44.035 -70.04 ;
        RECT -44.365 -71.565 -44.035 -71.235 ;
        RECT -44.365 -72.925 -44.035 -72.595 ;
        RECT -44.365 -74.285 -44.035 -73.955 ;
        RECT -44.365 -75.645 -44.035 -75.315 ;
        RECT -44.365 -77.005 -44.035 -76.675 ;
        RECT -44.365 -79.725 -44.035 -79.395 ;
        RECT -44.365 -80.91 -44.035 -80.58 ;
        RECT -44.365 -82.445 -44.035 -82.115 ;
        RECT -44.365 -83.805 -44.035 -83.475 ;
        RECT -44.365 -85.165 -44.035 -84.835 ;
        RECT -44.365 -87.885 -44.035 -87.555 ;
        RECT -44.365 -89.245 -44.035 -88.915 ;
        RECT -44.365 -93.325 -44.035 -92.995 ;
        RECT -44.365 -94.685 -44.035 -94.355 ;
        RECT -44.365 -96.045 -44.035 -95.715 ;
        RECT -44.365 -98.765 -44.035 -98.435 ;
        RECT -44.365 -100.125 -44.035 -99.795 ;
        RECT -44.365 -101.485 -44.035 -101.155 ;
        RECT -44.365 -102.845 -44.035 -102.515 ;
        RECT -44.365 -104.205 -44.035 -103.875 ;
        RECT -44.365 -105.565 -44.035 -105.235 ;
        RECT -44.365 -106.925 -44.035 -106.595 ;
        RECT -44.365 -108.285 -44.035 -107.955 ;
        RECT -44.365 -109.645 -44.035 -109.315 ;
        RECT -44.365 -111.005 -44.035 -110.675 ;
        RECT -44.365 -112.365 -44.035 -112.035 ;
        RECT -44.365 -113.725 -44.035 -113.395 ;
        RECT -44.365 -115.085 -44.035 -114.755 ;
        RECT -44.365 -116.445 -44.035 -116.115 ;
        RECT -44.365 -117.805 -44.035 -117.475 ;
        RECT -44.365 -119.165 -44.035 -118.835 ;
        RECT -44.365 -120.525 -44.035 -120.195 ;
        RECT -44.365 -121.885 -44.035 -121.555 ;
        RECT -44.365 -123.245 -44.035 -122.915 ;
        RECT -44.365 -124.605 -44.035 -124.275 ;
        RECT -44.365 -125.965 -44.035 -125.635 ;
        RECT -44.365 -127.325 -44.035 -126.995 ;
        RECT -44.365 -128.685 -44.035 -128.355 ;
        RECT -44.365 -130.045 -44.035 -129.715 ;
        RECT -44.365 -131.405 -44.035 -131.075 ;
        RECT -44.365 -132.765 -44.035 -132.435 ;
        RECT -44.365 -134.125 -44.035 -133.795 ;
        RECT -44.365 -135.485 -44.035 -135.155 ;
        RECT -44.365 -136.845 -44.035 -136.515 ;
        RECT -44.365 -138.205 -44.035 -137.875 ;
        RECT -44.365 -139.565 -44.035 -139.235 ;
        RECT -44.365 -140.925 -44.035 -140.595 ;
        RECT -44.365 -142.285 -44.035 -141.955 ;
        RECT -44.365 -143.645 -44.035 -143.315 ;
        RECT -44.365 -145.005 -44.035 -144.675 ;
        RECT -44.365 -146.365 -44.035 -146.035 ;
        RECT -44.365 -148.215 -44.035 -147.885 ;
        RECT -44.365 -149.085 -44.035 -148.755 ;
        RECT -44.365 -150.445 -44.035 -150.115 ;
        RECT -44.365 -154.525 -44.035 -154.195 ;
        RECT -44.365 -157.245 -44.035 -156.915 ;
        RECT -44.365 -162.89 -44.035 -161.76 ;
        RECT -44.36 -163.005 -44.04 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 14.115 -42.675 14.445 ;
        RECT -43.005 12.755 -42.675 13.085 ;
        RECT -43.005 11.395 -42.675 11.725 ;
        RECT -43.005 10.035 -42.675 10.365 ;
        RECT -43.005 8.675 -42.675 9.005 ;
        RECT -43.005 7.315 -42.675 7.645 ;
        RECT -43.005 5.955 -42.675 6.285 ;
        RECT -43.005 4.595 -42.675 4.925 ;
        RECT -43.005 3.235 -42.675 3.565 ;
        RECT -43.005 1.875 -42.675 2.205 ;
        RECT -43.005 0.515 -42.675 0.845 ;
        RECT -43.005 -0.845 -42.675 -0.515 ;
        RECT -43.005 -2.205 -42.675 -1.875 ;
        RECT -43.005 -3.565 -42.675 -3.235 ;
        RECT -43.005 -4.925 -42.675 -4.595 ;
        RECT -43.005 -7.645 -42.675 -7.315 ;
        RECT -43.005 -11.725 -42.675 -11.395 ;
        RECT -43.005 -13.085 -42.675 -12.755 ;
        RECT -43.005 -14.445 -42.675 -14.115 ;
        RECT -43.005 -15.805 -42.675 -15.475 ;
        RECT -43.005 -17.165 -42.675 -16.835 ;
        RECT -43.005 -19.885 -42.675 -19.555 ;
        RECT -43.005 -21.245 -42.675 -20.915 ;
        RECT -43.005 -22.605 -42.675 -22.275 ;
        RECT -43.005 -28.045 -42.675 -27.715 ;
        RECT -43.005 -29.405 -42.675 -29.075 ;
        RECT -43.005 -30.765 -42.675 -30.435 ;
        RECT -43.005 -32.125 -42.675 -31.795 ;
        RECT -43.005 -33.485 -42.675 -33.155 ;
        RECT -43.005 -34.845 -42.675 -34.515 ;
        RECT -43.005 -36.205 -42.675 -35.875 ;
        RECT -43.005 -37.565 -42.675 -37.235 ;
        RECT -43.005 -38.925 -42.675 -38.595 ;
        RECT -43.005 -40.285 -42.675 -39.955 ;
        RECT -43.005 -41.645 -42.675 -41.315 ;
        RECT -43.005 -43.005 -42.675 -42.675 ;
        RECT -43.005 -44.365 -42.675 -44.035 ;
        RECT -43.005 -45.725 -42.675 -45.395 ;
        RECT -43.005 -47.085 -42.675 -46.755 ;
        RECT -43.005 -48.445 -42.675 -48.115 ;
        RECT -43.005 -49.805 -42.675 -49.475 ;
        RECT -43.005 -51.165 -42.675 -50.835 ;
        RECT -43.005 -52.525 -42.675 -52.195 ;
        RECT -43.005 -53.885 -42.675 -53.555 ;
        RECT -43.005 -55.245 -42.675 -54.915 ;
        RECT -43.005 -56.605 -42.675 -56.275 ;
        RECT -43.005 -57.965 -42.675 -57.635 ;
        RECT -43.005 -59.325 -42.675 -58.995 ;
        RECT -43.005 -60.685 -42.675 -60.355 ;
        RECT -43.005 -62.045 -42.675 -61.715 ;
        RECT -43.005 -63.405 -42.675 -63.075 ;
        RECT -43.005 -64.765 -42.675 -64.435 ;
        RECT -43.005 -66.125 -42.675 -65.795 ;
        RECT -43.005 -67.485 -42.675 -67.155 ;
        RECT -43.005 -68.845 -42.675 -68.515 ;
        RECT -43.005 -70.37 -42.675 -70.04 ;
        RECT -43.005 -71.565 -42.675 -71.235 ;
        RECT -43.005 -72.925 -42.675 -72.595 ;
        RECT -43.005 -74.285 -42.675 -73.955 ;
        RECT -43.005 -75.645 -42.675 -75.315 ;
        RECT -43.005 -77.005 -42.675 -76.675 ;
        RECT -43.005 -79.725 -42.675 -79.395 ;
        RECT -43.005 -80.91 -42.675 -80.58 ;
        RECT -43.005 -82.445 -42.675 -82.115 ;
        RECT -43.005 -83.805 -42.675 -83.475 ;
        RECT -43.005 -85.165 -42.675 -84.835 ;
        RECT -43.005 -87.885 -42.675 -87.555 ;
        RECT -43.005 -89.245 -42.675 -88.915 ;
        RECT -43.005 -91.965 -42.675 -91.635 ;
        RECT -43.005 -93.325 -42.675 -92.995 ;
        RECT -43.005 -94.685 -42.675 -94.355 ;
        RECT -43.005 -96.045 -42.675 -95.715 ;
        RECT -43.005 -98.765 -42.675 -98.435 ;
        RECT -43.005 -100.125 -42.675 -99.795 ;
        RECT -43.005 -101.485 -42.675 -101.155 ;
        RECT -43.005 -102.845 -42.675 -102.515 ;
        RECT -43.005 -104.205 -42.675 -103.875 ;
        RECT -43.005 -105.565 -42.675 -105.235 ;
        RECT -43.005 -106.925 -42.675 -106.595 ;
        RECT -43.005 -108.285 -42.675 -107.955 ;
        RECT -43.005 -109.645 -42.675 -109.315 ;
        RECT -43.005 -111.005 -42.675 -110.675 ;
        RECT -43.005 -112.365 -42.675 -112.035 ;
        RECT -43.005 -113.725 -42.675 -113.395 ;
        RECT -43.005 -115.085 -42.675 -114.755 ;
        RECT -43.005 -116.445 -42.675 -116.115 ;
        RECT -43.005 -117.805 -42.675 -117.475 ;
        RECT -43.005 -119.165 -42.675 -118.835 ;
        RECT -43.005 -120.525 -42.675 -120.195 ;
        RECT -43.005 -121.885 -42.675 -121.555 ;
        RECT -43.005 -123.245 -42.675 -122.915 ;
        RECT -43.005 -124.605 -42.675 -124.275 ;
        RECT -43.005 -125.965 -42.675 -125.635 ;
        RECT -43.005 -127.325 -42.675 -126.995 ;
        RECT -43.005 -128.685 -42.675 -128.355 ;
        RECT -43.005 -130.045 -42.675 -129.715 ;
        RECT -43.005 -131.405 -42.675 -131.075 ;
        RECT -43.005 -132.765 -42.675 -132.435 ;
        RECT -43.005 -134.125 -42.675 -133.795 ;
        RECT -43.005 -135.485 -42.675 -135.155 ;
        RECT -43.005 -136.845 -42.675 -136.515 ;
        RECT -43.005 -138.205 -42.675 -137.875 ;
        RECT -43.005 -139.565 -42.675 -139.235 ;
        RECT -43.005 -140.925 -42.675 -140.595 ;
        RECT -43.005 -142.285 -42.675 -141.955 ;
        RECT -43.005 -143.645 -42.675 -143.315 ;
        RECT -43.005 -145.005 -42.675 -144.675 ;
        RECT -43.005 -146.365 -42.675 -146.035 ;
        RECT -43.005 -148.215 -42.675 -147.885 ;
        RECT -43.005 -149.085 -42.675 -148.755 ;
        RECT -43.005 -150.445 -42.675 -150.115 ;
        RECT -43.005 -151.805 -42.675 -151.475 ;
        RECT -43.005 -154.525 -42.675 -154.195 ;
        RECT -43.005 -157.245 -42.675 -156.915 ;
        RECT -43.005 -162.89 -42.675 -161.76 ;
        RECT -43 -163.005 -42.68 131.19 ;
        RECT -43.005 129.945 -42.675 131.075 ;
        RECT -43.005 125.635 -42.675 125.965 ;
        RECT -43.005 124.275 -42.675 124.605 ;
        RECT -43.005 122.915 -42.675 123.245 ;
        RECT -43.005 121.555 -42.675 121.885 ;
        RECT -43.005 120.195 -42.675 120.525 ;
        RECT -43.005 118.835 -42.675 119.165 ;
        RECT -43.005 117.475 -42.675 117.805 ;
        RECT -43.005 116.115 -42.675 116.445 ;
        RECT -43.005 114.755 -42.675 115.085 ;
        RECT -43.005 113.395 -42.675 113.725 ;
        RECT -43.005 112.035 -42.675 112.365 ;
        RECT -43.005 110.675 -42.675 111.005 ;
        RECT -43.005 109.315 -42.675 109.645 ;
        RECT -43.005 107.955 -42.675 108.285 ;
        RECT -43.005 106.595 -42.675 106.925 ;
        RECT -43.005 105.235 -42.675 105.565 ;
        RECT -43.005 103.875 -42.675 104.205 ;
        RECT -43.005 102.515 -42.675 102.845 ;
        RECT -43.005 101.155 -42.675 101.485 ;
        RECT -43.005 99.795 -42.675 100.125 ;
        RECT -43.005 98.435 -42.675 98.765 ;
        RECT -43.005 97.075 -42.675 97.405 ;
        RECT -43.005 95.715 -42.675 96.045 ;
        RECT -43.005 94.355 -42.675 94.685 ;
        RECT -43.005 92.995 -42.675 93.325 ;
        RECT -43.005 91.635 -42.675 91.965 ;
        RECT -43.005 90.275 -42.675 90.605 ;
        RECT -43.005 88.915 -42.675 89.245 ;
        RECT -43.005 87.555 -42.675 87.885 ;
        RECT -43.005 86.195 -42.675 86.525 ;
        RECT -43.005 84.835 -42.675 85.165 ;
        RECT -43.005 83.475 -42.675 83.805 ;
        RECT -43.005 82.115 -42.675 82.445 ;
        RECT -43.005 80.755 -42.675 81.085 ;
        RECT -43.005 79.395 -42.675 79.725 ;
        RECT -43.005 78.035 -42.675 78.365 ;
        RECT -43.005 76.675 -42.675 77.005 ;
        RECT -43.005 75.315 -42.675 75.645 ;
        RECT -43.005 73.955 -42.675 74.285 ;
        RECT -43.005 72.595 -42.675 72.925 ;
        RECT -43.005 71.235 -42.675 71.565 ;
        RECT -43.005 69.875 -42.675 70.205 ;
        RECT -43.005 68.515 -42.675 68.845 ;
        RECT -43.005 67.155 -42.675 67.485 ;
        RECT -43.005 65.795 -42.675 66.125 ;
        RECT -43.005 64.435 -42.675 64.765 ;
        RECT -43.005 63.075 -42.675 63.405 ;
        RECT -43.005 61.715 -42.675 62.045 ;
        RECT -43.005 60.355 -42.675 60.685 ;
        RECT -43.005 58.995 -42.675 59.325 ;
        RECT -43.005 57.635 -42.675 57.965 ;
        RECT -43.005 56.275 -42.675 56.605 ;
        RECT -43.005 54.915 -42.675 55.245 ;
        RECT -43.005 53.555 -42.675 53.885 ;
        RECT -43.005 52.195 -42.675 52.525 ;
        RECT -43.005 50.835 -42.675 51.165 ;
        RECT -43.005 49.475 -42.675 49.805 ;
        RECT -43.005 48.115 -42.675 48.445 ;
        RECT -43.005 46.755 -42.675 47.085 ;
        RECT -43.005 45.395 -42.675 45.725 ;
        RECT -43.005 44.035 -42.675 44.365 ;
        RECT -43.005 42.675 -42.675 43.005 ;
        RECT -43.005 41.315 -42.675 41.645 ;
        RECT -43.005 39.955 -42.675 40.285 ;
        RECT -43.005 38.595 -42.675 38.925 ;
        RECT -43.005 37.235 -42.675 37.565 ;
        RECT -43.005 35.875 -42.675 36.205 ;
        RECT -43.005 34.515 -42.675 34.845 ;
        RECT -43.005 33.155 -42.675 33.485 ;
        RECT -43.005 31.795 -42.675 32.125 ;
        RECT -43.005 30.435 -42.675 30.765 ;
        RECT -43.005 29.075 -42.675 29.405 ;
        RECT -43.005 27.715 -42.675 28.045 ;
        RECT -43.005 26.355 -42.675 26.685 ;
        RECT -43.005 24.995 -42.675 25.325 ;
        RECT -43.005 23.635 -42.675 23.965 ;
        RECT -43.005 22.275 -42.675 22.605 ;
        RECT -43.005 20.915 -42.675 21.245 ;
        RECT -43.005 19.555 -42.675 19.885 ;
        RECT -43.005 18.195 -42.675 18.525 ;
        RECT -43.005 16.835 -42.675 17.165 ;
        RECT -43.005 15.475 -42.675 15.805 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 129.945 -56.275 131.075 ;
        RECT -56.605 125.635 -56.275 125.965 ;
        RECT -56.605 124.275 -56.275 124.605 ;
        RECT -56.605 122.915 -56.275 123.245 ;
        RECT -56.605 121.555 -56.275 121.885 ;
        RECT -56.605 120.195 -56.275 120.525 ;
        RECT -56.605 118.835 -56.275 119.165 ;
        RECT -56.605 117.475 -56.275 117.805 ;
        RECT -56.605 116.115 -56.275 116.445 ;
        RECT -56.605 114.755 -56.275 115.085 ;
        RECT -56.605 113.395 -56.275 113.725 ;
        RECT -56.605 112.035 -56.275 112.365 ;
        RECT -56.605 110.675 -56.275 111.005 ;
        RECT -56.605 109.315 -56.275 109.645 ;
        RECT -56.605 107.955 -56.275 108.285 ;
        RECT -56.605 106.595 -56.275 106.925 ;
        RECT -56.605 105.235 -56.275 105.565 ;
        RECT -56.605 103.875 -56.275 104.205 ;
        RECT -56.605 102.515 -56.275 102.845 ;
        RECT -56.605 101.155 -56.275 101.485 ;
        RECT -56.605 99.795 -56.275 100.125 ;
        RECT -56.605 98.435 -56.275 98.765 ;
        RECT -56.605 97.075 -56.275 97.405 ;
        RECT -56.605 95.715 -56.275 96.045 ;
        RECT -56.605 94.355 -56.275 94.685 ;
        RECT -56.605 92.995 -56.275 93.325 ;
        RECT -56.605 91.635 -56.275 91.965 ;
        RECT -56.605 90.275 -56.275 90.605 ;
        RECT -56.605 88.915 -56.275 89.245 ;
        RECT -56.605 87.555 -56.275 87.885 ;
        RECT -56.605 86.195 -56.275 86.525 ;
        RECT -56.605 84.835 -56.275 85.165 ;
        RECT -56.605 83.475 -56.275 83.805 ;
        RECT -56.605 82.115 -56.275 82.445 ;
        RECT -56.605 80.755 -56.275 81.085 ;
        RECT -56.605 79.395 -56.275 79.725 ;
        RECT -56.605 78.035 -56.275 78.365 ;
        RECT -56.605 76.675 -56.275 77.005 ;
        RECT -56.605 75.315 -56.275 75.645 ;
        RECT -56.605 73.955 -56.275 74.285 ;
        RECT -56.605 71.64 -56.275 71.97 ;
        RECT -56.605 69.465 -56.275 69.795 ;
        RECT -56.605 68.615 -56.275 68.945 ;
        RECT -56.605 66.305 -56.275 66.635 ;
        RECT -56.605 65.455 -56.275 65.785 ;
        RECT -56.605 63.145 -56.275 63.475 ;
        RECT -56.605 62.295 -56.275 62.625 ;
        RECT -56.605 59.985 -56.275 60.315 ;
        RECT -56.605 59.135 -56.275 59.465 ;
        RECT -56.605 56.825 -56.275 57.155 ;
        RECT -56.605 55.975 -56.275 56.305 ;
        RECT -56.605 53.665 -56.275 53.995 ;
        RECT -56.605 52.815 -56.275 53.145 ;
        RECT -56.605 50.64 -56.275 50.97 ;
        RECT -56.605 48.115 -56.275 48.445 ;
        RECT -56.605 46.755 -56.275 47.085 ;
        RECT -56.605 45.395 -56.275 45.725 ;
        RECT -56.605 44.035 -56.275 44.365 ;
        RECT -56.605 42.675 -56.275 43.005 ;
        RECT -56.605 41.315 -56.275 41.645 ;
        RECT -56.605 39.955 -56.275 40.285 ;
        RECT -56.605 38.595 -56.275 38.925 ;
        RECT -56.605 37.235 -56.275 37.565 ;
        RECT -56.605 35.875 -56.275 36.205 ;
        RECT -56.605 34.515 -56.275 34.845 ;
        RECT -56.605 33.155 -56.275 33.485 ;
        RECT -56.605 31.795 -56.275 32.125 ;
        RECT -56.605 30.435 -56.275 30.765 ;
        RECT -56.605 29.075 -56.275 29.405 ;
        RECT -56.605 27.715 -56.275 28.045 ;
        RECT -56.605 26.355 -56.275 26.685 ;
        RECT -56.605 24.995 -56.275 25.325 ;
        RECT -56.605 23.635 -56.275 23.965 ;
        RECT -56.605 22.275 -56.275 22.605 ;
        RECT -56.605 20.915 -56.275 21.245 ;
        RECT -56.605 19.555 -56.275 19.885 ;
        RECT -56.605 18.195 -56.275 18.525 ;
        RECT -56.605 16.835 -56.275 17.165 ;
        RECT -56.605 15.475 -56.275 15.805 ;
        RECT -56.605 14.115 -56.275 14.445 ;
        RECT -56.605 12.755 -56.275 13.085 ;
        RECT -56.605 11.395 -56.275 11.725 ;
        RECT -56.605 10.035 -56.275 10.365 ;
        RECT -56.605 8.675 -56.275 9.005 ;
        RECT -56.605 7.315 -56.275 7.645 ;
        RECT -56.605 5.955 -56.275 6.285 ;
        RECT -56.605 4.595 -56.275 4.925 ;
        RECT -56.605 3.235 -56.275 3.565 ;
        RECT -56.605 1.875 -56.275 2.205 ;
        RECT -56.605 0.515 -56.275 0.845 ;
        RECT -56.605 -0.845 -56.275 -0.515 ;
        RECT -56.605 -2.205 -56.275 -1.875 ;
        RECT -56.605 -3.565 -56.275 -3.235 ;
        RECT -56.605 -4.925 -56.275 -4.595 ;
        RECT -56.605 -6.285 -56.275 -5.955 ;
        RECT -56.605 -7.645 -56.275 -7.315 ;
        RECT -56.605 -9.005 -56.275 -8.675 ;
        RECT -56.605 -10.365 -56.275 -10.035 ;
        RECT -56.605 -11.725 -56.275 -11.395 ;
        RECT -56.605 -13.085 -56.275 -12.755 ;
        RECT -56.605 -14.445 -56.275 -14.115 ;
        RECT -56.605 -15.805 -56.275 -15.475 ;
        RECT -56.605 -17.165 -56.275 -16.835 ;
        RECT -56.605 -18.525 -56.275 -18.195 ;
        RECT -56.605 -19.885 -56.275 -19.555 ;
        RECT -56.605 -21.245 -56.275 -20.915 ;
        RECT -56.605 -22.605 -56.275 -22.275 ;
        RECT -56.605 -23.965 -56.275 -23.635 ;
        RECT -56.605 -25.325 -56.275 -24.995 ;
        RECT -56.605 -26.685 -56.275 -26.355 ;
        RECT -56.605 -28.045 -56.275 -27.715 ;
        RECT -56.605 -29.405 -56.275 -29.075 ;
        RECT -56.605 -30.765 -56.275 -30.435 ;
        RECT -56.605 -32.125 -56.275 -31.795 ;
        RECT -56.605 -33.485 -56.275 -33.155 ;
        RECT -56.605 -34.845 -56.275 -34.515 ;
        RECT -56.605 -36.205 -56.275 -35.875 ;
        RECT -56.605 -37.565 -56.275 -37.235 ;
        RECT -56.605 -38.925 -56.275 -38.595 ;
        RECT -56.605 -40.285 -56.275 -39.955 ;
        RECT -56.605 -41.645 -56.275 -41.315 ;
        RECT -56.605 -43.005 -56.275 -42.675 ;
        RECT -56.605 -44.365 -56.275 -44.035 ;
        RECT -56.605 -45.725 -56.275 -45.395 ;
        RECT -56.605 -47.085 -56.275 -46.755 ;
        RECT -56.605 -48.445 -56.275 -48.115 ;
        RECT -56.605 -49.805 -56.275 -49.475 ;
        RECT -56.605 -51.165 -56.275 -50.835 ;
        RECT -56.605 -52.525 -56.275 -52.195 ;
        RECT -56.605 -53.885 -56.275 -53.555 ;
        RECT -56.605 -55.245 -56.275 -54.915 ;
        RECT -56.605 -56.605 -56.275 -56.275 ;
        RECT -56.605 -57.965 -56.275 -57.635 ;
        RECT -56.605 -59.325 -56.275 -58.995 ;
        RECT -56.605 -60.685 -56.275 -60.355 ;
        RECT -56.605 -62.045 -56.275 -61.715 ;
        RECT -56.605 -63.405 -56.275 -63.075 ;
        RECT -56.605 -64.765 -56.275 -64.435 ;
        RECT -56.605 -66.125 -56.275 -65.795 ;
        RECT -56.605 -67.485 -56.275 -67.155 ;
        RECT -56.605 -68.845 -56.275 -68.515 ;
        RECT -56.605 -71.565 -56.275 -71.235 ;
        RECT -56.605 -72.925 -56.275 -72.595 ;
        RECT -56.605 -74.285 -56.275 -73.955 ;
        RECT -56.605 -75.645 -56.275 -75.315 ;
        RECT -56.605 -77.005 -56.275 -76.675 ;
        RECT -56.605 -79.725 -56.275 -79.395 ;
        RECT -56.605 -82.445 -56.275 -82.115 ;
        RECT -56.605 -83.805 -56.275 -83.475 ;
        RECT -56.605 -85.165 -56.275 -84.835 ;
        RECT -56.605 -87.885 -56.275 -87.555 ;
        RECT -56.605 -89.245 -56.275 -88.915 ;
        RECT -56.6 -90.6 -56.28 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 -100.125 -56.275 -99.795 ;
        RECT -56.605 -101.485 -56.275 -101.155 ;
        RECT -56.605 -102.845 -56.275 -102.515 ;
        RECT -56.605 -104.205 -56.275 -103.875 ;
        RECT -56.605 -105.565 -56.275 -105.235 ;
        RECT -56.605 -106.925 -56.275 -106.595 ;
        RECT -56.605 -108.285 -56.275 -107.955 ;
        RECT -56.605 -109.645 -56.275 -109.315 ;
        RECT -56.605 -111.005 -56.275 -110.675 ;
        RECT -56.605 -112.365 -56.275 -112.035 ;
        RECT -56.605 -113.725 -56.275 -113.395 ;
        RECT -56.605 -115.085 -56.275 -114.755 ;
        RECT -56.605 -116.445 -56.275 -116.115 ;
        RECT -56.605 -117.805 -56.275 -117.475 ;
        RECT -56.605 -119.165 -56.275 -118.835 ;
        RECT -56.605 -120.525 -56.275 -120.195 ;
        RECT -56.605 -121.885 -56.275 -121.555 ;
        RECT -56.605 -123.245 -56.275 -122.915 ;
        RECT -56.605 -124.605 -56.275 -124.275 ;
        RECT -56.605 -125.965 -56.275 -125.635 ;
        RECT -56.605 -127.325 -56.275 -126.995 ;
        RECT -56.605 -128.685 -56.275 -128.355 ;
        RECT -56.605 -130.045 -56.275 -129.715 ;
        RECT -56.605 -131.405 -56.275 -131.075 ;
        RECT -56.605 -132.765 -56.275 -132.435 ;
        RECT -56.605 -134.125 -56.275 -133.795 ;
        RECT -56.605 -135.485 -56.275 -135.155 ;
        RECT -56.605 -136.845 -56.275 -136.515 ;
        RECT -56.605 -138.205 -56.275 -137.875 ;
        RECT -56.605 -139.565 -56.275 -139.235 ;
        RECT -56.605 -140.925 -56.275 -140.595 ;
        RECT -56.605 -142.285 -56.275 -141.955 ;
        RECT -56.605 -143.645 -56.275 -143.315 ;
        RECT -56.605 -145.005 -56.275 -144.675 ;
        RECT -56.605 -146.365 -56.275 -146.035 ;
        RECT -56.605 -148.215 -56.275 -147.885 ;
        RECT -56.605 -149.085 -56.275 -148.755 ;
        RECT -56.605 -150.445 -56.275 -150.115 ;
        RECT -56.605 -151.805 -56.275 -151.475 ;
        RECT -56.605 -153.165 -56.275 -152.835 ;
        RECT -56.605 -154.525 -56.275 -154.195 ;
        RECT -56.605 -157.245 -56.275 -156.915 ;
        RECT -56.605 -162.89 -56.275 -161.76 ;
        RECT -56.6 -163.005 -56.28 -99.795 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 129.945 -54.915 131.075 ;
        RECT -55.245 125.635 -54.915 125.965 ;
        RECT -55.245 124.275 -54.915 124.605 ;
        RECT -55.245 122.915 -54.915 123.245 ;
        RECT -55.245 121.555 -54.915 121.885 ;
        RECT -55.245 120.195 -54.915 120.525 ;
        RECT -55.245 118.835 -54.915 119.165 ;
        RECT -55.245 117.475 -54.915 117.805 ;
        RECT -55.245 116.115 -54.915 116.445 ;
        RECT -55.245 114.755 -54.915 115.085 ;
        RECT -55.245 113.395 -54.915 113.725 ;
        RECT -55.245 112.035 -54.915 112.365 ;
        RECT -55.245 110.675 -54.915 111.005 ;
        RECT -55.245 109.315 -54.915 109.645 ;
        RECT -55.245 107.955 -54.915 108.285 ;
        RECT -55.245 106.595 -54.915 106.925 ;
        RECT -55.245 105.235 -54.915 105.565 ;
        RECT -55.245 103.875 -54.915 104.205 ;
        RECT -55.245 102.515 -54.915 102.845 ;
        RECT -55.245 101.155 -54.915 101.485 ;
        RECT -55.245 99.795 -54.915 100.125 ;
        RECT -55.245 98.435 -54.915 98.765 ;
        RECT -55.245 97.075 -54.915 97.405 ;
        RECT -55.245 95.715 -54.915 96.045 ;
        RECT -55.245 94.355 -54.915 94.685 ;
        RECT -55.245 92.995 -54.915 93.325 ;
        RECT -55.245 91.635 -54.915 91.965 ;
        RECT -55.245 90.275 -54.915 90.605 ;
        RECT -55.245 88.915 -54.915 89.245 ;
        RECT -55.245 87.555 -54.915 87.885 ;
        RECT -55.245 86.195 -54.915 86.525 ;
        RECT -55.245 84.835 -54.915 85.165 ;
        RECT -55.245 83.475 -54.915 83.805 ;
        RECT -55.245 82.115 -54.915 82.445 ;
        RECT -55.245 80.755 -54.915 81.085 ;
        RECT -55.245 79.395 -54.915 79.725 ;
        RECT -55.245 78.035 -54.915 78.365 ;
        RECT -55.245 76.675 -54.915 77.005 ;
        RECT -55.245 75.315 -54.915 75.645 ;
        RECT -55.245 73.955 -54.915 74.285 ;
        RECT -55.245 71.64 -54.915 71.97 ;
        RECT -55.245 69.465 -54.915 69.795 ;
        RECT -55.245 68.615 -54.915 68.945 ;
        RECT -55.245 66.305 -54.915 66.635 ;
        RECT -55.245 65.455 -54.915 65.785 ;
        RECT -55.245 63.145 -54.915 63.475 ;
        RECT -55.245 62.295 -54.915 62.625 ;
        RECT -55.245 59.985 -54.915 60.315 ;
        RECT -55.245 59.135 -54.915 59.465 ;
        RECT -55.245 56.825 -54.915 57.155 ;
        RECT -55.245 55.975 -54.915 56.305 ;
        RECT -55.245 53.665 -54.915 53.995 ;
        RECT -55.245 52.815 -54.915 53.145 ;
        RECT -55.245 50.64 -54.915 50.97 ;
        RECT -55.245 48.115 -54.915 48.445 ;
        RECT -55.245 46.755 -54.915 47.085 ;
        RECT -55.245 45.395 -54.915 45.725 ;
        RECT -55.245 44.035 -54.915 44.365 ;
        RECT -55.245 42.675 -54.915 43.005 ;
        RECT -55.245 41.315 -54.915 41.645 ;
        RECT -55.245 39.955 -54.915 40.285 ;
        RECT -55.245 38.595 -54.915 38.925 ;
        RECT -55.24 38.595 -54.92 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 -11.725 -54.915 -11.395 ;
        RECT -55.245 -13.085 -54.915 -12.755 ;
        RECT -55.245 -14.445 -54.915 -14.115 ;
        RECT -55.245 -15.805 -54.915 -15.475 ;
        RECT -55.245 -17.165 -54.915 -16.835 ;
        RECT -55.245 -18.525 -54.915 -18.195 ;
        RECT -55.245 -19.885 -54.915 -19.555 ;
        RECT -55.245 -21.245 -54.915 -20.915 ;
        RECT -55.245 -22.605 -54.915 -22.275 ;
        RECT -55.245 -23.965 -54.915 -23.635 ;
        RECT -55.245 -25.325 -54.915 -24.995 ;
        RECT -55.245 -26.685 -54.915 -26.355 ;
        RECT -55.245 -28.045 -54.915 -27.715 ;
        RECT -55.245 -29.405 -54.915 -29.075 ;
        RECT -55.245 -30.765 -54.915 -30.435 ;
        RECT -55.245 -32.125 -54.915 -31.795 ;
        RECT -55.245 -33.485 -54.915 -33.155 ;
        RECT -55.245 -34.845 -54.915 -34.515 ;
        RECT -55.245 -36.205 -54.915 -35.875 ;
        RECT -55.245 -37.565 -54.915 -37.235 ;
        RECT -55.245 -38.925 -54.915 -38.595 ;
        RECT -55.245 -40.285 -54.915 -39.955 ;
        RECT -55.245 -41.645 -54.915 -41.315 ;
        RECT -55.245 -43.005 -54.915 -42.675 ;
        RECT -55.245 -44.365 -54.915 -44.035 ;
        RECT -55.245 -45.725 -54.915 -45.395 ;
        RECT -55.245 -47.085 -54.915 -46.755 ;
        RECT -55.245 -48.445 -54.915 -48.115 ;
        RECT -55.245 -49.805 -54.915 -49.475 ;
        RECT -55.245 -51.165 -54.915 -50.835 ;
        RECT -55.245 -52.525 -54.915 -52.195 ;
        RECT -55.245 -53.885 -54.915 -53.555 ;
        RECT -55.245 -55.245 -54.915 -54.915 ;
        RECT -55.245 -56.605 -54.915 -56.275 ;
        RECT -55.245 -57.965 -54.915 -57.635 ;
        RECT -55.245 -59.325 -54.915 -58.995 ;
        RECT -55.245 -60.685 -54.915 -60.355 ;
        RECT -55.245 -62.045 -54.915 -61.715 ;
        RECT -55.245 -63.405 -54.915 -63.075 ;
        RECT -55.245 -64.765 -54.915 -64.435 ;
        RECT -55.245 -66.125 -54.915 -65.795 ;
        RECT -55.245 -67.485 -54.915 -67.155 ;
        RECT -55.245 -68.845 -54.915 -68.515 ;
        RECT -55.245 -70.37 -54.915 -70.04 ;
        RECT -55.245 -71.565 -54.915 -71.235 ;
        RECT -55.245 -72.925 -54.915 -72.595 ;
        RECT -55.245 -74.285 -54.915 -73.955 ;
        RECT -55.245 -75.645 -54.915 -75.315 ;
        RECT -55.245 -77.005 -54.915 -76.675 ;
        RECT -55.245 -79.725 -54.915 -79.395 ;
        RECT -55.245 -80.91 -54.915 -80.58 ;
        RECT -55.245 -82.445 -54.915 -82.115 ;
        RECT -55.245 -83.805 -54.915 -83.475 ;
        RECT -55.245 -85.165 -54.915 -84.835 ;
        RECT -55.245 -87.885 -54.915 -87.555 ;
        RECT -55.245 -89.245 -54.915 -88.915 ;
        RECT -55.245 -93.325 -54.915 -92.995 ;
        RECT -55.245 -94.685 -54.915 -94.355 ;
        RECT -55.245 -96.045 -54.915 -95.715 ;
        RECT -55.245 -97.405 -54.915 -97.075 ;
        RECT -55.245 -98.765 -54.915 -98.435 ;
        RECT -55.245 -100.125 -54.915 -99.795 ;
        RECT -55.245 -101.485 -54.915 -101.155 ;
        RECT -55.245 -102.845 -54.915 -102.515 ;
        RECT -55.245 -104.205 -54.915 -103.875 ;
        RECT -55.245 -105.565 -54.915 -105.235 ;
        RECT -55.245 -106.925 -54.915 -106.595 ;
        RECT -55.245 -108.285 -54.915 -107.955 ;
        RECT -55.245 -109.645 -54.915 -109.315 ;
        RECT -55.245 -111.005 -54.915 -110.675 ;
        RECT -55.245 -112.365 -54.915 -112.035 ;
        RECT -55.245 -113.725 -54.915 -113.395 ;
        RECT -55.245 -115.085 -54.915 -114.755 ;
        RECT -55.245 -116.445 -54.915 -116.115 ;
        RECT -55.245 -117.805 -54.915 -117.475 ;
        RECT -55.245 -119.165 -54.915 -118.835 ;
        RECT -55.245 -120.525 -54.915 -120.195 ;
        RECT -55.245 -121.885 -54.915 -121.555 ;
        RECT -55.245 -123.245 -54.915 -122.915 ;
        RECT -55.245 -124.605 -54.915 -124.275 ;
        RECT -55.245 -125.965 -54.915 -125.635 ;
        RECT -55.245 -127.325 -54.915 -126.995 ;
        RECT -55.245 -128.685 -54.915 -128.355 ;
        RECT -55.245 -130.045 -54.915 -129.715 ;
        RECT -55.245 -131.405 -54.915 -131.075 ;
        RECT -55.245 -132.765 -54.915 -132.435 ;
        RECT -55.245 -134.125 -54.915 -133.795 ;
        RECT -55.245 -135.485 -54.915 -135.155 ;
        RECT -55.245 -136.845 -54.915 -136.515 ;
        RECT -55.245 -138.205 -54.915 -137.875 ;
        RECT -55.245 -139.565 -54.915 -139.235 ;
        RECT -55.245 -140.925 -54.915 -140.595 ;
        RECT -55.245 -142.285 -54.915 -141.955 ;
        RECT -55.245 -143.645 -54.915 -143.315 ;
        RECT -55.245 -145.005 -54.915 -144.675 ;
        RECT -55.245 -146.365 -54.915 -146.035 ;
        RECT -55.245 -148.215 -54.915 -147.885 ;
        RECT -55.245 -149.085 -54.915 -148.755 ;
        RECT -55.245 -150.445 -54.915 -150.115 ;
        RECT -55.245 -151.805 -54.915 -151.475 ;
        RECT -55.245 -153.165 -54.915 -152.835 ;
        RECT -55.245 -154.525 -54.915 -154.195 ;
        RECT -55.245 -157.245 -54.915 -156.915 ;
        RECT -55.245 -162.89 -54.915 -161.76 ;
        RECT -55.24 -163.005 -54.92 -11.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 129.945 -53.555 131.075 ;
        RECT -53.885 125.635 -53.555 125.965 ;
        RECT -53.885 124.275 -53.555 124.605 ;
        RECT -53.885 122.915 -53.555 123.245 ;
        RECT -53.885 121.555 -53.555 121.885 ;
        RECT -53.885 120.195 -53.555 120.525 ;
        RECT -53.885 118.835 -53.555 119.165 ;
        RECT -53.885 117.475 -53.555 117.805 ;
        RECT -53.885 116.115 -53.555 116.445 ;
        RECT -53.885 114.755 -53.555 115.085 ;
        RECT -53.885 113.395 -53.555 113.725 ;
        RECT -53.885 112.035 -53.555 112.365 ;
        RECT -53.885 110.675 -53.555 111.005 ;
        RECT -53.885 109.315 -53.555 109.645 ;
        RECT -53.885 107.955 -53.555 108.285 ;
        RECT -53.885 106.595 -53.555 106.925 ;
        RECT -53.885 105.235 -53.555 105.565 ;
        RECT -53.885 103.875 -53.555 104.205 ;
        RECT -53.885 102.515 -53.555 102.845 ;
        RECT -53.885 101.155 -53.555 101.485 ;
        RECT -53.885 99.795 -53.555 100.125 ;
        RECT -53.885 98.435 -53.555 98.765 ;
        RECT -53.885 97.075 -53.555 97.405 ;
        RECT -53.885 95.715 -53.555 96.045 ;
        RECT -53.885 94.355 -53.555 94.685 ;
        RECT -53.885 92.995 -53.555 93.325 ;
        RECT -53.885 91.635 -53.555 91.965 ;
        RECT -53.885 90.275 -53.555 90.605 ;
        RECT -53.885 88.915 -53.555 89.245 ;
        RECT -53.885 87.555 -53.555 87.885 ;
        RECT -53.885 86.195 -53.555 86.525 ;
        RECT -53.885 84.835 -53.555 85.165 ;
        RECT -53.885 83.475 -53.555 83.805 ;
        RECT -53.885 82.115 -53.555 82.445 ;
        RECT -53.885 80.755 -53.555 81.085 ;
        RECT -53.885 79.395 -53.555 79.725 ;
        RECT -53.885 78.035 -53.555 78.365 ;
        RECT -53.885 76.675 -53.555 77.005 ;
        RECT -53.885 75.315 -53.555 75.645 ;
        RECT -53.885 73.955 -53.555 74.285 ;
        RECT -53.88 73.28 -53.56 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 48.115 -53.555 48.445 ;
        RECT -53.885 46.755 -53.555 47.085 ;
        RECT -53.885 45.395 -53.555 45.725 ;
        RECT -53.885 44.035 -53.555 44.365 ;
        RECT -53.885 39.955 -53.555 40.285 ;
        RECT -53.885 38.595 -53.555 38.925 ;
        RECT -53.885 35.875 -53.555 36.205 ;
        RECT -53.885 34.515 -53.555 34.845 ;
        RECT -53.885 33.155 -53.555 33.485 ;
        RECT -53.885 31.795 -53.555 32.125 ;
        RECT -53.885 30.435 -53.555 30.765 ;
        RECT -53.885 29.075 -53.555 29.405 ;
        RECT -53.885 27.715 -53.555 28.045 ;
        RECT -53.885 26.355 -53.555 26.685 ;
        RECT -53.885 24.995 -53.555 25.325 ;
        RECT -53.885 23.635 -53.555 23.965 ;
        RECT -53.885 22.275 -53.555 22.605 ;
        RECT -53.885 20.915 -53.555 21.245 ;
        RECT -53.885 19.555 -53.555 19.885 ;
        RECT -53.885 18.195 -53.555 18.525 ;
        RECT -53.885 16.835 -53.555 17.165 ;
        RECT -53.885 15.475 -53.555 15.805 ;
        RECT -53.885 14.115 -53.555 14.445 ;
        RECT -53.885 12.755 -53.555 13.085 ;
        RECT -53.885 11.395 -53.555 11.725 ;
        RECT -53.885 10.035 -53.555 10.365 ;
        RECT -53.885 8.675 -53.555 9.005 ;
        RECT -53.885 7.315 -53.555 7.645 ;
        RECT -53.885 5.955 -53.555 6.285 ;
        RECT -53.885 4.595 -53.555 4.925 ;
        RECT -53.885 3.235 -53.555 3.565 ;
        RECT -53.885 1.875 -53.555 2.205 ;
        RECT -53.885 0.515 -53.555 0.845 ;
        RECT -53.885 -0.845 -53.555 -0.515 ;
        RECT -53.885 -2.205 -53.555 -1.875 ;
        RECT -53.885 -3.565 -53.555 -3.235 ;
        RECT -53.885 -4.925 -53.555 -4.595 ;
        RECT -53.885 -6.285 -53.555 -5.955 ;
        RECT -53.885 -7.645 -53.555 -7.315 ;
        RECT -53.885 -9.005 -53.555 -8.675 ;
        RECT -53.885 -10.365 -53.555 -10.035 ;
        RECT -53.885 -11.725 -53.555 -11.395 ;
        RECT -53.885 -13.085 -53.555 -12.755 ;
        RECT -53.885 -14.445 -53.555 -14.115 ;
        RECT -53.885 -15.805 -53.555 -15.475 ;
        RECT -53.885 -17.165 -53.555 -16.835 ;
        RECT -53.885 -18.525 -53.555 -18.195 ;
        RECT -53.885 -19.885 -53.555 -19.555 ;
        RECT -53.885 -21.245 -53.555 -20.915 ;
        RECT -53.885 -22.605 -53.555 -22.275 ;
        RECT -53.885 -23.965 -53.555 -23.635 ;
        RECT -53.885 -25.325 -53.555 -24.995 ;
        RECT -53.885 -26.685 -53.555 -26.355 ;
        RECT -53.885 -28.045 -53.555 -27.715 ;
        RECT -53.885 -29.405 -53.555 -29.075 ;
        RECT -53.885 -30.765 -53.555 -30.435 ;
        RECT -53.885 -32.125 -53.555 -31.795 ;
        RECT -53.885 -33.485 -53.555 -33.155 ;
        RECT -53.885 -34.845 -53.555 -34.515 ;
        RECT -53.885 -36.205 -53.555 -35.875 ;
        RECT -53.885 -37.565 -53.555 -37.235 ;
        RECT -53.885 -38.925 -53.555 -38.595 ;
        RECT -53.885 -40.285 -53.555 -39.955 ;
        RECT -53.885 -41.645 -53.555 -41.315 ;
        RECT -53.885 -43.005 -53.555 -42.675 ;
        RECT -53.885 -44.365 -53.555 -44.035 ;
        RECT -53.885 -45.725 -53.555 -45.395 ;
        RECT -53.885 -47.085 -53.555 -46.755 ;
        RECT -53.885 -48.445 -53.555 -48.115 ;
        RECT -53.885 -49.805 -53.555 -49.475 ;
        RECT -53.885 -51.165 -53.555 -50.835 ;
        RECT -53.885 -52.525 -53.555 -52.195 ;
        RECT -53.885 -53.885 -53.555 -53.555 ;
        RECT -53.885 -55.245 -53.555 -54.915 ;
        RECT -53.885 -56.605 -53.555 -56.275 ;
        RECT -53.885 -57.965 -53.555 -57.635 ;
        RECT -53.885 -59.325 -53.555 -58.995 ;
        RECT -53.885 -60.685 -53.555 -60.355 ;
        RECT -53.885 -62.045 -53.555 -61.715 ;
        RECT -53.885 -63.405 -53.555 -63.075 ;
        RECT -53.885 -64.765 -53.555 -64.435 ;
        RECT -53.885 -66.125 -53.555 -65.795 ;
        RECT -53.885 -67.485 -53.555 -67.155 ;
        RECT -53.885 -68.845 -53.555 -68.515 ;
        RECT -53.885 -70.37 -53.555 -70.04 ;
        RECT -53.885 -71.565 -53.555 -71.235 ;
        RECT -53.885 -72.925 -53.555 -72.595 ;
        RECT -53.885 -74.285 -53.555 -73.955 ;
        RECT -53.885 -75.645 -53.555 -75.315 ;
        RECT -53.885 -77.005 -53.555 -76.675 ;
        RECT -53.885 -79.725 -53.555 -79.395 ;
        RECT -53.885 -80.91 -53.555 -80.58 ;
        RECT -53.885 -82.445 -53.555 -82.115 ;
        RECT -53.885 -83.805 -53.555 -83.475 ;
        RECT -53.885 -85.165 -53.555 -84.835 ;
        RECT -53.885 -87.885 -53.555 -87.555 ;
        RECT -53.885 -89.245 -53.555 -88.915 ;
        RECT -53.88 -92.64 -53.56 49.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 -154.525 -53.555 -154.195 ;
        RECT -53.885 -157.245 -53.555 -156.915 ;
        RECT -53.885 -162.89 -53.555 -161.76 ;
        RECT -53.88 -163.005 -53.56 -152.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 129.945 -52.195 131.075 ;
        RECT -52.525 125.635 -52.195 125.965 ;
        RECT -52.525 124.275 -52.195 124.605 ;
        RECT -52.525 122.915 -52.195 123.245 ;
        RECT -52.525 121.555 -52.195 121.885 ;
        RECT -52.525 120.195 -52.195 120.525 ;
        RECT -52.525 118.835 -52.195 119.165 ;
        RECT -52.525 117.475 -52.195 117.805 ;
        RECT -52.525 116.115 -52.195 116.445 ;
        RECT -52.525 114.755 -52.195 115.085 ;
        RECT -52.525 113.395 -52.195 113.725 ;
        RECT -52.525 112.035 -52.195 112.365 ;
        RECT -52.525 110.675 -52.195 111.005 ;
        RECT -52.525 109.315 -52.195 109.645 ;
        RECT -52.525 107.955 -52.195 108.285 ;
        RECT -52.525 106.595 -52.195 106.925 ;
        RECT -52.525 105.235 -52.195 105.565 ;
        RECT -52.525 103.875 -52.195 104.205 ;
        RECT -52.525 102.515 -52.195 102.845 ;
        RECT -52.525 101.155 -52.195 101.485 ;
        RECT -52.525 99.795 -52.195 100.125 ;
        RECT -52.525 98.435 -52.195 98.765 ;
        RECT -52.525 97.075 -52.195 97.405 ;
        RECT -52.525 95.715 -52.195 96.045 ;
        RECT -52.525 94.355 -52.195 94.685 ;
        RECT -52.525 92.995 -52.195 93.325 ;
        RECT -52.525 91.635 -52.195 91.965 ;
        RECT -52.525 90.275 -52.195 90.605 ;
        RECT -52.525 88.915 -52.195 89.245 ;
        RECT -52.525 87.555 -52.195 87.885 ;
        RECT -52.525 86.195 -52.195 86.525 ;
        RECT -52.525 84.835 -52.195 85.165 ;
        RECT -52.525 83.475 -52.195 83.805 ;
        RECT -52.525 82.115 -52.195 82.445 ;
        RECT -52.525 80.755 -52.195 81.085 ;
        RECT -52.525 79.395 -52.195 79.725 ;
        RECT -52.525 78.035 -52.195 78.365 ;
        RECT -52.525 76.675 -52.195 77.005 ;
        RECT -52.525 75.315 -52.195 75.645 ;
        RECT -52.525 73.955 -52.195 74.285 ;
        RECT -52.52 73.28 -52.2 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 48.115 -52.195 48.445 ;
        RECT -52.525 46.755 -52.195 47.085 ;
        RECT -52.525 45.395 -52.195 45.725 ;
        RECT -52.525 44.035 -52.195 44.365 ;
        RECT -52.525 39.955 -52.195 40.285 ;
        RECT -52.525 38.595 -52.195 38.925 ;
        RECT -52.525 35.875 -52.195 36.205 ;
        RECT -52.525 34.515 -52.195 34.845 ;
        RECT -52.525 33.155 -52.195 33.485 ;
        RECT -52.525 31.795 -52.195 32.125 ;
        RECT -52.525 30.435 -52.195 30.765 ;
        RECT -52.525 29.075 -52.195 29.405 ;
        RECT -52.525 27.715 -52.195 28.045 ;
        RECT -52.525 26.355 -52.195 26.685 ;
        RECT -52.525 24.995 -52.195 25.325 ;
        RECT -52.525 23.635 -52.195 23.965 ;
        RECT -52.525 22.275 -52.195 22.605 ;
        RECT -52.525 20.915 -52.195 21.245 ;
        RECT -52.525 19.555 -52.195 19.885 ;
        RECT -52.525 18.195 -52.195 18.525 ;
        RECT -52.525 16.835 -52.195 17.165 ;
        RECT -52.525 15.475 -52.195 15.805 ;
        RECT -52.525 14.115 -52.195 14.445 ;
        RECT -52.525 12.755 -52.195 13.085 ;
        RECT -52.525 11.395 -52.195 11.725 ;
        RECT -52.525 10.035 -52.195 10.365 ;
        RECT -52.525 8.675 -52.195 9.005 ;
        RECT -52.525 7.315 -52.195 7.645 ;
        RECT -52.525 5.955 -52.195 6.285 ;
        RECT -52.525 4.595 -52.195 4.925 ;
        RECT -52.525 3.235 -52.195 3.565 ;
        RECT -52.525 1.875 -52.195 2.205 ;
        RECT -52.525 0.515 -52.195 0.845 ;
        RECT -52.525 -0.845 -52.195 -0.515 ;
        RECT -52.525 -2.205 -52.195 -1.875 ;
        RECT -52.525 -3.565 -52.195 -3.235 ;
        RECT -52.525 -4.925 -52.195 -4.595 ;
        RECT -52.525 -6.285 -52.195 -5.955 ;
        RECT -52.525 -7.645 -52.195 -7.315 ;
        RECT -52.525 -9.005 -52.195 -8.675 ;
        RECT -52.525 -10.365 -52.195 -10.035 ;
        RECT -52.525 -11.725 -52.195 -11.395 ;
        RECT -52.525 -13.085 -52.195 -12.755 ;
        RECT -52.525 -14.445 -52.195 -14.115 ;
        RECT -52.525 -15.805 -52.195 -15.475 ;
        RECT -52.525 -17.165 -52.195 -16.835 ;
        RECT -52.525 -18.525 -52.195 -18.195 ;
        RECT -52.525 -19.885 -52.195 -19.555 ;
        RECT -52.525 -21.245 -52.195 -20.915 ;
        RECT -52.525 -22.605 -52.195 -22.275 ;
        RECT -52.525 -25.325 -52.195 -24.995 ;
        RECT -52.525 -26.685 -52.195 -26.355 ;
        RECT -52.525 -28.045 -52.195 -27.715 ;
        RECT -52.525 -29.405 -52.195 -29.075 ;
        RECT -52.525 -30.765 -52.195 -30.435 ;
        RECT -52.525 -32.125 -52.195 -31.795 ;
        RECT -52.525 -33.485 -52.195 -33.155 ;
        RECT -52.525 -34.845 -52.195 -34.515 ;
        RECT -52.525 -36.205 -52.195 -35.875 ;
        RECT -52.525 -37.565 -52.195 -37.235 ;
        RECT -52.525 -38.925 -52.195 -38.595 ;
        RECT -52.525 -40.285 -52.195 -39.955 ;
        RECT -52.525 -41.645 -52.195 -41.315 ;
        RECT -52.525 -43.005 -52.195 -42.675 ;
        RECT -52.525 -44.365 -52.195 -44.035 ;
        RECT -52.525 -45.725 -52.195 -45.395 ;
        RECT -52.525 -47.085 -52.195 -46.755 ;
        RECT -52.525 -48.445 -52.195 -48.115 ;
        RECT -52.525 -49.805 -52.195 -49.475 ;
        RECT -52.525 -51.165 -52.195 -50.835 ;
        RECT -52.525 -52.525 -52.195 -52.195 ;
        RECT -52.525 -53.885 -52.195 -53.555 ;
        RECT -52.525 -55.245 -52.195 -54.915 ;
        RECT -52.525 -56.605 -52.195 -56.275 ;
        RECT -52.525 -57.965 -52.195 -57.635 ;
        RECT -52.525 -59.325 -52.195 -58.995 ;
        RECT -52.525 -60.685 -52.195 -60.355 ;
        RECT -52.525 -62.045 -52.195 -61.715 ;
        RECT -52.525 -63.405 -52.195 -63.075 ;
        RECT -52.525 -64.765 -52.195 -64.435 ;
        RECT -52.525 -66.125 -52.195 -65.795 ;
        RECT -52.525 -67.485 -52.195 -67.155 ;
        RECT -52.525 -68.845 -52.195 -68.515 ;
        RECT -52.525 -70.37 -52.195 -70.04 ;
        RECT -52.525 -71.565 -52.195 -71.235 ;
        RECT -52.525 -72.925 -52.195 -72.595 ;
        RECT -52.525 -74.285 -52.195 -73.955 ;
        RECT -52.525 -75.645 -52.195 -75.315 ;
        RECT -52.525 -77.005 -52.195 -76.675 ;
        RECT -52.525 -79.725 -52.195 -79.395 ;
        RECT -52.525 -80.91 -52.195 -80.58 ;
        RECT -52.525 -82.445 -52.195 -82.115 ;
        RECT -52.525 -83.805 -52.195 -83.475 ;
        RECT -52.525 -85.165 -52.195 -84.835 ;
        RECT -52.525 -87.885 -52.195 -87.555 ;
        RECT -52.525 -89.245 -52.195 -88.915 ;
        RECT -52.525 -91.965 -52.195 -91.635 ;
        RECT -52.525 -94.685 -52.195 -94.355 ;
        RECT -52.525 -96.045 -52.195 -95.715 ;
        RECT -52.525 -97.405 -52.195 -97.075 ;
        RECT -52.525 -98.765 -52.195 -98.435 ;
        RECT -52.525 -100.125 -52.195 -99.795 ;
        RECT -52.525 -101.485 -52.195 -101.155 ;
        RECT -52.525 -102.845 -52.195 -102.515 ;
        RECT -52.525 -104.205 -52.195 -103.875 ;
        RECT -52.525 -105.565 -52.195 -105.235 ;
        RECT -52.525 -106.925 -52.195 -106.595 ;
        RECT -52.525 -108.285 -52.195 -107.955 ;
        RECT -52.525 -109.645 -52.195 -109.315 ;
        RECT -52.525 -111.005 -52.195 -110.675 ;
        RECT -52.525 -112.365 -52.195 -112.035 ;
        RECT -52.525 -113.725 -52.195 -113.395 ;
        RECT -52.525 -115.085 -52.195 -114.755 ;
        RECT -52.525 -116.445 -52.195 -116.115 ;
        RECT -52.525 -117.805 -52.195 -117.475 ;
        RECT -52.525 -119.165 -52.195 -118.835 ;
        RECT -52.525 -120.525 -52.195 -120.195 ;
        RECT -52.525 -121.885 -52.195 -121.555 ;
        RECT -52.525 -123.245 -52.195 -122.915 ;
        RECT -52.525 -124.605 -52.195 -124.275 ;
        RECT -52.525 -125.965 -52.195 -125.635 ;
        RECT -52.525 -127.325 -52.195 -126.995 ;
        RECT -52.525 -128.685 -52.195 -128.355 ;
        RECT -52.525 -130.045 -52.195 -129.715 ;
        RECT -52.525 -131.405 -52.195 -131.075 ;
        RECT -52.525 -132.765 -52.195 -132.435 ;
        RECT -52.525 -134.125 -52.195 -133.795 ;
        RECT -52.525 -135.485 -52.195 -135.155 ;
        RECT -52.525 -136.845 -52.195 -136.515 ;
        RECT -52.525 -138.205 -52.195 -137.875 ;
        RECT -52.525 -139.565 -52.195 -139.235 ;
        RECT -52.525 -140.925 -52.195 -140.595 ;
        RECT -52.525 -142.285 -52.195 -141.955 ;
        RECT -52.525 -143.645 -52.195 -143.315 ;
        RECT -52.525 -145.005 -52.195 -144.675 ;
        RECT -52.525 -146.365 -52.195 -146.035 ;
        RECT -52.525 -148.215 -52.195 -147.885 ;
        RECT -52.525 -149.085 -52.195 -148.755 ;
        RECT -52.525 -150.445 -52.195 -150.115 ;
        RECT -52.525 -151.805 -52.195 -151.475 ;
        RECT -52.52 -151.805 -52.2 49.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 129.945 -50.835 131.075 ;
        RECT -51.165 125.635 -50.835 125.965 ;
        RECT -51.165 124.275 -50.835 124.605 ;
        RECT -51.165 122.915 -50.835 123.245 ;
        RECT -51.165 121.555 -50.835 121.885 ;
        RECT -51.165 120.195 -50.835 120.525 ;
        RECT -51.165 118.835 -50.835 119.165 ;
        RECT -51.165 117.475 -50.835 117.805 ;
        RECT -51.165 116.115 -50.835 116.445 ;
        RECT -51.165 114.755 -50.835 115.085 ;
        RECT -51.165 113.395 -50.835 113.725 ;
        RECT -51.165 112.035 -50.835 112.365 ;
        RECT -51.165 110.675 -50.835 111.005 ;
        RECT -51.165 109.315 -50.835 109.645 ;
        RECT -51.165 107.955 -50.835 108.285 ;
        RECT -51.165 106.595 -50.835 106.925 ;
        RECT -51.165 105.235 -50.835 105.565 ;
        RECT -51.165 103.875 -50.835 104.205 ;
        RECT -51.165 102.515 -50.835 102.845 ;
        RECT -51.165 101.155 -50.835 101.485 ;
        RECT -51.165 99.795 -50.835 100.125 ;
        RECT -51.165 98.435 -50.835 98.765 ;
        RECT -51.165 97.075 -50.835 97.405 ;
        RECT -51.165 95.715 -50.835 96.045 ;
        RECT -51.165 94.355 -50.835 94.685 ;
        RECT -51.165 92.995 -50.835 93.325 ;
        RECT -51.165 91.635 -50.835 91.965 ;
        RECT -51.165 90.275 -50.835 90.605 ;
        RECT -51.165 88.915 -50.835 89.245 ;
        RECT -51.165 87.555 -50.835 87.885 ;
        RECT -51.165 86.195 -50.835 86.525 ;
        RECT -51.165 84.835 -50.835 85.165 ;
        RECT -51.165 83.475 -50.835 83.805 ;
        RECT -51.165 82.115 -50.835 82.445 ;
        RECT -51.165 80.755 -50.835 81.085 ;
        RECT -51.165 79.395 -50.835 79.725 ;
        RECT -51.165 78.035 -50.835 78.365 ;
        RECT -51.165 76.675 -50.835 77.005 ;
        RECT -51.165 75.315 -50.835 75.645 ;
        RECT -51.165 73.955 -50.835 74.285 ;
        RECT -51.16 73.28 -50.84 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 19.555 -50.835 19.885 ;
        RECT -51.165 18.195 -50.835 18.525 ;
        RECT -51.165 16.835 -50.835 17.165 ;
        RECT -51.165 15.475 -50.835 15.805 ;
        RECT -51.165 14.115 -50.835 14.445 ;
        RECT -51.165 12.755 -50.835 13.085 ;
        RECT -51.165 11.395 -50.835 11.725 ;
        RECT -51.165 10.035 -50.835 10.365 ;
        RECT -51.165 8.675 -50.835 9.005 ;
        RECT -51.165 7.315 -50.835 7.645 ;
        RECT -51.165 5.955 -50.835 6.285 ;
        RECT -51.165 4.595 -50.835 4.925 ;
        RECT -51.165 3.235 -50.835 3.565 ;
        RECT -51.165 1.875 -50.835 2.205 ;
        RECT -51.165 0.515 -50.835 0.845 ;
        RECT -51.165 -0.845 -50.835 -0.515 ;
        RECT -51.165 -2.205 -50.835 -1.875 ;
        RECT -51.165 -3.565 -50.835 -3.235 ;
        RECT -51.165 -4.925 -50.835 -4.595 ;
        RECT -51.165 -6.285 -50.835 -5.955 ;
        RECT -51.165 -7.645 -50.835 -7.315 ;
        RECT -51.165 -9.005 -50.835 -8.675 ;
        RECT -51.165 -10.365 -50.835 -10.035 ;
        RECT -51.165 -11.725 -50.835 -11.395 ;
        RECT -51.165 -13.085 -50.835 -12.755 ;
        RECT -51.165 -14.445 -50.835 -14.115 ;
        RECT -51.165 -15.805 -50.835 -15.475 ;
        RECT -51.165 -17.165 -50.835 -16.835 ;
        RECT -51.165 -18.525 -50.835 -18.195 ;
        RECT -51.165 -19.885 -50.835 -19.555 ;
        RECT -51.165 -21.245 -50.835 -20.915 ;
        RECT -51.165 -22.605 -50.835 -22.275 ;
        RECT -51.165 -25.325 -50.835 -24.995 ;
        RECT -51.165 -26.685 -50.835 -26.355 ;
        RECT -51.165 -28.045 -50.835 -27.715 ;
        RECT -51.165 -29.405 -50.835 -29.075 ;
        RECT -51.165 -30.765 -50.835 -30.435 ;
        RECT -51.165 -32.125 -50.835 -31.795 ;
        RECT -51.165 -33.485 -50.835 -33.155 ;
        RECT -51.165 -34.845 -50.835 -34.515 ;
        RECT -51.165 -36.205 -50.835 -35.875 ;
        RECT -51.165 -37.565 -50.835 -37.235 ;
        RECT -51.165 -38.925 -50.835 -38.595 ;
        RECT -51.165 -40.285 -50.835 -39.955 ;
        RECT -51.165 -41.645 -50.835 -41.315 ;
        RECT -51.165 -43.005 -50.835 -42.675 ;
        RECT -51.165 -44.365 -50.835 -44.035 ;
        RECT -51.165 -45.725 -50.835 -45.395 ;
        RECT -51.165 -47.085 -50.835 -46.755 ;
        RECT -51.165 -48.445 -50.835 -48.115 ;
        RECT -51.165 -49.805 -50.835 -49.475 ;
        RECT -51.165 -51.165 -50.835 -50.835 ;
        RECT -51.165 -52.525 -50.835 -52.195 ;
        RECT -51.165 -53.885 -50.835 -53.555 ;
        RECT -51.165 -55.245 -50.835 -54.915 ;
        RECT -51.165 -56.605 -50.835 -56.275 ;
        RECT -51.165 -57.965 -50.835 -57.635 ;
        RECT -51.165 -59.325 -50.835 -58.995 ;
        RECT -51.165 -60.685 -50.835 -60.355 ;
        RECT -51.165 -62.045 -50.835 -61.715 ;
        RECT -51.165 -63.405 -50.835 -63.075 ;
        RECT -51.165 -64.765 -50.835 -64.435 ;
        RECT -51.165 -66.125 -50.835 -65.795 ;
        RECT -51.165 -67.485 -50.835 -67.155 ;
        RECT -51.165 -68.845 -50.835 -68.515 ;
        RECT -51.165 -70.37 -50.835 -70.04 ;
        RECT -51.165 -71.565 -50.835 -71.235 ;
        RECT -51.165 -72.925 -50.835 -72.595 ;
        RECT -51.165 -74.285 -50.835 -73.955 ;
        RECT -51.165 -75.645 -50.835 -75.315 ;
        RECT -51.165 -77.005 -50.835 -76.675 ;
        RECT -51.165 -79.725 -50.835 -79.395 ;
        RECT -51.165 -80.91 -50.835 -80.58 ;
        RECT -51.165 -82.445 -50.835 -82.115 ;
        RECT -51.165 -83.805 -50.835 -83.475 ;
        RECT -51.165 -85.165 -50.835 -84.835 ;
        RECT -51.165 -87.885 -50.835 -87.555 ;
        RECT -51.165 -89.245 -50.835 -88.915 ;
        RECT -51.165 -91.965 -50.835 -91.635 ;
        RECT -51.165 -94.685 -50.835 -94.355 ;
        RECT -51.165 -96.045 -50.835 -95.715 ;
        RECT -51.165 -97.405 -50.835 -97.075 ;
        RECT -51.165 -98.765 -50.835 -98.435 ;
        RECT -51.165 -100.125 -50.835 -99.795 ;
        RECT -51.165 -101.485 -50.835 -101.155 ;
        RECT -51.165 -102.845 -50.835 -102.515 ;
        RECT -51.165 -104.205 -50.835 -103.875 ;
        RECT -51.165 -105.565 -50.835 -105.235 ;
        RECT -51.165 -106.925 -50.835 -106.595 ;
        RECT -51.165 -108.285 -50.835 -107.955 ;
        RECT -51.165 -109.645 -50.835 -109.315 ;
        RECT -51.165 -111.005 -50.835 -110.675 ;
        RECT -51.165 -112.365 -50.835 -112.035 ;
        RECT -51.165 -113.725 -50.835 -113.395 ;
        RECT -51.165 -115.085 -50.835 -114.755 ;
        RECT -51.165 -116.445 -50.835 -116.115 ;
        RECT -51.165 -117.805 -50.835 -117.475 ;
        RECT -51.165 -119.165 -50.835 -118.835 ;
        RECT -51.165 -120.525 -50.835 -120.195 ;
        RECT -51.165 -121.885 -50.835 -121.555 ;
        RECT -51.165 -123.245 -50.835 -122.915 ;
        RECT -51.165 -124.605 -50.835 -124.275 ;
        RECT -51.165 -125.965 -50.835 -125.635 ;
        RECT -51.165 -127.325 -50.835 -126.995 ;
        RECT -51.165 -128.685 -50.835 -128.355 ;
        RECT -51.165 -130.045 -50.835 -129.715 ;
        RECT -51.165 -131.405 -50.835 -131.075 ;
        RECT -51.165 -132.765 -50.835 -132.435 ;
        RECT -51.165 -134.125 -50.835 -133.795 ;
        RECT -51.165 -135.485 -50.835 -135.155 ;
        RECT -51.165 -136.845 -50.835 -136.515 ;
        RECT -51.165 -138.205 -50.835 -137.875 ;
        RECT -51.165 -139.565 -50.835 -139.235 ;
        RECT -51.165 -140.925 -50.835 -140.595 ;
        RECT -51.165 -142.285 -50.835 -141.955 ;
        RECT -51.165 -143.645 -50.835 -143.315 ;
        RECT -51.165 -145.005 -50.835 -144.675 ;
        RECT -51.165 -146.365 -50.835 -146.035 ;
        RECT -51.165 -148.215 -50.835 -147.885 ;
        RECT -51.165 -149.085 -50.835 -148.755 ;
        RECT -51.165 -150.445 -50.835 -150.115 ;
        RECT -51.165 -154.525 -50.835 -154.195 ;
        RECT -51.165 -157.245 -50.835 -156.915 ;
        RECT -51.165 -162.89 -50.835 -161.76 ;
        RECT -51.16 -163.005 -50.84 49.12 ;
        RECT -51.165 48.115 -50.835 48.445 ;
        RECT -51.165 46.755 -50.835 47.085 ;
        RECT -51.165 45.395 -50.835 45.725 ;
        RECT -51.165 44.035 -50.835 44.365 ;
        RECT -51.165 39.955 -50.835 40.285 ;
        RECT -51.165 38.595 -50.835 38.925 ;
        RECT -51.165 35.875 -50.835 36.205 ;
        RECT -51.165 34.515 -50.835 34.845 ;
        RECT -51.165 33.155 -50.835 33.485 ;
        RECT -51.165 31.795 -50.835 32.125 ;
        RECT -51.165 30.435 -50.835 30.765 ;
        RECT -51.165 29.075 -50.835 29.405 ;
        RECT -51.165 27.715 -50.835 28.045 ;
        RECT -51.165 26.355 -50.835 26.685 ;
        RECT -51.165 24.995 -50.835 25.325 ;
        RECT -51.165 23.635 -50.835 23.965 ;
        RECT -51.165 22.275 -50.835 22.605 ;
        RECT -51.165 20.915 -50.835 21.245 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.405 129.945 -63.075 131.075 ;
        RECT -63.405 125.635 -63.075 125.965 ;
        RECT -63.405 124.275 -63.075 124.605 ;
        RECT -63.405 122.915 -63.075 123.245 ;
        RECT -63.405 121.555 -63.075 121.885 ;
        RECT -63.405 120.195 -63.075 120.525 ;
        RECT -63.405 118.835 -63.075 119.165 ;
        RECT -63.405 117.475 -63.075 117.805 ;
        RECT -63.405 116.115 -63.075 116.445 ;
        RECT -63.405 114.755 -63.075 115.085 ;
        RECT -63.405 113.395 -63.075 113.725 ;
        RECT -63.405 112.035 -63.075 112.365 ;
        RECT -63.405 110.675 -63.075 111.005 ;
        RECT -63.405 109.315 -63.075 109.645 ;
        RECT -63.405 107.955 -63.075 108.285 ;
        RECT -63.405 106.595 -63.075 106.925 ;
        RECT -63.405 105.235 -63.075 105.565 ;
        RECT -63.405 103.875 -63.075 104.205 ;
        RECT -63.405 102.515 -63.075 102.845 ;
        RECT -63.405 101.155 -63.075 101.485 ;
        RECT -63.405 99.795 -63.075 100.125 ;
        RECT -63.405 98.435 -63.075 98.765 ;
        RECT -63.405 97.075 -63.075 97.405 ;
        RECT -63.405 95.715 -63.075 96.045 ;
        RECT -63.405 94.355 -63.075 94.685 ;
        RECT -63.405 92.995 -63.075 93.325 ;
        RECT -63.405 91.635 -63.075 91.965 ;
        RECT -63.405 90.275 -63.075 90.605 ;
        RECT -63.405 88.915 -63.075 89.245 ;
        RECT -63.405 87.555 -63.075 87.885 ;
        RECT -63.405 86.195 -63.075 86.525 ;
        RECT -63.405 84.835 -63.075 85.165 ;
        RECT -63.405 83.475 -63.075 83.805 ;
        RECT -63.405 82.115 -63.075 82.445 ;
        RECT -63.405 80.755 -63.075 81.085 ;
        RECT -63.405 79.395 -63.075 79.725 ;
        RECT -63.405 78.035 -63.075 78.365 ;
        RECT -63.405 76.675 -63.075 77.005 ;
        RECT -63.405 75.315 -63.075 75.645 ;
        RECT -63.405 73.955 -63.075 74.285 ;
        RECT -63.405 72.595 -63.075 72.925 ;
        RECT -63.405 71.235 -63.075 71.565 ;
        RECT -63.405 69.875 -63.075 70.205 ;
        RECT -63.405 68.515 -63.075 68.845 ;
        RECT -63.405 67.155 -63.075 67.485 ;
        RECT -63.405 65.795 -63.075 66.125 ;
        RECT -63.405 64.435 -63.075 64.765 ;
        RECT -63.405 63.075 -63.075 63.405 ;
        RECT -63.405 61.715 -63.075 62.045 ;
        RECT -63.405 60.355 -63.075 60.685 ;
        RECT -63.405 58.995 -63.075 59.325 ;
        RECT -63.405 57.635 -63.075 57.965 ;
        RECT -63.405 56.275 -63.075 56.605 ;
        RECT -63.405 54.915 -63.075 55.245 ;
        RECT -63.405 53.555 -63.075 53.885 ;
        RECT -63.405 52.195 -63.075 52.525 ;
        RECT -63.405 50.835 -63.075 51.165 ;
        RECT -63.405 49.475 -63.075 49.805 ;
        RECT -63.405 48.115 -63.075 48.445 ;
        RECT -63.405 46.755 -63.075 47.085 ;
        RECT -63.405 45.395 -63.075 45.725 ;
        RECT -63.405 44.035 -63.075 44.365 ;
        RECT -63.405 42.675 -63.075 43.005 ;
        RECT -63.405 41.315 -63.075 41.645 ;
        RECT -63.405 39.955 -63.075 40.285 ;
        RECT -63.405 38.595 -63.075 38.925 ;
        RECT -63.405 37.235 -63.075 37.565 ;
        RECT -63.405 35.875 -63.075 36.205 ;
        RECT -63.405 34.515 -63.075 34.845 ;
        RECT -63.405 33.155 -63.075 33.485 ;
        RECT -63.405 31.795 -63.075 32.125 ;
        RECT -63.405 30.435 -63.075 30.765 ;
        RECT -63.405 29.075 -63.075 29.405 ;
        RECT -63.405 27.715 -63.075 28.045 ;
        RECT -63.405 26.355 -63.075 26.685 ;
        RECT -63.405 24.995 -63.075 25.325 ;
        RECT -63.405 23.635 -63.075 23.965 ;
        RECT -63.405 22.275 -63.075 22.605 ;
        RECT -63.405 20.915 -63.075 21.245 ;
        RECT -63.405 19.555 -63.075 19.885 ;
        RECT -63.405 18.195 -63.075 18.525 ;
        RECT -63.405 16.835 -63.075 17.165 ;
        RECT -63.405 15.475 -63.075 15.805 ;
        RECT -63.405 14.115 -63.075 14.445 ;
        RECT -63.405 12.755 -63.075 13.085 ;
        RECT -63.405 11.395 -63.075 11.725 ;
        RECT -63.405 10.035 -63.075 10.365 ;
        RECT -63.405 8.675 -63.075 9.005 ;
        RECT -63.405 7.315 -63.075 7.645 ;
        RECT -63.405 5.955 -63.075 6.285 ;
        RECT -63.405 4.595 -63.075 4.925 ;
        RECT -63.405 3.235 -63.075 3.565 ;
        RECT -63.405 1.875 -63.075 2.205 ;
        RECT -63.405 0.515 -63.075 0.845 ;
        RECT -63.405 -0.845 -63.075 -0.515 ;
        RECT -63.405 -2.205 -63.075 -1.875 ;
        RECT -63.405 -3.565 -63.075 -3.235 ;
        RECT -63.405 -4.925 -63.075 -4.595 ;
        RECT -63.405 -6.285 -63.075 -5.955 ;
        RECT -63.405 -7.645 -63.075 -7.315 ;
        RECT -63.405 -9.005 -63.075 -8.675 ;
        RECT -63.405 -10.365 -63.075 -10.035 ;
        RECT -63.405 -11.725 -63.075 -11.395 ;
        RECT -63.405 -13.085 -63.075 -12.755 ;
        RECT -63.405 -14.445 -63.075 -14.115 ;
        RECT -63.405 -15.805 -63.075 -15.475 ;
        RECT -63.405 -17.165 -63.075 -16.835 ;
        RECT -63.405 -18.525 -63.075 -18.195 ;
        RECT -63.405 -19.885 -63.075 -19.555 ;
        RECT -63.405 -21.245 -63.075 -20.915 ;
        RECT -63.405 -22.605 -63.075 -22.275 ;
        RECT -63.405 -23.965 -63.075 -23.635 ;
        RECT -63.405 -25.325 -63.075 -24.995 ;
        RECT -63.405 -26.685 -63.075 -26.355 ;
        RECT -63.405 -28.045 -63.075 -27.715 ;
        RECT -63.405 -29.405 -63.075 -29.075 ;
        RECT -63.405 -30.765 -63.075 -30.435 ;
        RECT -63.405 -32.125 -63.075 -31.795 ;
        RECT -63.405 -33.485 -63.075 -33.155 ;
        RECT -63.405 -34.845 -63.075 -34.515 ;
        RECT -63.405 -36.205 -63.075 -35.875 ;
        RECT -63.405 -37.565 -63.075 -37.235 ;
        RECT -63.405 -38.925 -63.075 -38.595 ;
        RECT -63.405 -40.285 -63.075 -39.955 ;
        RECT -63.405 -41.645 -63.075 -41.315 ;
        RECT -63.405 -43.005 -63.075 -42.675 ;
        RECT -63.405 -44.365 -63.075 -44.035 ;
        RECT -63.405 -45.725 -63.075 -45.395 ;
        RECT -63.405 -47.085 -63.075 -46.755 ;
        RECT -63.405 -48.445 -63.075 -48.115 ;
        RECT -63.405 -49.805 -63.075 -49.475 ;
        RECT -63.405 -51.165 -63.075 -50.835 ;
        RECT -63.405 -52.525 -63.075 -52.195 ;
        RECT -63.405 -53.885 -63.075 -53.555 ;
        RECT -63.405 -55.245 -63.075 -54.915 ;
        RECT -63.405 -56.605 -63.075 -56.275 ;
        RECT -63.405 -57.965 -63.075 -57.635 ;
        RECT -63.405 -59.325 -63.075 -58.995 ;
        RECT -63.405 -60.685 -63.075 -60.355 ;
        RECT -63.405 -62.045 -63.075 -61.715 ;
        RECT -63.405 -63.405 -63.075 -63.075 ;
        RECT -63.405 -64.765 -63.075 -64.435 ;
        RECT -63.405 -66.125 -63.075 -65.795 ;
        RECT -63.405 -67.485 -63.075 -67.155 ;
        RECT -63.405 -68.845 -63.075 -68.515 ;
        RECT -63.405 -70.205 -63.075 -69.875 ;
        RECT -63.405 -71.565 -63.075 -71.235 ;
        RECT -63.405 -72.925 -63.075 -72.595 ;
        RECT -63.405 -74.285 -63.075 -73.955 ;
        RECT -63.405 -75.645 -63.075 -75.315 ;
        RECT -63.405 -77.005 -63.075 -76.675 ;
        RECT -63.405 -78.365 -63.075 -78.035 ;
        RECT -63.405 -79.725 -63.075 -79.395 ;
        RECT -63.405 -81.085 -63.075 -80.755 ;
        RECT -63.405 -82.445 -63.075 -82.115 ;
        RECT -63.405 -83.805 -63.075 -83.475 ;
        RECT -63.405 -85.165 -63.075 -84.835 ;
        RECT -63.405 -86.525 -63.075 -86.195 ;
        RECT -63.405 -87.885 -63.075 -87.555 ;
        RECT -63.405 -89.245 -63.075 -88.915 ;
        RECT -63.405 -90.605 -63.075 -90.275 ;
        RECT -63.405 -91.965 -63.075 -91.635 ;
        RECT -63.405 -93.325 -63.075 -92.995 ;
        RECT -63.405 -94.685 -63.075 -94.355 ;
        RECT -63.405 -96.045 -63.075 -95.715 ;
        RECT -63.405 -97.405 -63.075 -97.075 ;
        RECT -63.405 -98.765 -63.075 -98.435 ;
        RECT -63.405 -100.125 -63.075 -99.795 ;
        RECT -63.405 -101.485 -63.075 -101.155 ;
        RECT -63.405 -102.845 -63.075 -102.515 ;
        RECT -63.405 -104.205 -63.075 -103.875 ;
        RECT -63.405 -105.565 -63.075 -105.235 ;
        RECT -63.405 -106.925 -63.075 -106.595 ;
        RECT -63.405 -108.285 -63.075 -107.955 ;
        RECT -63.405 -109.645 -63.075 -109.315 ;
        RECT -63.405 -111.005 -63.075 -110.675 ;
        RECT -63.405 -112.365 -63.075 -112.035 ;
        RECT -63.405 -113.725 -63.075 -113.395 ;
        RECT -63.405 -115.085 -63.075 -114.755 ;
        RECT -63.405 -116.445 -63.075 -116.115 ;
        RECT -63.405 -117.805 -63.075 -117.475 ;
        RECT -63.405 -119.165 -63.075 -118.835 ;
        RECT -63.405 -120.525 -63.075 -120.195 ;
        RECT -63.405 -121.885 -63.075 -121.555 ;
        RECT -63.405 -123.245 -63.075 -122.915 ;
        RECT -63.405 -124.605 -63.075 -124.275 ;
        RECT -63.405 -125.965 -63.075 -125.635 ;
        RECT -63.405 -127.325 -63.075 -126.995 ;
        RECT -63.405 -128.685 -63.075 -128.355 ;
        RECT -63.405 -130.045 -63.075 -129.715 ;
        RECT -63.405 -131.405 -63.075 -131.075 ;
        RECT -63.405 -132.765 -63.075 -132.435 ;
        RECT -63.405 -134.125 -63.075 -133.795 ;
        RECT -63.405 -135.485 -63.075 -135.155 ;
        RECT -63.405 -136.845 -63.075 -136.515 ;
        RECT -63.405 -138.205 -63.075 -137.875 ;
        RECT -63.405 -139.565 -63.075 -139.235 ;
        RECT -63.405 -140.925 -63.075 -140.595 ;
        RECT -63.405 -142.285 -63.075 -141.955 ;
        RECT -63.405 -143.645 -63.075 -143.315 ;
        RECT -63.405 -145.005 -63.075 -144.675 ;
        RECT -63.405 -146.365 -63.075 -146.035 ;
        RECT -63.405 -148.215 -63.075 -147.885 ;
        RECT -63.405 -149.085 -63.075 -148.755 ;
        RECT -63.405 -150.445 -63.075 -150.115 ;
        RECT -63.405 -153.165 -63.075 -152.835 ;
        RECT -63.405 -154.525 -63.075 -154.195 ;
        RECT -63.405 -157.245 -63.075 -156.915 ;
        RECT -63.405 -162.89 -63.075 -161.76 ;
        RECT -63.4 -163.005 -63.08 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.045 129.945 -61.715 131.075 ;
        RECT -62.045 125.635 -61.715 125.965 ;
        RECT -62.045 124.275 -61.715 124.605 ;
        RECT -62.045 122.915 -61.715 123.245 ;
        RECT -62.045 121.555 -61.715 121.885 ;
        RECT -62.045 120.195 -61.715 120.525 ;
        RECT -62.045 118.835 -61.715 119.165 ;
        RECT -62.045 117.475 -61.715 117.805 ;
        RECT -62.045 116.115 -61.715 116.445 ;
        RECT -62.045 114.755 -61.715 115.085 ;
        RECT -62.045 113.395 -61.715 113.725 ;
        RECT -62.045 112.035 -61.715 112.365 ;
        RECT -62.045 110.675 -61.715 111.005 ;
        RECT -62.045 109.315 -61.715 109.645 ;
        RECT -62.045 107.955 -61.715 108.285 ;
        RECT -62.045 106.595 -61.715 106.925 ;
        RECT -62.045 105.235 -61.715 105.565 ;
        RECT -62.045 103.875 -61.715 104.205 ;
        RECT -62.045 102.515 -61.715 102.845 ;
        RECT -62.045 101.155 -61.715 101.485 ;
        RECT -62.045 99.795 -61.715 100.125 ;
        RECT -62.045 98.435 -61.715 98.765 ;
        RECT -62.045 97.075 -61.715 97.405 ;
        RECT -62.045 95.715 -61.715 96.045 ;
        RECT -62.045 94.355 -61.715 94.685 ;
        RECT -62.045 92.995 -61.715 93.325 ;
        RECT -62.045 91.635 -61.715 91.965 ;
        RECT -62.045 90.275 -61.715 90.605 ;
        RECT -62.045 88.915 -61.715 89.245 ;
        RECT -62.045 87.555 -61.715 87.885 ;
        RECT -62.045 86.195 -61.715 86.525 ;
        RECT -62.045 84.835 -61.715 85.165 ;
        RECT -62.045 83.475 -61.715 83.805 ;
        RECT -62.045 82.115 -61.715 82.445 ;
        RECT -62.045 80.755 -61.715 81.085 ;
        RECT -62.045 79.395 -61.715 79.725 ;
        RECT -62.045 78.035 -61.715 78.365 ;
        RECT -62.045 76.675 -61.715 77.005 ;
        RECT -62.045 75.315 -61.715 75.645 ;
        RECT -62.045 73.955 -61.715 74.285 ;
        RECT -62.045 72.595 -61.715 72.925 ;
        RECT -62.045 71.235 -61.715 71.565 ;
        RECT -62.045 69.875 -61.715 70.205 ;
        RECT -62.045 68.515 -61.715 68.845 ;
        RECT -62.045 67.155 -61.715 67.485 ;
        RECT -62.045 65.795 -61.715 66.125 ;
        RECT -62.045 64.435 -61.715 64.765 ;
        RECT -62.045 63.075 -61.715 63.405 ;
        RECT -62.045 61.715 -61.715 62.045 ;
        RECT -62.045 60.355 -61.715 60.685 ;
        RECT -62.045 58.995 -61.715 59.325 ;
        RECT -62.045 57.635 -61.715 57.965 ;
        RECT -62.045 56.275 -61.715 56.605 ;
        RECT -62.045 54.915 -61.715 55.245 ;
        RECT -62.045 53.555 -61.715 53.885 ;
        RECT -62.045 52.195 -61.715 52.525 ;
        RECT -62.045 50.835 -61.715 51.165 ;
        RECT -62.045 49.475 -61.715 49.805 ;
        RECT -62.045 48.115 -61.715 48.445 ;
        RECT -62.045 46.755 -61.715 47.085 ;
        RECT -62.045 45.395 -61.715 45.725 ;
        RECT -62.045 44.035 -61.715 44.365 ;
        RECT -62.045 42.675 -61.715 43.005 ;
        RECT -62.045 41.315 -61.715 41.645 ;
        RECT -62.045 39.955 -61.715 40.285 ;
        RECT -62.045 38.595 -61.715 38.925 ;
        RECT -62.045 37.235 -61.715 37.565 ;
        RECT -62.045 35.875 -61.715 36.205 ;
        RECT -62.045 34.515 -61.715 34.845 ;
        RECT -62.045 33.155 -61.715 33.485 ;
        RECT -62.045 31.795 -61.715 32.125 ;
        RECT -62.045 30.435 -61.715 30.765 ;
        RECT -62.045 29.075 -61.715 29.405 ;
        RECT -62.045 27.715 -61.715 28.045 ;
        RECT -62.045 26.355 -61.715 26.685 ;
        RECT -62.045 24.995 -61.715 25.325 ;
        RECT -62.045 23.635 -61.715 23.965 ;
        RECT -62.045 22.275 -61.715 22.605 ;
        RECT -62.045 20.915 -61.715 21.245 ;
        RECT -62.045 19.555 -61.715 19.885 ;
        RECT -62.045 18.195 -61.715 18.525 ;
        RECT -62.045 16.835 -61.715 17.165 ;
        RECT -62.045 15.475 -61.715 15.805 ;
        RECT -62.045 14.115 -61.715 14.445 ;
        RECT -62.045 12.755 -61.715 13.085 ;
        RECT -62.045 11.395 -61.715 11.725 ;
        RECT -62.045 10.035 -61.715 10.365 ;
        RECT -62.045 8.675 -61.715 9.005 ;
        RECT -62.045 7.315 -61.715 7.645 ;
        RECT -62.045 5.955 -61.715 6.285 ;
        RECT -62.045 4.595 -61.715 4.925 ;
        RECT -62.045 3.235 -61.715 3.565 ;
        RECT -62.045 1.875 -61.715 2.205 ;
        RECT -62.045 0.515 -61.715 0.845 ;
        RECT -62.045 -0.845 -61.715 -0.515 ;
        RECT -62.045 -2.205 -61.715 -1.875 ;
        RECT -62.045 -3.565 -61.715 -3.235 ;
        RECT -62.045 -4.925 -61.715 -4.595 ;
        RECT -62.045 -6.285 -61.715 -5.955 ;
        RECT -62.045 -7.645 -61.715 -7.315 ;
        RECT -62.045 -9.005 -61.715 -8.675 ;
        RECT -62.045 -10.365 -61.715 -10.035 ;
        RECT -62.045 -11.725 -61.715 -11.395 ;
        RECT -62.045 -13.085 -61.715 -12.755 ;
        RECT -62.045 -14.445 -61.715 -14.115 ;
        RECT -62.045 -15.805 -61.715 -15.475 ;
        RECT -62.045 -17.165 -61.715 -16.835 ;
        RECT -62.045 -18.525 -61.715 -18.195 ;
        RECT -62.045 -19.885 -61.715 -19.555 ;
        RECT -62.045 -21.245 -61.715 -20.915 ;
        RECT -62.045 -22.605 -61.715 -22.275 ;
        RECT -62.045 -23.965 -61.715 -23.635 ;
        RECT -62.045 -25.325 -61.715 -24.995 ;
        RECT -62.045 -26.685 -61.715 -26.355 ;
        RECT -62.045 -28.045 -61.715 -27.715 ;
        RECT -62.045 -29.405 -61.715 -29.075 ;
        RECT -62.045 -30.765 -61.715 -30.435 ;
        RECT -62.045 -32.125 -61.715 -31.795 ;
        RECT -62.045 -33.485 -61.715 -33.155 ;
        RECT -62.045 -34.845 -61.715 -34.515 ;
        RECT -62.045 -36.205 -61.715 -35.875 ;
        RECT -62.045 -37.565 -61.715 -37.235 ;
        RECT -62.045 -38.925 -61.715 -38.595 ;
        RECT -62.045 -40.285 -61.715 -39.955 ;
        RECT -62.045 -41.645 -61.715 -41.315 ;
        RECT -62.045 -43.005 -61.715 -42.675 ;
        RECT -62.045 -44.365 -61.715 -44.035 ;
        RECT -62.045 -45.725 -61.715 -45.395 ;
        RECT -62.045 -47.085 -61.715 -46.755 ;
        RECT -62.045 -48.445 -61.715 -48.115 ;
        RECT -62.045 -49.805 -61.715 -49.475 ;
        RECT -62.045 -51.165 -61.715 -50.835 ;
        RECT -62.045 -52.525 -61.715 -52.195 ;
        RECT -62.045 -53.885 -61.715 -53.555 ;
        RECT -62.045 -55.245 -61.715 -54.915 ;
        RECT -62.045 -56.605 -61.715 -56.275 ;
        RECT -62.045 -57.965 -61.715 -57.635 ;
        RECT -62.045 -59.325 -61.715 -58.995 ;
        RECT -62.045 -60.685 -61.715 -60.355 ;
        RECT -62.045 -62.045 -61.715 -61.715 ;
        RECT -62.045 -63.405 -61.715 -63.075 ;
        RECT -62.045 -64.765 -61.715 -64.435 ;
        RECT -62.045 -66.125 -61.715 -65.795 ;
        RECT -62.045 -67.485 -61.715 -67.155 ;
        RECT -62.045 -68.845 -61.715 -68.515 ;
        RECT -62.045 -70.205 -61.715 -69.875 ;
        RECT -62.045 -71.565 -61.715 -71.235 ;
        RECT -62.045 -72.925 -61.715 -72.595 ;
        RECT -62.045 -74.285 -61.715 -73.955 ;
        RECT -62.045 -75.645 -61.715 -75.315 ;
        RECT -62.045 -77.005 -61.715 -76.675 ;
        RECT -62.045 -78.365 -61.715 -78.035 ;
        RECT -62.045 -79.725 -61.715 -79.395 ;
        RECT -62.045 -81.085 -61.715 -80.755 ;
        RECT -62.045 -82.445 -61.715 -82.115 ;
        RECT -62.045 -83.805 -61.715 -83.475 ;
        RECT -62.045 -85.165 -61.715 -84.835 ;
        RECT -62.045 -86.525 -61.715 -86.195 ;
        RECT -62.045 -87.885 -61.715 -87.555 ;
        RECT -62.045 -89.245 -61.715 -88.915 ;
        RECT -62.045 -90.605 -61.715 -90.275 ;
        RECT -62.045 -91.965 -61.715 -91.635 ;
        RECT -62.045 -93.325 -61.715 -92.995 ;
        RECT -62.045 -94.685 -61.715 -94.355 ;
        RECT -62.045 -96.045 -61.715 -95.715 ;
        RECT -62.045 -97.405 -61.715 -97.075 ;
        RECT -62.045 -98.765 -61.715 -98.435 ;
        RECT -62.045 -100.125 -61.715 -99.795 ;
        RECT -62.045 -101.485 -61.715 -101.155 ;
        RECT -62.045 -102.845 -61.715 -102.515 ;
        RECT -62.045 -104.205 -61.715 -103.875 ;
        RECT -62.045 -105.565 -61.715 -105.235 ;
        RECT -62.045 -106.925 -61.715 -106.595 ;
        RECT -62.045 -108.285 -61.715 -107.955 ;
        RECT -62.045 -109.645 -61.715 -109.315 ;
        RECT -62.045 -111.005 -61.715 -110.675 ;
        RECT -62.045 -112.365 -61.715 -112.035 ;
        RECT -62.045 -113.725 -61.715 -113.395 ;
        RECT -62.045 -115.085 -61.715 -114.755 ;
        RECT -62.045 -116.445 -61.715 -116.115 ;
        RECT -62.045 -117.805 -61.715 -117.475 ;
        RECT -62.045 -119.165 -61.715 -118.835 ;
        RECT -62.045 -120.525 -61.715 -120.195 ;
        RECT -62.045 -121.885 -61.715 -121.555 ;
        RECT -62.045 -123.245 -61.715 -122.915 ;
        RECT -62.045 -124.605 -61.715 -124.275 ;
        RECT -62.045 -125.965 -61.715 -125.635 ;
        RECT -62.045 -127.325 -61.715 -126.995 ;
        RECT -62.045 -128.685 -61.715 -128.355 ;
        RECT -62.045 -130.045 -61.715 -129.715 ;
        RECT -62.045 -131.405 -61.715 -131.075 ;
        RECT -62.045 -132.765 -61.715 -132.435 ;
        RECT -62.045 -134.125 -61.715 -133.795 ;
        RECT -62.045 -135.485 -61.715 -135.155 ;
        RECT -62.045 -136.845 -61.715 -136.515 ;
        RECT -62.045 -138.205 -61.715 -137.875 ;
        RECT -62.045 -139.565 -61.715 -139.235 ;
        RECT -62.045 -140.925 -61.715 -140.595 ;
        RECT -62.045 -142.285 -61.715 -141.955 ;
        RECT -62.045 -143.645 -61.715 -143.315 ;
        RECT -62.045 -145.005 -61.715 -144.675 ;
        RECT -62.045 -146.365 -61.715 -146.035 ;
        RECT -62.045 -148.215 -61.715 -147.885 ;
        RECT -62.045 -149.085 -61.715 -148.755 ;
        RECT -62.045 -150.445 -61.715 -150.115 ;
        RECT -62.045 -151.805 -61.715 -151.475 ;
        RECT -62.045 -153.165 -61.715 -152.835 ;
        RECT -62.045 -154.525 -61.715 -154.195 ;
        RECT -62.045 -157.245 -61.715 -156.915 ;
        RECT -62.045 -162.89 -61.715 -161.76 ;
        RECT -62.04 -163.005 -61.72 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 129.945 -60.355 131.075 ;
        RECT -60.685 125.635 -60.355 125.965 ;
        RECT -60.685 124.275 -60.355 124.605 ;
        RECT -60.685 122.915 -60.355 123.245 ;
        RECT -60.685 121.555 -60.355 121.885 ;
        RECT -60.685 120.195 -60.355 120.525 ;
        RECT -60.685 118.835 -60.355 119.165 ;
        RECT -60.685 117.475 -60.355 117.805 ;
        RECT -60.685 116.115 -60.355 116.445 ;
        RECT -60.685 114.755 -60.355 115.085 ;
        RECT -60.685 113.395 -60.355 113.725 ;
        RECT -60.685 112.035 -60.355 112.365 ;
        RECT -60.685 110.675 -60.355 111.005 ;
        RECT -60.685 109.315 -60.355 109.645 ;
        RECT -60.685 107.955 -60.355 108.285 ;
        RECT -60.685 106.595 -60.355 106.925 ;
        RECT -60.685 105.235 -60.355 105.565 ;
        RECT -60.685 103.875 -60.355 104.205 ;
        RECT -60.685 102.515 -60.355 102.845 ;
        RECT -60.685 101.155 -60.355 101.485 ;
        RECT -60.685 99.795 -60.355 100.125 ;
        RECT -60.685 98.435 -60.355 98.765 ;
        RECT -60.685 97.075 -60.355 97.405 ;
        RECT -60.685 95.715 -60.355 96.045 ;
        RECT -60.685 94.355 -60.355 94.685 ;
        RECT -60.685 92.995 -60.355 93.325 ;
        RECT -60.685 91.635 -60.355 91.965 ;
        RECT -60.685 90.275 -60.355 90.605 ;
        RECT -60.685 88.915 -60.355 89.245 ;
        RECT -60.685 87.555 -60.355 87.885 ;
        RECT -60.685 86.195 -60.355 86.525 ;
        RECT -60.685 84.835 -60.355 85.165 ;
        RECT -60.685 83.475 -60.355 83.805 ;
        RECT -60.685 82.115 -60.355 82.445 ;
        RECT -60.685 80.755 -60.355 81.085 ;
        RECT -60.685 79.395 -60.355 79.725 ;
        RECT -60.685 78.035 -60.355 78.365 ;
        RECT -60.685 76.675 -60.355 77.005 ;
        RECT -60.685 75.315 -60.355 75.645 ;
        RECT -60.685 73.955 -60.355 74.285 ;
        RECT -60.685 48.115 -60.355 48.445 ;
        RECT -60.685 46.755 -60.355 47.085 ;
        RECT -60.685 45.395 -60.355 45.725 ;
        RECT -60.685 44.035 -60.355 44.365 ;
        RECT -60.685 42.675 -60.355 43.005 ;
        RECT -60.685 41.315 -60.355 41.645 ;
        RECT -60.685 39.955 -60.355 40.285 ;
        RECT -60.685 38.595 -60.355 38.925 ;
        RECT -60.685 37.235 -60.355 37.565 ;
        RECT -60.685 35.875 -60.355 36.205 ;
        RECT -60.685 34.515 -60.355 34.845 ;
        RECT -60.685 33.155 -60.355 33.485 ;
        RECT -60.685 31.795 -60.355 32.125 ;
        RECT -60.685 30.435 -60.355 30.765 ;
        RECT -60.685 29.075 -60.355 29.405 ;
        RECT -60.685 27.715 -60.355 28.045 ;
        RECT -60.685 26.355 -60.355 26.685 ;
        RECT -60.685 24.995 -60.355 25.325 ;
        RECT -60.685 23.635 -60.355 23.965 ;
        RECT -60.685 22.275 -60.355 22.605 ;
        RECT -60.685 20.915 -60.355 21.245 ;
        RECT -60.685 19.555 -60.355 19.885 ;
        RECT -60.685 18.195 -60.355 18.525 ;
        RECT -60.685 16.835 -60.355 17.165 ;
        RECT -60.685 15.475 -60.355 15.805 ;
        RECT -60.685 14.115 -60.355 14.445 ;
        RECT -60.685 12.755 -60.355 13.085 ;
        RECT -60.685 11.395 -60.355 11.725 ;
        RECT -60.685 10.035 -60.355 10.365 ;
        RECT -60.685 8.675 -60.355 9.005 ;
        RECT -60.685 7.315 -60.355 7.645 ;
        RECT -60.685 5.955 -60.355 6.285 ;
        RECT -60.685 4.595 -60.355 4.925 ;
        RECT -60.685 3.235 -60.355 3.565 ;
        RECT -60.685 1.875 -60.355 2.205 ;
        RECT -60.685 0.515 -60.355 0.845 ;
        RECT -60.685 -0.845 -60.355 -0.515 ;
        RECT -60.685 -2.205 -60.355 -1.875 ;
        RECT -60.685 -3.565 -60.355 -3.235 ;
        RECT -60.685 -4.925 -60.355 -4.595 ;
        RECT -60.685 -6.285 -60.355 -5.955 ;
        RECT -60.685 -7.645 -60.355 -7.315 ;
        RECT -60.685 -9.005 -60.355 -8.675 ;
        RECT -60.685 -10.365 -60.355 -10.035 ;
        RECT -60.685 -11.725 -60.355 -11.395 ;
        RECT -60.685 -13.085 -60.355 -12.755 ;
        RECT -60.685 -14.445 -60.355 -14.115 ;
        RECT -60.685 -15.805 -60.355 -15.475 ;
        RECT -60.685 -17.165 -60.355 -16.835 ;
        RECT -60.685 -18.525 -60.355 -18.195 ;
        RECT -60.685 -19.885 -60.355 -19.555 ;
        RECT -60.685 -21.245 -60.355 -20.915 ;
        RECT -60.685 -22.605 -60.355 -22.275 ;
        RECT -60.685 -23.965 -60.355 -23.635 ;
        RECT -60.685 -25.325 -60.355 -24.995 ;
        RECT -60.685 -26.685 -60.355 -26.355 ;
        RECT -60.685 -28.045 -60.355 -27.715 ;
        RECT -60.685 -29.405 -60.355 -29.075 ;
        RECT -60.685 -30.765 -60.355 -30.435 ;
        RECT -60.685 -32.125 -60.355 -31.795 ;
        RECT -60.685 -33.485 -60.355 -33.155 ;
        RECT -60.685 -34.845 -60.355 -34.515 ;
        RECT -60.685 -36.205 -60.355 -35.875 ;
        RECT -60.685 -37.565 -60.355 -37.235 ;
        RECT -60.685 -38.925 -60.355 -38.595 ;
        RECT -60.685 -40.285 -60.355 -39.955 ;
        RECT -60.685 -41.645 -60.355 -41.315 ;
        RECT -60.685 -43.005 -60.355 -42.675 ;
        RECT -60.685 -44.365 -60.355 -44.035 ;
        RECT -60.685 -45.725 -60.355 -45.395 ;
        RECT -60.685 -47.085 -60.355 -46.755 ;
        RECT -60.685 -48.445 -60.355 -48.115 ;
        RECT -60.685 -49.805 -60.355 -49.475 ;
        RECT -60.685 -51.165 -60.355 -50.835 ;
        RECT -60.685 -52.525 -60.355 -52.195 ;
        RECT -60.685 -53.885 -60.355 -53.555 ;
        RECT -60.685 -55.245 -60.355 -54.915 ;
        RECT -60.685 -56.605 -60.355 -56.275 ;
        RECT -60.685 -57.965 -60.355 -57.635 ;
        RECT -60.685 -59.325 -60.355 -58.995 ;
        RECT -60.685 -60.685 -60.355 -60.355 ;
        RECT -60.685 -62.045 -60.355 -61.715 ;
        RECT -60.685 -63.405 -60.355 -63.075 ;
        RECT -60.685 -64.765 -60.355 -64.435 ;
        RECT -60.685 -66.125 -60.355 -65.795 ;
        RECT -60.685 -67.485 -60.355 -67.155 ;
        RECT -60.685 -68.845 -60.355 -68.515 ;
        RECT -60.685 -70.205 -60.355 -69.875 ;
        RECT -60.685 -71.565 -60.355 -71.235 ;
        RECT -60.685 -72.925 -60.355 -72.595 ;
        RECT -60.685 -74.285 -60.355 -73.955 ;
        RECT -60.685 -75.645 -60.355 -75.315 ;
        RECT -60.685 -77.005 -60.355 -76.675 ;
        RECT -60.685 -78.365 -60.355 -78.035 ;
        RECT -60.685 -79.725 -60.355 -79.395 ;
        RECT -60.685 -81.085 -60.355 -80.755 ;
        RECT -60.685 -82.445 -60.355 -82.115 ;
        RECT -60.685 -83.805 -60.355 -83.475 ;
        RECT -60.685 -85.165 -60.355 -84.835 ;
        RECT -60.685 -86.525 -60.355 -86.195 ;
        RECT -60.685 -87.885 -60.355 -87.555 ;
        RECT -60.685 -89.245 -60.355 -88.915 ;
        RECT -60.685 -90.605 -60.355 -90.275 ;
        RECT -60.685 -91.965 -60.355 -91.635 ;
        RECT -60.68 -91.965 -60.36 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 -154.525 -60.355 -154.195 ;
        RECT -60.685 -157.245 -60.355 -156.915 ;
        RECT -60.685 -162.89 -60.355 -161.76 ;
        RECT -60.68 -163.005 -60.36 -153.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.325 129.945 -58.995 131.075 ;
        RECT -59.325 125.635 -58.995 125.965 ;
        RECT -59.325 124.275 -58.995 124.605 ;
        RECT -59.325 122.915 -58.995 123.245 ;
        RECT -59.325 121.555 -58.995 121.885 ;
        RECT -59.325 120.195 -58.995 120.525 ;
        RECT -59.325 118.835 -58.995 119.165 ;
        RECT -59.325 117.475 -58.995 117.805 ;
        RECT -59.325 116.115 -58.995 116.445 ;
        RECT -59.325 114.755 -58.995 115.085 ;
        RECT -59.325 113.395 -58.995 113.725 ;
        RECT -59.325 112.035 -58.995 112.365 ;
        RECT -59.325 110.675 -58.995 111.005 ;
        RECT -59.325 109.315 -58.995 109.645 ;
        RECT -59.325 107.955 -58.995 108.285 ;
        RECT -59.325 106.595 -58.995 106.925 ;
        RECT -59.325 105.235 -58.995 105.565 ;
        RECT -59.325 103.875 -58.995 104.205 ;
        RECT -59.325 102.515 -58.995 102.845 ;
        RECT -59.325 101.155 -58.995 101.485 ;
        RECT -59.325 99.795 -58.995 100.125 ;
        RECT -59.325 98.435 -58.995 98.765 ;
        RECT -59.325 97.075 -58.995 97.405 ;
        RECT -59.325 95.715 -58.995 96.045 ;
        RECT -59.325 94.355 -58.995 94.685 ;
        RECT -59.325 92.995 -58.995 93.325 ;
        RECT -59.325 91.635 -58.995 91.965 ;
        RECT -59.325 90.275 -58.995 90.605 ;
        RECT -59.325 88.915 -58.995 89.245 ;
        RECT -59.325 87.555 -58.995 87.885 ;
        RECT -59.325 86.195 -58.995 86.525 ;
        RECT -59.325 84.835 -58.995 85.165 ;
        RECT -59.325 83.475 -58.995 83.805 ;
        RECT -59.325 82.115 -58.995 82.445 ;
        RECT -59.325 80.755 -58.995 81.085 ;
        RECT -59.325 79.395 -58.995 79.725 ;
        RECT -59.325 78.035 -58.995 78.365 ;
        RECT -59.325 76.675 -58.995 77.005 ;
        RECT -59.325 75.315 -58.995 75.645 ;
        RECT -59.325 73.955 -58.995 74.285 ;
        RECT -59.325 71.64 -58.995 71.97 ;
        RECT -59.325 69.465 -58.995 69.795 ;
        RECT -59.325 68.615 -58.995 68.945 ;
        RECT -59.325 66.305 -58.995 66.635 ;
        RECT -59.325 65.455 -58.995 65.785 ;
        RECT -59.325 63.145 -58.995 63.475 ;
        RECT -59.325 62.295 -58.995 62.625 ;
        RECT -59.325 59.985 -58.995 60.315 ;
        RECT -59.325 59.135 -58.995 59.465 ;
        RECT -59.325 56.825 -58.995 57.155 ;
        RECT -59.325 55.975 -58.995 56.305 ;
        RECT -59.325 53.665 -58.995 53.995 ;
        RECT -59.325 52.815 -58.995 53.145 ;
        RECT -59.325 50.64 -58.995 50.97 ;
        RECT -59.325 48.115 -58.995 48.445 ;
        RECT -59.325 46.755 -58.995 47.085 ;
        RECT -59.325 45.395 -58.995 45.725 ;
        RECT -59.325 44.035 -58.995 44.365 ;
        RECT -59.325 42.675 -58.995 43.005 ;
        RECT -59.325 41.315 -58.995 41.645 ;
        RECT -59.325 39.955 -58.995 40.285 ;
        RECT -59.325 38.595 -58.995 38.925 ;
        RECT -59.325 37.235 -58.995 37.565 ;
        RECT -59.325 35.875 -58.995 36.205 ;
        RECT -59.325 34.515 -58.995 34.845 ;
        RECT -59.325 33.155 -58.995 33.485 ;
        RECT -59.325 31.795 -58.995 32.125 ;
        RECT -59.325 30.435 -58.995 30.765 ;
        RECT -59.325 29.075 -58.995 29.405 ;
        RECT -59.325 27.715 -58.995 28.045 ;
        RECT -59.325 26.355 -58.995 26.685 ;
        RECT -59.325 24.995 -58.995 25.325 ;
        RECT -59.325 23.635 -58.995 23.965 ;
        RECT -59.325 22.275 -58.995 22.605 ;
        RECT -59.325 20.915 -58.995 21.245 ;
        RECT -59.325 19.555 -58.995 19.885 ;
        RECT -59.325 18.195 -58.995 18.525 ;
        RECT -59.325 16.835 -58.995 17.165 ;
        RECT -59.325 15.475 -58.995 15.805 ;
        RECT -59.325 14.115 -58.995 14.445 ;
        RECT -59.325 12.755 -58.995 13.085 ;
        RECT -59.325 11.395 -58.995 11.725 ;
        RECT -59.325 10.035 -58.995 10.365 ;
        RECT -59.325 8.675 -58.995 9.005 ;
        RECT -59.325 7.315 -58.995 7.645 ;
        RECT -59.325 5.955 -58.995 6.285 ;
        RECT -59.325 4.595 -58.995 4.925 ;
        RECT -59.325 3.235 -58.995 3.565 ;
        RECT -59.325 1.875 -58.995 2.205 ;
        RECT -59.325 0.515 -58.995 0.845 ;
        RECT -59.325 -0.845 -58.995 -0.515 ;
        RECT -59.325 -2.205 -58.995 -1.875 ;
        RECT -59.325 -3.565 -58.995 -3.235 ;
        RECT -59.325 -4.925 -58.995 -4.595 ;
        RECT -59.325 -6.285 -58.995 -5.955 ;
        RECT -59.325 -7.645 -58.995 -7.315 ;
        RECT -59.325 -9.005 -58.995 -8.675 ;
        RECT -59.325 -10.365 -58.995 -10.035 ;
        RECT -59.325 -11.725 -58.995 -11.395 ;
        RECT -59.325 -13.085 -58.995 -12.755 ;
        RECT -59.325 -14.445 -58.995 -14.115 ;
        RECT -59.325 -15.805 -58.995 -15.475 ;
        RECT -59.325 -17.165 -58.995 -16.835 ;
        RECT -59.325 -18.525 -58.995 -18.195 ;
        RECT -59.325 -19.885 -58.995 -19.555 ;
        RECT -59.325 -21.245 -58.995 -20.915 ;
        RECT -59.325 -22.605 -58.995 -22.275 ;
        RECT -59.325 -23.965 -58.995 -23.635 ;
        RECT -59.325 -25.325 -58.995 -24.995 ;
        RECT -59.325 -26.685 -58.995 -26.355 ;
        RECT -59.325 -28.045 -58.995 -27.715 ;
        RECT -59.325 -29.405 -58.995 -29.075 ;
        RECT -59.325 -30.765 -58.995 -30.435 ;
        RECT -59.325 -32.125 -58.995 -31.795 ;
        RECT -59.325 -33.485 -58.995 -33.155 ;
        RECT -59.325 -34.845 -58.995 -34.515 ;
        RECT -59.325 -36.205 -58.995 -35.875 ;
        RECT -59.325 -37.565 -58.995 -37.235 ;
        RECT -59.325 -38.925 -58.995 -38.595 ;
        RECT -59.325 -40.285 -58.995 -39.955 ;
        RECT -59.325 -41.645 -58.995 -41.315 ;
        RECT -59.325 -43.005 -58.995 -42.675 ;
        RECT -59.325 -44.365 -58.995 -44.035 ;
        RECT -59.325 -45.725 -58.995 -45.395 ;
        RECT -59.325 -47.085 -58.995 -46.755 ;
        RECT -59.325 -48.445 -58.995 -48.115 ;
        RECT -59.325 -49.805 -58.995 -49.475 ;
        RECT -59.325 -51.165 -58.995 -50.835 ;
        RECT -59.325 -52.525 -58.995 -52.195 ;
        RECT -59.325 -53.885 -58.995 -53.555 ;
        RECT -59.325 -55.245 -58.995 -54.915 ;
        RECT -59.325 -56.605 -58.995 -56.275 ;
        RECT -59.325 -57.965 -58.995 -57.635 ;
        RECT -59.325 -59.325 -58.995 -58.995 ;
        RECT -59.325 -60.685 -58.995 -60.355 ;
        RECT -59.325 -62.045 -58.995 -61.715 ;
        RECT -59.325 -63.405 -58.995 -63.075 ;
        RECT -59.325 -64.765 -58.995 -64.435 ;
        RECT -59.325 -66.125 -58.995 -65.795 ;
        RECT -59.325 -67.485 -58.995 -67.155 ;
        RECT -59.325 -68.845 -58.995 -68.515 ;
        RECT -59.325 -70.205 -58.995 -69.875 ;
        RECT -59.325 -71.565 -58.995 -71.235 ;
        RECT -59.325 -72.925 -58.995 -72.595 ;
        RECT -59.325 -74.285 -58.995 -73.955 ;
        RECT -59.325 -75.645 -58.995 -75.315 ;
        RECT -59.325 -77.005 -58.995 -76.675 ;
        RECT -59.325 -78.365 -58.995 -78.035 ;
        RECT -59.325 -79.725 -58.995 -79.395 ;
        RECT -59.325 -81.085 -58.995 -80.755 ;
        RECT -59.325 -82.445 -58.995 -82.115 ;
        RECT -59.325 -83.805 -58.995 -83.475 ;
        RECT -59.325 -85.165 -58.995 -84.835 ;
        RECT -59.325 -86.525 -58.995 -86.195 ;
        RECT -59.325 -87.885 -58.995 -87.555 ;
        RECT -59.325 -89.245 -58.995 -88.915 ;
        RECT -59.325 -90.605 -58.995 -90.275 ;
        RECT -59.325 -93.325 -58.995 -92.995 ;
        RECT -59.325 -94.685 -58.995 -94.355 ;
        RECT -59.325 -96.045 -58.995 -95.715 ;
        RECT -59.325 -97.405 -58.995 -97.075 ;
        RECT -59.325 -98.765 -58.995 -98.435 ;
        RECT -59.325 -100.125 -58.995 -99.795 ;
        RECT -59.325 -101.485 -58.995 -101.155 ;
        RECT -59.325 -102.845 -58.995 -102.515 ;
        RECT -59.325 -104.205 -58.995 -103.875 ;
        RECT -59.325 -105.565 -58.995 -105.235 ;
        RECT -59.325 -106.925 -58.995 -106.595 ;
        RECT -59.325 -108.285 -58.995 -107.955 ;
        RECT -59.325 -109.645 -58.995 -109.315 ;
        RECT -59.325 -111.005 -58.995 -110.675 ;
        RECT -59.325 -112.365 -58.995 -112.035 ;
        RECT -59.325 -113.725 -58.995 -113.395 ;
        RECT -59.325 -115.085 -58.995 -114.755 ;
        RECT -59.325 -116.445 -58.995 -116.115 ;
        RECT -59.325 -117.805 -58.995 -117.475 ;
        RECT -59.325 -119.165 -58.995 -118.835 ;
        RECT -59.325 -120.525 -58.995 -120.195 ;
        RECT -59.325 -121.885 -58.995 -121.555 ;
        RECT -59.325 -123.245 -58.995 -122.915 ;
        RECT -59.325 -124.605 -58.995 -124.275 ;
        RECT -59.325 -125.965 -58.995 -125.635 ;
        RECT -59.325 -127.325 -58.995 -126.995 ;
        RECT -59.325 -128.685 -58.995 -128.355 ;
        RECT -59.325 -130.045 -58.995 -129.715 ;
        RECT -59.325 -131.405 -58.995 -131.075 ;
        RECT -59.325 -132.765 -58.995 -132.435 ;
        RECT -59.325 -134.125 -58.995 -133.795 ;
        RECT -59.325 -135.485 -58.995 -135.155 ;
        RECT -59.325 -136.845 -58.995 -136.515 ;
        RECT -59.325 -138.205 -58.995 -137.875 ;
        RECT -59.325 -139.565 -58.995 -139.235 ;
        RECT -59.325 -140.925 -58.995 -140.595 ;
        RECT -59.325 -142.285 -58.995 -141.955 ;
        RECT -59.325 -143.645 -58.995 -143.315 ;
        RECT -59.325 -145.005 -58.995 -144.675 ;
        RECT -59.325 -146.365 -58.995 -146.035 ;
        RECT -59.325 -149.085 -58.995 -148.755 ;
        RECT -59.325 -150.445 -58.995 -150.115 ;
        RECT -59.325 -153.165 -58.995 -152.835 ;
        RECT -59.325 -154.525 -58.995 -154.195 ;
        RECT -59.325 -157.245 -58.995 -156.915 ;
        RECT -59.325 -162.89 -58.995 -161.76 ;
        RECT -59.32 -163.005 -59 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.965 -74.285 -57.635 -73.955 ;
        RECT -57.965 -75.645 -57.635 -75.315 ;
        RECT -57.965 -77.005 -57.635 -76.675 ;
        RECT -57.965 -78.365 -57.635 -78.035 ;
        RECT -57.965 -79.725 -57.635 -79.395 ;
        RECT -57.965 -81.085 -57.635 -80.755 ;
        RECT -57.965 -82.445 -57.635 -82.115 ;
        RECT -57.965 -83.805 -57.635 -83.475 ;
        RECT -57.965 -85.165 -57.635 -84.835 ;
        RECT -57.965 -86.525 -57.635 -86.195 ;
        RECT -57.965 -87.885 -57.635 -87.555 ;
        RECT -57.965 -89.245 -57.635 -88.915 ;
        RECT -57.965 -90.605 -57.635 -90.275 ;
        RECT -57.965 -93.325 -57.635 -92.995 ;
        RECT -57.965 -94.685 -57.635 -94.355 ;
        RECT -57.965 -96.045 -57.635 -95.715 ;
        RECT -57.965 -97.405 -57.635 -97.075 ;
        RECT -57.965 -98.765 -57.635 -98.435 ;
        RECT -57.965 -100.125 -57.635 -99.795 ;
        RECT -57.965 -101.485 -57.635 -101.155 ;
        RECT -57.965 -102.845 -57.635 -102.515 ;
        RECT -57.965 -104.205 -57.635 -103.875 ;
        RECT -57.965 -105.565 -57.635 -105.235 ;
        RECT -57.965 -106.925 -57.635 -106.595 ;
        RECT -57.965 -108.285 -57.635 -107.955 ;
        RECT -57.965 -109.645 -57.635 -109.315 ;
        RECT -57.965 -111.005 -57.635 -110.675 ;
        RECT -57.965 -112.365 -57.635 -112.035 ;
        RECT -57.965 -113.725 -57.635 -113.395 ;
        RECT -57.965 -115.085 -57.635 -114.755 ;
        RECT -57.965 -116.445 -57.635 -116.115 ;
        RECT -57.965 -117.805 -57.635 -117.475 ;
        RECT -57.965 -119.165 -57.635 -118.835 ;
        RECT -57.965 -120.525 -57.635 -120.195 ;
        RECT -57.965 -121.885 -57.635 -121.555 ;
        RECT -57.965 -123.245 -57.635 -122.915 ;
        RECT -57.965 -124.605 -57.635 -124.275 ;
        RECT -57.965 -125.965 -57.635 -125.635 ;
        RECT -57.965 -127.325 -57.635 -126.995 ;
        RECT -57.965 -128.685 -57.635 -128.355 ;
        RECT -57.965 -130.045 -57.635 -129.715 ;
        RECT -57.965 -131.405 -57.635 -131.075 ;
        RECT -57.965 -132.765 -57.635 -132.435 ;
        RECT -57.965 -134.125 -57.635 -133.795 ;
        RECT -57.965 -135.485 -57.635 -135.155 ;
        RECT -57.965 -136.845 -57.635 -136.515 ;
        RECT -57.965 -138.205 -57.635 -137.875 ;
        RECT -57.965 -139.565 -57.635 -139.235 ;
        RECT -57.965 -140.925 -57.635 -140.595 ;
        RECT -57.965 -142.285 -57.635 -141.955 ;
        RECT -57.965 -143.645 -57.635 -143.315 ;
        RECT -57.965 -145.005 -57.635 -144.675 ;
        RECT -57.965 -146.365 -57.635 -146.035 ;
        RECT -57.965 -148.215 -57.635 -147.885 ;
        RECT -57.965 -149.085 -57.635 -148.755 ;
        RECT -57.965 -150.445 -57.635 -150.115 ;
        RECT -57.965 -153.165 -57.635 -152.835 ;
        RECT -57.965 -154.525 -57.635 -154.195 ;
        RECT -57.965 -157.245 -57.635 -156.915 ;
        RECT -57.965 -162.89 -57.635 -161.76 ;
        RECT -57.96 -163.005 -57.64 131.19 ;
        RECT -57.965 129.945 -57.635 131.075 ;
        RECT -57.965 125.635 -57.635 125.965 ;
        RECT -57.965 124.275 -57.635 124.605 ;
        RECT -57.965 122.915 -57.635 123.245 ;
        RECT -57.965 121.555 -57.635 121.885 ;
        RECT -57.965 120.195 -57.635 120.525 ;
        RECT -57.965 118.835 -57.635 119.165 ;
        RECT -57.965 117.475 -57.635 117.805 ;
        RECT -57.965 116.115 -57.635 116.445 ;
        RECT -57.965 114.755 -57.635 115.085 ;
        RECT -57.965 113.395 -57.635 113.725 ;
        RECT -57.965 112.035 -57.635 112.365 ;
        RECT -57.965 110.675 -57.635 111.005 ;
        RECT -57.965 109.315 -57.635 109.645 ;
        RECT -57.965 107.955 -57.635 108.285 ;
        RECT -57.965 106.595 -57.635 106.925 ;
        RECT -57.965 105.235 -57.635 105.565 ;
        RECT -57.965 103.875 -57.635 104.205 ;
        RECT -57.965 102.515 -57.635 102.845 ;
        RECT -57.965 101.155 -57.635 101.485 ;
        RECT -57.965 99.795 -57.635 100.125 ;
        RECT -57.965 98.435 -57.635 98.765 ;
        RECT -57.965 97.075 -57.635 97.405 ;
        RECT -57.965 95.715 -57.635 96.045 ;
        RECT -57.965 94.355 -57.635 94.685 ;
        RECT -57.965 92.995 -57.635 93.325 ;
        RECT -57.965 91.635 -57.635 91.965 ;
        RECT -57.965 90.275 -57.635 90.605 ;
        RECT -57.965 88.915 -57.635 89.245 ;
        RECT -57.965 87.555 -57.635 87.885 ;
        RECT -57.965 86.195 -57.635 86.525 ;
        RECT -57.965 84.835 -57.635 85.165 ;
        RECT -57.965 83.475 -57.635 83.805 ;
        RECT -57.965 82.115 -57.635 82.445 ;
        RECT -57.965 80.755 -57.635 81.085 ;
        RECT -57.965 79.395 -57.635 79.725 ;
        RECT -57.965 78.035 -57.635 78.365 ;
        RECT -57.965 76.675 -57.635 77.005 ;
        RECT -57.965 75.315 -57.635 75.645 ;
        RECT -57.965 73.955 -57.635 74.285 ;
        RECT -57.965 71.64 -57.635 71.97 ;
        RECT -57.965 69.465 -57.635 69.795 ;
        RECT -57.965 68.615 -57.635 68.945 ;
        RECT -57.965 66.305 -57.635 66.635 ;
        RECT -57.965 65.455 -57.635 65.785 ;
        RECT -57.965 63.145 -57.635 63.475 ;
        RECT -57.965 62.295 -57.635 62.625 ;
        RECT -57.965 59.985 -57.635 60.315 ;
        RECT -57.965 59.135 -57.635 59.465 ;
        RECT -57.965 56.825 -57.635 57.155 ;
        RECT -57.965 55.975 -57.635 56.305 ;
        RECT -57.965 53.665 -57.635 53.995 ;
        RECT -57.965 52.815 -57.635 53.145 ;
        RECT -57.965 50.64 -57.635 50.97 ;
        RECT -57.965 48.115 -57.635 48.445 ;
        RECT -57.965 46.755 -57.635 47.085 ;
        RECT -57.965 45.395 -57.635 45.725 ;
        RECT -57.965 44.035 -57.635 44.365 ;
        RECT -57.965 42.675 -57.635 43.005 ;
        RECT -57.965 41.315 -57.635 41.645 ;
        RECT -57.965 39.955 -57.635 40.285 ;
        RECT -57.965 38.595 -57.635 38.925 ;
        RECT -57.965 37.235 -57.635 37.565 ;
        RECT -57.965 35.875 -57.635 36.205 ;
        RECT -57.965 34.515 -57.635 34.845 ;
        RECT -57.965 33.155 -57.635 33.485 ;
        RECT -57.965 31.795 -57.635 32.125 ;
        RECT -57.965 30.435 -57.635 30.765 ;
        RECT -57.965 29.075 -57.635 29.405 ;
        RECT -57.965 27.715 -57.635 28.045 ;
        RECT -57.965 26.355 -57.635 26.685 ;
        RECT -57.965 24.995 -57.635 25.325 ;
        RECT -57.965 23.635 -57.635 23.965 ;
        RECT -57.965 22.275 -57.635 22.605 ;
        RECT -57.965 20.915 -57.635 21.245 ;
        RECT -57.965 19.555 -57.635 19.885 ;
        RECT -57.965 18.195 -57.635 18.525 ;
        RECT -57.965 16.835 -57.635 17.165 ;
        RECT -57.965 15.475 -57.635 15.805 ;
        RECT -57.965 14.115 -57.635 14.445 ;
        RECT -57.965 12.755 -57.635 13.085 ;
        RECT -57.965 11.395 -57.635 11.725 ;
        RECT -57.965 10.035 -57.635 10.365 ;
        RECT -57.965 8.675 -57.635 9.005 ;
        RECT -57.965 7.315 -57.635 7.645 ;
        RECT -57.965 5.955 -57.635 6.285 ;
        RECT -57.965 4.595 -57.635 4.925 ;
        RECT -57.965 3.235 -57.635 3.565 ;
        RECT -57.965 1.875 -57.635 2.205 ;
        RECT -57.965 0.515 -57.635 0.845 ;
        RECT -57.965 -0.845 -57.635 -0.515 ;
        RECT -57.965 -2.205 -57.635 -1.875 ;
        RECT -57.965 -3.565 -57.635 -3.235 ;
        RECT -57.965 -4.925 -57.635 -4.595 ;
        RECT -57.965 -6.285 -57.635 -5.955 ;
        RECT -57.965 -7.645 -57.635 -7.315 ;
        RECT -57.965 -9.005 -57.635 -8.675 ;
        RECT -57.965 -10.365 -57.635 -10.035 ;
        RECT -57.965 -11.725 -57.635 -11.395 ;
        RECT -57.965 -13.085 -57.635 -12.755 ;
        RECT -57.965 -14.445 -57.635 -14.115 ;
        RECT -57.965 -15.805 -57.635 -15.475 ;
        RECT -57.965 -17.165 -57.635 -16.835 ;
        RECT -57.965 -18.525 -57.635 -18.195 ;
        RECT -57.965 -19.885 -57.635 -19.555 ;
        RECT -57.965 -21.245 -57.635 -20.915 ;
        RECT -57.965 -22.605 -57.635 -22.275 ;
        RECT -57.965 -23.965 -57.635 -23.635 ;
        RECT -57.965 -25.325 -57.635 -24.995 ;
        RECT -57.965 -26.685 -57.635 -26.355 ;
        RECT -57.965 -28.045 -57.635 -27.715 ;
        RECT -57.965 -29.405 -57.635 -29.075 ;
        RECT -57.965 -30.765 -57.635 -30.435 ;
        RECT -57.965 -32.125 -57.635 -31.795 ;
        RECT -57.965 -33.485 -57.635 -33.155 ;
        RECT -57.965 -34.845 -57.635 -34.515 ;
        RECT -57.965 -36.205 -57.635 -35.875 ;
        RECT -57.965 -37.565 -57.635 -37.235 ;
        RECT -57.965 -38.925 -57.635 -38.595 ;
        RECT -57.965 -40.285 -57.635 -39.955 ;
        RECT -57.965 -41.645 -57.635 -41.315 ;
        RECT -57.965 -43.005 -57.635 -42.675 ;
        RECT -57.965 -44.365 -57.635 -44.035 ;
        RECT -57.965 -45.725 -57.635 -45.395 ;
        RECT -57.965 -47.085 -57.635 -46.755 ;
        RECT -57.965 -48.445 -57.635 -48.115 ;
        RECT -57.965 -49.805 -57.635 -49.475 ;
        RECT -57.965 -51.165 -57.635 -50.835 ;
        RECT -57.965 -52.525 -57.635 -52.195 ;
        RECT -57.965 -53.885 -57.635 -53.555 ;
        RECT -57.965 -55.245 -57.635 -54.915 ;
        RECT -57.965 -56.605 -57.635 -56.275 ;
        RECT -57.965 -57.965 -57.635 -57.635 ;
        RECT -57.965 -59.325 -57.635 -58.995 ;
        RECT -57.965 -60.685 -57.635 -60.355 ;
        RECT -57.965 -62.045 -57.635 -61.715 ;
        RECT -57.965 -63.405 -57.635 -63.075 ;
        RECT -57.965 -64.765 -57.635 -64.435 ;
        RECT -57.965 -66.125 -57.635 -65.795 ;
        RECT -57.965 -67.485 -57.635 -67.155 ;
        RECT -57.965 -68.845 -57.635 -68.515 ;
        RECT -57.965 -70.205 -57.635 -69.875 ;
        RECT -57.965 -71.565 -57.635 -71.235 ;
        RECT -57.965 -72.925 -57.635 -72.595 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.485 129.945 -67.155 131.075 ;
        RECT -67.485 125.635 -67.155 125.965 ;
        RECT -67.485 124.275 -67.155 124.605 ;
        RECT -67.485 122.915 -67.155 123.245 ;
        RECT -67.485 121.555 -67.155 121.885 ;
        RECT -67.485 120.195 -67.155 120.525 ;
        RECT -67.485 118.835 -67.155 119.165 ;
        RECT -67.485 117.475 -67.155 117.805 ;
        RECT -67.485 116.115 -67.155 116.445 ;
        RECT -67.485 114.755 -67.155 115.085 ;
        RECT -67.485 113.395 -67.155 113.725 ;
        RECT -67.485 112.035 -67.155 112.365 ;
        RECT -67.485 110.675 -67.155 111.005 ;
        RECT -67.485 109.315 -67.155 109.645 ;
        RECT -67.485 107.955 -67.155 108.285 ;
        RECT -67.485 106.595 -67.155 106.925 ;
        RECT -67.485 105.235 -67.155 105.565 ;
        RECT -67.485 103.875 -67.155 104.205 ;
        RECT -67.485 102.515 -67.155 102.845 ;
        RECT -67.485 101.155 -67.155 101.485 ;
        RECT -67.485 99.795 -67.155 100.125 ;
        RECT -67.485 98.435 -67.155 98.765 ;
        RECT -67.485 97.075 -67.155 97.405 ;
        RECT -67.485 95.715 -67.155 96.045 ;
        RECT -67.485 94.355 -67.155 94.685 ;
        RECT -67.485 92.995 -67.155 93.325 ;
        RECT -67.485 91.635 -67.155 91.965 ;
        RECT -67.485 90.275 -67.155 90.605 ;
        RECT -67.485 88.915 -67.155 89.245 ;
        RECT -67.485 87.555 -67.155 87.885 ;
        RECT -67.485 86.195 -67.155 86.525 ;
        RECT -67.485 84.835 -67.155 85.165 ;
        RECT -67.485 83.475 -67.155 83.805 ;
        RECT -67.485 82.115 -67.155 82.445 ;
        RECT -67.485 80.755 -67.155 81.085 ;
        RECT -67.485 79.395 -67.155 79.725 ;
        RECT -67.485 78.035 -67.155 78.365 ;
        RECT -67.485 76.675 -67.155 77.005 ;
        RECT -67.485 75.315 -67.155 75.645 ;
        RECT -67.485 73.955 -67.155 74.285 ;
        RECT -67.485 72.595 -67.155 72.925 ;
        RECT -67.485 71.235 -67.155 71.565 ;
        RECT -67.485 69.875 -67.155 70.205 ;
        RECT -67.485 68.515 -67.155 68.845 ;
        RECT -67.485 67.155 -67.155 67.485 ;
        RECT -67.485 65.795 -67.155 66.125 ;
        RECT -67.485 64.435 -67.155 64.765 ;
        RECT -67.485 63.075 -67.155 63.405 ;
        RECT -67.485 61.715 -67.155 62.045 ;
        RECT -67.485 60.355 -67.155 60.685 ;
        RECT -67.485 58.995 -67.155 59.325 ;
        RECT -67.485 57.635 -67.155 57.965 ;
        RECT -67.485 56.275 -67.155 56.605 ;
        RECT -67.485 54.915 -67.155 55.245 ;
        RECT -67.485 53.555 -67.155 53.885 ;
        RECT -67.485 52.195 -67.155 52.525 ;
        RECT -67.485 50.835 -67.155 51.165 ;
        RECT -67.485 49.475 -67.155 49.805 ;
        RECT -67.485 48.115 -67.155 48.445 ;
        RECT -67.485 46.755 -67.155 47.085 ;
        RECT -67.485 45.395 -67.155 45.725 ;
        RECT -67.485 44.035 -67.155 44.365 ;
        RECT -67.485 42.675 -67.155 43.005 ;
        RECT -67.485 41.315 -67.155 41.645 ;
        RECT -67.485 39.955 -67.155 40.285 ;
        RECT -67.485 38.595 -67.155 38.925 ;
        RECT -67.485 37.235 -67.155 37.565 ;
        RECT -67.485 35.875 -67.155 36.205 ;
        RECT -67.485 34.515 -67.155 34.845 ;
        RECT -67.485 33.155 -67.155 33.485 ;
        RECT -67.485 31.795 -67.155 32.125 ;
        RECT -67.485 30.435 -67.155 30.765 ;
        RECT -67.485 29.075 -67.155 29.405 ;
        RECT -67.485 27.715 -67.155 28.045 ;
        RECT -67.485 26.355 -67.155 26.685 ;
        RECT -67.485 24.995 -67.155 25.325 ;
        RECT -67.485 23.635 -67.155 23.965 ;
        RECT -67.485 22.275 -67.155 22.605 ;
        RECT -67.485 20.915 -67.155 21.245 ;
        RECT -67.485 19.555 -67.155 19.885 ;
        RECT -67.485 18.195 -67.155 18.525 ;
        RECT -67.485 16.835 -67.155 17.165 ;
        RECT -67.485 15.475 -67.155 15.805 ;
        RECT -67.485 14.115 -67.155 14.445 ;
        RECT -67.485 12.755 -67.155 13.085 ;
        RECT -67.485 11.395 -67.155 11.725 ;
        RECT -67.485 10.035 -67.155 10.365 ;
        RECT -67.485 8.675 -67.155 9.005 ;
        RECT -67.485 7.315 -67.155 7.645 ;
        RECT -67.485 5.955 -67.155 6.285 ;
        RECT -67.485 4.595 -67.155 4.925 ;
        RECT -67.485 3.235 -67.155 3.565 ;
        RECT -67.485 1.875 -67.155 2.205 ;
        RECT -67.485 0.515 -67.155 0.845 ;
        RECT -67.485 -0.845 -67.155 -0.515 ;
        RECT -67.485 -2.205 -67.155 -1.875 ;
        RECT -67.485 -3.565 -67.155 -3.235 ;
        RECT -67.485 -4.925 -67.155 -4.595 ;
        RECT -67.485 -6.285 -67.155 -5.955 ;
        RECT -67.485 -7.645 -67.155 -7.315 ;
        RECT -67.485 -9.005 -67.155 -8.675 ;
        RECT -67.485 -10.365 -67.155 -10.035 ;
        RECT -67.485 -11.725 -67.155 -11.395 ;
        RECT -67.485 -13.085 -67.155 -12.755 ;
        RECT -67.485 -14.445 -67.155 -14.115 ;
        RECT -67.485 -15.805 -67.155 -15.475 ;
        RECT -67.485 -17.165 -67.155 -16.835 ;
        RECT -67.485 -18.525 -67.155 -18.195 ;
        RECT -67.485 -19.885 -67.155 -19.555 ;
        RECT -67.485 -21.245 -67.155 -20.915 ;
        RECT -67.485 -22.605 -67.155 -22.275 ;
        RECT -67.485 -23.965 -67.155 -23.635 ;
        RECT -67.485 -25.325 -67.155 -24.995 ;
        RECT -67.485 -26.685 -67.155 -26.355 ;
        RECT -67.485 -28.045 -67.155 -27.715 ;
        RECT -67.485 -29.405 -67.155 -29.075 ;
        RECT -67.485 -30.765 -67.155 -30.435 ;
        RECT -67.485 -32.125 -67.155 -31.795 ;
        RECT -67.485 -33.485 -67.155 -33.155 ;
        RECT -67.485 -34.845 -67.155 -34.515 ;
        RECT -67.485 -36.205 -67.155 -35.875 ;
        RECT -67.485 -37.565 -67.155 -37.235 ;
        RECT -67.485 -38.925 -67.155 -38.595 ;
        RECT -67.485 -40.285 -67.155 -39.955 ;
        RECT -67.485 -41.645 -67.155 -41.315 ;
        RECT -67.485 -43.005 -67.155 -42.675 ;
        RECT -67.485 -44.365 -67.155 -44.035 ;
        RECT -67.485 -45.725 -67.155 -45.395 ;
        RECT -67.485 -47.085 -67.155 -46.755 ;
        RECT -67.485 -48.445 -67.155 -48.115 ;
        RECT -67.485 -49.805 -67.155 -49.475 ;
        RECT -67.485 -51.165 -67.155 -50.835 ;
        RECT -67.485 -52.525 -67.155 -52.195 ;
        RECT -67.485 -53.885 -67.155 -53.555 ;
        RECT -67.485 -55.245 -67.155 -54.915 ;
        RECT -67.485 -56.605 -67.155 -56.275 ;
        RECT -67.485 -57.965 -67.155 -57.635 ;
        RECT -67.485 -59.325 -67.155 -58.995 ;
        RECT -67.485 -60.685 -67.155 -60.355 ;
        RECT -67.485 -62.045 -67.155 -61.715 ;
        RECT -67.485 -63.405 -67.155 -63.075 ;
        RECT -67.485 -64.765 -67.155 -64.435 ;
        RECT -67.485 -66.125 -67.155 -65.795 ;
        RECT -67.485 -67.485 -67.155 -67.155 ;
        RECT -67.485 -68.845 -67.155 -68.515 ;
        RECT -67.485 -70.205 -67.155 -69.875 ;
        RECT -67.485 -71.565 -67.155 -71.235 ;
        RECT -67.485 -72.925 -67.155 -72.595 ;
        RECT -67.485 -74.285 -67.155 -73.955 ;
        RECT -67.485 -75.645 -67.155 -75.315 ;
        RECT -67.485 -77.005 -67.155 -76.675 ;
        RECT -67.485 -78.365 -67.155 -78.035 ;
        RECT -67.485 -79.725 -67.155 -79.395 ;
        RECT -67.485 -81.085 -67.155 -80.755 ;
        RECT -67.485 -82.445 -67.155 -82.115 ;
        RECT -67.485 -83.805 -67.155 -83.475 ;
        RECT -67.485 -85.165 -67.155 -84.835 ;
        RECT -67.485 -86.525 -67.155 -86.195 ;
        RECT -67.485 -87.885 -67.155 -87.555 ;
        RECT -67.485 -89.245 -67.155 -88.915 ;
        RECT -67.485 -90.605 -67.155 -90.275 ;
        RECT -67.485 -91.965 -67.155 -91.635 ;
        RECT -67.485 -93.325 -67.155 -92.995 ;
        RECT -67.485 -94.685 -67.155 -94.355 ;
        RECT -67.485 -96.045 -67.155 -95.715 ;
        RECT -67.485 -97.405 -67.155 -97.075 ;
        RECT -67.485 -98.765 -67.155 -98.435 ;
        RECT -67.485 -100.125 -67.155 -99.795 ;
        RECT -67.485 -101.485 -67.155 -101.155 ;
        RECT -67.485 -102.845 -67.155 -102.515 ;
        RECT -67.485 -104.205 -67.155 -103.875 ;
        RECT -67.485 -105.565 -67.155 -105.235 ;
        RECT -67.485 -106.925 -67.155 -106.595 ;
        RECT -67.485 -108.285 -67.155 -107.955 ;
        RECT -67.485 -109.645 -67.155 -109.315 ;
        RECT -67.485 -111.005 -67.155 -110.675 ;
        RECT -67.485 -112.365 -67.155 -112.035 ;
        RECT -67.485 -113.725 -67.155 -113.395 ;
        RECT -67.485 -115.085 -67.155 -114.755 ;
        RECT -67.485 -116.445 -67.155 -116.115 ;
        RECT -67.485 -117.805 -67.155 -117.475 ;
        RECT -67.485 -119.165 -67.155 -118.835 ;
        RECT -67.485 -120.525 -67.155 -120.195 ;
        RECT -67.485 -121.885 -67.155 -121.555 ;
        RECT -67.485 -123.245 -67.155 -122.915 ;
        RECT -67.485 -124.605 -67.155 -124.275 ;
        RECT -67.485 -125.965 -67.155 -125.635 ;
        RECT -67.485 -127.325 -67.155 -126.995 ;
        RECT -67.485 -128.685 -67.155 -128.355 ;
        RECT -67.485 -130.045 -67.155 -129.715 ;
        RECT -67.485 -131.405 -67.155 -131.075 ;
        RECT -67.485 -132.765 -67.155 -132.435 ;
        RECT -67.485 -134.125 -67.155 -133.795 ;
        RECT -67.485 -135.485 -67.155 -135.155 ;
        RECT -67.485 -136.845 -67.155 -136.515 ;
        RECT -67.485 -138.205 -67.155 -137.875 ;
        RECT -67.485 -139.565 -67.155 -139.235 ;
        RECT -67.485 -140.925 -67.155 -140.595 ;
        RECT -67.485 -142.285 -67.155 -141.955 ;
        RECT -67.485 -143.645 -67.155 -143.315 ;
        RECT -67.485 -145.005 -67.155 -144.675 ;
        RECT -67.485 -146.365 -67.155 -146.035 ;
        RECT -67.485 -147.725 -67.155 -147.395 ;
        RECT -67.485 -149.085 -67.155 -148.755 ;
        RECT -67.485 -150.445 -67.155 -150.115 ;
        RECT -67.485 -151.805 -67.155 -151.475 ;
        RECT -67.485 -153.165 -67.155 -152.835 ;
        RECT -67.485 -154.525 -67.155 -154.195 ;
        RECT -67.485 -155.885 -67.155 -155.555 ;
        RECT -67.485 -157.245 -67.155 -156.915 ;
        RECT -67.485 -162.89 -67.155 -161.76 ;
        RECT -67.48 -163.005 -67.16 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.125 129.945 -65.795 131.075 ;
        RECT -66.125 125.635 -65.795 125.965 ;
        RECT -66.125 124.275 -65.795 124.605 ;
        RECT -66.125 122.915 -65.795 123.245 ;
        RECT -66.125 121.555 -65.795 121.885 ;
        RECT -66.125 120.195 -65.795 120.525 ;
        RECT -66.125 118.835 -65.795 119.165 ;
        RECT -66.125 117.475 -65.795 117.805 ;
        RECT -66.125 116.115 -65.795 116.445 ;
        RECT -66.125 114.755 -65.795 115.085 ;
        RECT -66.125 113.395 -65.795 113.725 ;
        RECT -66.125 112.035 -65.795 112.365 ;
        RECT -66.125 110.675 -65.795 111.005 ;
        RECT -66.125 109.315 -65.795 109.645 ;
        RECT -66.125 107.955 -65.795 108.285 ;
        RECT -66.125 106.595 -65.795 106.925 ;
        RECT -66.125 105.235 -65.795 105.565 ;
        RECT -66.125 103.875 -65.795 104.205 ;
        RECT -66.125 102.515 -65.795 102.845 ;
        RECT -66.125 101.155 -65.795 101.485 ;
        RECT -66.125 99.795 -65.795 100.125 ;
        RECT -66.125 98.435 -65.795 98.765 ;
        RECT -66.125 97.075 -65.795 97.405 ;
        RECT -66.125 95.715 -65.795 96.045 ;
        RECT -66.125 94.355 -65.795 94.685 ;
        RECT -66.125 92.995 -65.795 93.325 ;
        RECT -66.125 91.635 -65.795 91.965 ;
        RECT -66.125 90.275 -65.795 90.605 ;
        RECT -66.125 88.915 -65.795 89.245 ;
        RECT -66.125 87.555 -65.795 87.885 ;
        RECT -66.125 86.195 -65.795 86.525 ;
        RECT -66.125 84.835 -65.795 85.165 ;
        RECT -66.125 83.475 -65.795 83.805 ;
        RECT -66.125 82.115 -65.795 82.445 ;
        RECT -66.125 80.755 -65.795 81.085 ;
        RECT -66.125 79.395 -65.795 79.725 ;
        RECT -66.125 78.035 -65.795 78.365 ;
        RECT -66.125 76.675 -65.795 77.005 ;
        RECT -66.125 75.315 -65.795 75.645 ;
        RECT -66.125 73.955 -65.795 74.285 ;
        RECT -66.125 72.595 -65.795 72.925 ;
        RECT -66.125 71.235 -65.795 71.565 ;
        RECT -66.125 69.875 -65.795 70.205 ;
        RECT -66.125 68.515 -65.795 68.845 ;
        RECT -66.125 67.155 -65.795 67.485 ;
        RECT -66.125 65.795 -65.795 66.125 ;
        RECT -66.125 64.435 -65.795 64.765 ;
        RECT -66.125 63.075 -65.795 63.405 ;
        RECT -66.125 61.715 -65.795 62.045 ;
        RECT -66.125 60.355 -65.795 60.685 ;
        RECT -66.125 58.995 -65.795 59.325 ;
        RECT -66.125 57.635 -65.795 57.965 ;
        RECT -66.125 56.275 -65.795 56.605 ;
        RECT -66.125 54.915 -65.795 55.245 ;
        RECT -66.125 53.555 -65.795 53.885 ;
        RECT -66.125 52.195 -65.795 52.525 ;
        RECT -66.125 50.835 -65.795 51.165 ;
        RECT -66.125 49.475 -65.795 49.805 ;
        RECT -66.125 48.115 -65.795 48.445 ;
        RECT -66.125 46.755 -65.795 47.085 ;
        RECT -66.125 45.395 -65.795 45.725 ;
        RECT -66.125 44.035 -65.795 44.365 ;
        RECT -66.125 42.675 -65.795 43.005 ;
        RECT -66.125 41.315 -65.795 41.645 ;
        RECT -66.125 39.955 -65.795 40.285 ;
        RECT -66.125 38.595 -65.795 38.925 ;
        RECT -66.125 37.235 -65.795 37.565 ;
        RECT -66.125 35.875 -65.795 36.205 ;
        RECT -66.125 34.515 -65.795 34.845 ;
        RECT -66.125 33.155 -65.795 33.485 ;
        RECT -66.125 31.795 -65.795 32.125 ;
        RECT -66.125 30.435 -65.795 30.765 ;
        RECT -66.125 29.075 -65.795 29.405 ;
        RECT -66.125 27.715 -65.795 28.045 ;
        RECT -66.125 26.355 -65.795 26.685 ;
        RECT -66.125 24.995 -65.795 25.325 ;
        RECT -66.125 23.635 -65.795 23.965 ;
        RECT -66.125 22.275 -65.795 22.605 ;
        RECT -66.125 20.915 -65.795 21.245 ;
        RECT -66.125 19.555 -65.795 19.885 ;
        RECT -66.125 18.195 -65.795 18.525 ;
        RECT -66.125 16.835 -65.795 17.165 ;
        RECT -66.125 15.475 -65.795 15.805 ;
        RECT -66.125 14.115 -65.795 14.445 ;
        RECT -66.125 12.755 -65.795 13.085 ;
        RECT -66.125 11.395 -65.795 11.725 ;
        RECT -66.125 10.035 -65.795 10.365 ;
        RECT -66.125 8.675 -65.795 9.005 ;
        RECT -66.125 7.315 -65.795 7.645 ;
        RECT -66.125 5.955 -65.795 6.285 ;
        RECT -66.125 4.595 -65.795 4.925 ;
        RECT -66.125 3.235 -65.795 3.565 ;
        RECT -66.125 1.875 -65.795 2.205 ;
        RECT -66.125 0.515 -65.795 0.845 ;
        RECT -66.125 -0.845 -65.795 -0.515 ;
        RECT -66.125 -2.205 -65.795 -1.875 ;
        RECT -66.125 -3.565 -65.795 -3.235 ;
        RECT -66.125 -4.925 -65.795 -4.595 ;
        RECT -66.125 -6.285 -65.795 -5.955 ;
        RECT -66.125 -7.645 -65.795 -7.315 ;
        RECT -66.125 -9.005 -65.795 -8.675 ;
        RECT -66.125 -10.365 -65.795 -10.035 ;
        RECT -66.125 -11.725 -65.795 -11.395 ;
        RECT -66.125 -13.085 -65.795 -12.755 ;
        RECT -66.125 -14.445 -65.795 -14.115 ;
        RECT -66.125 -15.805 -65.795 -15.475 ;
        RECT -66.125 -17.165 -65.795 -16.835 ;
        RECT -66.125 -18.525 -65.795 -18.195 ;
        RECT -66.125 -19.885 -65.795 -19.555 ;
        RECT -66.125 -21.245 -65.795 -20.915 ;
        RECT -66.125 -22.605 -65.795 -22.275 ;
        RECT -66.125 -23.965 -65.795 -23.635 ;
        RECT -66.125 -25.325 -65.795 -24.995 ;
        RECT -66.125 -26.685 -65.795 -26.355 ;
        RECT -66.125 -28.045 -65.795 -27.715 ;
        RECT -66.125 -29.405 -65.795 -29.075 ;
        RECT -66.125 -30.765 -65.795 -30.435 ;
        RECT -66.125 -32.125 -65.795 -31.795 ;
        RECT -66.125 -33.485 -65.795 -33.155 ;
        RECT -66.125 -34.845 -65.795 -34.515 ;
        RECT -66.125 -36.205 -65.795 -35.875 ;
        RECT -66.125 -37.565 -65.795 -37.235 ;
        RECT -66.125 -38.925 -65.795 -38.595 ;
        RECT -66.125 -40.285 -65.795 -39.955 ;
        RECT -66.125 -41.645 -65.795 -41.315 ;
        RECT -66.125 -43.005 -65.795 -42.675 ;
        RECT -66.125 -44.365 -65.795 -44.035 ;
        RECT -66.125 -45.725 -65.795 -45.395 ;
        RECT -66.125 -47.085 -65.795 -46.755 ;
        RECT -66.125 -48.445 -65.795 -48.115 ;
        RECT -66.125 -49.805 -65.795 -49.475 ;
        RECT -66.125 -51.165 -65.795 -50.835 ;
        RECT -66.125 -52.525 -65.795 -52.195 ;
        RECT -66.125 -53.885 -65.795 -53.555 ;
        RECT -66.125 -55.245 -65.795 -54.915 ;
        RECT -66.125 -56.605 -65.795 -56.275 ;
        RECT -66.125 -57.965 -65.795 -57.635 ;
        RECT -66.125 -59.325 -65.795 -58.995 ;
        RECT -66.125 -60.685 -65.795 -60.355 ;
        RECT -66.125 -62.045 -65.795 -61.715 ;
        RECT -66.125 -63.405 -65.795 -63.075 ;
        RECT -66.125 -64.765 -65.795 -64.435 ;
        RECT -66.125 -66.125 -65.795 -65.795 ;
        RECT -66.125 -67.485 -65.795 -67.155 ;
        RECT -66.125 -68.845 -65.795 -68.515 ;
        RECT -66.125 -70.205 -65.795 -69.875 ;
        RECT -66.125 -71.565 -65.795 -71.235 ;
        RECT -66.125 -72.925 -65.795 -72.595 ;
        RECT -66.125 -74.285 -65.795 -73.955 ;
        RECT -66.125 -75.645 -65.795 -75.315 ;
        RECT -66.125 -77.005 -65.795 -76.675 ;
        RECT -66.125 -78.365 -65.795 -78.035 ;
        RECT -66.125 -79.725 -65.795 -79.395 ;
        RECT -66.125 -81.085 -65.795 -80.755 ;
        RECT -66.125 -82.445 -65.795 -82.115 ;
        RECT -66.125 -83.805 -65.795 -83.475 ;
        RECT -66.125 -85.165 -65.795 -84.835 ;
        RECT -66.125 -86.525 -65.795 -86.195 ;
        RECT -66.125 -87.885 -65.795 -87.555 ;
        RECT -66.125 -89.245 -65.795 -88.915 ;
        RECT -66.125 -90.605 -65.795 -90.275 ;
        RECT -66.125 -91.965 -65.795 -91.635 ;
        RECT -66.125 -93.325 -65.795 -92.995 ;
        RECT -66.125 -94.685 -65.795 -94.355 ;
        RECT -66.125 -96.045 -65.795 -95.715 ;
        RECT -66.125 -97.405 -65.795 -97.075 ;
        RECT -66.125 -98.765 -65.795 -98.435 ;
        RECT -66.125 -100.125 -65.795 -99.795 ;
        RECT -66.125 -101.485 -65.795 -101.155 ;
        RECT -66.125 -102.845 -65.795 -102.515 ;
        RECT -66.125 -104.205 -65.795 -103.875 ;
        RECT -66.125 -105.565 -65.795 -105.235 ;
        RECT -66.125 -106.925 -65.795 -106.595 ;
        RECT -66.125 -108.285 -65.795 -107.955 ;
        RECT -66.125 -109.645 -65.795 -109.315 ;
        RECT -66.125 -111.005 -65.795 -110.675 ;
        RECT -66.125 -112.365 -65.795 -112.035 ;
        RECT -66.125 -113.725 -65.795 -113.395 ;
        RECT -66.125 -115.085 -65.795 -114.755 ;
        RECT -66.125 -116.445 -65.795 -116.115 ;
        RECT -66.125 -117.805 -65.795 -117.475 ;
        RECT -66.125 -119.165 -65.795 -118.835 ;
        RECT -66.125 -120.525 -65.795 -120.195 ;
        RECT -66.125 -121.885 -65.795 -121.555 ;
        RECT -66.125 -123.245 -65.795 -122.915 ;
        RECT -66.125 -124.605 -65.795 -124.275 ;
        RECT -66.125 -125.965 -65.795 -125.635 ;
        RECT -66.125 -127.325 -65.795 -126.995 ;
        RECT -66.125 -128.685 -65.795 -128.355 ;
        RECT -66.125 -130.045 -65.795 -129.715 ;
        RECT -66.125 -131.405 -65.795 -131.075 ;
        RECT -66.125 -132.765 -65.795 -132.435 ;
        RECT -66.125 -134.125 -65.795 -133.795 ;
        RECT -66.125 -135.485 -65.795 -135.155 ;
        RECT -66.125 -136.845 -65.795 -136.515 ;
        RECT -66.125 -138.205 -65.795 -137.875 ;
        RECT -66.125 -139.565 -65.795 -139.235 ;
        RECT -66.125 -140.925 -65.795 -140.595 ;
        RECT -66.125 -142.285 -65.795 -141.955 ;
        RECT -66.125 -143.645 -65.795 -143.315 ;
        RECT -66.125 -145.005 -65.795 -144.675 ;
        RECT -66.125 -146.365 -65.795 -146.035 ;
        RECT -66.125 -147.725 -65.795 -147.395 ;
        RECT -66.125 -149.085 -65.795 -148.755 ;
        RECT -66.125 -150.445 -65.795 -150.115 ;
        RECT -66.125 -151.805 -65.795 -151.475 ;
        RECT -66.125 -153.165 -65.795 -152.835 ;
        RECT -66.125 -154.525 -65.795 -154.195 ;
        RECT -66.125 -155.885 -65.795 -155.555 ;
        RECT -66.125 -157.245 -65.795 -156.915 ;
        RECT -66.125 -162.89 -65.795 -161.76 ;
        RECT -66.12 -163.005 -65.8 131.19 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.765 -97.405 -64.435 -97.075 ;
        RECT -64.765 -98.765 -64.435 -98.435 ;
        RECT -64.765 -100.125 -64.435 -99.795 ;
        RECT -64.765 -101.485 -64.435 -101.155 ;
        RECT -64.765 -102.845 -64.435 -102.515 ;
        RECT -64.765 -104.205 -64.435 -103.875 ;
        RECT -64.765 -105.565 -64.435 -105.235 ;
        RECT -64.765 -106.925 -64.435 -106.595 ;
        RECT -64.765 -108.285 -64.435 -107.955 ;
        RECT -64.765 -109.645 -64.435 -109.315 ;
        RECT -64.765 -111.005 -64.435 -110.675 ;
        RECT -64.765 -112.365 -64.435 -112.035 ;
        RECT -64.765 -113.725 -64.435 -113.395 ;
        RECT -64.765 -115.085 -64.435 -114.755 ;
        RECT -64.765 -116.445 -64.435 -116.115 ;
        RECT -64.765 -117.805 -64.435 -117.475 ;
        RECT -64.765 -119.165 -64.435 -118.835 ;
        RECT -64.765 -120.525 -64.435 -120.195 ;
        RECT -64.765 -121.885 -64.435 -121.555 ;
        RECT -64.765 -123.245 -64.435 -122.915 ;
        RECT -64.765 -124.605 -64.435 -124.275 ;
        RECT -64.765 -125.965 -64.435 -125.635 ;
        RECT -64.765 -127.325 -64.435 -126.995 ;
        RECT -64.765 -128.685 -64.435 -128.355 ;
        RECT -64.765 -130.045 -64.435 -129.715 ;
        RECT -64.765 -131.405 -64.435 -131.075 ;
        RECT -64.765 -132.765 -64.435 -132.435 ;
        RECT -64.765 -134.125 -64.435 -133.795 ;
        RECT -64.765 -135.485 -64.435 -135.155 ;
        RECT -64.765 -136.845 -64.435 -136.515 ;
        RECT -64.765 -138.205 -64.435 -137.875 ;
        RECT -64.765 -139.565 -64.435 -139.235 ;
        RECT -64.765 -140.925 -64.435 -140.595 ;
        RECT -64.765 -142.285 -64.435 -141.955 ;
        RECT -64.765 -143.645 -64.435 -143.315 ;
        RECT -64.765 -145.005 -64.435 -144.675 ;
        RECT -64.765 -146.365 -64.435 -146.035 ;
        RECT -64.765 -148.215 -64.435 -147.885 ;
        RECT -64.765 -149.085 -64.435 -148.755 ;
        RECT -64.765 -150.445 -64.435 -150.115 ;
        RECT -64.765 -151.805 -64.435 -151.475 ;
        RECT -64.76 -151.805 -64.44 131.19 ;
        RECT -64.765 129.945 -64.435 131.075 ;
        RECT -64.765 125.635 -64.435 125.965 ;
        RECT -64.765 124.275 -64.435 124.605 ;
        RECT -64.765 122.915 -64.435 123.245 ;
        RECT -64.765 121.555 -64.435 121.885 ;
        RECT -64.765 120.195 -64.435 120.525 ;
        RECT -64.765 118.835 -64.435 119.165 ;
        RECT -64.765 117.475 -64.435 117.805 ;
        RECT -64.765 116.115 -64.435 116.445 ;
        RECT -64.765 114.755 -64.435 115.085 ;
        RECT -64.765 113.395 -64.435 113.725 ;
        RECT -64.765 112.035 -64.435 112.365 ;
        RECT -64.765 110.675 -64.435 111.005 ;
        RECT -64.765 109.315 -64.435 109.645 ;
        RECT -64.765 107.955 -64.435 108.285 ;
        RECT -64.765 106.595 -64.435 106.925 ;
        RECT -64.765 105.235 -64.435 105.565 ;
        RECT -64.765 103.875 -64.435 104.205 ;
        RECT -64.765 102.515 -64.435 102.845 ;
        RECT -64.765 101.155 -64.435 101.485 ;
        RECT -64.765 99.795 -64.435 100.125 ;
        RECT -64.765 98.435 -64.435 98.765 ;
        RECT -64.765 97.075 -64.435 97.405 ;
        RECT -64.765 95.715 -64.435 96.045 ;
        RECT -64.765 94.355 -64.435 94.685 ;
        RECT -64.765 92.995 -64.435 93.325 ;
        RECT -64.765 91.635 -64.435 91.965 ;
        RECT -64.765 90.275 -64.435 90.605 ;
        RECT -64.765 88.915 -64.435 89.245 ;
        RECT -64.765 87.555 -64.435 87.885 ;
        RECT -64.765 86.195 -64.435 86.525 ;
        RECT -64.765 84.835 -64.435 85.165 ;
        RECT -64.765 83.475 -64.435 83.805 ;
        RECT -64.765 82.115 -64.435 82.445 ;
        RECT -64.765 80.755 -64.435 81.085 ;
        RECT -64.765 79.395 -64.435 79.725 ;
        RECT -64.765 78.035 -64.435 78.365 ;
        RECT -64.765 76.675 -64.435 77.005 ;
        RECT -64.765 75.315 -64.435 75.645 ;
        RECT -64.765 73.955 -64.435 74.285 ;
        RECT -64.765 72.595 -64.435 72.925 ;
        RECT -64.765 71.235 -64.435 71.565 ;
        RECT -64.765 69.875 -64.435 70.205 ;
        RECT -64.765 68.515 -64.435 68.845 ;
        RECT -64.765 67.155 -64.435 67.485 ;
        RECT -64.765 65.795 -64.435 66.125 ;
        RECT -64.765 64.435 -64.435 64.765 ;
        RECT -64.765 63.075 -64.435 63.405 ;
        RECT -64.765 61.715 -64.435 62.045 ;
        RECT -64.765 60.355 -64.435 60.685 ;
        RECT -64.765 58.995 -64.435 59.325 ;
        RECT -64.765 57.635 -64.435 57.965 ;
        RECT -64.765 56.275 -64.435 56.605 ;
        RECT -64.765 54.915 -64.435 55.245 ;
        RECT -64.765 53.555 -64.435 53.885 ;
        RECT -64.765 52.195 -64.435 52.525 ;
        RECT -64.765 50.835 -64.435 51.165 ;
        RECT -64.765 49.475 -64.435 49.805 ;
        RECT -64.765 48.115 -64.435 48.445 ;
        RECT -64.765 46.755 -64.435 47.085 ;
        RECT -64.765 45.395 -64.435 45.725 ;
        RECT -64.765 44.035 -64.435 44.365 ;
        RECT -64.765 42.675 -64.435 43.005 ;
        RECT -64.765 41.315 -64.435 41.645 ;
        RECT -64.765 39.955 -64.435 40.285 ;
        RECT -64.765 38.595 -64.435 38.925 ;
        RECT -64.765 37.235 -64.435 37.565 ;
        RECT -64.765 35.875 -64.435 36.205 ;
        RECT -64.765 34.515 -64.435 34.845 ;
        RECT -64.765 33.155 -64.435 33.485 ;
        RECT -64.765 31.795 -64.435 32.125 ;
        RECT -64.765 30.435 -64.435 30.765 ;
        RECT -64.765 29.075 -64.435 29.405 ;
        RECT -64.765 27.715 -64.435 28.045 ;
        RECT -64.765 26.355 -64.435 26.685 ;
        RECT -64.765 24.995 -64.435 25.325 ;
        RECT -64.765 23.635 -64.435 23.965 ;
        RECT -64.765 22.275 -64.435 22.605 ;
        RECT -64.765 20.915 -64.435 21.245 ;
        RECT -64.765 19.555 -64.435 19.885 ;
        RECT -64.765 18.195 -64.435 18.525 ;
        RECT -64.765 16.835 -64.435 17.165 ;
        RECT -64.765 15.475 -64.435 15.805 ;
        RECT -64.765 14.115 -64.435 14.445 ;
        RECT -64.765 12.755 -64.435 13.085 ;
        RECT -64.765 11.395 -64.435 11.725 ;
        RECT -64.765 10.035 -64.435 10.365 ;
        RECT -64.765 8.675 -64.435 9.005 ;
        RECT -64.765 7.315 -64.435 7.645 ;
        RECT -64.765 5.955 -64.435 6.285 ;
        RECT -64.765 4.595 -64.435 4.925 ;
        RECT -64.765 3.235 -64.435 3.565 ;
        RECT -64.765 1.875 -64.435 2.205 ;
        RECT -64.765 0.515 -64.435 0.845 ;
        RECT -64.765 -0.845 -64.435 -0.515 ;
        RECT -64.765 -2.205 -64.435 -1.875 ;
        RECT -64.765 -3.565 -64.435 -3.235 ;
        RECT -64.765 -4.925 -64.435 -4.595 ;
        RECT -64.765 -6.285 -64.435 -5.955 ;
        RECT -64.765 -7.645 -64.435 -7.315 ;
        RECT -64.765 -9.005 -64.435 -8.675 ;
        RECT -64.765 -10.365 -64.435 -10.035 ;
        RECT -64.765 -11.725 -64.435 -11.395 ;
        RECT -64.765 -13.085 -64.435 -12.755 ;
        RECT -64.765 -14.445 -64.435 -14.115 ;
        RECT -64.765 -15.805 -64.435 -15.475 ;
        RECT -64.765 -17.165 -64.435 -16.835 ;
        RECT -64.765 -18.525 -64.435 -18.195 ;
        RECT -64.765 -19.885 -64.435 -19.555 ;
        RECT -64.765 -21.245 -64.435 -20.915 ;
        RECT -64.765 -22.605 -64.435 -22.275 ;
        RECT -64.765 -23.965 -64.435 -23.635 ;
        RECT -64.765 -25.325 -64.435 -24.995 ;
        RECT -64.765 -26.685 -64.435 -26.355 ;
        RECT -64.765 -28.045 -64.435 -27.715 ;
        RECT -64.765 -29.405 -64.435 -29.075 ;
        RECT -64.765 -30.765 -64.435 -30.435 ;
        RECT -64.765 -32.125 -64.435 -31.795 ;
        RECT -64.765 -33.485 -64.435 -33.155 ;
        RECT -64.765 -34.845 -64.435 -34.515 ;
        RECT -64.765 -36.205 -64.435 -35.875 ;
        RECT -64.765 -37.565 -64.435 -37.235 ;
        RECT -64.765 -38.925 -64.435 -38.595 ;
        RECT -64.765 -40.285 -64.435 -39.955 ;
        RECT -64.765 -41.645 -64.435 -41.315 ;
        RECT -64.765 -43.005 -64.435 -42.675 ;
        RECT -64.765 -44.365 -64.435 -44.035 ;
        RECT -64.765 -45.725 -64.435 -45.395 ;
        RECT -64.765 -47.085 -64.435 -46.755 ;
        RECT -64.765 -48.445 -64.435 -48.115 ;
        RECT -64.765 -49.805 -64.435 -49.475 ;
        RECT -64.765 -51.165 -64.435 -50.835 ;
        RECT -64.765 -52.525 -64.435 -52.195 ;
        RECT -64.765 -53.885 -64.435 -53.555 ;
        RECT -64.765 -55.245 -64.435 -54.915 ;
        RECT -64.765 -56.605 -64.435 -56.275 ;
        RECT -64.765 -57.965 -64.435 -57.635 ;
        RECT -64.765 -59.325 -64.435 -58.995 ;
        RECT -64.765 -60.685 -64.435 -60.355 ;
        RECT -64.765 -62.045 -64.435 -61.715 ;
        RECT -64.765 -63.405 -64.435 -63.075 ;
        RECT -64.765 -64.765 -64.435 -64.435 ;
        RECT -64.765 -66.125 -64.435 -65.795 ;
        RECT -64.765 -67.485 -64.435 -67.155 ;
        RECT -64.765 -68.845 -64.435 -68.515 ;
        RECT -64.765 -70.205 -64.435 -69.875 ;
        RECT -64.765 -71.565 -64.435 -71.235 ;
        RECT -64.765 -72.925 -64.435 -72.595 ;
        RECT -64.765 -74.285 -64.435 -73.955 ;
        RECT -64.765 -75.645 -64.435 -75.315 ;
        RECT -64.765 -77.005 -64.435 -76.675 ;
        RECT -64.765 -78.365 -64.435 -78.035 ;
        RECT -64.765 -79.725 -64.435 -79.395 ;
        RECT -64.765 -81.085 -64.435 -80.755 ;
        RECT -64.765 -82.445 -64.435 -82.115 ;
        RECT -64.765 -83.805 -64.435 -83.475 ;
        RECT -64.765 -85.165 -64.435 -84.835 ;
        RECT -64.765 -86.525 -64.435 -86.195 ;
        RECT -64.765 -87.885 -64.435 -87.555 ;
        RECT -64.765 -89.245 -64.435 -88.915 ;
        RECT -64.765 -90.605 -64.435 -90.275 ;
        RECT -64.765 -91.965 -64.435 -91.635 ;
        RECT -64.765 -93.325 -64.435 -92.995 ;
        RECT -64.765 -94.685 -64.435 -94.355 ;
        RECT -64.765 -96.045 -64.435 -95.715 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 197.86 -94.075 198.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 127.225 198.725 128.355 ;
        RECT 198.395 124.955 198.725 125.285 ;
        RECT 198.395 123.595 198.725 123.925 ;
        RECT 198.4 123.595 198.72 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 -95.365 198.725 -95.035 ;
        RECT 198.395 -96.725 198.725 -96.395 ;
        RECT 198.395 -98.085 198.725 -97.755 ;
        RECT 198.395 -99.445 198.725 -99.115 ;
        RECT 198.395 -100.805 198.725 -100.475 ;
        RECT 198.395 -102.165 198.725 -101.835 ;
        RECT 198.395 -103.525 198.725 -103.195 ;
        RECT 198.395 -104.885 198.725 -104.555 ;
        RECT 198.395 -106.245 198.725 -105.915 ;
        RECT 198.395 -107.605 198.725 -107.275 ;
        RECT 198.395 -108.965 198.725 -108.635 ;
        RECT 198.395 -110.325 198.725 -109.995 ;
        RECT 198.395 -111.685 198.725 -111.355 ;
        RECT 198.395 -113.045 198.725 -112.715 ;
        RECT 198.395 -114.405 198.725 -114.075 ;
        RECT 198.395 -115.765 198.725 -115.435 ;
        RECT 198.395 -117.125 198.725 -116.795 ;
        RECT 198.395 -118.485 198.725 -118.155 ;
        RECT 198.395 -119.845 198.725 -119.515 ;
        RECT 198.395 -121.205 198.725 -120.875 ;
        RECT 198.395 -122.565 198.725 -122.235 ;
        RECT 198.395 -123.925 198.725 -123.595 ;
        RECT 198.395 -125.285 198.725 -124.955 ;
        RECT 198.395 -126.645 198.725 -126.315 ;
        RECT 198.395 -128.005 198.725 -127.675 ;
        RECT 198.395 -129.365 198.725 -129.035 ;
        RECT 198.395 -130.725 198.725 -130.395 ;
        RECT 198.395 -132.085 198.725 -131.755 ;
        RECT 198.395 -133.445 198.725 -133.115 ;
        RECT 198.395 -134.805 198.725 -134.475 ;
        RECT 198.395 -136.165 198.725 -135.835 ;
        RECT 198.395 -137.525 198.725 -137.195 ;
        RECT 198.395 -138.885 198.725 -138.555 ;
        RECT 198.395 -140.245 198.725 -139.915 ;
        RECT 198.395 -141.605 198.725 -141.275 ;
        RECT 198.395 -142.965 198.725 -142.635 ;
        RECT 198.395 -144.325 198.725 -143.995 ;
        RECT 198.395 -145.685 198.725 -145.355 ;
        RECT 198.395 -147.045 198.725 -146.715 ;
        RECT 198.395 -148.405 198.725 -148.075 ;
        RECT 198.395 -149.765 198.725 -149.435 ;
        RECT 198.395 -151.125 198.725 -150.795 ;
        RECT 198.395 -152.485 198.725 -152.155 ;
        RECT 198.395 -153.845 198.725 -153.515 ;
        RECT 198.395 -155.205 198.725 -154.875 ;
        RECT 198.395 -156.565 198.725 -156.235 ;
        RECT 198.395 -157.925 198.725 -157.595 ;
        RECT 198.395 -160.17 198.725 -159.04 ;
        RECT 198.4 -160.285 198.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 127.225 200.085 128.355 ;
        RECT 199.755 124.955 200.085 125.285 ;
        RECT 199.755 123.595 200.085 123.925 ;
        RECT 199.76 123.595 200.08 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 -1.525 200.085 -1.195 ;
        RECT 199.755 -2.885 200.085 -2.555 ;
        RECT 199.76 -3.56 200.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 -91.285 200.085 -90.955 ;
        RECT 199.755 -92.645 200.085 -92.315 ;
        RECT 199.755 -94.005 200.085 -93.675 ;
        RECT 199.755 -95.365 200.085 -95.035 ;
        RECT 199.755 -96.725 200.085 -96.395 ;
        RECT 199.755 -98.085 200.085 -97.755 ;
        RECT 199.755 -99.445 200.085 -99.115 ;
        RECT 199.755 -100.805 200.085 -100.475 ;
        RECT 199.755 -102.165 200.085 -101.835 ;
        RECT 199.755 -103.525 200.085 -103.195 ;
        RECT 199.755 -104.885 200.085 -104.555 ;
        RECT 199.755 -106.245 200.085 -105.915 ;
        RECT 199.755 -107.605 200.085 -107.275 ;
        RECT 199.755 -108.965 200.085 -108.635 ;
        RECT 199.755 -110.325 200.085 -109.995 ;
        RECT 199.755 -111.685 200.085 -111.355 ;
        RECT 199.755 -113.045 200.085 -112.715 ;
        RECT 199.755 -114.405 200.085 -114.075 ;
        RECT 199.755 -115.765 200.085 -115.435 ;
        RECT 199.755 -117.125 200.085 -116.795 ;
        RECT 199.755 -118.485 200.085 -118.155 ;
        RECT 199.755 -119.845 200.085 -119.515 ;
        RECT 199.755 -121.205 200.085 -120.875 ;
        RECT 199.755 -122.565 200.085 -122.235 ;
        RECT 199.755 -123.925 200.085 -123.595 ;
        RECT 199.755 -125.285 200.085 -124.955 ;
        RECT 199.755 -126.645 200.085 -126.315 ;
        RECT 199.755 -128.005 200.085 -127.675 ;
        RECT 199.755 -129.365 200.085 -129.035 ;
        RECT 199.755 -130.725 200.085 -130.395 ;
        RECT 199.755 -132.085 200.085 -131.755 ;
        RECT 199.755 -133.445 200.085 -133.115 ;
        RECT 199.755 -134.805 200.085 -134.475 ;
        RECT 199.755 -136.165 200.085 -135.835 ;
        RECT 199.755 -137.525 200.085 -137.195 ;
        RECT 199.755 -138.885 200.085 -138.555 ;
        RECT 199.755 -140.245 200.085 -139.915 ;
        RECT 199.755 -141.605 200.085 -141.275 ;
        RECT 199.755 -142.965 200.085 -142.635 ;
        RECT 199.755 -144.325 200.085 -143.995 ;
        RECT 199.755 -145.685 200.085 -145.355 ;
        RECT 199.755 -147.045 200.085 -146.715 ;
        RECT 199.755 -148.405 200.085 -148.075 ;
        RECT 199.755 -149.765 200.085 -149.435 ;
        RECT 199.755 -151.125 200.085 -150.795 ;
        RECT 199.755 -152.485 200.085 -152.155 ;
        RECT 199.755 -153.845 200.085 -153.515 ;
        RECT 199.755 -155.205 200.085 -154.875 ;
        RECT 199.755 -156.565 200.085 -156.235 ;
        RECT 199.755 -157.925 200.085 -157.595 ;
        RECT 199.755 -160.17 200.085 -159.04 ;
        RECT 199.76 -160.285 200.08 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 127.225 201.445 128.355 ;
        RECT 201.115 124.955 201.445 125.285 ;
        RECT 201.115 123.595 201.445 123.925 ;
        RECT 201.12 123.595 201.44 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -1.525 201.445 -1.195 ;
        RECT 201.115 -2.885 201.445 -2.555 ;
        RECT 201.12 -3.56 201.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -91.285 201.445 -90.955 ;
        RECT 201.115 -92.645 201.445 -92.315 ;
        RECT 201.115 -94.005 201.445 -93.675 ;
        RECT 201.115 -95.365 201.445 -95.035 ;
        RECT 201.115 -96.725 201.445 -96.395 ;
        RECT 201.115 -98.085 201.445 -97.755 ;
        RECT 201.115 -99.445 201.445 -99.115 ;
        RECT 201.115 -100.805 201.445 -100.475 ;
        RECT 201.115 -102.165 201.445 -101.835 ;
        RECT 201.115 -103.525 201.445 -103.195 ;
        RECT 201.115 -104.885 201.445 -104.555 ;
        RECT 201.115 -106.245 201.445 -105.915 ;
        RECT 201.115 -107.605 201.445 -107.275 ;
        RECT 201.115 -108.965 201.445 -108.635 ;
        RECT 201.115 -110.325 201.445 -109.995 ;
        RECT 201.115 -111.685 201.445 -111.355 ;
        RECT 201.115 -113.045 201.445 -112.715 ;
        RECT 201.115 -114.405 201.445 -114.075 ;
        RECT 201.115 -115.765 201.445 -115.435 ;
        RECT 201.115 -117.125 201.445 -116.795 ;
        RECT 201.115 -118.485 201.445 -118.155 ;
        RECT 201.115 -119.845 201.445 -119.515 ;
        RECT 201.115 -121.205 201.445 -120.875 ;
        RECT 201.115 -122.565 201.445 -122.235 ;
        RECT 201.115 -123.925 201.445 -123.595 ;
        RECT 201.115 -125.285 201.445 -124.955 ;
        RECT 201.115 -126.645 201.445 -126.315 ;
        RECT 201.115 -128.005 201.445 -127.675 ;
        RECT 201.115 -129.365 201.445 -129.035 ;
        RECT 201.115 -130.725 201.445 -130.395 ;
        RECT 201.115 -132.085 201.445 -131.755 ;
        RECT 201.115 -133.445 201.445 -133.115 ;
        RECT 201.115 -134.805 201.445 -134.475 ;
        RECT 201.115 -136.165 201.445 -135.835 ;
        RECT 201.115 -137.525 201.445 -137.195 ;
        RECT 201.115 -138.885 201.445 -138.555 ;
        RECT 201.115 -140.245 201.445 -139.915 ;
        RECT 201.115 -141.605 201.445 -141.275 ;
        RECT 201.115 -142.965 201.445 -142.635 ;
        RECT 201.115 -144.325 201.445 -143.995 ;
        RECT 201.115 -145.685 201.445 -145.355 ;
        RECT 201.115 -147.045 201.445 -146.715 ;
        RECT 201.115 -148.405 201.445 -148.075 ;
        RECT 201.115 -149.765 201.445 -149.435 ;
        RECT 201.115 -151.125 201.445 -150.795 ;
        RECT 201.115 -152.485 201.445 -152.155 ;
        RECT 201.115 -153.845 201.445 -153.515 ;
        RECT 201.115 -155.205 201.445 -154.875 ;
        RECT 201.115 -156.565 201.445 -156.235 ;
        RECT 201.115 -157.925 201.445 -157.595 ;
        RECT 201.115 -160.17 201.445 -159.04 ;
        RECT 201.12 -160.285 201.44 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 127.225 202.805 128.355 ;
        RECT 202.475 124.955 202.805 125.285 ;
        RECT 202.475 123.595 202.805 123.925 ;
        RECT 202.475 122.215 202.805 122.545 ;
        RECT 202.475 120.165 202.805 120.495 ;
        RECT 202.475 118.235 202.805 118.565 ;
        RECT 202.475 116.395 202.805 116.725 ;
        RECT 202.475 114.905 202.805 115.235 ;
        RECT 202.475 113.235 202.805 113.565 ;
        RECT 202.475 111.745 202.805 112.075 ;
        RECT 202.475 110.075 202.805 110.405 ;
        RECT 202.475 108.585 202.805 108.915 ;
        RECT 202.475 106.915 202.805 107.245 ;
        RECT 202.475 105.425 202.805 105.755 ;
        RECT 202.475 104.015 202.805 104.345 ;
        RECT 202.475 102.175 202.805 102.505 ;
        RECT 202.475 100.685 202.805 101.015 ;
        RECT 202.475 99.015 202.805 99.345 ;
        RECT 202.475 97.525 202.805 97.855 ;
        RECT 202.475 95.855 202.805 96.185 ;
        RECT 202.475 94.365 202.805 94.695 ;
        RECT 202.475 92.695 202.805 93.025 ;
        RECT 202.475 91.205 202.805 91.535 ;
        RECT 202.475 89.795 202.805 90.125 ;
        RECT 202.475 87.955 202.805 88.285 ;
        RECT 202.475 86.465 202.805 86.795 ;
        RECT 202.475 84.795 202.805 85.125 ;
        RECT 202.475 83.305 202.805 83.635 ;
        RECT 202.475 81.635 202.805 81.965 ;
        RECT 202.475 80.145 202.805 80.475 ;
        RECT 202.475 78.475 202.805 78.805 ;
        RECT 202.475 76.985 202.805 77.315 ;
        RECT 202.475 75.575 202.805 75.905 ;
        RECT 202.475 73.735 202.805 74.065 ;
        RECT 202.475 72.245 202.805 72.575 ;
        RECT 202.475 70.575 202.805 70.905 ;
        RECT 202.475 69.085 202.805 69.415 ;
        RECT 202.475 67.415 202.805 67.745 ;
        RECT 202.475 65.925 202.805 66.255 ;
        RECT 202.475 64.255 202.805 64.585 ;
        RECT 202.475 62.765 202.805 63.095 ;
        RECT 202.475 61.355 202.805 61.685 ;
        RECT 202.475 59.515 202.805 59.845 ;
        RECT 202.475 58.025 202.805 58.355 ;
        RECT 202.475 56.355 202.805 56.685 ;
        RECT 202.475 54.865 202.805 55.195 ;
        RECT 202.475 53.195 202.805 53.525 ;
        RECT 202.475 51.705 202.805 52.035 ;
        RECT 202.475 50.035 202.805 50.365 ;
        RECT 202.475 48.545 202.805 48.875 ;
        RECT 202.475 47.135 202.805 47.465 ;
        RECT 202.475 45.295 202.805 45.625 ;
        RECT 202.475 43.805 202.805 44.135 ;
        RECT 202.475 42.135 202.805 42.465 ;
        RECT 202.475 40.645 202.805 40.975 ;
        RECT 202.475 38.975 202.805 39.305 ;
        RECT 202.475 37.485 202.805 37.815 ;
        RECT 202.475 35.815 202.805 36.145 ;
        RECT 202.475 34.325 202.805 34.655 ;
        RECT 202.475 32.915 202.805 33.245 ;
        RECT 202.475 31.075 202.805 31.405 ;
        RECT 202.475 29.585 202.805 29.915 ;
        RECT 202.475 27.915 202.805 28.245 ;
        RECT 202.475 26.425 202.805 26.755 ;
        RECT 202.475 24.755 202.805 25.085 ;
        RECT 202.475 23.265 202.805 23.595 ;
        RECT 202.475 21.595 202.805 21.925 ;
        RECT 202.475 20.105 202.805 20.435 ;
        RECT 202.475 18.695 202.805 19.025 ;
        RECT 202.475 16.855 202.805 17.185 ;
        RECT 202.475 15.365 202.805 15.695 ;
        RECT 202.475 13.695 202.805 14.025 ;
        RECT 202.475 12.205 202.805 12.535 ;
        RECT 202.475 10.535 202.805 10.865 ;
        RECT 202.475 9.045 202.805 9.375 ;
        RECT 202.475 7.375 202.805 7.705 ;
        RECT 202.475 5.885 202.805 6.215 ;
        RECT 202.475 4.475 202.805 4.805 ;
        RECT 202.475 2.115 202.805 2.445 ;
        RECT 202.475 0.06 202.805 0.39 ;
        RECT 202.475 -1.525 202.805 -1.195 ;
        RECT 202.475 -2.885 202.805 -2.555 ;
        RECT 202.475 -4.245 202.805 -3.915 ;
        RECT 202.475 -5.605 202.805 -5.275 ;
        RECT 202.475 -6.965 202.805 -6.635 ;
        RECT 202.475 -8.325 202.805 -7.995 ;
        RECT 202.475 -9.685 202.805 -9.355 ;
        RECT 202.475 -11.045 202.805 -10.715 ;
        RECT 202.475 -12.405 202.805 -12.075 ;
        RECT 202.475 -13.765 202.805 -13.435 ;
        RECT 202.475 -15.125 202.805 -14.795 ;
        RECT 202.475 -16.485 202.805 -16.155 ;
        RECT 202.475 -17.845 202.805 -17.515 ;
        RECT 202.475 -19.205 202.805 -18.875 ;
        RECT 202.475 -20.565 202.805 -20.235 ;
        RECT 202.475 -21.925 202.805 -21.595 ;
        RECT 202.475 -23.285 202.805 -22.955 ;
        RECT 202.475 -24.645 202.805 -24.315 ;
        RECT 202.475 -26.005 202.805 -25.675 ;
        RECT 202.475 -27.365 202.805 -27.035 ;
        RECT 202.475 -28.725 202.805 -28.395 ;
        RECT 202.475 -30.085 202.805 -29.755 ;
        RECT 202.475 -31.445 202.805 -31.115 ;
        RECT 202.475 -32.805 202.805 -32.475 ;
        RECT 202.475 -34.165 202.805 -33.835 ;
        RECT 202.475 -35.525 202.805 -35.195 ;
        RECT 202.475 -36.885 202.805 -36.555 ;
        RECT 202.475 -38.245 202.805 -37.915 ;
        RECT 202.475 -39.605 202.805 -39.275 ;
        RECT 202.475 -40.965 202.805 -40.635 ;
        RECT 202.475 -42.325 202.805 -41.995 ;
        RECT 202.475 -43.685 202.805 -43.355 ;
        RECT 202.475 -45.045 202.805 -44.715 ;
        RECT 202.475 -46.405 202.805 -46.075 ;
        RECT 202.475 -47.765 202.805 -47.435 ;
        RECT 202.475 -49.125 202.805 -48.795 ;
        RECT 202.475 -50.485 202.805 -50.155 ;
        RECT 202.475 -51.845 202.805 -51.515 ;
        RECT 202.475 -53.205 202.805 -52.875 ;
        RECT 202.475 -54.565 202.805 -54.235 ;
        RECT 202.475 -55.925 202.805 -55.595 ;
        RECT 202.475 -57.285 202.805 -56.955 ;
        RECT 202.475 -58.645 202.805 -58.315 ;
        RECT 202.475 -60.005 202.805 -59.675 ;
        RECT 202.475 -61.365 202.805 -61.035 ;
        RECT 202.475 -62.725 202.805 -62.395 ;
        RECT 202.475 -64.085 202.805 -63.755 ;
        RECT 202.475 -65.445 202.805 -65.115 ;
        RECT 202.475 -66.805 202.805 -66.475 ;
        RECT 202.475 -68.165 202.805 -67.835 ;
        RECT 202.475 -69.525 202.805 -69.195 ;
        RECT 202.475 -70.885 202.805 -70.555 ;
        RECT 202.475 -72.245 202.805 -71.915 ;
        RECT 202.475 -73.605 202.805 -73.275 ;
        RECT 202.475 -74.965 202.805 -74.635 ;
        RECT 202.475 -76.325 202.805 -75.995 ;
        RECT 202.475 -77.685 202.805 -77.355 ;
        RECT 202.475 -79.045 202.805 -78.715 ;
        RECT 202.475 -80.405 202.805 -80.075 ;
        RECT 202.475 -81.765 202.805 -81.435 ;
        RECT 202.475 -83.125 202.805 -82.795 ;
        RECT 202.475 -84.485 202.805 -84.155 ;
        RECT 202.475 -85.845 202.805 -85.515 ;
        RECT 202.475 -87.205 202.805 -86.875 ;
        RECT 202.475 -88.565 202.805 -88.235 ;
        RECT 202.475 -89.925 202.805 -89.595 ;
        RECT 202.475 -91.285 202.805 -90.955 ;
        RECT 202.475 -92.645 202.805 -92.315 ;
        RECT 202.475 -94.005 202.805 -93.675 ;
        RECT 202.475 -95.365 202.805 -95.035 ;
        RECT 202.475 -96.725 202.805 -96.395 ;
        RECT 202.475 -98.085 202.805 -97.755 ;
        RECT 202.475 -99.445 202.805 -99.115 ;
        RECT 202.475 -100.805 202.805 -100.475 ;
        RECT 202.475 -102.165 202.805 -101.835 ;
        RECT 202.475 -103.525 202.805 -103.195 ;
        RECT 202.475 -104.885 202.805 -104.555 ;
        RECT 202.475 -106.245 202.805 -105.915 ;
        RECT 202.475 -107.605 202.805 -107.275 ;
        RECT 202.475 -108.965 202.805 -108.635 ;
        RECT 202.475 -110.325 202.805 -109.995 ;
        RECT 202.475 -111.685 202.805 -111.355 ;
        RECT 202.475 -113.045 202.805 -112.715 ;
        RECT 202.475 -114.405 202.805 -114.075 ;
        RECT 202.475 -115.765 202.805 -115.435 ;
        RECT 202.475 -117.125 202.805 -116.795 ;
        RECT 202.475 -118.485 202.805 -118.155 ;
        RECT 202.475 -119.845 202.805 -119.515 ;
        RECT 202.475 -121.205 202.805 -120.875 ;
        RECT 202.475 -122.565 202.805 -122.235 ;
        RECT 202.475 -123.925 202.805 -123.595 ;
        RECT 202.475 -125.285 202.805 -124.955 ;
        RECT 202.475 -126.645 202.805 -126.315 ;
        RECT 202.475 -128.005 202.805 -127.675 ;
        RECT 202.475 -129.365 202.805 -129.035 ;
        RECT 202.475 -130.725 202.805 -130.395 ;
        RECT 202.475 -132.085 202.805 -131.755 ;
        RECT 202.475 -133.445 202.805 -133.115 ;
        RECT 202.475 -134.805 202.805 -134.475 ;
        RECT 202.475 -136.165 202.805 -135.835 ;
        RECT 202.475 -137.525 202.805 -137.195 ;
        RECT 202.475 -138.885 202.805 -138.555 ;
        RECT 202.475 -140.245 202.805 -139.915 ;
        RECT 202.475 -141.605 202.805 -141.275 ;
        RECT 202.475 -142.965 202.805 -142.635 ;
        RECT 202.475 -144.325 202.805 -143.995 ;
        RECT 202.475 -145.685 202.805 -145.355 ;
        RECT 202.475 -147.045 202.805 -146.715 ;
        RECT 202.475 -148.405 202.805 -148.075 ;
        RECT 202.475 -149.765 202.805 -149.435 ;
        RECT 202.475 -151.125 202.805 -150.795 ;
        RECT 202.475 -152.485 202.805 -152.155 ;
        RECT 202.475 -153.845 202.805 -153.515 ;
        RECT 202.475 -155.205 202.805 -154.875 ;
        RECT 202.475 -156.565 202.805 -156.235 ;
        RECT 202.475 -157.925 202.805 -157.595 ;
        RECT 202.475 -160.17 202.805 -159.04 ;
        RECT 202.48 -160.285 202.8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 127.225 204.165 128.355 ;
        RECT 203.835 124.955 204.165 125.285 ;
        RECT 203.835 123.595 204.165 123.925 ;
        RECT 203.835 122.215 204.165 122.545 ;
        RECT 203.835 120.165 204.165 120.495 ;
        RECT 203.835 118.235 204.165 118.565 ;
        RECT 203.835 116.395 204.165 116.725 ;
        RECT 203.835 114.905 204.165 115.235 ;
        RECT 203.835 113.235 204.165 113.565 ;
        RECT 203.835 111.745 204.165 112.075 ;
        RECT 203.835 110.075 204.165 110.405 ;
        RECT 203.835 108.585 204.165 108.915 ;
        RECT 203.835 106.915 204.165 107.245 ;
        RECT 203.835 105.425 204.165 105.755 ;
        RECT 203.835 104.015 204.165 104.345 ;
        RECT 203.835 102.175 204.165 102.505 ;
        RECT 203.835 100.685 204.165 101.015 ;
        RECT 203.835 99.015 204.165 99.345 ;
        RECT 203.835 97.525 204.165 97.855 ;
        RECT 203.835 95.855 204.165 96.185 ;
        RECT 203.835 94.365 204.165 94.695 ;
        RECT 203.835 92.695 204.165 93.025 ;
        RECT 203.835 91.205 204.165 91.535 ;
        RECT 203.835 89.795 204.165 90.125 ;
        RECT 203.835 87.955 204.165 88.285 ;
        RECT 203.835 86.465 204.165 86.795 ;
        RECT 203.835 84.795 204.165 85.125 ;
        RECT 203.835 83.305 204.165 83.635 ;
        RECT 203.835 81.635 204.165 81.965 ;
        RECT 203.835 80.145 204.165 80.475 ;
        RECT 203.835 78.475 204.165 78.805 ;
        RECT 203.835 76.985 204.165 77.315 ;
        RECT 203.835 75.575 204.165 75.905 ;
        RECT 203.835 73.735 204.165 74.065 ;
        RECT 203.835 72.245 204.165 72.575 ;
        RECT 203.835 70.575 204.165 70.905 ;
        RECT 203.835 69.085 204.165 69.415 ;
        RECT 203.835 67.415 204.165 67.745 ;
        RECT 203.835 65.925 204.165 66.255 ;
        RECT 203.835 64.255 204.165 64.585 ;
        RECT 203.835 62.765 204.165 63.095 ;
        RECT 203.835 61.355 204.165 61.685 ;
        RECT 203.835 59.515 204.165 59.845 ;
        RECT 203.835 58.025 204.165 58.355 ;
        RECT 203.835 56.355 204.165 56.685 ;
        RECT 203.835 54.865 204.165 55.195 ;
        RECT 203.835 53.195 204.165 53.525 ;
        RECT 203.835 51.705 204.165 52.035 ;
        RECT 203.835 50.035 204.165 50.365 ;
        RECT 203.835 48.545 204.165 48.875 ;
        RECT 203.835 47.135 204.165 47.465 ;
        RECT 203.835 45.295 204.165 45.625 ;
        RECT 203.835 43.805 204.165 44.135 ;
        RECT 203.835 42.135 204.165 42.465 ;
        RECT 203.835 40.645 204.165 40.975 ;
        RECT 203.835 38.975 204.165 39.305 ;
        RECT 203.835 37.485 204.165 37.815 ;
        RECT 203.835 35.815 204.165 36.145 ;
        RECT 203.835 34.325 204.165 34.655 ;
        RECT 203.835 32.915 204.165 33.245 ;
        RECT 203.835 31.075 204.165 31.405 ;
        RECT 203.835 29.585 204.165 29.915 ;
        RECT 203.835 27.915 204.165 28.245 ;
        RECT 203.835 26.425 204.165 26.755 ;
        RECT 203.835 24.755 204.165 25.085 ;
        RECT 203.835 23.265 204.165 23.595 ;
        RECT 203.835 21.595 204.165 21.925 ;
        RECT 203.835 20.105 204.165 20.435 ;
        RECT 203.835 18.695 204.165 19.025 ;
        RECT 203.835 16.855 204.165 17.185 ;
        RECT 203.835 15.365 204.165 15.695 ;
        RECT 203.835 13.695 204.165 14.025 ;
        RECT 203.835 12.205 204.165 12.535 ;
        RECT 203.835 10.535 204.165 10.865 ;
        RECT 203.835 9.045 204.165 9.375 ;
        RECT 203.835 7.375 204.165 7.705 ;
        RECT 203.835 5.885 204.165 6.215 ;
        RECT 203.835 4.475 204.165 4.805 ;
        RECT 203.835 2.115 204.165 2.445 ;
        RECT 203.835 0.06 204.165 0.39 ;
        RECT 203.835 -1.525 204.165 -1.195 ;
        RECT 203.835 -2.885 204.165 -2.555 ;
        RECT 203.835 -4.245 204.165 -3.915 ;
        RECT 203.835 -5.605 204.165 -5.275 ;
        RECT 203.835 -6.965 204.165 -6.635 ;
        RECT 203.835 -8.325 204.165 -7.995 ;
        RECT 203.835 -9.685 204.165 -9.355 ;
        RECT 203.835 -11.045 204.165 -10.715 ;
        RECT 203.835 -12.405 204.165 -12.075 ;
        RECT 203.835 -13.765 204.165 -13.435 ;
        RECT 203.835 -15.125 204.165 -14.795 ;
        RECT 203.835 -16.485 204.165 -16.155 ;
        RECT 203.835 -17.845 204.165 -17.515 ;
        RECT 203.835 -19.205 204.165 -18.875 ;
        RECT 203.835 -20.565 204.165 -20.235 ;
        RECT 203.835 -21.925 204.165 -21.595 ;
        RECT 203.835 -23.285 204.165 -22.955 ;
        RECT 203.835 -24.645 204.165 -24.315 ;
        RECT 203.835 -26.005 204.165 -25.675 ;
        RECT 203.835 -27.365 204.165 -27.035 ;
        RECT 203.835 -28.725 204.165 -28.395 ;
        RECT 203.835 -30.085 204.165 -29.755 ;
        RECT 203.835 -31.445 204.165 -31.115 ;
        RECT 203.835 -32.805 204.165 -32.475 ;
        RECT 203.835 -34.165 204.165 -33.835 ;
        RECT 203.835 -35.525 204.165 -35.195 ;
        RECT 203.835 -36.885 204.165 -36.555 ;
        RECT 203.835 -38.245 204.165 -37.915 ;
        RECT 203.835 -39.605 204.165 -39.275 ;
        RECT 203.835 -40.965 204.165 -40.635 ;
        RECT 203.835 -42.325 204.165 -41.995 ;
        RECT 203.835 -43.685 204.165 -43.355 ;
        RECT 203.835 -45.045 204.165 -44.715 ;
        RECT 203.835 -46.405 204.165 -46.075 ;
        RECT 203.835 -47.765 204.165 -47.435 ;
        RECT 203.835 -49.125 204.165 -48.795 ;
        RECT 203.835 -50.485 204.165 -50.155 ;
        RECT 203.835 -51.845 204.165 -51.515 ;
        RECT 203.835 -53.205 204.165 -52.875 ;
        RECT 203.835 -54.565 204.165 -54.235 ;
        RECT 203.835 -55.925 204.165 -55.595 ;
        RECT 203.835 -57.285 204.165 -56.955 ;
        RECT 203.835 -58.645 204.165 -58.315 ;
        RECT 203.835 -60.005 204.165 -59.675 ;
        RECT 203.835 -61.365 204.165 -61.035 ;
        RECT 203.835 -62.725 204.165 -62.395 ;
        RECT 203.835 -64.085 204.165 -63.755 ;
        RECT 203.835 -65.445 204.165 -65.115 ;
        RECT 203.835 -66.805 204.165 -66.475 ;
        RECT 203.835 -68.165 204.165 -67.835 ;
        RECT 203.835 -69.525 204.165 -69.195 ;
        RECT 203.835 -70.885 204.165 -70.555 ;
        RECT 203.835 -72.245 204.165 -71.915 ;
        RECT 203.835 -73.605 204.165 -73.275 ;
        RECT 203.835 -74.965 204.165 -74.635 ;
        RECT 203.835 -76.325 204.165 -75.995 ;
        RECT 203.835 -77.685 204.165 -77.355 ;
        RECT 203.835 -79.045 204.165 -78.715 ;
        RECT 203.835 -80.405 204.165 -80.075 ;
        RECT 203.835 -81.765 204.165 -81.435 ;
        RECT 203.835 -83.125 204.165 -82.795 ;
        RECT 203.835 -84.485 204.165 -84.155 ;
        RECT 203.835 -85.845 204.165 -85.515 ;
        RECT 203.835 -87.205 204.165 -86.875 ;
        RECT 203.835 -88.565 204.165 -88.235 ;
        RECT 203.835 -89.925 204.165 -89.595 ;
        RECT 203.835 -91.285 204.165 -90.955 ;
        RECT 203.835 -92.645 204.165 -92.315 ;
        RECT 203.835 -94.005 204.165 -93.675 ;
        RECT 203.835 -95.365 204.165 -95.035 ;
        RECT 203.835 -96.725 204.165 -96.395 ;
        RECT 203.835 -98.085 204.165 -97.755 ;
        RECT 203.835 -99.445 204.165 -99.115 ;
        RECT 203.835 -100.805 204.165 -100.475 ;
        RECT 203.835 -102.165 204.165 -101.835 ;
        RECT 203.835 -103.525 204.165 -103.195 ;
        RECT 203.835 -104.885 204.165 -104.555 ;
        RECT 203.835 -106.245 204.165 -105.915 ;
        RECT 203.835 -107.605 204.165 -107.275 ;
        RECT 203.835 -108.965 204.165 -108.635 ;
        RECT 203.835 -110.325 204.165 -109.995 ;
        RECT 203.835 -111.685 204.165 -111.355 ;
        RECT 203.835 -113.045 204.165 -112.715 ;
        RECT 203.835 -114.405 204.165 -114.075 ;
        RECT 203.835 -115.765 204.165 -115.435 ;
        RECT 203.835 -117.125 204.165 -116.795 ;
        RECT 203.835 -118.485 204.165 -118.155 ;
        RECT 203.835 -119.845 204.165 -119.515 ;
        RECT 203.835 -121.205 204.165 -120.875 ;
        RECT 203.835 -122.565 204.165 -122.235 ;
        RECT 203.835 -123.925 204.165 -123.595 ;
        RECT 203.835 -125.285 204.165 -124.955 ;
        RECT 203.835 -126.645 204.165 -126.315 ;
        RECT 203.835 -128.005 204.165 -127.675 ;
        RECT 203.835 -129.365 204.165 -129.035 ;
        RECT 203.835 -130.725 204.165 -130.395 ;
        RECT 203.835 -132.085 204.165 -131.755 ;
        RECT 203.835 -133.445 204.165 -133.115 ;
        RECT 203.835 -134.805 204.165 -134.475 ;
        RECT 203.835 -136.165 204.165 -135.835 ;
        RECT 203.835 -137.525 204.165 -137.195 ;
        RECT 203.835 -138.885 204.165 -138.555 ;
        RECT 203.835 -140.245 204.165 -139.915 ;
        RECT 203.835 -141.605 204.165 -141.275 ;
        RECT 203.835 -142.965 204.165 -142.635 ;
        RECT 203.835 -144.325 204.165 -143.995 ;
        RECT 203.835 -145.685 204.165 -145.355 ;
        RECT 203.835 -147.045 204.165 -146.715 ;
        RECT 203.835 -148.405 204.165 -148.075 ;
        RECT 203.835 -149.765 204.165 -149.435 ;
        RECT 203.835 -151.125 204.165 -150.795 ;
        RECT 203.835 -152.485 204.165 -152.155 ;
        RECT 203.835 -153.845 204.165 -153.515 ;
        RECT 203.835 -155.205 204.165 -154.875 ;
        RECT 203.835 -156.565 204.165 -156.235 ;
        RECT 203.835 -157.925 204.165 -157.595 ;
        RECT 203.835 -160.17 204.165 -159.04 ;
        RECT 203.84 -160.285 204.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 127.225 205.525 128.355 ;
        RECT 205.195 124.955 205.525 125.285 ;
        RECT 205.195 123.595 205.525 123.925 ;
        RECT 205.195 122.215 205.525 122.545 ;
        RECT 205.195 120.165 205.525 120.495 ;
        RECT 205.195 118.235 205.525 118.565 ;
        RECT 205.195 116.395 205.525 116.725 ;
        RECT 205.195 114.905 205.525 115.235 ;
        RECT 205.195 113.235 205.525 113.565 ;
        RECT 205.195 111.745 205.525 112.075 ;
        RECT 205.195 110.075 205.525 110.405 ;
        RECT 205.195 108.585 205.525 108.915 ;
        RECT 205.195 106.915 205.525 107.245 ;
        RECT 205.195 105.425 205.525 105.755 ;
        RECT 205.195 104.015 205.525 104.345 ;
        RECT 205.195 102.175 205.525 102.505 ;
        RECT 205.195 100.685 205.525 101.015 ;
        RECT 205.195 99.015 205.525 99.345 ;
        RECT 205.195 97.525 205.525 97.855 ;
        RECT 205.195 95.855 205.525 96.185 ;
        RECT 205.195 94.365 205.525 94.695 ;
        RECT 205.195 92.695 205.525 93.025 ;
        RECT 205.195 91.205 205.525 91.535 ;
        RECT 205.195 89.795 205.525 90.125 ;
        RECT 205.195 87.955 205.525 88.285 ;
        RECT 205.195 86.465 205.525 86.795 ;
        RECT 205.195 84.795 205.525 85.125 ;
        RECT 205.195 83.305 205.525 83.635 ;
        RECT 205.195 81.635 205.525 81.965 ;
        RECT 205.195 80.145 205.525 80.475 ;
        RECT 205.195 78.475 205.525 78.805 ;
        RECT 205.195 76.985 205.525 77.315 ;
        RECT 205.195 75.575 205.525 75.905 ;
        RECT 205.195 73.735 205.525 74.065 ;
        RECT 205.195 72.245 205.525 72.575 ;
        RECT 205.195 70.575 205.525 70.905 ;
        RECT 205.195 69.085 205.525 69.415 ;
        RECT 205.195 67.415 205.525 67.745 ;
        RECT 205.195 65.925 205.525 66.255 ;
        RECT 205.195 64.255 205.525 64.585 ;
        RECT 205.195 62.765 205.525 63.095 ;
        RECT 205.195 61.355 205.525 61.685 ;
        RECT 205.195 59.515 205.525 59.845 ;
        RECT 205.195 58.025 205.525 58.355 ;
        RECT 205.195 56.355 205.525 56.685 ;
        RECT 205.195 54.865 205.525 55.195 ;
        RECT 205.195 53.195 205.525 53.525 ;
        RECT 205.195 51.705 205.525 52.035 ;
        RECT 205.195 50.035 205.525 50.365 ;
        RECT 205.195 48.545 205.525 48.875 ;
        RECT 205.195 47.135 205.525 47.465 ;
        RECT 205.195 45.295 205.525 45.625 ;
        RECT 205.195 43.805 205.525 44.135 ;
        RECT 205.195 42.135 205.525 42.465 ;
        RECT 205.195 40.645 205.525 40.975 ;
        RECT 205.195 38.975 205.525 39.305 ;
        RECT 205.195 37.485 205.525 37.815 ;
        RECT 205.195 35.815 205.525 36.145 ;
        RECT 205.195 34.325 205.525 34.655 ;
        RECT 205.195 32.915 205.525 33.245 ;
        RECT 205.195 31.075 205.525 31.405 ;
        RECT 205.195 29.585 205.525 29.915 ;
        RECT 205.195 27.915 205.525 28.245 ;
        RECT 205.195 26.425 205.525 26.755 ;
        RECT 205.195 24.755 205.525 25.085 ;
        RECT 205.195 23.265 205.525 23.595 ;
        RECT 205.195 21.595 205.525 21.925 ;
        RECT 205.195 20.105 205.525 20.435 ;
        RECT 205.195 18.695 205.525 19.025 ;
        RECT 205.195 16.855 205.525 17.185 ;
        RECT 205.195 15.365 205.525 15.695 ;
        RECT 205.195 13.695 205.525 14.025 ;
        RECT 205.195 12.205 205.525 12.535 ;
        RECT 205.195 10.535 205.525 10.865 ;
        RECT 205.195 9.045 205.525 9.375 ;
        RECT 205.195 7.375 205.525 7.705 ;
        RECT 205.195 5.885 205.525 6.215 ;
        RECT 205.195 4.475 205.525 4.805 ;
        RECT 205.195 2.115 205.525 2.445 ;
        RECT 205.195 0.06 205.525 0.39 ;
        RECT 205.195 -1.525 205.525 -1.195 ;
        RECT 205.195 -2.885 205.525 -2.555 ;
        RECT 205.195 -4.245 205.525 -3.915 ;
        RECT 205.195 -5.605 205.525 -5.275 ;
        RECT 205.195 -6.965 205.525 -6.635 ;
        RECT 205.195 -8.325 205.525 -7.995 ;
        RECT 205.195 -9.685 205.525 -9.355 ;
        RECT 205.195 -11.045 205.525 -10.715 ;
        RECT 205.195 -12.405 205.525 -12.075 ;
        RECT 205.195 -13.765 205.525 -13.435 ;
        RECT 205.195 -15.125 205.525 -14.795 ;
        RECT 205.195 -16.485 205.525 -16.155 ;
        RECT 205.195 -17.845 205.525 -17.515 ;
        RECT 205.195 -19.205 205.525 -18.875 ;
        RECT 205.195 -20.565 205.525 -20.235 ;
        RECT 205.195 -21.925 205.525 -21.595 ;
        RECT 205.195 -23.285 205.525 -22.955 ;
        RECT 205.195 -24.645 205.525 -24.315 ;
        RECT 205.195 -26.005 205.525 -25.675 ;
        RECT 205.195 -27.365 205.525 -27.035 ;
        RECT 205.195 -28.725 205.525 -28.395 ;
        RECT 205.195 -30.085 205.525 -29.755 ;
        RECT 205.195 -31.445 205.525 -31.115 ;
        RECT 205.195 -32.805 205.525 -32.475 ;
        RECT 205.195 -34.165 205.525 -33.835 ;
        RECT 205.195 -35.525 205.525 -35.195 ;
        RECT 205.195 -36.885 205.525 -36.555 ;
        RECT 205.195 -38.245 205.525 -37.915 ;
        RECT 205.195 -39.605 205.525 -39.275 ;
        RECT 205.195 -40.965 205.525 -40.635 ;
        RECT 205.195 -42.325 205.525 -41.995 ;
        RECT 205.195 -43.685 205.525 -43.355 ;
        RECT 205.195 -45.045 205.525 -44.715 ;
        RECT 205.195 -46.405 205.525 -46.075 ;
        RECT 205.195 -47.765 205.525 -47.435 ;
        RECT 205.195 -49.125 205.525 -48.795 ;
        RECT 205.195 -50.485 205.525 -50.155 ;
        RECT 205.195 -51.845 205.525 -51.515 ;
        RECT 205.195 -53.205 205.525 -52.875 ;
        RECT 205.195 -54.565 205.525 -54.235 ;
        RECT 205.195 -55.925 205.525 -55.595 ;
        RECT 205.195 -57.285 205.525 -56.955 ;
        RECT 205.195 -58.645 205.525 -58.315 ;
        RECT 205.195 -60.005 205.525 -59.675 ;
        RECT 205.195 -61.365 205.525 -61.035 ;
        RECT 205.195 -62.725 205.525 -62.395 ;
        RECT 205.195 -64.085 205.525 -63.755 ;
        RECT 205.195 -65.445 205.525 -65.115 ;
        RECT 205.195 -66.805 205.525 -66.475 ;
        RECT 205.195 -68.165 205.525 -67.835 ;
        RECT 205.195 -69.525 205.525 -69.195 ;
        RECT 205.195 -70.885 205.525 -70.555 ;
        RECT 205.195 -72.245 205.525 -71.915 ;
        RECT 205.195 -73.605 205.525 -73.275 ;
        RECT 205.195 -74.965 205.525 -74.635 ;
        RECT 205.195 -76.325 205.525 -75.995 ;
        RECT 205.195 -77.685 205.525 -77.355 ;
        RECT 205.195 -79.045 205.525 -78.715 ;
        RECT 205.195 -80.405 205.525 -80.075 ;
        RECT 205.195 -81.765 205.525 -81.435 ;
        RECT 205.195 -83.125 205.525 -82.795 ;
        RECT 205.195 -84.485 205.525 -84.155 ;
        RECT 205.195 -85.845 205.525 -85.515 ;
        RECT 205.195 -87.205 205.525 -86.875 ;
        RECT 205.195 -88.565 205.525 -88.235 ;
        RECT 205.195 -89.925 205.525 -89.595 ;
        RECT 205.195 -91.285 205.525 -90.955 ;
        RECT 205.195 -92.645 205.525 -92.315 ;
        RECT 205.195 -94.005 205.525 -93.675 ;
        RECT 205.195 -95.365 205.525 -95.035 ;
        RECT 205.195 -96.725 205.525 -96.395 ;
        RECT 205.195 -98.085 205.525 -97.755 ;
        RECT 205.195 -99.445 205.525 -99.115 ;
        RECT 205.195 -100.805 205.525 -100.475 ;
        RECT 205.195 -102.165 205.525 -101.835 ;
        RECT 205.195 -103.525 205.525 -103.195 ;
        RECT 205.195 -104.885 205.525 -104.555 ;
        RECT 205.195 -106.245 205.525 -105.915 ;
        RECT 205.195 -107.605 205.525 -107.275 ;
        RECT 205.195 -108.965 205.525 -108.635 ;
        RECT 205.195 -110.325 205.525 -109.995 ;
        RECT 205.195 -111.685 205.525 -111.355 ;
        RECT 205.195 -113.045 205.525 -112.715 ;
        RECT 205.195 -114.405 205.525 -114.075 ;
        RECT 205.195 -115.765 205.525 -115.435 ;
        RECT 205.195 -117.125 205.525 -116.795 ;
        RECT 205.195 -118.485 205.525 -118.155 ;
        RECT 205.195 -119.845 205.525 -119.515 ;
        RECT 205.195 -121.205 205.525 -120.875 ;
        RECT 205.195 -122.565 205.525 -122.235 ;
        RECT 205.195 -123.925 205.525 -123.595 ;
        RECT 205.195 -125.285 205.525 -124.955 ;
        RECT 205.195 -126.645 205.525 -126.315 ;
        RECT 205.195 -128.005 205.525 -127.675 ;
        RECT 205.195 -129.365 205.525 -129.035 ;
        RECT 205.195 -130.725 205.525 -130.395 ;
        RECT 205.195 -132.085 205.525 -131.755 ;
        RECT 205.195 -133.445 205.525 -133.115 ;
        RECT 205.195 -134.805 205.525 -134.475 ;
        RECT 205.195 -136.165 205.525 -135.835 ;
        RECT 205.195 -137.525 205.525 -137.195 ;
        RECT 205.195 -138.885 205.525 -138.555 ;
        RECT 205.195 -140.245 205.525 -139.915 ;
        RECT 205.195 -141.605 205.525 -141.275 ;
        RECT 205.195 -142.965 205.525 -142.635 ;
        RECT 205.195 -144.325 205.525 -143.995 ;
        RECT 205.195 -145.685 205.525 -145.355 ;
        RECT 205.195 -147.045 205.525 -146.715 ;
        RECT 205.195 -148.405 205.525 -148.075 ;
        RECT 205.195 -149.765 205.525 -149.435 ;
        RECT 205.195 -151.125 205.525 -150.795 ;
        RECT 205.195 -152.485 205.525 -152.155 ;
        RECT 205.195 -153.845 205.525 -153.515 ;
        RECT 205.195 -155.205 205.525 -154.875 ;
        RECT 205.195 -156.565 205.525 -156.235 ;
        RECT 205.195 -157.925 205.525 -157.595 ;
        RECT 205.195 -160.17 205.525 -159.04 ;
        RECT 205.2 -160.285 205.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 127.225 206.885 128.355 ;
        RECT 206.555 124.955 206.885 125.285 ;
        RECT 206.555 123.595 206.885 123.925 ;
        RECT 206.555 122.215 206.885 122.545 ;
        RECT 206.555 120.165 206.885 120.495 ;
        RECT 206.555 118.235 206.885 118.565 ;
        RECT 206.555 116.395 206.885 116.725 ;
        RECT 206.555 114.905 206.885 115.235 ;
        RECT 206.555 113.235 206.885 113.565 ;
        RECT 206.555 111.745 206.885 112.075 ;
        RECT 206.555 110.075 206.885 110.405 ;
        RECT 206.555 108.585 206.885 108.915 ;
        RECT 206.555 106.915 206.885 107.245 ;
        RECT 206.555 105.425 206.885 105.755 ;
        RECT 206.555 104.015 206.885 104.345 ;
        RECT 206.555 102.175 206.885 102.505 ;
        RECT 206.555 100.685 206.885 101.015 ;
        RECT 206.555 99.015 206.885 99.345 ;
        RECT 206.555 97.525 206.885 97.855 ;
        RECT 206.555 95.855 206.885 96.185 ;
        RECT 206.555 94.365 206.885 94.695 ;
        RECT 206.555 92.695 206.885 93.025 ;
        RECT 206.555 91.205 206.885 91.535 ;
        RECT 206.555 89.795 206.885 90.125 ;
        RECT 206.555 87.955 206.885 88.285 ;
        RECT 206.555 86.465 206.885 86.795 ;
        RECT 206.555 84.795 206.885 85.125 ;
        RECT 206.555 83.305 206.885 83.635 ;
        RECT 206.555 81.635 206.885 81.965 ;
        RECT 206.555 80.145 206.885 80.475 ;
        RECT 206.555 78.475 206.885 78.805 ;
        RECT 206.555 76.985 206.885 77.315 ;
        RECT 206.555 75.575 206.885 75.905 ;
        RECT 206.555 73.735 206.885 74.065 ;
        RECT 206.555 72.245 206.885 72.575 ;
        RECT 206.555 70.575 206.885 70.905 ;
        RECT 206.555 69.085 206.885 69.415 ;
        RECT 206.555 67.415 206.885 67.745 ;
        RECT 206.555 65.925 206.885 66.255 ;
        RECT 206.555 64.255 206.885 64.585 ;
        RECT 206.555 62.765 206.885 63.095 ;
        RECT 206.555 61.355 206.885 61.685 ;
        RECT 206.555 59.515 206.885 59.845 ;
        RECT 206.555 58.025 206.885 58.355 ;
        RECT 206.555 56.355 206.885 56.685 ;
        RECT 206.555 54.865 206.885 55.195 ;
        RECT 206.555 53.195 206.885 53.525 ;
        RECT 206.555 51.705 206.885 52.035 ;
        RECT 206.555 50.035 206.885 50.365 ;
        RECT 206.555 48.545 206.885 48.875 ;
        RECT 206.555 47.135 206.885 47.465 ;
        RECT 206.555 45.295 206.885 45.625 ;
        RECT 206.555 43.805 206.885 44.135 ;
        RECT 206.555 42.135 206.885 42.465 ;
        RECT 206.555 40.645 206.885 40.975 ;
        RECT 206.555 38.975 206.885 39.305 ;
        RECT 206.555 37.485 206.885 37.815 ;
        RECT 206.555 35.815 206.885 36.145 ;
        RECT 206.555 34.325 206.885 34.655 ;
        RECT 206.555 32.915 206.885 33.245 ;
        RECT 206.555 31.075 206.885 31.405 ;
        RECT 206.555 29.585 206.885 29.915 ;
        RECT 206.555 27.915 206.885 28.245 ;
        RECT 206.555 26.425 206.885 26.755 ;
        RECT 206.555 24.755 206.885 25.085 ;
        RECT 206.555 23.265 206.885 23.595 ;
        RECT 206.555 21.595 206.885 21.925 ;
        RECT 206.555 20.105 206.885 20.435 ;
        RECT 206.555 18.695 206.885 19.025 ;
        RECT 206.555 16.855 206.885 17.185 ;
        RECT 206.555 15.365 206.885 15.695 ;
        RECT 206.555 13.695 206.885 14.025 ;
        RECT 206.555 12.205 206.885 12.535 ;
        RECT 206.555 10.535 206.885 10.865 ;
        RECT 206.555 9.045 206.885 9.375 ;
        RECT 206.555 7.375 206.885 7.705 ;
        RECT 206.555 5.885 206.885 6.215 ;
        RECT 206.555 4.475 206.885 4.805 ;
        RECT 206.555 2.115 206.885 2.445 ;
        RECT 206.555 0.06 206.885 0.39 ;
        RECT 206.555 -1.525 206.885 -1.195 ;
        RECT 206.555 -2.885 206.885 -2.555 ;
        RECT 206.555 -4.245 206.885 -3.915 ;
        RECT 206.555 -5.605 206.885 -5.275 ;
        RECT 206.555 -6.965 206.885 -6.635 ;
        RECT 206.555 -8.325 206.885 -7.995 ;
        RECT 206.555 -9.685 206.885 -9.355 ;
        RECT 206.555 -11.045 206.885 -10.715 ;
        RECT 206.555 -12.405 206.885 -12.075 ;
        RECT 206.555 -13.765 206.885 -13.435 ;
        RECT 206.555 -15.125 206.885 -14.795 ;
        RECT 206.555 -16.485 206.885 -16.155 ;
        RECT 206.555 -17.845 206.885 -17.515 ;
        RECT 206.555 -19.205 206.885 -18.875 ;
        RECT 206.555 -20.565 206.885 -20.235 ;
        RECT 206.555 -21.925 206.885 -21.595 ;
        RECT 206.555 -23.285 206.885 -22.955 ;
        RECT 206.555 -24.645 206.885 -24.315 ;
        RECT 206.555 -26.005 206.885 -25.675 ;
        RECT 206.555 -27.365 206.885 -27.035 ;
        RECT 206.555 -28.725 206.885 -28.395 ;
        RECT 206.555 -30.085 206.885 -29.755 ;
        RECT 206.555 -31.445 206.885 -31.115 ;
        RECT 206.555 -32.805 206.885 -32.475 ;
        RECT 206.555 -34.165 206.885 -33.835 ;
        RECT 206.555 -35.525 206.885 -35.195 ;
        RECT 206.555 -36.885 206.885 -36.555 ;
        RECT 206.555 -38.245 206.885 -37.915 ;
        RECT 206.555 -39.605 206.885 -39.275 ;
        RECT 206.555 -40.965 206.885 -40.635 ;
        RECT 206.555 -42.325 206.885 -41.995 ;
        RECT 206.555 -43.685 206.885 -43.355 ;
        RECT 206.555 -45.045 206.885 -44.715 ;
        RECT 206.555 -46.405 206.885 -46.075 ;
        RECT 206.555 -47.765 206.885 -47.435 ;
        RECT 206.555 -49.125 206.885 -48.795 ;
        RECT 206.555 -50.485 206.885 -50.155 ;
        RECT 206.555 -51.845 206.885 -51.515 ;
        RECT 206.555 -53.205 206.885 -52.875 ;
        RECT 206.555 -54.565 206.885 -54.235 ;
        RECT 206.555 -55.925 206.885 -55.595 ;
        RECT 206.555 -57.285 206.885 -56.955 ;
        RECT 206.555 -58.645 206.885 -58.315 ;
        RECT 206.555 -60.005 206.885 -59.675 ;
        RECT 206.555 -61.365 206.885 -61.035 ;
        RECT 206.555 -62.725 206.885 -62.395 ;
        RECT 206.555 -64.085 206.885 -63.755 ;
        RECT 206.555 -65.445 206.885 -65.115 ;
        RECT 206.555 -66.805 206.885 -66.475 ;
        RECT 206.555 -68.165 206.885 -67.835 ;
        RECT 206.555 -69.525 206.885 -69.195 ;
        RECT 206.555 -70.885 206.885 -70.555 ;
        RECT 206.555 -72.245 206.885 -71.915 ;
        RECT 206.555 -73.605 206.885 -73.275 ;
        RECT 206.555 -74.965 206.885 -74.635 ;
        RECT 206.555 -76.325 206.885 -75.995 ;
        RECT 206.555 -77.685 206.885 -77.355 ;
        RECT 206.555 -79.045 206.885 -78.715 ;
        RECT 206.555 -80.405 206.885 -80.075 ;
        RECT 206.555 -81.765 206.885 -81.435 ;
        RECT 206.555 -83.125 206.885 -82.795 ;
        RECT 206.555 -84.485 206.885 -84.155 ;
        RECT 206.555 -85.845 206.885 -85.515 ;
        RECT 206.555 -87.205 206.885 -86.875 ;
        RECT 206.555 -88.565 206.885 -88.235 ;
        RECT 206.555 -89.925 206.885 -89.595 ;
        RECT 206.555 -91.285 206.885 -90.955 ;
        RECT 206.555 -92.645 206.885 -92.315 ;
        RECT 206.555 -94.005 206.885 -93.675 ;
        RECT 206.555 -95.365 206.885 -95.035 ;
        RECT 206.555 -96.725 206.885 -96.395 ;
        RECT 206.555 -98.085 206.885 -97.755 ;
        RECT 206.555 -99.445 206.885 -99.115 ;
        RECT 206.555 -100.805 206.885 -100.475 ;
        RECT 206.555 -102.165 206.885 -101.835 ;
        RECT 206.555 -103.525 206.885 -103.195 ;
        RECT 206.555 -104.885 206.885 -104.555 ;
        RECT 206.555 -106.245 206.885 -105.915 ;
        RECT 206.555 -107.605 206.885 -107.275 ;
        RECT 206.555 -108.965 206.885 -108.635 ;
        RECT 206.555 -110.325 206.885 -109.995 ;
        RECT 206.555 -111.685 206.885 -111.355 ;
        RECT 206.555 -113.045 206.885 -112.715 ;
        RECT 206.555 -114.405 206.885 -114.075 ;
        RECT 206.555 -115.765 206.885 -115.435 ;
        RECT 206.555 -117.125 206.885 -116.795 ;
        RECT 206.555 -118.485 206.885 -118.155 ;
        RECT 206.555 -119.845 206.885 -119.515 ;
        RECT 206.555 -121.205 206.885 -120.875 ;
        RECT 206.555 -122.565 206.885 -122.235 ;
        RECT 206.555 -123.925 206.885 -123.595 ;
        RECT 206.555 -125.285 206.885 -124.955 ;
        RECT 206.555 -126.645 206.885 -126.315 ;
        RECT 206.555 -128.005 206.885 -127.675 ;
        RECT 206.555 -129.365 206.885 -129.035 ;
        RECT 206.555 -130.725 206.885 -130.395 ;
        RECT 206.555 -132.085 206.885 -131.755 ;
        RECT 206.555 -133.445 206.885 -133.115 ;
        RECT 206.555 -134.805 206.885 -134.475 ;
        RECT 206.555 -136.165 206.885 -135.835 ;
        RECT 206.555 -137.525 206.885 -137.195 ;
        RECT 206.555 -138.885 206.885 -138.555 ;
        RECT 206.555 -140.245 206.885 -139.915 ;
        RECT 206.555 -141.605 206.885 -141.275 ;
        RECT 206.555 -142.965 206.885 -142.635 ;
        RECT 206.555 -144.325 206.885 -143.995 ;
        RECT 206.555 -145.685 206.885 -145.355 ;
        RECT 206.555 -147.045 206.885 -146.715 ;
        RECT 206.555 -148.405 206.885 -148.075 ;
        RECT 206.555 -149.765 206.885 -149.435 ;
        RECT 206.555 -151.125 206.885 -150.795 ;
        RECT 206.555 -152.485 206.885 -152.155 ;
        RECT 206.555 -153.845 206.885 -153.515 ;
        RECT 206.555 -155.205 206.885 -154.875 ;
        RECT 206.555 -156.565 206.885 -156.235 ;
        RECT 206.555 -157.925 206.885 -157.595 ;
        RECT 206.555 -160.17 206.885 -159.04 ;
        RECT 206.56 -160.285 206.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 127.225 160.645 128.355 ;
        RECT 160.315 124.955 160.645 125.285 ;
        RECT 160.315 123.595 160.645 123.925 ;
        RECT 160.32 123.595 160.64 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -1.525 160.645 -1.195 ;
        RECT 160.315 -2.885 160.645 -2.555 ;
        RECT 160.32 -3.56 160.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -91.285 160.645 -90.955 ;
        RECT 160.315 -92.645 160.645 -92.315 ;
        RECT 160.315 -94.005 160.645 -93.675 ;
        RECT 160.315 -95.365 160.645 -95.035 ;
        RECT 160.315 -96.725 160.645 -96.395 ;
        RECT 160.315 -98.085 160.645 -97.755 ;
        RECT 160.315 -99.445 160.645 -99.115 ;
        RECT 160.315 -100.805 160.645 -100.475 ;
        RECT 160.315 -102.165 160.645 -101.835 ;
        RECT 160.315 -103.525 160.645 -103.195 ;
        RECT 160.315 -104.885 160.645 -104.555 ;
        RECT 160.315 -106.245 160.645 -105.915 ;
        RECT 160.315 -107.605 160.645 -107.275 ;
        RECT 160.315 -108.965 160.645 -108.635 ;
        RECT 160.315 -110.325 160.645 -109.995 ;
        RECT 160.315 -111.685 160.645 -111.355 ;
        RECT 160.315 -113.045 160.645 -112.715 ;
        RECT 160.315 -114.405 160.645 -114.075 ;
        RECT 160.315 -115.765 160.645 -115.435 ;
        RECT 160.315 -117.125 160.645 -116.795 ;
        RECT 160.315 -118.485 160.645 -118.155 ;
        RECT 160.315 -119.845 160.645 -119.515 ;
        RECT 160.315 -121.205 160.645 -120.875 ;
        RECT 160.315 -122.565 160.645 -122.235 ;
        RECT 160.315 -123.925 160.645 -123.595 ;
        RECT 160.315 -125.285 160.645 -124.955 ;
        RECT 160.315 -126.645 160.645 -126.315 ;
        RECT 160.315 -128.005 160.645 -127.675 ;
        RECT 160.315 -129.365 160.645 -129.035 ;
        RECT 160.315 -130.725 160.645 -130.395 ;
        RECT 160.315 -132.085 160.645 -131.755 ;
        RECT 160.315 -133.445 160.645 -133.115 ;
        RECT 160.315 -134.805 160.645 -134.475 ;
        RECT 160.315 -136.165 160.645 -135.835 ;
        RECT 160.315 -137.525 160.645 -137.195 ;
        RECT 160.315 -138.885 160.645 -138.555 ;
        RECT 160.315 -140.245 160.645 -139.915 ;
        RECT 160.315 -141.605 160.645 -141.275 ;
        RECT 160.315 -142.965 160.645 -142.635 ;
        RECT 160.315 -144.325 160.645 -143.995 ;
        RECT 160.315 -145.685 160.645 -145.355 ;
        RECT 160.315 -147.045 160.645 -146.715 ;
        RECT 160.315 -148.405 160.645 -148.075 ;
        RECT 160.315 -149.765 160.645 -149.435 ;
        RECT 160.315 -151.125 160.645 -150.795 ;
        RECT 160.315 -152.485 160.645 -152.155 ;
        RECT 160.315 -153.845 160.645 -153.515 ;
        RECT 160.315 -155.205 160.645 -154.875 ;
        RECT 160.315 -156.565 160.645 -156.235 ;
        RECT 160.315 -157.925 160.645 -157.595 ;
        RECT 160.315 -160.17 160.645 -159.04 ;
        RECT 160.32 -160.285 160.64 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 127.225 162.005 128.355 ;
        RECT 161.675 124.955 162.005 125.285 ;
        RECT 161.675 123.595 162.005 123.925 ;
        RECT 161.68 123.595 162 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 -95.365 162.005 -95.035 ;
        RECT 161.675 -96.725 162.005 -96.395 ;
        RECT 161.675 -98.085 162.005 -97.755 ;
        RECT 161.675 -99.445 162.005 -99.115 ;
        RECT 161.675 -100.805 162.005 -100.475 ;
        RECT 161.675 -102.165 162.005 -101.835 ;
        RECT 161.675 -103.525 162.005 -103.195 ;
        RECT 161.675 -104.885 162.005 -104.555 ;
        RECT 161.675 -106.245 162.005 -105.915 ;
        RECT 161.675 -107.605 162.005 -107.275 ;
        RECT 161.675 -108.965 162.005 -108.635 ;
        RECT 161.675 -110.325 162.005 -109.995 ;
        RECT 161.675 -111.685 162.005 -111.355 ;
        RECT 161.675 -113.045 162.005 -112.715 ;
        RECT 161.675 -114.405 162.005 -114.075 ;
        RECT 161.675 -115.765 162.005 -115.435 ;
        RECT 161.675 -117.125 162.005 -116.795 ;
        RECT 161.675 -118.485 162.005 -118.155 ;
        RECT 161.675 -119.845 162.005 -119.515 ;
        RECT 161.675 -121.205 162.005 -120.875 ;
        RECT 161.675 -122.565 162.005 -122.235 ;
        RECT 161.675 -123.925 162.005 -123.595 ;
        RECT 161.675 -125.285 162.005 -124.955 ;
        RECT 161.675 -126.645 162.005 -126.315 ;
        RECT 161.675 -128.005 162.005 -127.675 ;
        RECT 161.675 -129.365 162.005 -129.035 ;
        RECT 161.675 -130.725 162.005 -130.395 ;
        RECT 161.675 -132.085 162.005 -131.755 ;
        RECT 161.675 -133.445 162.005 -133.115 ;
        RECT 161.675 -134.805 162.005 -134.475 ;
        RECT 161.675 -136.165 162.005 -135.835 ;
        RECT 161.675 -137.525 162.005 -137.195 ;
        RECT 161.675 -138.885 162.005 -138.555 ;
        RECT 161.675 -140.245 162.005 -139.915 ;
        RECT 161.675 -141.605 162.005 -141.275 ;
        RECT 161.675 -142.965 162.005 -142.635 ;
        RECT 161.675 -144.325 162.005 -143.995 ;
        RECT 161.675 -145.685 162.005 -145.355 ;
        RECT 161.675 -147.045 162.005 -146.715 ;
        RECT 161.675 -148.405 162.005 -148.075 ;
        RECT 161.675 -149.765 162.005 -149.435 ;
        RECT 161.675 -151.125 162.005 -150.795 ;
        RECT 161.675 -152.485 162.005 -152.155 ;
        RECT 161.675 -153.845 162.005 -153.515 ;
        RECT 161.675 -155.205 162.005 -154.875 ;
        RECT 161.675 -156.565 162.005 -156.235 ;
        RECT 161.675 -157.925 162.005 -157.595 ;
        RECT 161.675 -160.17 162.005 -159.04 ;
        RECT 161.68 -160.285 162 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.91 -94.075 162.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 127.225 163.365 128.355 ;
        RECT 163.035 124.955 163.365 125.285 ;
        RECT 163.035 123.595 163.365 123.925 ;
        RECT 163.04 123.595 163.36 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 -1.525 163.365 -1.195 ;
        RECT 163.035 -2.885 163.365 -2.555 ;
        RECT 163.04 -3.56 163.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 127.225 164.725 128.355 ;
        RECT 164.395 124.955 164.725 125.285 ;
        RECT 164.395 123.595 164.725 123.925 ;
        RECT 164.4 123.595 164.72 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 -1.525 164.725 -1.195 ;
        RECT 164.395 -2.885 164.725 -2.555 ;
        RECT 164.4 -3.56 164.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 127.225 166.085 128.355 ;
        RECT 165.755 124.955 166.085 125.285 ;
        RECT 165.755 123.595 166.085 123.925 ;
        RECT 165.76 123.595 166.08 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 -1.525 166.085 -1.195 ;
        RECT 165.755 -2.885 166.085 -2.555 ;
        RECT 165.76 -3.56 166.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 -91.285 166.085 -90.955 ;
        RECT 165.755 -92.645 166.085 -92.315 ;
        RECT 165.755 -94.005 166.085 -93.675 ;
        RECT 165.755 -95.365 166.085 -95.035 ;
        RECT 165.755 -96.725 166.085 -96.395 ;
        RECT 165.755 -98.085 166.085 -97.755 ;
        RECT 165.755 -99.445 166.085 -99.115 ;
        RECT 165.755 -100.805 166.085 -100.475 ;
        RECT 165.755 -102.165 166.085 -101.835 ;
        RECT 165.755 -103.525 166.085 -103.195 ;
        RECT 165.755 -104.885 166.085 -104.555 ;
        RECT 165.755 -106.245 166.085 -105.915 ;
        RECT 165.755 -107.605 166.085 -107.275 ;
        RECT 165.755 -108.965 166.085 -108.635 ;
        RECT 165.755 -110.325 166.085 -109.995 ;
        RECT 165.755 -111.685 166.085 -111.355 ;
        RECT 165.755 -113.045 166.085 -112.715 ;
        RECT 165.755 -114.405 166.085 -114.075 ;
        RECT 165.755 -115.765 166.085 -115.435 ;
        RECT 165.755 -117.125 166.085 -116.795 ;
        RECT 165.755 -118.485 166.085 -118.155 ;
        RECT 165.755 -119.845 166.085 -119.515 ;
        RECT 165.755 -121.205 166.085 -120.875 ;
        RECT 165.755 -122.565 166.085 -122.235 ;
        RECT 165.755 -123.925 166.085 -123.595 ;
        RECT 165.755 -125.285 166.085 -124.955 ;
        RECT 165.755 -126.645 166.085 -126.315 ;
        RECT 165.755 -128.005 166.085 -127.675 ;
        RECT 165.755 -129.365 166.085 -129.035 ;
        RECT 165.755 -130.725 166.085 -130.395 ;
        RECT 165.755 -132.085 166.085 -131.755 ;
        RECT 165.755 -133.445 166.085 -133.115 ;
        RECT 165.755 -134.805 166.085 -134.475 ;
        RECT 165.755 -136.165 166.085 -135.835 ;
        RECT 165.755 -137.525 166.085 -137.195 ;
        RECT 165.755 -138.885 166.085 -138.555 ;
        RECT 165.755 -140.245 166.085 -139.915 ;
        RECT 165.755 -141.605 166.085 -141.275 ;
        RECT 165.755 -142.965 166.085 -142.635 ;
        RECT 165.755 -144.325 166.085 -143.995 ;
        RECT 165.755 -145.685 166.085 -145.355 ;
        RECT 165.755 -147.045 166.085 -146.715 ;
        RECT 165.755 -148.405 166.085 -148.075 ;
        RECT 165.755 -149.765 166.085 -149.435 ;
        RECT 165.755 -151.125 166.085 -150.795 ;
        RECT 165.755 -152.485 166.085 -152.155 ;
        RECT 165.755 -153.845 166.085 -153.515 ;
        RECT 165.755 -155.205 166.085 -154.875 ;
        RECT 165.755 -156.565 166.085 -156.235 ;
        RECT 165.755 -157.925 166.085 -157.595 ;
        RECT 165.755 -160.17 166.085 -159.04 ;
        RECT 165.76 -160.285 166.08 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 127.225 167.445 128.355 ;
        RECT 167.115 124.955 167.445 125.285 ;
        RECT 167.115 123.595 167.445 123.925 ;
        RECT 167.12 123.595 167.44 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 -95.365 167.445 -95.035 ;
        RECT 167.115 -96.725 167.445 -96.395 ;
        RECT 167.115 -98.085 167.445 -97.755 ;
        RECT 167.115 -99.445 167.445 -99.115 ;
        RECT 167.115 -100.805 167.445 -100.475 ;
        RECT 167.115 -102.165 167.445 -101.835 ;
        RECT 167.115 -103.525 167.445 -103.195 ;
        RECT 167.115 -104.885 167.445 -104.555 ;
        RECT 167.115 -106.245 167.445 -105.915 ;
        RECT 167.115 -107.605 167.445 -107.275 ;
        RECT 167.115 -108.965 167.445 -108.635 ;
        RECT 167.115 -110.325 167.445 -109.995 ;
        RECT 167.115 -111.685 167.445 -111.355 ;
        RECT 167.115 -113.045 167.445 -112.715 ;
        RECT 167.115 -114.405 167.445 -114.075 ;
        RECT 167.115 -115.765 167.445 -115.435 ;
        RECT 167.115 -117.125 167.445 -116.795 ;
        RECT 167.115 -118.485 167.445 -118.155 ;
        RECT 167.115 -119.845 167.445 -119.515 ;
        RECT 167.115 -121.205 167.445 -120.875 ;
        RECT 167.115 -122.565 167.445 -122.235 ;
        RECT 167.115 -123.925 167.445 -123.595 ;
        RECT 167.115 -125.285 167.445 -124.955 ;
        RECT 167.115 -126.645 167.445 -126.315 ;
        RECT 167.115 -128.005 167.445 -127.675 ;
        RECT 167.115 -129.365 167.445 -129.035 ;
        RECT 167.115 -130.725 167.445 -130.395 ;
        RECT 167.115 -132.085 167.445 -131.755 ;
        RECT 167.115 -133.445 167.445 -133.115 ;
        RECT 167.115 -134.805 167.445 -134.475 ;
        RECT 167.115 -136.165 167.445 -135.835 ;
        RECT 167.115 -137.525 167.445 -137.195 ;
        RECT 167.115 -138.885 167.445 -138.555 ;
        RECT 167.115 -140.245 167.445 -139.915 ;
        RECT 167.115 -141.605 167.445 -141.275 ;
        RECT 167.115 -142.965 167.445 -142.635 ;
        RECT 167.115 -144.325 167.445 -143.995 ;
        RECT 167.115 -145.685 167.445 -145.355 ;
        RECT 167.115 -147.045 167.445 -146.715 ;
        RECT 167.115 -148.405 167.445 -148.075 ;
        RECT 167.115 -149.765 167.445 -149.435 ;
        RECT 167.115 -151.125 167.445 -150.795 ;
        RECT 167.115 -152.485 167.445 -152.155 ;
        RECT 167.115 -153.845 167.445 -153.515 ;
        RECT 167.115 -155.205 167.445 -154.875 ;
        RECT 167.115 -156.565 167.445 -156.235 ;
        RECT 167.115 -157.925 167.445 -157.595 ;
        RECT 167.115 -160.17 167.445 -159.04 ;
        RECT 167.12 -160.285 167.44 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.01 -94.075 168.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 127.225 168.805 128.355 ;
        RECT 168.475 124.955 168.805 125.285 ;
        RECT 168.475 123.595 168.805 123.925 ;
        RECT 168.48 123.595 168.8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 127.225 170.165 128.355 ;
        RECT 169.835 124.955 170.165 125.285 ;
        RECT 169.835 123.595 170.165 123.925 ;
        RECT 169.84 123.595 170.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 -1.525 170.165 -1.195 ;
        RECT 169.835 -2.885 170.165 -2.555 ;
        RECT 169.84 -3.56 170.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 127.225 171.525 128.355 ;
        RECT 171.195 124.955 171.525 125.285 ;
        RECT 171.195 123.595 171.525 123.925 ;
        RECT 171.2 123.595 171.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -1.525 171.525 -1.195 ;
        RECT 171.195 -2.885 171.525 -2.555 ;
        RECT 171.2 -3.56 171.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -91.285 171.525 -90.955 ;
        RECT 171.195 -92.645 171.525 -92.315 ;
        RECT 171.195 -94.005 171.525 -93.675 ;
        RECT 171.195 -95.365 171.525 -95.035 ;
        RECT 171.195 -96.725 171.525 -96.395 ;
        RECT 171.195 -98.085 171.525 -97.755 ;
        RECT 171.195 -99.445 171.525 -99.115 ;
        RECT 171.195 -100.805 171.525 -100.475 ;
        RECT 171.195 -102.165 171.525 -101.835 ;
        RECT 171.195 -103.525 171.525 -103.195 ;
        RECT 171.195 -104.885 171.525 -104.555 ;
        RECT 171.195 -106.245 171.525 -105.915 ;
        RECT 171.195 -107.605 171.525 -107.275 ;
        RECT 171.195 -108.965 171.525 -108.635 ;
        RECT 171.195 -110.325 171.525 -109.995 ;
        RECT 171.195 -111.685 171.525 -111.355 ;
        RECT 171.195 -113.045 171.525 -112.715 ;
        RECT 171.195 -114.405 171.525 -114.075 ;
        RECT 171.195 -115.765 171.525 -115.435 ;
        RECT 171.195 -117.125 171.525 -116.795 ;
        RECT 171.195 -118.485 171.525 -118.155 ;
        RECT 171.195 -119.845 171.525 -119.515 ;
        RECT 171.195 -121.205 171.525 -120.875 ;
        RECT 171.195 -122.565 171.525 -122.235 ;
        RECT 171.195 -123.925 171.525 -123.595 ;
        RECT 171.195 -125.285 171.525 -124.955 ;
        RECT 171.195 -126.645 171.525 -126.315 ;
        RECT 171.195 -128.005 171.525 -127.675 ;
        RECT 171.195 -129.365 171.525 -129.035 ;
        RECT 171.195 -130.725 171.525 -130.395 ;
        RECT 171.195 -132.085 171.525 -131.755 ;
        RECT 171.195 -133.445 171.525 -133.115 ;
        RECT 171.195 -134.805 171.525 -134.475 ;
        RECT 171.195 -136.165 171.525 -135.835 ;
        RECT 171.195 -137.525 171.525 -137.195 ;
        RECT 171.195 -138.885 171.525 -138.555 ;
        RECT 171.195 -140.245 171.525 -139.915 ;
        RECT 171.195 -141.605 171.525 -141.275 ;
        RECT 171.195 -142.965 171.525 -142.635 ;
        RECT 171.195 -144.325 171.525 -143.995 ;
        RECT 171.195 -145.685 171.525 -145.355 ;
        RECT 171.195 -147.045 171.525 -146.715 ;
        RECT 171.195 -148.405 171.525 -148.075 ;
        RECT 171.195 -149.765 171.525 -149.435 ;
        RECT 171.195 -151.125 171.525 -150.795 ;
        RECT 171.195 -152.485 171.525 -152.155 ;
        RECT 171.195 -153.845 171.525 -153.515 ;
        RECT 171.195 -155.205 171.525 -154.875 ;
        RECT 171.195 -156.565 171.525 -156.235 ;
        RECT 171.195 -157.925 171.525 -157.595 ;
        RECT 171.195 -160.17 171.525 -159.04 ;
        RECT 171.2 -160.285 171.52 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 127.225 172.885 128.355 ;
        RECT 172.555 124.955 172.885 125.285 ;
        RECT 172.555 123.595 172.885 123.925 ;
        RECT 172.56 123.595 172.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -1.525 172.885 -1.195 ;
        RECT 172.555 -2.885 172.885 -2.555 ;
        RECT 172.56 -3.56 172.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -91.285 172.885 -90.955 ;
        RECT 172.555 -92.645 172.885 -92.315 ;
        RECT 172.555 -94.005 172.885 -93.675 ;
        RECT 172.555 -95.365 172.885 -95.035 ;
        RECT 172.555 -96.725 172.885 -96.395 ;
        RECT 172.555 -98.085 172.885 -97.755 ;
        RECT 172.555 -99.445 172.885 -99.115 ;
        RECT 172.555 -100.805 172.885 -100.475 ;
        RECT 172.555 -102.165 172.885 -101.835 ;
        RECT 172.555 -103.525 172.885 -103.195 ;
        RECT 172.555 -104.885 172.885 -104.555 ;
        RECT 172.555 -106.245 172.885 -105.915 ;
        RECT 172.555 -107.605 172.885 -107.275 ;
        RECT 172.555 -108.965 172.885 -108.635 ;
        RECT 172.555 -110.325 172.885 -109.995 ;
        RECT 172.555 -111.685 172.885 -111.355 ;
        RECT 172.555 -113.045 172.885 -112.715 ;
        RECT 172.555 -114.405 172.885 -114.075 ;
        RECT 172.555 -115.765 172.885 -115.435 ;
        RECT 172.555 -117.125 172.885 -116.795 ;
        RECT 172.555 -118.485 172.885 -118.155 ;
        RECT 172.555 -119.845 172.885 -119.515 ;
        RECT 172.555 -121.205 172.885 -120.875 ;
        RECT 172.555 -122.565 172.885 -122.235 ;
        RECT 172.555 -123.925 172.885 -123.595 ;
        RECT 172.555 -125.285 172.885 -124.955 ;
        RECT 172.555 -126.645 172.885 -126.315 ;
        RECT 172.555 -128.005 172.885 -127.675 ;
        RECT 172.555 -129.365 172.885 -129.035 ;
        RECT 172.555 -130.725 172.885 -130.395 ;
        RECT 172.555 -132.085 172.885 -131.755 ;
        RECT 172.555 -133.445 172.885 -133.115 ;
        RECT 172.555 -134.805 172.885 -134.475 ;
        RECT 172.555 -136.165 172.885 -135.835 ;
        RECT 172.555 -137.525 172.885 -137.195 ;
        RECT 172.555 -138.885 172.885 -138.555 ;
        RECT 172.555 -140.245 172.885 -139.915 ;
        RECT 172.555 -141.605 172.885 -141.275 ;
        RECT 172.555 -142.965 172.885 -142.635 ;
        RECT 172.555 -144.325 172.885 -143.995 ;
        RECT 172.555 -145.685 172.885 -145.355 ;
        RECT 172.555 -147.045 172.885 -146.715 ;
        RECT 172.555 -148.405 172.885 -148.075 ;
        RECT 172.555 -149.765 172.885 -149.435 ;
        RECT 172.555 -151.125 172.885 -150.795 ;
        RECT 172.555 -152.485 172.885 -152.155 ;
        RECT 172.555 -153.845 172.885 -153.515 ;
        RECT 172.555 -155.205 172.885 -154.875 ;
        RECT 172.555 -156.565 172.885 -156.235 ;
        RECT 172.555 -157.925 172.885 -157.595 ;
        RECT 172.555 -160.17 172.885 -159.04 ;
        RECT 172.56 -160.285 172.88 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 127.225 174.245 128.355 ;
        RECT 173.915 124.955 174.245 125.285 ;
        RECT 173.915 123.595 174.245 123.925 ;
        RECT 173.92 123.595 174.24 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 -95.365 174.245 -95.035 ;
        RECT 173.915 -96.725 174.245 -96.395 ;
        RECT 173.915 -98.085 174.245 -97.755 ;
        RECT 173.915 -99.445 174.245 -99.115 ;
        RECT 173.915 -100.805 174.245 -100.475 ;
        RECT 173.915 -102.165 174.245 -101.835 ;
        RECT 173.915 -103.525 174.245 -103.195 ;
        RECT 173.915 -104.885 174.245 -104.555 ;
        RECT 173.915 -106.245 174.245 -105.915 ;
        RECT 173.915 -107.605 174.245 -107.275 ;
        RECT 173.915 -108.965 174.245 -108.635 ;
        RECT 173.915 -110.325 174.245 -109.995 ;
        RECT 173.915 -111.685 174.245 -111.355 ;
        RECT 173.915 -113.045 174.245 -112.715 ;
        RECT 173.915 -114.405 174.245 -114.075 ;
        RECT 173.915 -115.765 174.245 -115.435 ;
        RECT 173.915 -117.125 174.245 -116.795 ;
        RECT 173.915 -118.485 174.245 -118.155 ;
        RECT 173.915 -119.845 174.245 -119.515 ;
        RECT 173.915 -121.205 174.245 -120.875 ;
        RECT 173.915 -122.565 174.245 -122.235 ;
        RECT 173.915 -123.925 174.245 -123.595 ;
        RECT 173.915 -125.285 174.245 -124.955 ;
        RECT 173.915 -126.645 174.245 -126.315 ;
        RECT 173.915 -128.005 174.245 -127.675 ;
        RECT 173.915 -129.365 174.245 -129.035 ;
        RECT 173.915 -130.725 174.245 -130.395 ;
        RECT 173.915 -132.085 174.245 -131.755 ;
        RECT 173.915 -133.445 174.245 -133.115 ;
        RECT 173.915 -134.805 174.245 -134.475 ;
        RECT 173.915 -136.165 174.245 -135.835 ;
        RECT 173.915 -137.525 174.245 -137.195 ;
        RECT 173.915 -138.885 174.245 -138.555 ;
        RECT 173.915 -140.245 174.245 -139.915 ;
        RECT 173.915 -141.605 174.245 -141.275 ;
        RECT 173.915 -142.965 174.245 -142.635 ;
        RECT 173.915 -144.325 174.245 -143.995 ;
        RECT 173.915 -145.685 174.245 -145.355 ;
        RECT 173.915 -147.045 174.245 -146.715 ;
        RECT 173.915 -148.405 174.245 -148.075 ;
        RECT 173.915 -149.765 174.245 -149.435 ;
        RECT 173.915 -151.125 174.245 -150.795 ;
        RECT 173.915 -152.485 174.245 -152.155 ;
        RECT 173.915 -153.845 174.245 -153.515 ;
        RECT 173.915 -155.205 174.245 -154.875 ;
        RECT 173.915 -156.565 174.245 -156.235 ;
        RECT 173.915 -157.925 174.245 -157.595 ;
        RECT 173.915 -160.17 174.245 -159.04 ;
        RECT 173.92 -160.285 174.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.11 -94.075 174.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 127.225 175.605 128.355 ;
        RECT 175.275 124.955 175.605 125.285 ;
        RECT 175.275 123.595 175.605 123.925 ;
        RECT 175.28 123.595 175.6 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -1.525 175.605 -1.195 ;
        RECT 175.275 -2.885 175.605 -2.555 ;
        RECT 175.28 -3.56 175.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 127.225 176.965 128.355 ;
        RECT 176.635 124.955 176.965 125.285 ;
        RECT 176.635 123.595 176.965 123.925 ;
        RECT 176.64 123.595 176.96 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 -1.525 176.965 -1.195 ;
        RECT 176.635 -2.885 176.965 -2.555 ;
        RECT 176.64 -3.56 176.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 127.225 178.325 128.355 ;
        RECT 177.995 124.955 178.325 125.285 ;
        RECT 177.995 123.595 178.325 123.925 ;
        RECT 178 123.595 178.32 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 -1.525 178.325 -1.195 ;
        RECT 177.995 -2.885 178.325 -2.555 ;
        RECT 178 -3.56 178.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 -91.285 178.325 -90.955 ;
        RECT 177.995 -92.645 178.325 -92.315 ;
        RECT 177.995 -94.005 178.325 -93.675 ;
        RECT 177.995 -95.365 178.325 -95.035 ;
        RECT 177.995 -96.725 178.325 -96.395 ;
        RECT 177.995 -98.085 178.325 -97.755 ;
        RECT 177.995 -99.445 178.325 -99.115 ;
        RECT 177.995 -100.805 178.325 -100.475 ;
        RECT 177.995 -102.165 178.325 -101.835 ;
        RECT 177.995 -103.525 178.325 -103.195 ;
        RECT 177.995 -104.885 178.325 -104.555 ;
        RECT 177.995 -106.245 178.325 -105.915 ;
        RECT 177.995 -107.605 178.325 -107.275 ;
        RECT 177.995 -108.965 178.325 -108.635 ;
        RECT 177.995 -110.325 178.325 -109.995 ;
        RECT 177.995 -111.685 178.325 -111.355 ;
        RECT 177.995 -113.045 178.325 -112.715 ;
        RECT 177.995 -114.405 178.325 -114.075 ;
        RECT 177.995 -115.765 178.325 -115.435 ;
        RECT 177.995 -117.125 178.325 -116.795 ;
        RECT 177.995 -118.485 178.325 -118.155 ;
        RECT 177.995 -119.845 178.325 -119.515 ;
        RECT 177.995 -121.205 178.325 -120.875 ;
        RECT 177.995 -122.565 178.325 -122.235 ;
        RECT 177.995 -123.925 178.325 -123.595 ;
        RECT 177.995 -125.285 178.325 -124.955 ;
        RECT 177.995 -126.645 178.325 -126.315 ;
        RECT 177.995 -128.005 178.325 -127.675 ;
        RECT 177.995 -129.365 178.325 -129.035 ;
        RECT 177.995 -130.725 178.325 -130.395 ;
        RECT 177.995 -132.085 178.325 -131.755 ;
        RECT 177.995 -133.445 178.325 -133.115 ;
        RECT 177.995 -134.805 178.325 -134.475 ;
        RECT 177.995 -136.165 178.325 -135.835 ;
        RECT 177.995 -137.525 178.325 -137.195 ;
        RECT 177.995 -138.885 178.325 -138.555 ;
        RECT 177.995 -140.245 178.325 -139.915 ;
        RECT 177.995 -141.605 178.325 -141.275 ;
        RECT 177.995 -142.965 178.325 -142.635 ;
        RECT 177.995 -144.325 178.325 -143.995 ;
        RECT 177.995 -145.685 178.325 -145.355 ;
        RECT 177.995 -147.045 178.325 -146.715 ;
        RECT 177.995 -148.405 178.325 -148.075 ;
        RECT 177.995 -149.765 178.325 -149.435 ;
        RECT 177.995 -151.125 178.325 -150.795 ;
        RECT 177.995 -152.485 178.325 -152.155 ;
        RECT 177.995 -153.845 178.325 -153.515 ;
        RECT 177.995 -155.205 178.325 -154.875 ;
        RECT 177.995 -156.565 178.325 -156.235 ;
        RECT 177.995 -157.925 178.325 -157.595 ;
        RECT 177.995 -160.17 178.325 -159.04 ;
        RECT 178 -160.285 178.32 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 127.225 179.685 128.355 ;
        RECT 179.355 124.955 179.685 125.285 ;
        RECT 179.355 123.595 179.685 123.925 ;
        RECT 179.36 123.595 179.68 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 -95.365 179.685 -95.035 ;
        RECT 179.355 -96.725 179.685 -96.395 ;
        RECT 179.355 -98.085 179.685 -97.755 ;
        RECT 179.355 -99.445 179.685 -99.115 ;
        RECT 179.355 -100.805 179.685 -100.475 ;
        RECT 179.355 -102.165 179.685 -101.835 ;
        RECT 179.355 -103.525 179.685 -103.195 ;
        RECT 179.355 -104.885 179.685 -104.555 ;
        RECT 179.355 -106.245 179.685 -105.915 ;
        RECT 179.355 -107.605 179.685 -107.275 ;
        RECT 179.355 -108.965 179.685 -108.635 ;
        RECT 179.355 -110.325 179.685 -109.995 ;
        RECT 179.355 -111.685 179.685 -111.355 ;
        RECT 179.355 -113.045 179.685 -112.715 ;
        RECT 179.355 -114.405 179.685 -114.075 ;
        RECT 179.355 -115.765 179.685 -115.435 ;
        RECT 179.355 -117.125 179.685 -116.795 ;
        RECT 179.355 -118.485 179.685 -118.155 ;
        RECT 179.355 -119.845 179.685 -119.515 ;
        RECT 179.355 -121.205 179.685 -120.875 ;
        RECT 179.355 -122.565 179.685 -122.235 ;
        RECT 179.355 -123.925 179.685 -123.595 ;
        RECT 179.355 -125.285 179.685 -124.955 ;
        RECT 179.355 -126.645 179.685 -126.315 ;
        RECT 179.355 -128.005 179.685 -127.675 ;
        RECT 179.355 -129.365 179.685 -129.035 ;
        RECT 179.355 -130.725 179.685 -130.395 ;
        RECT 179.355 -132.085 179.685 -131.755 ;
        RECT 179.355 -133.445 179.685 -133.115 ;
        RECT 179.355 -134.805 179.685 -134.475 ;
        RECT 179.355 -136.165 179.685 -135.835 ;
        RECT 179.355 -137.525 179.685 -137.195 ;
        RECT 179.355 -138.885 179.685 -138.555 ;
        RECT 179.355 -140.245 179.685 -139.915 ;
        RECT 179.355 -141.605 179.685 -141.275 ;
        RECT 179.355 -142.965 179.685 -142.635 ;
        RECT 179.355 -144.325 179.685 -143.995 ;
        RECT 179.355 -145.685 179.685 -145.355 ;
        RECT 179.355 -147.045 179.685 -146.715 ;
        RECT 179.355 -148.405 179.685 -148.075 ;
        RECT 179.355 -149.765 179.685 -149.435 ;
        RECT 179.355 -151.125 179.685 -150.795 ;
        RECT 179.355 -152.485 179.685 -152.155 ;
        RECT 179.355 -153.845 179.685 -153.515 ;
        RECT 179.355 -155.205 179.685 -154.875 ;
        RECT 179.355 -156.565 179.685 -156.235 ;
        RECT 179.355 -157.925 179.685 -157.595 ;
        RECT 179.355 -160.17 179.685 -159.04 ;
        RECT 179.36 -160.285 179.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.21 -94.075 180.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 127.225 181.045 128.355 ;
        RECT 180.715 124.955 181.045 125.285 ;
        RECT 180.715 123.595 181.045 123.925 ;
        RECT 180.72 123.595 181.04 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 127.225 182.405 128.355 ;
        RECT 182.075 124.955 182.405 125.285 ;
        RECT 182.075 123.595 182.405 123.925 ;
        RECT 182.08 123.595 182.4 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 -1.525 182.405 -1.195 ;
        RECT 182.075 -2.885 182.405 -2.555 ;
        RECT 182.08 -3.56 182.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 127.225 183.765 128.355 ;
        RECT 183.435 124.955 183.765 125.285 ;
        RECT 183.435 123.595 183.765 123.925 ;
        RECT 183.44 123.595 183.76 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -1.525 183.765 -1.195 ;
        RECT 183.435 -2.885 183.765 -2.555 ;
        RECT 183.44 -3.56 183.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -91.285 183.765 -90.955 ;
        RECT 183.435 -92.645 183.765 -92.315 ;
        RECT 183.435 -94.005 183.765 -93.675 ;
        RECT 183.435 -95.365 183.765 -95.035 ;
        RECT 183.435 -96.725 183.765 -96.395 ;
        RECT 183.435 -98.085 183.765 -97.755 ;
        RECT 183.435 -99.445 183.765 -99.115 ;
        RECT 183.435 -100.805 183.765 -100.475 ;
        RECT 183.435 -102.165 183.765 -101.835 ;
        RECT 183.435 -103.525 183.765 -103.195 ;
        RECT 183.435 -104.885 183.765 -104.555 ;
        RECT 183.435 -106.245 183.765 -105.915 ;
        RECT 183.435 -107.605 183.765 -107.275 ;
        RECT 183.435 -108.965 183.765 -108.635 ;
        RECT 183.435 -110.325 183.765 -109.995 ;
        RECT 183.435 -111.685 183.765 -111.355 ;
        RECT 183.435 -113.045 183.765 -112.715 ;
        RECT 183.435 -114.405 183.765 -114.075 ;
        RECT 183.435 -115.765 183.765 -115.435 ;
        RECT 183.435 -117.125 183.765 -116.795 ;
        RECT 183.435 -118.485 183.765 -118.155 ;
        RECT 183.435 -119.845 183.765 -119.515 ;
        RECT 183.435 -121.205 183.765 -120.875 ;
        RECT 183.435 -122.565 183.765 -122.235 ;
        RECT 183.435 -123.925 183.765 -123.595 ;
        RECT 183.435 -125.285 183.765 -124.955 ;
        RECT 183.435 -126.645 183.765 -126.315 ;
        RECT 183.435 -128.005 183.765 -127.675 ;
        RECT 183.435 -129.365 183.765 -129.035 ;
        RECT 183.435 -130.725 183.765 -130.395 ;
        RECT 183.435 -132.085 183.765 -131.755 ;
        RECT 183.435 -133.445 183.765 -133.115 ;
        RECT 183.435 -134.805 183.765 -134.475 ;
        RECT 183.435 -136.165 183.765 -135.835 ;
        RECT 183.435 -137.525 183.765 -137.195 ;
        RECT 183.435 -138.885 183.765 -138.555 ;
        RECT 183.435 -140.245 183.765 -139.915 ;
        RECT 183.435 -141.605 183.765 -141.275 ;
        RECT 183.435 -142.965 183.765 -142.635 ;
        RECT 183.435 -144.325 183.765 -143.995 ;
        RECT 183.435 -145.685 183.765 -145.355 ;
        RECT 183.435 -147.045 183.765 -146.715 ;
        RECT 183.435 -148.405 183.765 -148.075 ;
        RECT 183.435 -149.765 183.765 -149.435 ;
        RECT 183.435 -151.125 183.765 -150.795 ;
        RECT 183.435 -152.485 183.765 -152.155 ;
        RECT 183.435 -153.845 183.765 -153.515 ;
        RECT 183.435 -155.205 183.765 -154.875 ;
        RECT 183.435 -156.565 183.765 -156.235 ;
        RECT 183.435 -157.925 183.765 -157.595 ;
        RECT 183.435 -160.17 183.765 -159.04 ;
        RECT 183.44 -160.285 183.76 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 127.225 185.125 128.355 ;
        RECT 184.795 124.955 185.125 125.285 ;
        RECT 184.795 123.595 185.125 123.925 ;
        RECT 184.8 123.595 185.12 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -1.525 185.125 -1.195 ;
        RECT 184.795 -2.885 185.125 -2.555 ;
        RECT 184.8 -3.56 185.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -91.285 185.125 -90.955 ;
        RECT 184.795 -92.645 185.125 -92.315 ;
        RECT 184.795 -94.005 185.125 -93.675 ;
        RECT 184.795 -95.365 185.125 -95.035 ;
        RECT 184.795 -96.725 185.125 -96.395 ;
        RECT 184.795 -98.085 185.125 -97.755 ;
        RECT 184.795 -99.445 185.125 -99.115 ;
        RECT 184.795 -100.805 185.125 -100.475 ;
        RECT 184.795 -102.165 185.125 -101.835 ;
        RECT 184.795 -103.525 185.125 -103.195 ;
        RECT 184.795 -104.885 185.125 -104.555 ;
        RECT 184.795 -106.245 185.125 -105.915 ;
        RECT 184.795 -107.605 185.125 -107.275 ;
        RECT 184.795 -108.965 185.125 -108.635 ;
        RECT 184.795 -110.325 185.125 -109.995 ;
        RECT 184.795 -111.685 185.125 -111.355 ;
        RECT 184.795 -113.045 185.125 -112.715 ;
        RECT 184.795 -114.405 185.125 -114.075 ;
        RECT 184.795 -115.765 185.125 -115.435 ;
        RECT 184.795 -117.125 185.125 -116.795 ;
        RECT 184.795 -118.485 185.125 -118.155 ;
        RECT 184.795 -119.845 185.125 -119.515 ;
        RECT 184.795 -121.205 185.125 -120.875 ;
        RECT 184.795 -122.565 185.125 -122.235 ;
        RECT 184.795 -123.925 185.125 -123.595 ;
        RECT 184.795 -125.285 185.125 -124.955 ;
        RECT 184.795 -126.645 185.125 -126.315 ;
        RECT 184.795 -128.005 185.125 -127.675 ;
        RECT 184.795 -129.365 185.125 -129.035 ;
        RECT 184.795 -130.725 185.125 -130.395 ;
        RECT 184.795 -132.085 185.125 -131.755 ;
        RECT 184.795 -133.445 185.125 -133.115 ;
        RECT 184.795 -134.805 185.125 -134.475 ;
        RECT 184.795 -136.165 185.125 -135.835 ;
        RECT 184.795 -137.525 185.125 -137.195 ;
        RECT 184.795 -138.885 185.125 -138.555 ;
        RECT 184.795 -140.245 185.125 -139.915 ;
        RECT 184.795 -141.605 185.125 -141.275 ;
        RECT 184.795 -142.965 185.125 -142.635 ;
        RECT 184.795 -144.325 185.125 -143.995 ;
        RECT 184.795 -145.685 185.125 -145.355 ;
        RECT 184.795 -147.045 185.125 -146.715 ;
        RECT 184.795 -148.405 185.125 -148.075 ;
        RECT 184.795 -149.765 185.125 -149.435 ;
        RECT 184.795 -151.125 185.125 -150.795 ;
        RECT 184.795 -152.485 185.125 -152.155 ;
        RECT 184.795 -153.845 185.125 -153.515 ;
        RECT 184.795 -155.205 185.125 -154.875 ;
        RECT 184.795 -156.565 185.125 -156.235 ;
        RECT 184.795 -157.925 185.125 -157.595 ;
        RECT 184.795 -160.17 185.125 -159.04 ;
        RECT 184.8 -160.285 185.12 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 127.225 186.485 128.355 ;
        RECT 186.155 124.955 186.485 125.285 ;
        RECT 186.155 123.595 186.485 123.925 ;
        RECT 186.16 123.595 186.48 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 -95.365 186.485 -95.035 ;
        RECT 186.155 -96.725 186.485 -96.395 ;
        RECT 186.155 -98.085 186.485 -97.755 ;
        RECT 186.155 -99.445 186.485 -99.115 ;
        RECT 186.155 -100.805 186.485 -100.475 ;
        RECT 186.155 -102.165 186.485 -101.835 ;
        RECT 186.155 -103.525 186.485 -103.195 ;
        RECT 186.155 -104.885 186.485 -104.555 ;
        RECT 186.155 -106.245 186.485 -105.915 ;
        RECT 186.155 -107.605 186.485 -107.275 ;
        RECT 186.155 -108.965 186.485 -108.635 ;
        RECT 186.155 -110.325 186.485 -109.995 ;
        RECT 186.155 -111.685 186.485 -111.355 ;
        RECT 186.155 -113.045 186.485 -112.715 ;
        RECT 186.155 -114.405 186.485 -114.075 ;
        RECT 186.155 -115.765 186.485 -115.435 ;
        RECT 186.155 -117.125 186.485 -116.795 ;
        RECT 186.155 -118.485 186.485 -118.155 ;
        RECT 186.155 -119.845 186.485 -119.515 ;
        RECT 186.155 -121.205 186.485 -120.875 ;
        RECT 186.155 -122.565 186.485 -122.235 ;
        RECT 186.155 -123.925 186.485 -123.595 ;
        RECT 186.155 -125.285 186.485 -124.955 ;
        RECT 186.155 -126.645 186.485 -126.315 ;
        RECT 186.155 -128.005 186.485 -127.675 ;
        RECT 186.155 -129.365 186.485 -129.035 ;
        RECT 186.155 -130.725 186.485 -130.395 ;
        RECT 186.155 -132.085 186.485 -131.755 ;
        RECT 186.155 -133.445 186.485 -133.115 ;
        RECT 186.155 -134.805 186.485 -134.475 ;
        RECT 186.155 -136.165 186.485 -135.835 ;
        RECT 186.155 -137.525 186.485 -137.195 ;
        RECT 186.155 -138.885 186.485 -138.555 ;
        RECT 186.155 -140.245 186.485 -139.915 ;
        RECT 186.155 -141.605 186.485 -141.275 ;
        RECT 186.155 -142.965 186.485 -142.635 ;
        RECT 186.155 -144.325 186.485 -143.995 ;
        RECT 186.155 -145.685 186.485 -145.355 ;
        RECT 186.155 -147.045 186.485 -146.715 ;
        RECT 186.155 -148.405 186.485 -148.075 ;
        RECT 186.155 -149.765 186.485 -149.435 ;
        RECT 186.155 -151.125 186.485 -150.795 ;
        RECT 186.155 -152.485 186.485 -152.155 ;
        RECT 186.155 -153.845 186.485 -153.515 ;
        RECT 186.155 -155.205 186.485 -154.875 ;
        RECT 186.155 -156.565 186.485 -156.235 ;
        RECT 186.155 -157.925 186.485 -157.595 ;
        RECT 186.155 -160.17 186.485 -159.04 ;
        RECT 186.16 -160.285 186.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.31 -94.075 186.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 127.225 187.845 128.355 ;
        RECT 187.515 124.955 187.845 125.285 ;
        RECT 187.515 123.595 187.845 123.925 ;
        RECT 187.52 123.595 187.84 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 -1.525 187.845 -1.195 ;
        RECT 187.515 -2.885 187.845 -2.555 ;
        RECT 187.52 -3.56 187.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 127.225 189.205 128.355 ;
        RECT 188.875 124.955 189.205 125.285 ;
        RECT 188.875 123.595 189.205 123.925 ;
        RECT 188.88 123.595 189.2 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 -1.525 189.205 -1.195 ;
        RECT 188.875 -2.885 189.205 -2.555 ;
        RECT 188.88 -3.56 189.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 127.225 190.565 128.355 ;
        RECT 190.235 124.955 190.565 125.285 ;
        RECT 190.235 123.595 190.565 123.925 ;
        RECT 190.24 123.595 190.56 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 -1.525 190.565 -1.195 ;
        RECT 190.235 -2.885 190.565 -2.555 ;
        RECT 190.24 -3.56 190.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 -91.285 190.565 -90.955 ;
        RECT 190.235 -92.645 190.565 -92.315 ;
        RECT 190.235 -94.005 190.565 -93.675 ;
        RECT 190.235 -95.365 190.565 -95.035 ;
        RECT 190.235 -96.725 190.565 -96.395 ;
        RECT 190.235 -98.085 190.565 -97.755 ;
        RECT 190.235 -99.445 190.565 -99.115 ;
        RECT 190.235 -100.805 190.565 -100.475 ;
        RECT 190.235 -102.165 190.565 -101.835 ;
        RECT 190.235 -103.525 190.565 -103.195 ;
        RECT 190.235 -104.885 190.565 -104.555 ;
        RECT 190.235 -106.245 190.565 -105.915 ;
        RECT 190.235 -107.605 190.565 -107.275 ;
        RECT 190.235 -108.965 190.565 -108.635 ;
        RECT 190.235 -110.325 190.565 -109.995 ;
        RECT 190.235 -111.685 190.565 -111.355 ;
        RECT 190.235 -113.045 190.565 -112.715 ;
        RECT 190.235 -114.405 190.565 -114.075 ;
        RECT 190.235 -115.765 190.565 -115.435 ;
        RECT 190.235 -117.125 190.565 -116.795 ;
        RECT 190.235 -118.485 190.565 -118.155 ;
        RECT 190.235 -119.845 190.565 -119.515 ;
        RECT 190.235 -121.205 190.565 -120.875 ;
        RECT 190.235 -122.565 190.565 -122.235 ;
        RECT 190.235 -123.925 190.565 -123.595 ;
        RECT 190.235 -125.285 190.565 -124.955 ;
        RECT 190.235 -126.645 190.565 -126.315 ;
        RECT 190.235 -128.005 190.565 -127.675 ;
        RECT 190.235 -129.365 190.565 -129.035 ;
        RECT 190.235 -130.725 190.565 -130.395 ;
        RECT 190.235 -132.085 190.565 -131.755 ;
        RECT 190.235 -133.445 190.565 -133.115 ;
        RECT 190.235 -134.805 190.565 -134.475 ;
        RECT 190.235 -136.165 190.565 -135.835 ;
        RECT 190.235 -137.525 190.565 -137.195 ;
        RECT 190.235 -138.885 190.565 -138.555 ;
        RECT 190.235 -140.245 190.565 -139.915 ;
        RECT 190.235 -141.605 190.565 -141.275 ;
        RECT 190.235 -142.965 190.565 -142.635 ;
        RECT 190.235 -144.325 190.565 -143.995 ;
        RECT 190.235 -145.685 190.565 -145.355 ;
        RECT 190.235 -147.045 190.565 -146.715 ;
        RECT 190.235 -148.405 190.565 -148.075 ;
        RECT 190.235 -149.765 190.565 -149.435 ;
        RECT 190.235 -151.125 190.565 -150.795 ;
        RECT 190.235 -152.485 190.565 -152.155 ;
        RECT 190.235 -153.845 190.565 -153.515 ;
        RECT 190.235 -155.205 190.565 -154.875 ;
        RECT 190.235 -156.565 190.565 -156.235 ;
        RECT 190.235 -157.925 190.565 -157.595 ;
        RECT 190.235 -160.17 190.565 -159.04 ;
        RECT 190.24 -160.285 190.56 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 127.225 191.925 128.355 ;
        RECT 191.595 124.955 191.925 125.285 ;
        RECT 191.595 123.595 191.925 123.925 ;
        RECT 191.6 123.595 191.92 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 -95.365 191.925 -95.035 ;
        RECT 191.595 -96.725 191.925 -96.395 ;
        RECT 191.595 -98.085 191.925 -97.755 ;
        RECT 191.595 -99.445 191.925 -99.115 ;
        RECT 191.595 -100.805 191.925 -100.475 ;
        RECT 191.595 -102.165 191.925 -101.835 ;
        RECT 191.595 -103.525 191.925 -103.195 ;
        RECT 191.595 -104.885 191.925 -104.555 ;
        RECT 191.595 -106.245 191.925 -105.915 ;
        RECT 191.595 -107.605 191.925 -107.275 ;
        RECT 191.595 -108.965 191.925 -108.635 ;
        RECT 191.595 -110.325 191.925 -109.995 ;
        RECT 191.595 -111.685 191.925 -111.355 ;
        RECT 191.595 -113.045 191.925 -112.715 ;
        RECT 191.595 -114.405 191.925 -114.075 ;
        RECT 191.595 -115.765 191.925 -115.435 ;
        RECT 191.595 -117.125 191.925 -116.795 ;
        RECT 191.595 -118.485 191.925 -118.155 ;
        RECT 191.595 -119.845 191.925 -119.515 ;
        RECT 191.595 -121.205 191.925 -120.875 ;
        RECT 191.595 -122.565 191.925 -122.235 ;
        RECT 191.595 -123.925 191.925 -123.595 ;
        RECT 191.595 -125.285 191.925 -124.955 ;
        RECT 191.595 -126.645 191.925 -126.315 ;
        RECT 191.595 -128.005 191.925 -127.675 ;
        RECT 191.595 -129.365 191.925 -129.035 ;
        RECT 191.595 -130.725 191.925 -130.395 ;
        RECT 191.595 -132.085 191.925 -131.755 ;
        RECT 191.595 -133.445 191.925 -133.115 ;
        RECT 191.595 -134.805 191.925 -134.475 ;
        RECT 191.595 -136.165 191.925 -135.835 ;
        RECT 191.595 -137.525 191.925 -137.195 ;
        RECT 191.595 -138.885 191.925 -138.555 ;
        RECT 191.595 -140.245 191.925 -139.915 ;
        RECT 191.595 -141.605 191.925 -141.275 ;
        RECT 191.595 -142.965 191.925 -142.635 ;
        RECT 191.595 -144.325 191.925 -143.995 ;
        RECT 191.595 -145.685 191.925 -145.355 ;
        RECT 191.595 -147.045 191.925 -146.715 ;
        RECT 191.595 -148.405 191.925 -148.075 ;
        RECT 191.595 -149.765 191.925 -149.435 ;
        RECT 191.595 -151.125 191.925 -150.795 ;
        RECT 191.595 -152.485 191.925 -152.155 ;
        RECT 191.595 -153.845 191.925 -153.515 ;
        RECT 191.595 -155.205 191.925 -154.875 ;
        RECT 191.595 -156.565 191.925 -156.235 ;
        RECT 191.595 -157.925 191.925 -157.595 ;
        RECT 191.595 -160.17 191.925 -159.04 ;
        RECT 191.6 -160.285 191.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.41 -94.075 192.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 127.225 193.285 128.355 ;
        RECT 192.955 124.955 193.285 125.285 ;
        RECT 192.955 123.595 193.285 123.925 ;
        RECT 192.96 123.595 193.28 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 127.225 194.645 128.355 ;
        RECT 194.315 124.955 194.645 125.285 ;
        RECT 194.315 123.595 194.645 123.925 ;
        RECT 194.32 123.595 194.64 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 -1.525 194.645 -1.195 ;
        RECT 194.315 -2.885 194.645 -2.555 ;
        RECT 194.32 -3.56 194.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 127.225 196.005 128.355 ;
        RECT 195.675 124.955 196.005 125.285 ;
        RECT 195.675 123.595 196.005 123.925 ;
        RECT 195.68 123.595 196 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -1.525 196.005 -1.195 ;
        RECT 195.675 -2.885 196.005 -2.555 ;
        RECT 195.68 -3.56 196 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -91.285 196.005 -90.955 ;
        RECT 195.675 -92.645 196.005 -92.315 ;
        RECT 195.675 -94.005 196.005 -93.675 ;
        RECT 195.675 -95.365 196.005 -95.035 ;
        RECT 195.675 -96.725 196.005 -96.395 ;
        RECT 195.675 -98.085 196.005 -97.755 ;
        RECT 195.675 -99.445 196.005 -99.115 ;
        RECT 195.675 -100.805 196.005 -100.475 ;
        RECT 195.675 -102.165 196.005 -101.835 ;
        RECT 195.675 -103.525 196.005 -103.195 ;
        RECT 195.675 -104.885 196.005 -104.555 ;
        RECT 195.675 -106.245 196.005 -105.915 ;
        RECT 195.675 -107.605 196.005 -107.275 ;
        RECT 195.675 -108.965 196.005 -108.635 ;
        RECT 195.675 -110.325 196.005 -109.995 ;
        RECT 195.675 -111.685 196.005 -111.355 ;
        RECT 195.675 -113.045 196.005 -112.715 ;
        RECT 195.675 -114.405 196.005 -114.075 ;
        RECT 195.675 -115.765 196.005 -115.435 ;
        RECT 195.675 -117.125 196.005 -116.795 ;
        RECT 195.675 -118.485 196.005 -118.155 ;
        RECT 195.675 -119.845 196.005 -119.515 ;
        RECT 195.675 -121.205 196.005 -120.875 ;
        RECT 195.675 -122.565 196.005 -122.235 ;
        RECT 195.675 -123.925 196.005 -123.595 ;
        RECT 195.675 -125.285 196.005 -124.955 ;
        RECT 195.675 -126.645 196.005 -126.315 ;
        RECT 195.675 -128.005 196.005 -127.675 ;
        RECT 195.675 -129.365 196.005 -129.035 ;
        RECT 195.675 -130.725 196.005 -130.395 ;
        RECT 195.675 -132.085 196.005 -131.755 ;
        RECT 195.675 -133.445 196.005 -133.115 ;
        RECT 195.675 -134.805 196.005 -134.475 ;
        RECT 195.675 -136.165 196.005 -135.835 ;
        RECT 195.675 -137.525 196.005 -137.195 ;
        RECT 195.675 -138.885 196.005 -138.555 ;
        RECT 195.675 -140.245 196.005 -139.915 ;
        RECT 195.675 -141.605 196.005 -141.275 ;
        RECT 195.675 -142.965 196.005 -142.635 ;
        RECT 195.675 -144.325 196.005 -143.995 ;
        RECT 195.675 -145.685 196.005 -145.355 ;
        RECT 195.675 -147.045 196.005 -146.715 ;
        RECT 195.675 -148.405 196.005 -148.075 ;
        RECT 195.675 -149.765 196.005 -149.435 ;
        RECT 195.675 -151.125 196.005 -150.795 ;
        RECT 195.675 -152.485 196.005 -152.155 ;
        RECT 195.675 -153.845 196.005 -153.515 ;
        RECT 195.675 -155.205 196.005 -154.875 ;
        RECT 195.675 -156.565 196.005 -156.235 ;
        RECT 195.675 -157.925 196.005 -157.595 ;
        RECT 195.675 -160.17 196.005 -159.04 ;
        RECT 195.68 -160.285 196 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 127.225 197.365 128.355 ;
        RECT 197.035 124.955 197.365 125.285 ;
        RECT 197.035 123.595 197.365 123.925 ;
        RECT 197.04 123.595 197.36 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -1.525 197.365 -1.195 ;
        RECT 197.035 -2.885 197.365 -2.555 ;
        RECT 197.04 -3.56 197.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -140.245 197.365 -139.915 ;
        RECT 197.035 -141.605 197.365 -141.275 ;
        RECT 197.035 -142.965 197.365 -142.635 ;
        RECT 197.035 -144.325 197.365 -143.995 ;
        RECT 197.035 -145.685 197.365 -145.355 ;
        RECT 197.035 -147.045 197.365 -146.715 ;
        RECT 197.035 -148.405 197.365 -148.075 ;
        RECT 197.035 -149.765 197.365 -149.435 ;
        RECT 197.035 -151.125 197.365 -150.795 ;
        RECT 197.035 -152.485 197.365 -152.155 ;
        RECT 197.035 -153.845 197.365 -153.515 ;
        RECT 197.035 -155.205 197.365 -154.875 ;
        RECT 197.035 -156.565 197.365 -156.235 ;
        RECT 197.035 -157.925 197.365 -157.595 ;
        RECT 197.035 -160.17 197.365 -159.04 ;
        RECT 197.04 -160.285 197.36 -90.955 ;
        RECT 197.035 -91.285 197.365 -90.955 ;
        RECT 197.035 -92.645 197.365 -92.315 ;
        RECT 197.035 -94.005 197.365 -93.675 ;
        RECT 197.035 -95.365 197.365 -95.035 ;
        RECT 197.035 -96.725 197.365 -96.395 ;
        RECT 197.035 -98.085 197.365 -97.755 ;
        RECT 197.035 -99.445 197.365 -99.115 ;
        RECT 197.035 -100.805 197.365 -100.475 ;
        RECT 197.035 -102.165 197.365 -101.835 ;
        RECT 197.035 -103.525 197.365 -103.195 ;
        RECT 197.035 -104.885 197.365 -104.555 ;
        RECT 197.035 -106.245 197.365 -105.915 ;
        RECT 197.035 -107.605 197.365 -107.275 ;
        RECT 197.035 -108.965 197.365 -108.635 ;
        RECT 197.035 -110.325 197.365 -109.995 ;
        RECT 197.035 -111.685 197.365 -111.355 ;
        RECT 197.035 -113.045 197.365 -112.715 ;
        RECT 197.035 -114.405 197.365 -114.075 ;
        RECT 197.035 -115.765 197.365 -115.435 ;
        RECT 197.035 -117.125 197.365 -116.795 ;
        RECT 197.035 -118.485 197.365 -118.155 ;
        RECT 197.035 -119.845 197.365 -119.515 ;
        RECT 197.035 -121.205 197.365 -120.875 ;
        RECT 197.035 -122.565 197.365 -122.235 ;
        RECT 197.035 -123.925 197.365 -123.595 ;
        RECT 197.035 -125.285 197.365 -124.955 ;
        RECT 197.035 -126.645 197.365 -126.315 ;
        RECT 197.035 -128.005 197.365 -127.675 ;
        RECT 197.035 -129.365 197.365 -129.035 ;
        RECT 197.035 -130.725 197.365 -130.395 ;
        RECT 197.035 -132.085 197.365 -131.755 ;
        RECT 197.035 -133.445 197.365 -133.115 ;
        RECT 197.035 -134.805 197.365 -134.475 ;
        RECT 197.035 -136.165 197.365 -135.835 ;
        RECT 197.035 -137.525 197.365 -137.195 ;
        RECT 197.035 -138.885 197.365 -138.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.11 -94.075 113.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 127.225 114.405 128.355 ;
        RECT 114.075 124.955 114.405 125.285 ;
        RECT 114.075 123.595 114.405 123.925 ;
        RECT 114.08 123.595 114.4 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 -1.525 114.405 -1.195 ;
        RECT 114.075 -2.885 114.405 -2.555 ;
        RECT 114.08 -3.56 114.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 127.225 115.765 128.355 ;
        RECT 115.435 124.955 115.765 125.285 ;
        RECT 115.435 123.595 115.765 123.925 ;
        RECT 115.44 123.595 115.76 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 -1.525 115.765 -1.195 ;
        RECT 115.435 -2.885 115.765 -2.555 ;
        RECT 115.44 -3.56 115.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 127.225 117.125 128.355 ;
        RECT 116.795 124.955 117.125 125.285 ;
        RECT 116.795 123.595 117.125 123.925 ;
        RECT 116.8 123.595 117.12 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -1.525 117.125 -1.195 ;
        RECT 116.795 -2.885 117.125 -2.555 ;
        RECT 116.8 -3.56 117.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -91.285 117.125 -90.955 ;
        RECT 116.795 -92.645 117.125 -92.315 ;
        RECT 116.795 -94.005 117.125 -93.675 ;
        RECT 116.795 -95.365 117.125 -95.035 ;
        RECT 116.795 -96.725 117.125 -96.395 ;
        RECT 116.795 -98.085 117.125 -97.755 ;
        RECT 116.795 -99.445 117.125 -99.115 ;
        RECT 116.795 -100.805 117.125 -100.475 ;
        RECT 116.795 -102.165 117.125 -101.835 ;
        RECT 116.795 -103.525 117.125 -103.195 ;
        RECT 116.795 -104.885 117.125 -104.555 ;
        RECT 116.795 -106.245 117.125 -105.915 ;
        RECT 116.795 -107.605 117.125 -107.275 ;
        RECT 116.795 -108.965 117.125 -108.635 ;
        RECT 116.795 -110.325 117.125 -109.995 ;
        RECT 116.795 -111.685 117.125 -111.355 ;
        RECT 116.795 -113.045 117.125 -112.715 ;
        RECT 116.795 -114.405 117.125 -114.075 ;
        RECT 116.795 -115.765 117.125 -115.435 ;
        RECT 116.795 -117.125 117.125 -116.795 ;
        RECT 116.795 -118.485 117.125 -118.155 ;
        RECT 116.795 -119.845 117.125 -119.515 ;
        RECT 116.795 -121.205 117.125 -120.875 ;
        RECT 116.795 -122.565 117.125 -122.235 ;
        RECT 116.795 -123.925 117.125 -123.595 ;
        RECT 116.795 -125.285 117.125 -124.955 ;
        RECT 116.795 -126.645 117.125 -126.315 ;
        RECT 116.795 -128.005 117.125 -127.675 ;
        RECT 116.795 -129.365 117.125 -129.035 ;
        RECT 116.795 -130.725 117.125 -130.395 ;
        RECT 116.795 -132.085 117.125 -131.755 ;
        RECT 116.795 -133.445 117.125 -133.115 ;
        RECT 116.795 -134.805 117.125 -134.475 ;
        RECT 116.795 -136.165 117.125 -135.835 ;
        RECT 116.795 -137.525 117.125 -137.195 ;
        RECT 116.795 -138.885 117.125 -138.555 ;
        RECT 116.795 -140.245 117.125 -139.915 ;
        RECT 116.795 -141.605 117.125 -141.275 ;
        RECT 116.795 -142.965 117.125 -142.635 ;
        RECT 116.795 -144.325 117.125 -143.995 ;
        RECT 116.795 -145.685 117.125 -145.355 ;
        RECT 116.795 -147.045 117.125 -146.715 ;
        RECT 116.795 -148.405 117.125 -148.075 ;
        RECT 116.795 -149.765 117.125 -149.435 ;
        RECT 116.795 -151.125 117.125 -150.795 ;
        RECT 116.795 -152.485 117.125 -152.155 ;
        RECT 116.795 -153.845 117.125 -153.515 ;
        RECT 116.795 -155.205 117.125 -154.875 ;
        RECT 116.795 -156.565 117.125 -156.235 ;
        RECT 116.795 -157.925 117.125 -157.595 ;
        RECT 116.795 -160.17 117.125 -159.04 ;
        RECT 116.8 -160.285 117.12 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 127.225 118.485 128.355 ;
        RECT 118.155 124.955 118.485 125.285 ;
        RECT 118.155 123.595 118.485 123.925 ;
        RECT 118.16 123.595 118.48 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 -95.365 118.485 -95.035 ;
        RECT 118.155 -96.725 118.485 -96.395 ;
        RECT 118.155 -98.085 118.485 -97.755 ;
        RECT 118.155 -99.445 118.485 -99.115 ;
        RECT 118.155 -100.805 118.485 -100.475 ;
        RECT 118.155 -102.165 118.485 -101.835 ;
        RECT 118.155 -103.525 118.485 -103.195 ;
        RECT 118.155 -104.885 118.485 -104.555 ;
        RECT 118.155 -106.245 118.485 -105.915 ;
        RECT 118.155 -107.605 118.485 -107.275 ;
        RECT 118.155 -108.965 118.485 -108.635 ;
        RECT 118.155 -110.325 118.485 -109.995 ;
        RECT 118.155 -111.685 118.485 -111.355 ;
        RECT 118.155 -113.045 118.485 -112.715 ;
        RECT 118.155 -114.405 118.485 -114.075 ;
        RECT 118.155 -115.765 118.485 -115.435 ;
        RECT 118.155 -117.125 118.485 -116.795 ;
        RECT 118.155 -118.485 118.485 -118.155 ;
        RECT 118.155 -119.845 118.485 -119.515 ;
        RECT 118.155 -121.205 118.485 -120.875 ;
        RECT 118.155 -122.565 118.485 -122.235 ;
        RECT 118.155 -123.925 118.485 -123.595 ;
        RECT 118.155 -125.285 118.485 -124.955 ;
        RECT 118.155 -126.645 118.485 -126.315 ;
        RECT 118.155 -128.005 118.485 -127.675 ;
        RECT 118.155 -129.365 118.485 -129.035 ;
        RECT 118.155 -130.725 118.485 -130.395 ;
        RECT 118.155 -132.085 118.485 -131.755 ;
        RECT 118.155 -133.445 118.485 -133.115 ;
        RECT 118.155 -134.805 118.485 -134.475 ;
        RECT 118.155 -136.165 118.485 -135.835 ;
        RECT 118.155 -137.525 118.485 -137.195 ;
        RECT 118.155 -138.885 118.485 -138.555 ;
        RECT 118.155 -140.245 118.485 -139.915 ;
        RECT 118.155 -141.605 118.485 -141.275 ;
        RECT 118.155 -142.965 118.485 -142.635 ;
        RECT 118.155 -144.325 118.485 -143.995 ;
        RECT 118.155 -145.685 118.485 -145.355 ;
        RECT 118.155 -147.045 118.485 -146.715 ;
        RECT 118.155 -148.405 118.485 -148.075 ;
        RECT 118.155 -149.765 118.485 -149.435 ;
        RECT 118.155 -151.125 118.485 -150.795 ;
        RECT 118.155 -152.485 118.485 -152.155 ;
        RECT 118.155 -153.845 118.485 -153.515 ;
        RECT 118.155 -155.205 118.485 -154.875 ;
        RECT 118.155 -156.565 118.485 -156.235 ;
        RECT 118.155 -157.925 118.485 -157.595 ;
        RECT 118.155 -160.17 118.485 -159.04 ;
        RECT 118.16 -160.285 118.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.21 -94.075 119.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 127.225 119.845 128.355 ;
        RECT 119.515 124.955 119.845 125.285 ;
        RECT 119.515 123.595 119.845 123.925 ;
        RECT 119.52 123.595 119.84 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 127.225 121.205 128.355 ;
        RECT 120.875 124.955 121.205 125.285 ;
        RECT 120.875 123.595 121.205 123.925 ;
        RECT 120.88 123.595 121.2 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 -1.525 121.205 -1.195 ;
        RECT 120.875 -2.885 121.205 -2.555 ;
        RECT 120.88 -3.56 121.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 127.225 122.565 128.355 ;
        RECT 122.235 124.955 122.565 125.285 ;
        RECT 122.235 123.595 122.565 123.925 ;
        RECT 122.24 123.595 122.56 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 -1.525 122.565 -1.195 ;
        RECT 122.235 -2.885 122.565 -2.555 ;
        RECT 122.24 -3.56 122.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 127.225 123.925 128.355 ;
        RECT 123.595 124.955 123.925 125.285 ;
        RECT 123.595 123.595 123.925 123.925 ;
        RECT 123.6 123.595 123.92 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 -1.525 123.925 -1.195 ;
        RECT 123.595 -2.885 123.925 -2.555 ;
        RECT 123.6 -3.56 123.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 -91.285 123.925 -90.955 ;
        RECT 123.595 -92.645 123.925 -92.315 ;
        RECT 123.595 -94.005 123.925 -93.675 ;
        RECT 123.595 -95.365 123.925 -95.035 ;
        RECT 123.595 -96.725 123.925 -96.395 ;
        RECT 123.595 -98.085 123.925 -97.755 ;
        RECT 123.595 -99.445 123.925 -99.115 ;
        RECT 123.595 -100.805 123.925 -100.475 ;
        RECT 123.595 -102.165 123.925 -101.835 ;
        RECT 123.595 -103.525 123.925 -103.195 ;
        RECT 123.595 -104.885 123.925 -104.555 ;
        RECT 123.595 -106.245 123.925 -105.915 ;
        RECT 123.595 -107.605 123.925 -107.275 ;
        RECT 123.595 -108.965 123.925 -108.635 ;
        RECT 123.595 -110.325 123.925 -109.995 ;
        RECT 123.595 -111.685 123.925 -111.355 ;
        RECT 123.595 -113.045 123.925 -112.715 ;
        RECT 123.595 -114.405 123.925 -114.075 ;
        RECT 123.595 -115.765 123.925 -115.435 ;
        RECT 123.595 -117.125 123.925 -116.795 ;
        RECT 123.595 -118.485 123.925 -118.155 ;
        RECT 123.595 -119.845 123.925 -119.515 ;
        RECT 123.595 -121.205 123.925 -120.875 ;
        RECT 123.595 -122.565 123.925 -122.235 ;
        RECT 123.595 -123.925 123.925 -123.595 ;
        RECT 123.595 -125.285 123.925 -124.955 ;
        RECT 123.595 -126.645 123.925 -126.315 ;
        RECT 123.595 -128.005 123.925 -127.675 ;
        RECT 123.595 -129.365 123.925 -129.035 ;
        RECT 123.595 -130.725 123.925 -130.395 ;
        RECT 123.595 -132.085 123.925 -131.755 ;
        RECT 123.595 -133.445 123.925 -133.115 ;
        RECT 123.595 -134.805 123.925 -134.475 ;
        RECT 123.595 -136.165 123.925 -135.835 ;
        RECT 123.595 -137.525 123.925 -137.195 ;
        RECT 123.595 -138.885 123.925 -138.555 ;
        RECT 123.595 -140.245 123.925 -139.915 ;
        RECT 123.595 -141.605 123.925 -141.275 ;
        RECT 123.595 -142.965 123.925 -142.635 ;
        RECT 123.595 -144.325 123.925 -143.995 ;
        RECT 123.595 -145.685 123.925 -145.355 ;
        RECT 123.595 -147.045 123.925 -146.715 ;
        RECT 123.595 -148.405 123.925 -148.075 ;
        RECT 123.595 -149.765 123.925 -149.435 ;
        RECT 123.595 -151.125 123.925 -150.795 ;
        RECT 123.595 -152.485 123.925 -152.155 ;
        RECT 123.595 -153.845 123.925 -153.515 ;
        RECT 123.595 -155.205 123.925 -154.875 ;
        RECT 123.595 -156.565 123.925 -156.235 ;
        RECT 123.595 -157.925 123.925 -157.595 ;
        RECT 123.595 -160.17 123.925 -159.04 ;
        RECT 123.6 -160.285 123.92 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 127.225 125.285 128.355 ;
        RECT 124.955 124.955 125.285 125.285 ;
        RECT 124.955 123.595 125.285 123.925 ;
        RECT 124.96 123.595 125.28 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 -95.365 125.285 -95.035 ;
        RECT 124.955 -96.725 125.285 -96.395 ;
        RECT 124.955 -98.085 125.285 -97.755 ;
        RECT 124.955 -99.445 125.285 -99.115 ;
        RECT 124.955 -100.805 125.285 -100.475 ;
        RECT 124.955 -102.165 125.285 -101.835 ;
        RECT 124.955 -103.525 125.285 -103.195 ;
        RECT 124.955 -104.885 125.285 -104.555 ;
        RECT 124.955 -106.245 125.285 -105.915 ;
        RECT 124.955 -107.605 125.285 -107.275 ;
        RECT 124.955 -108.965 125.285 -108.635 ;
        RECT 124.955 -110.325 125.285 -109.995 ;
        RECT 124.955 -111.685 125.285 -111.355 ;
        RECT 124.955 -113.045 125.285 -112.715 ;
        RECT 124.955 -114.405 125.285 -114.075 ;
        RECT 124.955 -115.765 125.285 -115.435 ;
        RECT 124.955 -117.125 125.285 -116.795 ;
        RECT 124.955 -118.485 125.285 -118.155 ;
        RECT 124.955 -119.845 125.285 -119.515 ;
        RECT 124.955 -121.205 125.285 -120.875 ;
        RECT 124.955 -122.565 125.285 -122.235 ;
        RECT 124.955 -123.925 125.285 -123.595 ;
        RECT 124.955 -125.285 125.285 -124.955 ;
        RECT 124.955 -126.645 125.285 -126.315 ;
        RECT 124.955 -128.005 125.285 -127.675 ;
        RECT 124.955 -129.365 125.285 -129.035 ;
        RECT 124.955 -130.725 125.285 -130.395 ;
        RECT 124.955 -132.085 125.285 -131.755 ;
        RECT 124.955 -133.445 125.285 -133.115 ;
        RECT 124.955 -134.805 125.285 -134.475 ;
        RECT 124.955 -136.165 125.285 -135.835 ;
        RECT 124.955 -137.525 125.285 -137.195 ;
        RECT 124.955 -138.885 125.285 -138.555 ;
        RECT 124.955 -140.245 125.285 -139.915 ;
        RECT 124.955 -141.605 125.285 -141.275 ;
        RECT 124.955 -142.965 125.285 -142.635 ;
        RECT 124.955 -144.325 125.285 -143.995 ;
        RECT 124.955 -145.685 125.285 -145.355 ;
        RECT 124.955 -147.045 125.285 -146.715 ;
        RECT 124.955 -148.405 125.285 -148.075 ;
        RECT 124.955 -149.765 125.285 -149.435 ;
        RECT 124.955 -151.125 125.285 -150.795 ;
        RECT 124.955 -152.485 125.285 -152.155 ;
        RECT 124.955 -153.845 125.285 -153.515 ;
        RECT 124.955 -155.205 125.285 -154.875 ;
        RECT 124.955 -156.565 125.285 -156.235 ;
        RECT 124.955 -157.925 125.285 -157.595 ;
        RECT 124.955 -160.17 125.285 -159.04 ;
        RECT 124.96 -160.285 125.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.31 -94.075 125.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 127.225 126.645 128.355 ;
        RECT 126.315 124.955 126.645 125.285 ;
        RECT 126.315 123.595 126.645 123.925 ;
        RECT 126.32 123.595 126.64 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 -1.525 126.645 -1.195 ;
        RECT 126.315 -2.885 126.645 -2.555 ;
        RECT 126.32 -3.56 126.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 127.225 128.005 128.355 ;
        RECT 127.675 124.955 128.005 125.285 ;
        RECT 127.675 123.595 128.005 123.925 ;
        RECT 127.68 123.595 128 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 -1.525 128.005 -1.195 ;
        RECT 127.675 -2.885 128.005 -2.555 ;
        RECT 127.68 -3.56 128 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 127.225 129.365 128.355 ;
        RECT 129.035 124.955 129.365 125.285 ;
        RECT 129.035 123.595 129.365 123.925 ;
        RECT 129.04 123.595 129.36 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -1.525 129.365 -1.195 ;
        RECT 129.035 -2.885 129.365 -2.555 ;
        RECT 129.04 -3.56 129.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -91.285 129.365 -90.955 ;
        RECT 129.035 -92.645 129.365 -92.315 ;
        RECT 129.035 -94.005 129.365 -93.675 ;
        RECT 129.035 -95.365 129.365 -95.035 ;
        RECT 129.035 -96.725 129.365 -96.395 ;
        RECT 129.035 -98.085 129.365 -97.755 ;
        RECT 129.035 -99.445 129.365 -99.115 ;
        RECT 129.035 -100.805 129.365 -100.475 ;
        RECT 129.035 -102.165 129.365 -101.835 ;
        RECT 129.035 -103.525 129.365 -103.195 ;
        RECT 129.035 -104.885 129.365 -104.555 ;
        RECT 129.035 -106.245 129.365 -105.915 ;
        RECT 129.035 -107.605 129.365 -107.275 ;
        RECT 129.035 -108.965 129.365 -108.635 ;
        RECT 129.035 -110.325 129.365 -109.995 ;
        RECT 129.035 -111.685 129.365 -111.355 ;
        RECT 129.035 -113.045 129.365 -112.715 ;
        RECT 129.035 -114.405 129.365 -114.075 ;
        RECT 129.035 -115.765 129.365 -115.435 ;
        RECT 129.035 -117.125 129.365 -116.795 ;
        RECT 129.035 -118.485 129.365 -118.155 ;
        RECT 129.035 -119.845 129.365 -119.515 ;
        RECT 129.035 -121.205 129.365 -120.875 ;
        RECT 129.035 -122.565 129.365 -122.235 ;
        RECT 129.035 -123.925 129.365 -123.595 ;
        RECT 129.035 -125.285 129.365 -124.955 ;
        RECT 129.035 -126.645 129.365 -126.315 ;
        RECT 129.035 -128.005 129.365 -127.675 ;
        RECT 129.035 -129.365 129.365 -129.035 ;
        RECT 129.035 -130.725 129.365 -130.395 ;
        RECT 129.035 -132.085 129.365 -131.755 ;
        RECT 129.035 -133.445 129.365 -133.115 ;
        RECT 129.035 -134.805 129.365 -134.475 ;
        RECT 129.035 -136.165 129.365 -135.835 ;
        RECT 129.035 -137.525 129.365 -137.195 ;
        RECT 129.035 -138.885 129.365 -138.555 ;
        RECT 129.035 -140.245 129.365 -139.915 ;
        RECT 129.035 -141.605 129.365 -141.275 ;
        RECT 129.035 -142.965 129.365 -142.635 ;
        RECT 129.035 -144.325 129.365 -143.995 ;
        RECT 129.035 -145.685 129.365 -145.355 ;
        RECT 129.035 -147.045 129.365 -146.715 ;
        RECT 129.035 -148.405 129.365 -148.075 ;
        RECT 129.035 -149.765 129.365 -149.435 ;
        RECT 129.035 -151.125 129.365 -150.795 ;
        RECT 129.035 -152.485 129.365 -152.155 ;
        RECT 129.035 -153.845 129.365 -153.515 ;
        RECT 129.035 -155.205 129.365 -154.875 ;
        RECT 129.035 -156.565 129.365 -156.235 ;
        RECT 129.035 -157.925 129.365 -157.595 ;
        RECT 129.035 -160.17 129.365 -159.04 ;
        RECT 129.04 -160.285 129.36 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 127.225 130.725 128.355 ;
        RECT 130.395 124.955 130.725 125.285 ;
        RECT 130.395 123.595 130.725 123.925 ;
        RECT 130.4 123.595 130.72 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 -95.365 130.725 -95.035 ;
        RECT 130.395 -96.725 130.725 -96.395 ;
        RECT 130.395 -98.085 130.725 -97.755 ;
        RECT 130.395 -99.445 130.725 -99.115 ;
        RECT 130.395 -100.805 130.725 -100.475 ;
        RECT 130.395 -102.165 130.725 -101.835 ;
        RECT 130.395 -103.525 130.725 -103.195 ;
        RECT 130.395 -104.885 130.725 -104.555 ;
        RECT 130.395 -106.245 130.725 -105.915 ;
        RECT 130.395 -107.605 130.725 -107.275 ;
        RECT 130.395 -108.965 130.725 -108.635 ;
        RECT 130.395 -110.325 130.725 -109.995 ;
        RECT 130.395 -111.685 130.725 -111.355 ;
        RECT 130.395 -113.045 130.725 -112.715 ;
        RECT 130.395 -114.405 130.725 -114.075 ;
        RECT 130.395 -115.765 130.725 -115.435 ;
        RECT 130.395 -117.125 130.725 -116.795 ;
        RECT 130.395 -118.485 130.725 -118.155 ;
        RECT 130.395 -119.845 130.725 -119.515 ;
        RECT 130.395 -121.205 130.725 -120.875 ;
        RECT 130.395 -122.565 130.725 -122.235 ;
        RECT 130.395 -123.925 130.725 -123.595 ;
        RECT 130.395 -125.285 130.725 -124.955 ;
        RECT 130.395 -126.645 130.725 -126.315 ;
        RECT 130.395 -128.005 130.725 -127.675 ;
        RECT 130.395 -129.365 130.725 -129.035 ;
        RECT 130.395 -130.725 130.725 -130.395 ;
        RECT 130.395 -132.085 130.725 -131.755 ;
        RECT 130.395 -133.445 130.725 -133.115 ;
        RECT 130.395 -134.805 130.725 -134.475 ;
        RECT 130.395 -136.165 130.725 -135.835 ;
        RECT 130.395 -137.525 130.725 -137.195 ;
        RECT 130.395 -138.885 130.725 -138.555 ;
        RECT 130.395 -140.245 130.725 -139.915 ;
        RECT 130.395 -141.605 130.725 -141.275 ;
        RECT 130.395 -142.965 130.725 -142.635 ;
        RECT 130.395 -144.325 130.725 -143.995 ;
        RECT 130.395 -145.685 130.725 -145.355 ;
        RECT 130.395 -147.045 130.725 -146.715 ;
        RECT 130.395 -148.405 130.725 -148.075 ;
        RECT 130.395 -149.765 130.725 -149.435 ;
        RECT 130.395 -151.125 130.725 -150.795 ;
        RECT 130.395 -152.485 130.725 -152.155 ;
        RECT 130.395 -153.845 130.725 -153.515 ;
        RECT 130.395 -155.205 130.725 -154.875 ;
        RECT 130.395 -156.565 130.725 -156.235 ;
        RECT 130.395 -157.925 130.725 -157.595 ;
        RECT 130.395 -160.17 130.725 -159.04 ;
        RECT 130.4 -160.285 130.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.41 -94.075 131.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 127.225 132.085 128.355 ;
        RECT 131.755 124.955 132.085 125.285 ;
        RECT 131.755 123.595 132.085 123.925 ;
        RECT 131.76 123.595 132.08 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 127.225 133.445 128.355 ;
        RECT 133.115 124.955 133.445 125.285 ;
        RECT 133.115 123.595 133.445 123.925 ;
        RECT 133.12 123.595 133.44 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 -1.525 133.445 -1.195 ;
        RECT 133.115 -2.885 133.445 -2.555 ;
        RECT 133.12 -3.56 133.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 127.225 134.805 128.355 ;
        RECT 134.475 124.955 134.805 125.285 ;
        RECT 134.475 123.595 134.805 123.925 ;
        RECT 134.48 123.595 134.8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 -1.525 134.805 -1.195 ;
        RECT 134.475 -2.885 134.805 -2.555 ;
        RECT 134.48 -3.56 134.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 -91.285 134.805 -90.955 ;
        RECT 134.475 -92.645 134.805 -92.315 ;
        RECT 134.475 -94.005 134.805 -93.675 ;
        RECT 134.475 -95.365 134.805 -95.035 ;
        RECT 134.475 -96.725 134.805 -96.395 ;
        RECT 134.475 -98.085 134.805 -97.755 ;
        RECT 134.475 -99.445 134.805 -99.115 ;
        RECT 134.475 -100.805 134.805 -100.475 ;
        RECT 134.475 -102.165 134.805 -101.835 ;
        RECT 134.475 -103.525 134.805 -103.195 ;
        RECT 134.475 -104.885 134.805 -104.555 ;
        RECT 134.475 -106.245 134.805 -105.915 ;
        RECT 134.475 -107.605 134.805 -107.275 ;
        RECT 134.475 -108.965 134.805 -108.635 ;
        RECT 134.475 -110.325 134.805 -109.995 ;
        RECT 134.475 -111.685 134.805 -111.355 ;
        RECT 134.475 -113.045 134.805 -112.715 ;
        RECT 134.475 -114.405 134.805 -114.075 ;
        RECT 134.475 -115.765 134.805 -115.435 ;
        RECT 134.475 -117.125 134.805 -116.795 ;
        RECT 134.475 -118.485 134.805 -118.155 ;
        RECT 134.475 -119.845 134.805 -119.515 ;
        RECT 134.475 -121.205 134.805 -120.875 ;
        RECT 134.475 -122.565 134.805 -122.235 ;
        RECT 134.475 -123.925 134.805 -123.595 ;
        RECT 134.475 -125.285 134.805 -124.955 ;
        RECT 134.475 -126.645 134.805 -126.315 ;
        RECT 134.475 -128.005 134.805 -127.675 ;
        RECT 134.475 -129.365 134.805 -129.035 ;
        RECT 134.475 -130.725 134.805 -130.395 ;
        RECT 134.475 -132.085 134.805 -131.755 ;
        RECT 134.475 -133.445 134.805 -133.115 ;
        RECT 134.475 -134.805 134.805 -134.475 ;
        RECT 134.475 -136.165 134.805 -135.835 ;
        RECT 134.475 -137.525 134.805 -137.195 ;
        RECT 134.475 -138.885 134.805 -138.555 ;
        RECT 134.475 -140.245 134.805 -139.915 ;
        RECT 134.475 -141.605 134.805 -141.275 ;
        RECT 134.475 -142.965 134.805 -142.635 ;
        RECT 134.475 -144.325 134.805 -143.995 ;
        RECT 134.475 -145.685 134.805 -145.355 ;
        RECT 134.475 -147.045 134.805 -146.715 ;
        RECT 134.475 -148.405 134.805 -148.075 ;
        RECT 134.475 -149.765 134.805 -149.435 ;
        RECT 134.475 -151.125 134.805 -150.795 ;
        RECT 134.475 -152.485 134.805 -152.155 ;
        RECT 134.475 -153.845 134.805 -153.515 ;
        RECT 134.475 -155.205 134.805 -154.875 ;
        RECT 134.475 -156.565 134.805 -156.235 ;
        RECT 134.475 -157.925 134.805 -157.595 ;
        RECT 134.475 -160.17 134.805 -159.04 ;
        RECT 134.48 -160.285 134.8 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 127.225 136.165 128.355 ;
        RECT 135.835 124.955 136.165 125.285 ;
        RECT 135.835 123.595 136.165 123.925 ;
        RECT 135.84 123.595 136.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 -1.525 136.165 -1.195 ;
        RECT 135.835 -2.885 136.165 -2.555 ;
        RECT 135.84 -3.56 136.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 -91.285 136.165 -90.955 ;
        RECT 135.835 -92.645 136.165 -92.315 ;
        RECT 135.835 -94.005 136.165 -93.675 ;
        RECT 135.835 -95.365 136.165 -95.035 ;
        RECT 135.835 -96.725 136.165 -96.395 ;
        RECT 135.835 -98.085 136.165 -97.755 ;
        RECT 135.835 -99.445 136.165 -99.115 ;
        RECT 135.835 -100.805 136.165 -100.475 ;
        RECT 135.835 -102.165 136.165 -101.835 ;
        RECT 135.835 -103.525 136.165 -103.195 ;
        RECT 135.835 -104.885 136.165 -104.555 ;
        RECT 135.835 -106.245 136.165 -105.915 ;
        RECT 135.835 -107.605 136.165 -107.275 ;
        RECT 135.835 -108.965 136.165 -108.635 ;
        RECT 135.835 -110.325 136.165 -109.995 ;
        RECT 135.835 -111.685 136.165 -111.355 ;
        RECT 135.835 -113.045 136.165 -112.715 ;
        RECT 135.835 -114.405 136.165 -114.075 ;
        RECT 135.835 -115.765 136.165 -115.435 ;
        RECT 135.835 -117.125 136.165 -116.795 ;
        RECT 135.835 -118.485 136.165 -118.155 ;
        RECT 135.835 -119.845 136.165 -119.515 ;
        RECT 135.835 -121.205 136.165 -120.875 ;
        RECT 135.835 -122.565 136.165 -122.235 ;
        RECT 135.835 -123.925 136.165 -123.595 ;
        RECT 135.835 -125.285 136.165 -124.955 ;
        RECT 135.835 -126.645 136.165 -126.315 ;
        RECT 135.835 -128.005 136.165 -127.675 ;
        RECT 135.835 -129.365 136.165 -129.035 ;
        RECT 135.835 -130.725 136.165 -130.395 ;
        RECT 135.835 -132.085 136.165 -131.755 ;
        RECT 135.835 -133.445 136.165 -133.115 ;
        RECT 135.835 -134.805 136.165 -134.475 ;
        RECT 135.835 -136.165 136.165 -135.835 ;
        RECT 135.835 -137.525 136.165 -137.195 ;
        RECT 135.835 -138.885 136.165 -138.555 ;
        RECT 135.835 -140.245 136.165 -139.915 ;
        RECT 135.835 -141.605 136.165 -141.275 ;
        RECT 135.835 -142.965 136.165 -142.635 ;
        RECT 135.835 -144.325 136.165 -143.995 ;
        RECT 135.835 -145.685 136.165 -145.355 ;
        RECT 135.835 -147.045 136.165 -146.715 ;
        RECT 135.835 -148.405 136.165 -148.075 ;
        RECT 135.835 -149.765 136.165 -149.435 ;
        RECT 135.835 -151.125 136.165 -150.795 ;
        RECT 135.835 -152.485 136.165 -152.155 ;
        RECT 135.835 -153.845 136.165 -153.515 ;
        RECT 135.835 -155.205 136.165 -154.875 ;
        RECT 135.835 -156.565 136.165 -156.235 ;
        RECT 135.835 -157.925 136.165 -157.595 ;
        RECT 135.835 -160.17 136.165 -159.04 ;
        RECT 135.84 -160.285 136.16 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 127.225 137.525 128.355 ;
        RECT 137.195 124.955 137.525 125.285 ;
        RECT 137.195 123.595 137.525 123.925 ;
        RECT 137.2 123.595 137.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 -95.365 137.525 -95.035 ;
        RECT 137.195 -96.725 137.525 -96.395 ;
        RECT 137.195 -98.085 137.525 -97.755 ;
        RECT 137.195 -99.445 137.525 -99.115 ;
        RECT 137.195 -100.805 137.525 -100.475 ;
        RECT 137.195 -102.165 137.525 -101.835 ;
        RECT 137.195 -103.525 137.525 -103.195 ;
        RECT 137.195 -104.885 137.525 -104.555 ;
        RECT 137.195 -106.245 137.525 -105.915 ;
        RECT 137.195 -107.605 137.525 -107.275 ;
        RECT 137.195 -108.965 137.525 -108.635 ;
        RECT 137.195 -110.325 137.525 -109.995 ;
        RECT 137.195 -111.685 137.525 -111.355 ;
        RECT 137.195 -113.045 137.525 -112.715 ;
        RECT 137.195 -114.405 137.525 -114.075 ;
        RECT 137.195 -115.765 137.525 -115.435 ;
        RECT 137.195 -117.125 137.525 -116.795 ;
        RECT 137.195 -118.485 137.525 -118.155 ;
        RECT 137.195 -119.845 137.525 -119.515 ;
        RECT 137.195 -121.205 137.525 -120.875 ;
        RECT 137.195 -122.565 137.525 -122.235 ;
        RECT 137.195 -123.925 137.525 -123.595 ;
        RECT 137.195 -125.285 137.525 -124.955 ;
        RECT 137.195 -126.645 137.525 -126.315 ;
        RECT 137.195 -128.005 137.525 -127.675 ;
        RECT 137.195 -129.365 137.525 -129.035 ;
        RECT 137.195 -130.725 137.525 -130.395 ;
        RECT 137.195 -132.085 137.525 -131.755 ;
        RECT 137.195 -133.445 137.525 -133.115 ;
        RECT 137.195 -134.805 137.525 -134.475 ;
        RECT 137.195 -136.165 137.525 -135.835 ;
        RECT 137.195 -137.525 137.525 -137.195 ;
        RECT 137.195 -138.885 137.525 -138.555 ;
        RECT 137.195 -140.245 137.525 -139.915 ;
        RECT 137.195 -141.605 137.525 -141.275 ;
        RECT 137.195 -142.965 137.525 -142.635 ;
        RECT 137.195 -144.325 137.525 -143.995 ;
        RECT 137.195 -145.685 137.525 -145.355 ;
        RECT 137.195 -147.045 137.525 -146.715 ;
        RECT 137.195 -148.405 137.525 -148.075 ;
        RECT 137.195 -149.765 137.525 -149.435 ;
        RECT 137.195 -151.125 137.525 -150.795 ;
        RECT 137.195 -152.485 137.525 -152.155 ;
        RECT 137.195 -153.845 137.525 -153.515 ;
        RECT 137.195 -155.205 137.525 -154.875 ;
        RECT 137.195 -156.565 137.525 -156.235 ;
        RECT 137.195 -157.925 137.525 -157.595 ;
        RECT 137.195 -160.17 137.525 -159.04 ;
        RECT 137.2 -160.285 137.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.51 -94.075 137.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 127.225 138.885 128.355 ;
        RECT 138.555 124.955 138.885 125.285 ;
        RECT 138.555 123.595 138.885 123.925 ;
        RECT 138.56 123.595 138.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 -1.525 138.885 -1.195 ;
        RECT 138.555 -2.885 138.885 -2.555 ;
        RECT 138.56 -3.56 138.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 127.225 140.245 128.355 ;
        RECT 139.915 124.955 140.245 125.285 ;
        RECT 139.915 123.595 140.245 123.925 ;
        RECT 139.92 123.595 140.24 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 -1.525 140.245 -1.195 ;
        RECT 139.915 -2.885 140.245 -2.555 ;
        RECT 139.92 -3.56 140.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 127.225 141.605 128.355 ;
        RECT 141.275 124.955 141.605 125.285 ;
        RECT 141.275 123.595 141.605 123.925 ;
        RECT 141.28 123.595 141.6 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -1.525 141.605 -1.195 ;
        RECT 141.275 -2.885 141.605 -2.555 ;
        RECT 141.28 -3.56 141.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -91.285 141.605 -90.955 ;
        RECT 141.275 -92.645 141.605 -92.315 ;
        RECT 141.275 -94.005 141.605 -93.675 ;
        RECT 141.275 -95.365 141.605 -95.035 ;
        RECT 141.275 -96.725 141.605 -96.395 ;
        RECT 141.275 -98.085 141.605 -97.755 ;
        RECT 141.275 -99.445 141.605 -99.115 ;
        RECT 141.275 -100.805 141.605 -100.475 ;
        RECT 141.275 -102.165 141.605 -101.835 ;
        RECT 141.275 -103.525 141.605 -103.195 ;
        RECT 141.275 -104.885 141.605 -104.555 ;
        RECT 141.275 -106.245 141.605 -105.915 ;
        RECT 141.275 -107.605 141.605 -107.275 ;
        RECT 141.275 -108.965 141.605 -108.635 ;
        RECT 141.275 -110.325 141.605 -109.995 ;
        RECT 141.275 -111.685 141.605 -111.355 ;
        RECT 141.275 -113.045 141.605 -112.715 ;
        RECT 141.275 -114.405 141.605 -114.075 ;
        RECT 141.275 -115.765 141.605 -115.435 ;
        RECT 141.275 -117.125 141.605 -116.795 ;
        RECT 141.275 -118.485 141.605 -118.155 ;
        RECT 141.275 -119.845 141.605 -119.515 ;
        RECT 141.275 -121.205 141.605 -120.875 ;
        RECT 141.275 -122.565 141.605 -122.235 ;
        RECT 141.275 -123.925 141.605 -123.595 ;
        RECT 141.275 -125.285 141.605 -124.955 ;
        RECT 141.275 -126.645 141.605 -126.315 ;
        RECT 141.275 -128.005 141.605 -127.675 ;
        RECT 141.275 -129.365 141.605 -129.035 ;
        RECT 141.275 -130.725 141.605 -130.395 ;
        RECT 141.275 -132.085 141.605 -131.755 ;
        RECT 141.275 -133.445 141.605 -133.115 ;
        RECT 141.275 -134.805 141.605 -134.475 ;
        RECT 141.275 -136.165 141.605 -135.835 ;
        RECT 141.275 -137.525 141.605 -137.195 ;
        RECT 141.275 -138.885 141.605 -138.555 ;
        RECT 141.275 -140.245 141.605 -139.915 ;
        RECT 141.275 -141.605 141.605 -141.275 ;
        RECT 141.275 -142.965 141.605 -142.635 ;
        RECT 141.275 -144.325 141.605 -143.995 ;
        RECT 141.275 -145.685 141.605 -145.355 ;
        RECT 141.275 -147.045 141.605 -146.715 ;
        RECT 141.275 -148.405 141.605 -148.075 ;
        RECT 141.275 -149.765 141.605 -149.435 ;
        RECT 141.275 -151.125 141.605 -150.795 ;
        RECT 141.275 -152.485 141.605 -152.155 ;
        RECT 141.275 -153.845 141.605 -153.515 ;
        RECT 141.275 -155.205 141.605 -154.875 ;
        RECT 141.275 -156.565 141.605 -156.235 ;
        RECT 141.275 -157.925 141.605 -157.595 ;
        RECT 141.275 -160.17 141.605 -159.04 ;
        RECT 141.28 -160.285 141.6 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 127.225 142.965 128.355 ;
        RECT 142.635 124.955 142.965 125.285 ;
        RECT 142.635 123.595 142.965 123.925 ;
        RECT 142.64 123.595 142.96 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 -95.365 142.965 -95.035 ;
        RECT 142.635 -96.725 142.965 -96.395 ;
        RECT 142.635 -98.085 142.965 -97.755 ;
        RECT 142.635 -99.445 142.965 -99.115 ;
        RECT 142.635 -100.805 142.965 -100.475 ;
        RECT 142.635 -102.165 142.965 -101.835 ;
        RECT 142.635 -103.525 142.965 -103.195 ;
        RECT 142.635 -104.885 142.965 -104.555 ;
        RECT 142.635 -106.245 142.965 -105.915 ;
        RECT 142.635 -107.605 142.965 -107.275 ;
        RECT 142.635 -108.965 142.965 -108.635 ;
        RECT 142.635 -110.325 142.965 -109.995 ;
        RECT 142.635 -111.685 142.965 -111.355 ;
        RECT 142.635 -113.045 142.965 -112.715 ;
        RECT 142.635 -114.405 142.965 -114.075 ;
        RECT 142.635 -115.765 142.965 -115.435 ;
        RECT 142.635 -117.125 142.965 -116.795 ;
        RECT 142.635 -118.485 142.965 -118.155 ;
        RECT 142.635 -119.845 142.965 -119.515 ;
        RECT 142.635 -121.205 142.965 -120.875 ;
        RECT 142.635 -122.565 142.965 -122.235 ;
        RECT 142.635 -123.925 142.965 -123.595 ;
        RECT 142.635 -125.285 142.965 -124.955 ;
        RECT 142.635 -126.645 142.965 -126.315 ;
        RECT 142.635 -128.005 142.965 -127.675 ;
        RECT 142.635 -129.365 142.965 -129.035 ;
        RECT 142.635 -130.725 142.965 -130.395 ;
        RECT 142.635 -132.085 142.965 -131.755 ;
        RECT 142.635 -133.445 142.965 -133.115 ;
        RECT 142.635 -134.805 142.965 -134.475 ;
        RECT 142.635 -136.165 142.965 -135.835 ;
        RECT 142.635 -137.525 142.965 -137.195 ;
        RECT 142.635 -138.885 142.965 -138.555 ;
        RECT 142.635 -140.245 142.965 -139.915 ;
        RECT 142.635 -141.605 142.965 -141.275 ;
        RECT 142.635 -142.965 142.965 -142.635 ;
        RECT 142.635 -144.325 142.965 -143.995 ;
        RECT 142.635 -145.685 142.965 -145.355 ;
        RECT 142.635 -147.045 142.965 -146.715 ;
        RECT 142.635 -148.405 142.965 -148.075 ;
        RECT 142.635 -149.765 142.965 -149.435 ;
        RECT 142.635 -151.125 142.965 -150.795 ;
        RECT 142.635 -152.485 142.965 -152.155 ;
        RECT 142.635 -153.845 142.965 -153.515 ;
        RECT 142.635 -155.205 142.965 -154.875 ;
        RECT 142.635 -156.565 142.965 -156.235 ;
        RECT 142.635 -157.925 142.965 -157.595 ;
        RECT 142.635 -160.17 142.965 -159.04 ;
        RECT 142.64 -160.285 142.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.61 -94.075 143.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 127.225 144.325 128.355 ;
        RECT 143.995 124.955 144.325 125.285 ;
        RECT 143.995 123.595 144.325 123.925 ;
        RECT 144 123.595 144.32 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 127.225 145.685 128.355 ;
        RECT 145.355 124.955 145.685 125.285 ;
        RECT 145.355 123.595 145.685 123.925 ;
        RECT 145.36 123.595 145.68 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 -1.525 145.685 -1.195 ;
        RECT 145.355 -2.885 145.685 -2.555 ;
        RECT 145.36 -3.56 145.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 127.225 147.045 128.355 ;
        RECT 146.715 124.955 147.045 125.285 ;
        RECT 146.715 123.595 147.045 123.925 ;
        RECT 146.72 123.595 147.04 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 -1.525 147.045 -1.195 ;
        RECT 146.715 -2.885 147.045 -2.555 ;
        RECT 146.72 -3.56 147.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 -91.285 147.045 -90.955 ;
        RECT 146.715 -92.645 147.045 -92.315 ;
        RECT 146.715 -94.005 147.045 -93.675 ;
        RECT 146.715 -95.365 147.045 -95.035 ;
        RECT 146.715 -96.725 147.045 -96.395 ;
        RECT 146.715 -98.085 147.045 -97.755 ;
        RECT 146.715 -99.445 147.045 -99.115 ;
        RECT 146.715 -100.805 147.045 -100.475 ;
        RECT 146.715 -102.165 147.045 -101.835 ;
        RECT 146.715 -103.525 147.045 -103.195 ;
        RECT 146.715 -104.885 147.045 -104.555 ;
        RECT 146.715 -106.245 147.045 -105.915 ;
        RECT 146.715 -107.605 147.045 -107.275 ;
        RECT 146.715 -108.965 147.045 -108.635 ;
        RECT 146.715 -110.325 147.045 -109.995 ;
        RECT 146.715 -111.685 147.045 -111.355 ;
        RECT 146.715 -113.045 147.045 -112.715 ;
        RECT 146.715 -114.405 147.045 -114.075 ;
        RECT 146.715 -115.765 147.045 -115.435 ;
        RECT 146.715 -117.125 147.045 -116.795 ;
        RECT 146.715 -118.485 147.045 -118.155 ;
        RECT 146.715 -119.845 147.045 -119.515 ;
        RECT 146.715 -121.205 147.045 -120.875 ;
        RECT 146.715 -122.565 147.045 -122.235 ;
        RECT 146.715 -123.925 147.045 -123.595 ;
        RECT 146.715 -125.285 147.045 -124.955 ;
        RECT 146.715 -126.645 147.045 -126.315 ;
        RECT 146.715 -128.005 147.045 -127.675 ;
        RECT 146.715 -129.365 147.045 -129.035 ;
        RECT 146.715 -130.725 147.045 -130.395 ;
        RECT 146.715 -132.085 147.045 -131.755 ;
        RECT 146.715 -133.445 147.045 -133.115 ;
        RECT 146.715 -134.805 147.045 -134.475 ;
        RECT 146.715 -136.165 147.045 -135.835 ;
        RECT 146.715 -137.525 147.045 -137.195 ;
        RECT 146.715 -138.885 147.045 -138.555 ;
        RECT 146.715 -140.245 147.045 -139.915 ;
        RECT 146.715 -141.605 147.045 -141.275 ;
        RECT 146.715 -142.965 147.045 -142.635 ;
        RECT 146.715 -144.325 147.045 -143.995 ;
        RECT 146.715 -145.685 147.045 -145.355 ;
        RECT 146.715 -147.045 147.045 -146.715 ;
        RECT 146.715 -148.405 147.045 -148.075 ;
        RECT 146.715 -149.765 147.045 -149.435 ;
        RECT 146.715 -151.125 147.045 -150.795 ;
        RECT 146.715 -152.485 147.045 -152.155 ;
        RECT 146.715 -153.845 147.045 -153.515 ;
        RECT 146.715 -155.205 147.045 -154.875 ;
        RECT 146.715 -156.565 147.045 -156.235 ;
        RECT 146.715 -157.925 147.045 -157.595 ;
        RECT 146.715 -160.17 147.045 -159.04 ;
        RECT 146.72 -160.285 147.04 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 127.225 148.405 128.355 ;
        RECT 148.075 124.955 148.405 125.285 ;
        RECT 148.075 123.595 148.405 123.925 ;
        RECT 148.08 123.595 148.4 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -1.525 148.405 -1.195 ;
        RECT 148.075 -2.885 148.405 -2.555 ;
        RECT 148.08 -3.56 148.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -91.285 148.405 -90.955 ;
        RECT 148.075 -92.645 148.405 -92.315 ;
        RECT 148.075 -94.005 148.405 -93.675 ;
        RECT 148.075 -95.365 148.405 -95.035 ;
        RECT 148.075 -96.725 148.405 -96.395 ;
        RECT 148.075 -98.085 148.405 -97.755 ;
        RECT 148.075 -99.445 148.405 -99.115 ;
        RECT 148.075 -100.805 148.405 -100.475 ;
        RECT 148.075 -102.165 148.405 -101.835 ;
        RECT 148.075 -103.525 148.405 -103.195 ;
        RECT 148.075 -104.885 148.405 -104.555 ;
        RECT 148.075 -106.245 148.405 -105.915 ;
        RECT 148.075 -107.605 148.405 -107.275 ;
        RECT 148.075 -108.965 148.405 -108.635 ;
        RECT 148.075 -110.325 148.405 -109.995 ;
        RECT 148.075 -111.685 148.405 -111.355 ;
        RECT 148.075 -113.045 148.405 -112.715 ;
        RECT 148.075 -114.405 148.405 -114.075 ;
        RECT 148.075 -115.765 148.405 -115.435 ;
        RECT 148.075 -117.125 148.405 -116.795 ;
        RECT 148.075 -118.485 148.405 -118.155 ;
        RECT 148.075 -119.845 148.405 -119.515 ;
        RECT 148.075 -121.205 148.405 -120.875 ;
        RECT 148.075 -122.565 148.405 -122.235 ;
        RECT 148.075 -123.925 148.405 -123.595 ;
        RECT 148.075 -125.285 148.405 -124.955 ;
        RECT 148.075 -126.645 148.405 -126.315 ;
        RECT 148.075 -128.005 148.405 -127.675 ;
        RECT 148.075 -129.365 148.405 -129.035 ;
        RECT 148.075 -130.725 148.405 -130.395 ;
        RECT 148.075 -132.085 148.405 -131.755 ;
        RECT 148.075 -133.445 148.405 -133.115 ;
        RECT 148.075 -134.805 148.405 -134.475 ;
        RECT 148.075 -136.165 148.405 -135.835 ;
        RECT 148.075 -137.525 148.405 -137.195 ;
        RECT 148.075 -138.885 148.405 -138.555 ;
        RECT 148.075 -140.245 148.405 -139.915 ;
        RECT 148.075 -141.605 148.405 -141.275 ;
        RECT 148.075 -142.965 148.405 -142.635 ;
        RECT 148.075 -144.325 148.405 -143.995 ;
        RECT 148.075 -145.685 148.405 -145.355 ;
        RECT 148.075 -147.045 148.405 -146.715 ;
        RECT 148.075 -148.405 148.405 -148.075 ;
        RECT 148.075 -149.765 148.405 -149.435 ;
        RECT 148.075 -151.125 148.405 -150.795 ;
        RECT 148.075 -152.485 148.405 -152.155 ;
        RECT 148.075 -153.845 148.405 -153.515 ;
        RECT 148.075 -155.205 148.405 -154.875 ;
        RECT 148.075 -156.565 148.405 -156.235 ;
        RECT 148.075 -157.925 148.405 -157.595 ;
        RECT 148.075 -160.17 148.405 -159.04 ;
        RECT 148.08 -160.285 148.4 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 127.225 149.765 128.355 ;
        RECT 149.435 124.955 149.765 125.285 ;
        RECT 149.435 123.595 149.765 123.925 ;
        RECT 149.44 123.595 149.76 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 -95.365 149.765 -95.035 ;
        RECT 149.435 -96.725 149.765 -96.395 ;
        RECT 149.435 -98.085 149.765 -97.755 ;
        RECT 149.435 -99.445 149.765 -99.115 ;
        RECT 149.435 -100.805 149.765 -100.475 ;
        RECT 149.435 -102.165 149.765 -101.835 ;
        RECT 149.435 -103.525 149.765 -103.195 ;
        RECT 149.435 -104.885 149.765 -104.555 ;
        RECT 149.435 -106.245 149.765 -105.915 ;
        RECT 149.435 -107.605 149.765 -107.275 ;
        RECT 149.435 -108.965 149.765 -108.635 ;
        RECT 149.435 -110.325 149.765 -109.995 ;
        RECT 149.435 -111.685 149.765 -111.355 ;
        RECT 149.435 -113.045 149.765 -112.715 ;
        RECT 149.435 -114.405 149.765 -114.075 ;
        RECT 149.435 -115.765 149.765 -115.435 ;
        RECT 149.435 -117.125 149.765 -116.795 ;
        RECT 149.435 -118.485 149.765 -118.155 ;
        RECT 149.435 -119.845 149.765 -119.515 ;
        RECT 149.435 -121.205 149.765 -120.875 ;
        RECT 149.435 -122.565 149.765 -122.235 ;
        RECT 149.435 -123.925 149.765 -123.595 ;
        RECT 149.435 -125.285 149.765 -124.955 ;
        RECT 149.435 -126.645 149.765 -126.315 ;
        RECT 149.435 -128.005 149.765 -127.675 ;
        RECT 149.435 -129.365 149.765 -129.035 ;
        RECT 149.435 -130.725 149.765 -130.395 ;
        RECT 149.435 -132.085 149.765 -131.755 ;
        RECT 149.435 -133.445 149.765 -133.115 ;
        RECT 149.435 -134.805 149.765 -134.475 ;
        RECT 149.435 -136.165 149.765 -135.835 ;
        RECT 149.435 -137.525 149.765 -137.195 ;
        RECT 149.435 -138.885 149.765 -138.555 ;
        RECT 149.435 -140.245 149.765 -139.915 ;
        RECT 149.435 -141.605 149.765 -141.275 ;
        RECT 149.435 -142.965 149.765 -142.635 ;
        RECT 149.435 -144.325 149.765 -143.995 ;
        RECT 149.435 -145.685 149.765 -145.355 ;
        RECT 149.435 -147.045 149.765 -146.715 ;
        RECT 149.435 -148.405 149.765 -148.075 ;
        RECT 149.435 -149.765 149.765 -149.435 ;
        RECT 149.435 -151.125 149.765 -150.795 ;
        RECT 149.435 -152.485 149.765 -152.155 ;
        RECT 149.435 -153.845 149.765 -153.515 ;
        RECT 149.435 -155.205 149.765 -154.875 ;
        RECT 149.435 -156.565 149.765 -156.235 ;
        RECT 149.435 -157.925 149.765 -157.595 ;
        RECT 149.435 -160.17 149.765 -159.04 ;
        RECT 149.44 -160.285 149.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.71 -94.075 150.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 127.225 151.125 128.355 ;
        RECT 150.795 124.955 151.125 125.285 ;
        RECT 150.795 123.595 151.125 123.925 ;
        RECT 150.8 123.595 151.12 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 -1.525 151.125 -1.195 ;
        RECT 150.795 -2.885 151.125 -2.555 ;
        RECT 150.8 -3.56 151.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 127.225 152.485 128.355 ;
        RECT 152.155 124.955 152.485 125.285 ;
        RECT 152.155 123.595 152.485 123.925 ;
        RECT 152.16 123.595 152.48 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 -1.525 152.485 -1.195 ;
        RECT 152.155 -2.885 152.485 -2.555 ;
        RECT 152.16 -3.56 152.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 127.225 153.845 128.355 ;
        RECT 153.515 124.955 153.845 125.285 ;
        RECT 153.515 123.595 153.845 123.925 ;
        RECT 153.52 123.595 153.84 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 -1.525 153.845 -1.195 ;
        RECT 153.515 -2.885 153.845 -2.555 ;
        RECT 153.52 -3.56 153.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 127.225 155.205 128.355 ;
        RECT 154.875 124.955 155.205 125.285 ;
        RECT 154.875 123.595 155.205 123.925 ;
        RECT 154.88 123.595 155.2 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 -95.365 155.205 -95.035 ;
        RECT 154.875 -96.725 155.205 -96.395 ;
        RECT 154.875 -98.085 155.205 -97.755 ;
        RECT 154.875 -99.445 155.205 -99.115 ;
        RECT 154.875 -100.805 155.205 -100.475 ;
        RECT 154.875 -102.165 155.205 -101.835 ;
        RECT 154.875 -103.525 155.205 -103.195 ;
        RECT 154.875 -104.885 155.205 -104.555 ;
        RECT 154.875 -106.245 155.205 -105.915 ;
        RECT 154.875 -107.605 155.205 -107.275 ;
        RECT 154.875 -108.965 155.205 -108.635 ;
        RECT 154.875 -110.325 155.205 -109.995 ;
        RECT 154.875 -111.685 155.205 -111.355 ;
        RECT 154.875 -113.045 155.205 -112.715 ;
        RECT 154.875 -114.405 155.205 -114.075 ;
        RECT 154.875 -115.765 155.205 -115.435 ;
        RECT 154.875 -117.125 155.205 -116.795 ;
        RECT 154.875 -118.485 155.205 -118.155 ;
        RECT 154.875 -119.845 155.205 -119.515 ;
        RECT 154.875 -121.205 155.205 -120.875 ;
        RECT 154.875 -122.565 155.205 -122.235 ;
        RECT 154.875 -123.925 155.205 -123.595 ;
        RECT 154.875 -125.285 155.205 -124.955 ;
        RECT 154.875 -126.645 155.205 -126.315 ;
        RECT 154.875 -128.005 155.205 -127.675 ;
        RECT 154.875 -129.365 155.205 -129.035 ;
        RECT 154.875 -130.725 155.205 -130.395 ;
        RECT 154.875 -132.085 155.205 -131.755 ;
        RECT 154.875 -133.445 155.205 -133.115 ;
        RECT 154.875 -134.805 155.205 -134.475 ;
        RECT 154.875 -136.165 155.205 -135.835 ;
        RECT 154.875 -137.525 155.205 -137.195 ;
        RECT 154.875 -138.885 155.205 -138.555 ;
        RECT 154.875 -140.245 155.205 -139.915 ;
        RECT 154.875 -141.605 155.205 -141.275 ;
        RECT 154.875 -142.965 155.205 -142.635 ;
        RECT 154.875 -144.325 155.205 -143.995 ;
        RECT 154.875 -145.685 155.205 -145.355 ;
        RECT 154.875 -147.045 155.205 -146.715 ;
        RECT 154.875 -148.405 155.205 -148.075 ;
        RECT 154.875 -149.765 155.205 -149.435 ;
        RECT 154.875 -151.125 155.205 -150.795 ;
        RECT 154.875 -152.485 155.205 -152.155 ;
        RECT 154.875 -153.845 155.205 -153.515 ;
        RECT 154.875 -155.205 155.205 -154.875 ;
        RECT 154.875 -156.565 155.205 -156.235 ;
        RECT 154.875 -157.925 155.205 -157.595 ;
        RECT 154.875 -160.17 155.205 -159.04 ;
        RECT 154.88 -160.285 155.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.81 -94.075 156.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.235 127.225 156.565 128.355 ;
        RECT 156.235 124.955 156.565 125.285 ;
        RECT 156.235 123.595 156.565 123.925 ;
        RECT 156.24 123.595 156.56 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 127.225 157.925 128.355 ;
        RECT 157.595 124.955 157.925 125.285 ;
        RECT 157.595 123.595 157.925 123.925 ;
        RECT 157.6 123.595 157.92 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 -1.525 157.925 -1.195 ;
        RECT 157.595 -2.885 157.925 -2.555 ;
        RECT 157.6 -3.56 157.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 127.225 159.285 128.355 ;
        RECT 158.955 124.955 159.285 125.285 ;
        RECT 158.955 123.595 159.285 123.925 ;
        RECT 158.96 123.595 159.28 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -1.525 159.285 -1.195 ;
        RECT 158.955 -2.885 159.285 -2.555 ;
        RECT 158.96 -3.56 159.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -155.205 159.285 -154.875 ;
        RECT 158.955 -156.565 159.285 -156.235 ;
        RECT 158.955 -157.925 159.285 -157.595 ;
        RECT 158.955 -160.17 159.285 -159.04 ;
        RECT 158.96 -160.285 159.28 -90.955 ;
        RECT 158.955 -91.285 159.285 -90.955 ;
        RECT 158.955 -92.645 159.285 -92.315 ;
        RECT 158.955 -94.005 159.285 -93.675 ;
        RECT 158.955 -95.365 159.285 -95.035 ;
        RECT 158.955 -96.725 159.285 -96.395 ;
        RECT 158.955 -98.085 159.285 -97.755 ;
        RECT 158.955 -99.445 159.285 -99.115 ;
        RECT 158.955 -100.805 159.285 -100.475 ;
        RECT 158.955 -102.165 159.285 -101.835 ;
        RECT 158.955 -103.525 159.285 -103.195 ;
        RECT 158.955 -104.885 159.285 -104.555 ;
        RECT 158.955 -106.245 159.285 -105.915 ;
        RECT 158.955 -107.605 159.285 -107.275 ;
        RECT 158.955 -108.965 159.285 -108.635 ;
        RECT 158.955 -110.325 159.285 -109.995 ;
        RECT 158.955 -111.685 159.285 -111.355 ;
        RECT 158.955 -113.045 159.285 -112.715 ;
        RECT 158.955 -114.405 159.285 -114.075 ;
        RECT 158.955 -115.765 159.285 -115.435 ;
        RECT 158.955 -117.125 159.285 -116.795 ;
        RECT 158.955 -118.485 159.285 -118.155 ;
        RECT 158.955 -119.845 159.285 -119.515 ;
        RECT 158.955 -121.205 159.285 -120.875 ;
        RECT 158.955 -122.565 159.285 -122.235 ;
        RECT 158.955 -123.925 159.285 -123.595 ;
        RECT 158.955 -125.285 159.285 -124.955 ;
        RECT 158.955 -126.645 159.285 -126.315 ;
        RECT 158.955 -128.005 159.285 -127.675 ;
        RECT 158.955 -129.365 159.285 -129.035 ;
        RECT 158.955 -130.725 159.285 -130.395 ;
        RECT 158.955 -132.085 159.285 -131.755 ;
        RECT 158.955 -133.445 159.285 -133.115 ;
        RECT 158.955 -134.805 159.285 -134.475 ;
        RECT 158.955 -136.165 159.285 -135.835 ;
        RECT 158.955 -137.525 159.285 -137.195 ;
        RECT 158.955 -138.885 159.285 -138.555 ;
        RECT 158.955 -140.245 159.285 -139.915 ;
        RECT 158.955 -141.605 159.285 -141.275 ;
        RECT 158.955 -142.965 159.285 -142.635 ;
        RECT 158.955 -144.325 159.285 -143.995 ;
        RECT 158.955 -145.685 159.285 -145.355 ;
        RECT 158.955 -147.045 159.285 -146.715 ;
        RECT 158.955 -148.405 159.285 -148.075 ;
        RECT 158.955 -149.765 159.285 -149.435 ;
        RECT 158.955 -151.125 159.285 -150.795 ;
        RECT 158.955 -152.485 159.285 -152.155 ;
        RECT 158.955 -153.845 159.285 -153.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.41 -94.075 70.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 127.225 70.885 128.355 ;
        RECT 70.555 124.955 70.885 125.285 ;
        RECT 70.555 123.595 70.885 123.925 ;
        RECT 70.56 123.595 70.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 127.225 72.245 128.355 ;
        RECT 71.915 124.955 72.245 125.285 ;
        RECT 71.915 123.595 72.245 123.925 ;
        RECT 71.92 123.595 72.24 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -1.525 72.245 -1.195 ;
        RECT 71.915 -2.885 72.245 -2.555 ;
        RECT 71.92 -3.56 72.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -91.285 72.245 -90.955 ;
        RECT 71.915 -92.645 72.245 -92.315 ;
        RECT 71.915 -94.005 72.245 -93.675 ;
        RECT 71.915 -95.365 72.245 -95.035 ;
        RECT 71.915 -96.725 72.245 -96.395 ;
        RECT 71.915 -98.085 72.245 -97.755 ;
        RECT 71.915 -99.445 72.245 -99.115 ;
        RECT 71.915 -100.805 72.245 -100.475 ;
        RECT 71.915 -102.165 72.245 -101.835 ;
        RECT 71.915 -103.525 72.245 -103.195 ;
        RECT 71.915 -104.885 72.245 -104.555 ;
        RECT 71.915 -106.245 72.245 -105.915 ;
        RECT 71.915 -107.605 72.245 -107.275 ;
        RECT 71.915 -108.965 72.245 -108.635 ;
        RECT 71.915 -110.325 72.245 -109.995 ;
        RECT 71.915 -111.685 72.245 -111.355 ;
        RECT 71.915 -113.045 72.245 -112.715 ;
        RECT 71.915 -114.405 72.245 -114.075 ;
        RECT 71.915 -115.765 72.245 -115.435 ;
        RECT 71.915 -117.125 72.245 -116.795 ;
        RECT 71.915 -118.485 72.245 -118.155 ;
        RECT 71.915 -119.845 72.245 -119.515 ;
        RECT 71.915 -121.205 72.245 -120.875 ;
        RECT 71.915 -122.565 72.245 -122.235 ;
        RECT 71.915 -123.925 72.245 -123.595 ;
        RECT 71.915 -125.285 72.245 -124.955 ;
        RECT 71.915 -126.645 72.245 -126.315 ;
        RECT 71.915 -128.005 72.245 -127.675 ;
        RECT 71.915 -129.365 72.245 -129.035 ;
        RECT 71.915 -130.725 72.245 -130.395 ;
        RECT 71.915 -132.085 72.245 -131.755 ;
        RECT 71.915 -133.445 72.245 -133.115 ;
        RECT 71.915 -134.805 72.245 -134.475 ;
        RECT 71.915 -136.165 72.245 -135.835 ;
        RECT 71.915 -137.525 72.245 -137.195 ;
        RECT 71.915 -138.885 72.245 -138.555 ;
        RECT 71.915 -140.245 72.245 -139.915 ;
        RECT 71.915 -141.605 72.245 -141.275 ;
        RECT 71.915 -142.965 72.245 -142.635 ;
        RECT 71.915 -144.325 72.245 -143.995 ;
        RECT 71.915 -145.685 72.245 -145.355 ;
        RECT 71.915 -147.045 72.245 -146.715 ;
        RECT 71.915 -148.405 72.245 -148.075 ;
        RECT 71.915 -149.765 72.245 -149.435 ;
        RECT 71.915 -151.125 72.245 -150.795 ;
        RECT 71.915 -152.485 72.245 -152.155 ;
        RECT 71.915 -153.845 72.245 -153.515 ;
        RECT 71.915 -155.205 72.245 -154.875 ;
        RECT 71.915 -156.565 72.245 -156.235 ;
        RECT 71.915 -157.925 72.245 -157.595 ;
        RECT 71.915 -160.17 72.245 -159.04 ;
        RECT 71.92 -160.285 72.24 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 127.225 73.605 128.355 ;
        RECT 73.275 124.955 73.605 125.285 ;
        RECT 73.275 123.595 73.605 123.925 ;
        RECT 73.28 123.595 73.6 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 -1.525 73.605 -1.195 ;
        RECT 73.275 -2.885 73.605 -2.555 ;
        RECT 73.28 -3.56 73.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 127.225 74.965 128.355 ;
        RECT 74.635 124.955 74.965 125.285 ;
        RECT 74.635 123.595 74.965 123.925 ;
        RECT 74.64 123.595 74.96 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -1.525 74.965 -1.195 ;
        RECT 74.635 -2.885 74.965 -2.555 ;
        RECT 74.64 -3.56 74.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -91.285 74.965 -90.955 ;
        RECT 74.635 -92.645 74.965 -92.315 ;
        RECT 74.635 -94.005 74.965 -93.675 ;
        RECT 74.635 -95.365 74.965 -95.035 ;
        RECT 74.635 -96.725 74.965 -96.395 ;
        RECT 74.635 -98.085 74.965 -97.755 ;
        RECT 74.635 -99.445 74.965 -99.115 ;
        RECT 74.635 -100.805 74.965 -100.475 ;
        RECT 74.635 -102.165 74.965 -101.835 ;
        RECT 74.635 -103.525 74.965 -103.195 ;
        RECT 74.635 -104.885 74.965 -104.555 ;
        RECT 74.635 -106.245 74.965 -105.915 ;
        RECT 74.635 -107.605 74.965 -107.275 ;
        RECT 74.635 -108.965 74.965 -108.635 ;
        RECT 74.635 -110.325 74.965 -109.995 ;
        RECT 74.635 -111.685 74.965 -111.355 ;
        RECT 74.635 -113.045 74.965 -112.715 ;
        RECT 74.635 -114.405 74.965 -114.075 ;
        RECT 74.635 -115.765 74.965 -115.435 ;
        RECT 74.635 -117.125 74.965 -116.795 ;
        RECT 74.635 -118.485 74.965 -118.155 ;
        RECT 74.635 -119.845 74.965 -119.515 ;
        RECT 74.635 -121.205 74.965 -120.875 ;
        RECT 74.635 -122.565 74.965 -122.235 ;
        RECT 74.635 -123.925 74.965 -123.595 ;
        RECT 74.635 -125.285 74.965 -124.955 ;
        RECT 74.635 -126.645 74.965 -126.315 ;
        RECT 74.635 -128.005 74.965 -127.675 ;
        RECT 74.635 -129.365 74.965 -129.035 ;
        RECT 74.635 -130.725 74.965 -130.395 ;
        RECT 74.635 -132.085 74.965 -131.755 ;
        RECT 74.635 -133.445 74.965 -133.115 ;
        RECT 74.635 -134.805 74.965 -134.475 ;
        RECT 74.635 -136.165 74.965 -135.835 ;
        RECT 74.635 -137.525 74.965 -137.195 ;
        RECT 74.635 -138.885 74.965 -138.555 ;
        RECT 74.635 -140.245 74.965 -139.915 ;
        RECT 74.635 -141.605 74.965 -141.275 ;
        RECT 74.635 -142.965 74.965 -142.635 ;
        RECT 74.635 -144.325 74.965 -143.995 ;
        RECT 74.635 -145.685 74.965 -145.355 ;
        RECT 74.635 -147.045 74.965 -146.715 ;
        RECT 74.635 -148.405 74.965 -148.075 ;
        RECT 74.635 -149.765 74.965 -149.435 ;
        RECT 74.635 -151.125 74.965 -150.795 ;
        RECT 74.635 -152.485 74.965 -152.155 ;
        RECT 74.635 -153.845 74.965 -153.515 ;
        RECT 74.635 -155.205 74.965 -154.875 ;
        RECT 74.635 -156.565 74.965 -156.235 ;
        RECT 74.635 -157.925 74.965 -157.595 ;
        RECT 74.635 -160.17 74.965 -159.04 ;
        RECT 74.64 -160.285 74.96 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 127.225 76.325 128.355 ;
        RECT 75.995 124.955 76.325 125.285 ;
        RECT 75.995 123.595 76.325 123.925 ;
        RECT 76 123.595 76.32 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 -95.365 76.325 -95.035 ;
        RECT 75.995 -96.725 76.325 -96.395 ;
        RECT 75.995 -98.085 76.325 -97.755 ;
        RECT 75.995 -99.445 76.325 -99.115 ;
        RECT 75.995 -100.805 76.325 -100.475 ;
        RECT 75.995 -102.165 76.325 -101.835 ;
        RECT 75.995 -103.525 76.325 -103.195 ;
        RECT 75.995 -104.885 76.325 -104.555 ;
        RECT 75.995 -106.245 76.325 -105.915 ;
        RECT 75.995 -107.605 76.325 -107.275 ;
        RECT 75.995 -108.965 76.325 -108.635 ;
        RECT 75.995 -110.325 76.325 -109.995 ;
        RECT 75.995 -111.685 76.325 -111.355 ;
        RECT 75.995 -113.045 76.325 -112.715 ;
        RECT 75.995 -114.405 76.325 -114.075 ;
        RECT 75.995 -115.765 76.325 -115.435 ;
        RECT 75.995 -117.125 76.325 -116.795 ;
        RECT 75.995 -118.485 76.325 -118.155 ;
        RECT 75.995 -119.845 76.325 -119.515 ;
        RECT 75.995 -121.205 76.325 -120.875 ;
        RECT 75.995 -122.565 76.325 -122.235 ;
        RECT 75.995 -123.925 76.325 -123.595 ;
        RECT 75.995 -125.285 76.325 -124.955 ;
        RECT 75.995 -126.645 76.325 -126.315 ;
        RECT 75.995 -128.005 76.325 -127.675 ;
        RECT 75.995 -129.365 76.325 -129.035 ;
        RECT 75.995 -130.725 76.325 -130.395 ;
        RECT 75.995 -132.085 76.325 -131.755 ;
        RECT 75.995 -133.445 76.325 -133.115 ;
        RECT 75.995 -134.805 76.325 -134.475 ;
        RECT 75.995 -136.165 76.325 -135.835 ;
        RECT 75.995 -137.525 76.325 -137.195 ;
        RECT 75.995 -138.885 76.325 -138.555 ;
        RECT 75.995 -140.245 76.325 -139.915 ;
        RECT 75.995 -141.605 76.325 -141.275 ;
        RECT 75.995 -142.965 76.325 -142.635 ;
        RECT 75.995 -144.325 76.325 -143.995 ;
        RECT 75.995 -145.685 76.325 -145.355 ;
        RECT 75.995 -147.045 76.325 -146.715 ;
        RECT 75.995 -148.405 76.325 -148.075 ;
        RECT 75.995 -149.765 76.325 -149.435 ;
        RECT 75.995 -151.125 76.325 -150.795 ;
        RECT 75.995 -152.485 76.325 -152.155 ;
        RECT 75.995 -153.845 76.325 -153.515 ;
        RECT 75.995 -155.205 76.325 -154.875 ;
        RECT 75.995 -156.565 76.325 -156.235 ;
        RECT 75.995 -157.925 76.325 -157.595 ;
        RECT 75.995 -160.17 76.325 -159.04 ;
        RECT 76 -160.285 76.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.51 -94.075 76.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 127.225 77.685 128.355 ;
        RECT 77.355 124.955 77.685 125.285 ;
        RECT 77.355 123.595 77.685 123.925 ;
        RECT 77.36 123.595 77.68 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 -1.525 77.685 -1.195 ;
        RECT 77.355 -2.885 77.685 -2.555 ;
        RECT 77.36 -3.56 77.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 127.225 79.045 128.355 ;
        RECT 78.715 124.955 79.045 125.285 ;
        RECT 78.715 123.595 79.045 123.925 ;
        RECT 78.72 123.595 79.04 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 -1.525 79.045 -1.195 ;
        RECT 78.715 -2.885 79.045 -2.555 ;
        RECT 78.72 -3.56 79.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 127.225 80.405 128.355 ;
        RECT 80.075 124.955 80.405 125.285 ;
        RECT 80.075 123.595 80.405 123.925 ;
        RECT 80.08 123.595 80.4 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 -1.525 80.405 -1.195 ;
        RECT 80.075 -2.885 80.405 -2.555 ;
        RECT 80.08 -3.56 80.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 -91.285 80.405 -90.955 ;
        RECT 80.075 -92.645 80.405 -92.315 ;
        RECT 80.075 -94.005 80.405 -93.675 ;
        RECT 80.075 -95.365 80.405 -95.035 ;
        RECT 80.075 -96.725 80.405 -96.395 ;
        RECT 80.075 -98.085 80.405 -97.755 ;
        RECT 80.075 -99.445 80.405 -99.115 ;
        RECT 80.075 -100.805 80.405 -100.475 ;
        RECT 80.075 -102.165 80.405 -101.835 ;
        RECT 80.075 -103.525 80.405 -103.195 ;
        RECT 80.075 -104.885 80.405 -104.555 ;
        RECT 80.075 -106.245 80.405 -105.915 ;
        RECT 80.075 -107.605 80.405 -107.275 ;
        RECT 80.075 -108.965 80.405 -108.635 ;
        RECT 80.075 -110.325 80.405 -109.995 ;
        RECT 80.075 -111.685 80.405 -111.355 ;
        RECT 80.075 -113.045 80.405 -112.715 ;
        RECT 80.075 -114.405 80.405 -114.075 ;
        RECT 80.075 -115.765 80.405 -115.435 ;
        RECT 80.075 -117.125 80.405 -116.795 ;
        RECT 80.075 -118.485 80.405 -118.155 ;
        RECT 80.075 -119.845 80.405 -119.515 ;
        RECT 80.075 -121.205 80.405 -120.875 ;
        RECT 80.075 -122.565 80.405 -122.235 ;
        RECT 80.075 -123.925 80.405 -123.595 ;
        RECT 80.075 -125.285 80.405 -124.955 ;
        RECT 80.075 -126.645 80.405 -126.315 ;
        RECT 80.075 -128.005 80.405 -127.675 ;
        RECT 80.075 -129.365 80.405 -129.035 ;
        RECT 80.075 -130.725 80.405 -130.395 ;
        RECT 80.075 -132.085 80.405 -131.755 ;
        RECT 80.075 -133.445 80.405 -133.115 ;
        RECT 80.075 -134.805 80.405 -134.475 ;
        RECT 80.075 -136.165 80.405 -135.835 ;
        RECT 80.075 -137.525 80.405 -137.195 ;
        RECT 80.075 -138.885 80.405 -138.555 ;
        RECT 80.075 -140.245 80.405 -139.915 ;
        RECT 80.075 -141.605 80.405 -141.275 ;
        RECT 80.075 -142.965 80.405 -142.635 ;
        RECT 80.075 -144.325 80.405 -143.995 ;
        RECT 80.075 -145.685 80.405 -145.355 ;
        RECT 80.075 -147.045 80.405 -146.715 ;
        RECT 80.075 -148.405 80.405 -148.075 ;
        RECT 80.075 -149.765 80.405 -149.435 ;
        RECT 80.075 -151.125 80.405 -150.795 ;
        RECT 80.075 -152.485 80.405 -152.155 ;
        RECT 80.075 -153.845 80.405 -153.515 ;
        RECT 80.075 -155.205 80.405 -154.875 ;
        RECT 80.075 -156.565 80.405 -156.235 ;
        RECT 80.075 -157.925 80.405 -157.595 ;
        RECT 80.075 -160.17 80.405 -159.04 ;
        RECT 80.08 -160.285 80.4 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 127.225 81.765 128.355 ;
        RECT 81.435 124.955 81.765 125.285 ;
        RECT 81.435 123.595 81.765 123.925 ;
        RECT 81.44 123.595 81.76 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 -95.365 81.765 -95.035 ;
        RECT 81.435 -96.725 81.765 -96.395 ;
        RECT 81.435 -98.085 81.765 -97.755 ;
        RECT 81.435 -99.445 81.765 -99.115 ;
        RECT 81.435 -100.805 81.765 -100.475 ;
        RECT 81.435 -102.165 81.765 -101.835 ;
        RECT 81.435 -103.525 81.765 -103.195 ;
        RECT 81.435 -104.885 81.765 -104.555 ;
        RECT 81.435 -106.245 81.765 -105.915 ;
        RECT 81.435 -107.605 81.765 -107.275 ;
        RECT 81.435 -108.965 81.765 -108.635 ;
        RECT 81.435 -110.325 81.765 -109.995 ;
        RECT 81.435 -111.685 81.765 -111.355 ;
        RECT 81.435 -113.045 81.765 -112.715 ;
        RECT 81.435 -114.405 81.765 -114.075 ;
        RECT 81.435 -115.765 81.765 -115.435 ;
        RECT 81.435 -117.125 81.765 -116.795 ;
        RECT 81.435 -118.485 81.765 -118.155 ;
        RECT 81.435 -119.845 81.765 -119.515 ;
        RECT 81.435 -121.205 81.765 -120.875 ;
        RECT 81.435 -122.565 81.765 -122.235 ;
        RECT 81.435 -123.925 81.765 -123.595 ;
        RECT 81.435 -125.285 81.765 -124.955 ;
        RECT 81.435 -126.645 81.765 -126.315 ;
        RECT 81.435 -128.005 81.765 -127.675 ;
        RECT 81.435 -129.365 81.765 -129.035 ;
        RECT 81.435 -130.725 81.765 -130.395 ;
        RECT 81.435 -132.085 81.765 -131.755 ;
        RECT 81.435 -133.445 81.765 -133.115 ;
        RECT 81.435 -134.805 81.765 -134.475 ;
        RECT 81.435 -136.165 81.765 -135.835 ;
        RECT 81.435 -137.525 81.765 -137.195 ;
        RECT 81.435 -138.885 81.765 -138.555 ;
        RECT 81.435 -140.245 81.765 -139.915 ;
        RECT 81.435 -141.605 81.765 -141.275 ;
        RECT 81.435 -142.965 81.765 -142.635 ;
        RECT 81.435 -144.325 81.765 -143.995 ;
        RECT 81.435 -145.685 81.765 -145.355 ;
        RECT 81.435 -147.045 81.765 -146.715 ;
        RECT 81.435 -148.405 81.765 -148.075 ;
        RECT 81.435 -149.765 81.765 -149.435 ;
        RECT 81.435 -151.125 81.765 -150.795 ;
        RECT 81.435 -152.485 81.765 -152.155 ;
        RECT 81.435 -153.845 81.765 -153.515 ;
        RECT 81.435 -155.205 81.765 -154.875 ;
        RECT 81.435 -156.565 81.765 -156.235 ;
        RECT 81.435 -157.925 81.765 -157.595 ;
        RECT 81.435 -160.17 81.765 -159.04 ;
        RECT 81.44 -160.285 81.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.61 -94.075 82.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 127.225 83.125 128.355 ;
        RECT 82.795 124.955 83.125 125.285 ;
        RECT 82.795 123.595 83.125 123.925 ;
        RECT 82.8 123.595 83.12 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 127.225 84.485 128.355 ;
        RECT 84.155 124.955 84.485 125.285 ;
        RECT 84.155 123.595 84.485 123.925 ;
        RECT 84.16 123.595 84.48 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -1.525 84.485 -1.195 ;
        RECT 84.155 -2.885 84.485 -2.555 ;
        RECT 84.16 -3.56 84.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -91.285 84.485 -90.955 ;
        RECT 84.155 -92.645 84.485 -92.315 ;
        RECT 84.155 -94.005 84.485 -93.675 ;
        RECT 84.155 -95.365 84.485 -95.035 ;
        RECT 84.155 -96.725 84.485 -96.395 ;
        RECT 84.155 -98.085 84.485 -97.755 ;
        RECT 84.155 -99.445 84.485 -99.115 ;
        RECT 84.155 -100.805 84.485 -100.475 ;
        RECT 84.155 -102.165 84.485 -101.835 ;
        RECT 84.155 -103.525 84.485 -103.195 ;
        RECT 84.155 -104.885 84.485 -104.555 ;
        RECT 84.155 -106.245 84.485 -105.915 ;
        RECT 84.155 -107.605 84.485 -107.275 ;
        RECT 84.155 -108.965 84.485 -108.635 ;
        RECT 84.155 -110.325 84.485 -109.995 ;
        RECT 84.155 -111.685 84.485 -111.355 ;
        RECT 84.155 -113.045 84.485 -112.715 ;
        RECT 84.155 -114.405 84.485 -114.075 ;
        RECT 84.155 -115.765 84.485 -115.435 ;
        RECT 84.155 -117.125 84.485 -116.795 ;
        RECT 84.155 -118.485 84.485 -118.155 ;
        RECT 84.155 -119.845 84.485 -119.515 ;
        RECT 84.155 -121.205 84.485 -120.875 ;
        RECT 84.155 -122.565 84.485 -122.235 ;
        RECT 84.155 -123.925 84.485 -123.595 ;
        RECT 84.155 -125.285 84.485 -124.955 ;
        RECT 84.155 -126.645 84.485 -126.315 ;
        RECT 84.155 -128.005 84.485 -127.675 ;
        RECT 84.155 -129.365 84.485 -129.035 ;
        RECT 84.155 -130.725 84.485 -130.395 ;
        RECT 84.155 -132.085 84.485 -131.755 ;
        RECT 84.155 -133.445 84.485 -133.115 ;
        RECT 84.155 -134.805 84.485 -134.475 ;
        RECT 84.155 -136.165 84.485 -135.835 ;
        RECT 84.155 -137.525 84.485 -137.195 ;
        RECT 84.155 -138.885 84.485 -138.555 ;
        RECT 84.155 -140.245 84.485 -139.915 ;
        RECT 84.155 -141.605 84.485 -141.275 ;
        RECT 84.155 -142.965 84.485 -142.635 ;
        RECT 84.155 -144.325 84.485 -143.995 ;
        RECT 84.155 -145.685 84.485 -145.355 ;
        RECT 84.155 -147.045 84.485 -146.715 ;
        RECT 84.155 -148.405 84.485 -148.075 ;
        RECT 84.155 -149.765 84.485 -149.435 ;
        RECT 84.155 -151.125 84.485 -150.795 ;
        RECT 84.155 -152.485 84.485 -152.155 ;
        RECT 84.155 -153.845 84.485 -153.515 ;
        RECT 84.155 -155.205 84.485 -154.875 ;
        RECT 84.155 -156.565 84.485 -156.235 ;
        RECT 84.155 -157.925 84.485 -157.595 ;
        RECT 84.155 -160.17 84.485 -159.04 ;
        RECT 84.16 -160.285 84.48 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 127.225 85.845 128.355 ;
        RECT 85.515 124.955 85.845 125.285 ;
        RECT 85.515 123.595 85.845 123.925 ;
        RECT 85.52 123.595 85.84 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 -1.525 85.845 -1.195 ;
        RECT 85.515 -2.885 85.845 -2.555 ;
        RECT 85.52 -3.56 85.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 127.225 87.205 128.355 ;
        RECT 86.875 124.955 87.205 125.285 ;
        RECT 86.875 123.595 87.205 123.925 ;
        RECT 86.88 123.595 87.2 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -1.525 87.205 -1.195 ;
        RECT 86.875 -2.885 87.205 -2.555 ;
        RECT 86.88 -3.56 87.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -91.285 87.205 -90.955 ;
        RECT 86.875 -92.645 87.205 -92.315 ;
        RECT 86.875 -94.005 87.205 -93.675 ;
        RECT 86.875 -95.365 87.205 -95.035 ;
        RECT 86.875 -96.725 87.205 -96.395 ;
        RECT 86.875 -98.085 87.205 -97.755 ;
        RECT 86.875 -99.445 87.205 -99.115 ;
        RECT 86.875 -100.805 87.205 -100.475 ;
        RECT 86.875 -102.165 87.205 -101.835 ;
        RECT 86.875 -103.525 87.205 -103.195 ;
        RECT 86.875 -104.885 87.205 -104.555 ;
        RECT 86.875 -106.245 87.205 -105.915 ;
        RECT 86.875 -107.605 87.205 -107.275 ;
        RECT 86.875 -108.965 87.205 -108.635 ;
        RECT 86.875 -110.325 87.205 -109.995 ;
        RECT 86.875 -111.685 87.205 -111.355 ;
        RECT 86.875 -113.045 87.205 -112.715 ;
        RECT 86.875 -114.405 87.205 -114.075 ;
        RECT 86.875 -115.765 87.205 -115.435 ;
        RECT 86.875 -117.125 87.205 -116.795 ;
        RECT 86.875 -118.485 87.205 -118.155 ;
        RECT 86.875 -119.845 87.205 -119.515 ;
        RECT 86.875 -121.205 87.205 -120.875 ;
        RECT 86.875 -122.565 87.205 -122.235 ;
        RECT 86.875 -123.925 87.205 -123.595 ;
        RECT 86.875 -125.285 87.205 -124.955 ;
        RECT 86.875 -126.645 87.205 -126.315 ;
        RECT 86.875 -128.005 87.205 -127.675 ;
        RECT 86.875 -129.365 87.205 -129.035 ;
        RECT 86.875 -130.725 87.205 -130.395 ;
        RECT 86.875 -132.085 87.205 -131.755 ;
        RECT 86.875 -133.445 87.205 -133.115 ;
        RECT 86.875 -134.805 87.205 -134.475 ;
        RECT 86.875 -136.165 87.205 -135.835 ;
        RECT 86.875 -137.525 87.205 -137.195 ;
        RECT 86.875 -138.885 87.205 -138.555 ;
        RECT 86.875 -140.245 87.205 -139.915 ;
        RECT 86.875 -141.605 87.205 -141.275 ;
        RECT 86.875 -142.965 87.205 -142.635 ;
        RECT 86.875 -144.325 87.205 -143.995 ;
        RECT 86.875 -145.685 87.205 -145.355 ;
        RECT 86.875 -147.045 87.205 -146.715 ;
        RECT 86.875 -148.405 87.205 -148.075 ;
        RECT 86.875 -149.765 87.205 -149.435 ;
        RECT 86.875 -151.125 87.205 -150.795 ;
        RECT 86.875 -152.485 87.205 -152.155 ;
        RECT 86.875 -153.845 87.205 -153.515 ;
        RECT 86.875 -155.205 87.205 -154.875 ;
        RECT 86.875 -156.565 87.205 -156.235 ;
        RECT 86.875 -157.925 87.205 -157.595 ;
        RECT 86.875 -160.17 87.205 -159.04 ;
        RECT 86.88 -160.285 87.2 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 127.225 88.565 128.355 ;
        RECT 88.235 124.955 88.565 125.285 ;
        RECT 88.235 123.595 88.565 123.925 ;
        RECT 88.24 123.595 88.56 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 -95.365 88.565 -95.035 ;
        RECT 88.235 -96.725 88.565 -96.395 ;
        RECT 88.235 -98.085 88.565 -97.755 ;
        RECT 88.235 -99.445 88.565 -99.115 ;
        RECT 88.235 -100.805 88.565 -100.475 ;
        RECT 88.235 -102.165 88.565 -101.835 ;
        RECT 88.235 -103.525 88.565 -103.195 ;
        RECT 88.235 -104.885 88.565 -104.555 ;
        RECT 88.235 -106.245 88.565 -105.915 ;
        RECT 88.235 -107.605 88.565 -107.275 ;
        RECT 88.235 -108.965 88.565 -108.635 ;
        RECT 88.235 -110.325 88.565 -109.995 ;
        RECT 88.235 -111.685 88.565 -111.355 ;
        RECT 88.235 -113.045 88.565 -112.715 ;
        RECT 88.235 -114.405 88.565 -114.075 ;
        RECT 88.235 -115.765 88.565 -115.435 ;
        RECT 88.235 -117.125 88.565 -116.795 ;
        RECT 88.235 -118.485 88.565 -118.155 ;
        RECT 88.235 -119.845 88.565 -119.515 ;
        RECT 88.235 -121.205 88.565 -120.875 ;
        RECT 88.235 -122.565 88.565 -122.235 ;
        RECT 88.235 -123.925 88.565 -123.595 ;
        RECT 88.235 -125.285 88.565 -124.955 ;
        RECT 88.235 -126.645 88.565 -126.315 ;
        RECT 88.235 -128.005 88.565 -127.675 ;
        RECT 88.235 -129.365 88.565 -129.035 ;
        RECT 88.235 -130.725 88.565 -130.395 ;
        RECT 88.235 -132.085 88.565 -131.755 ;
        RECT 88.235 -133.445 88.565 -133.115 ;
        RECT 88.235 -134.805 88.565 -134.475 ;
        RECT 88.235 -136.165 88.565 -135.835 ;
        RECT 88.235 -137.525 88.565 -137.195 ;
        RECT 88.235 -138.885 88.565 -138.555 ;
        RECT 88.235 -140.245 88.565 -139.915 ;
        RECT 88.235 -141.605 88.565 -141.275 ;
        RECT 88.235 -142.965 88.565 -142.635 ;
        RECT 88.235 -144.325 88.565 -143.995 ;
        RECT 88.235 -145.685 88.565 -145.355 ;
        RECT 88.235 -147.045 88.565 -146.715 ;
        RECT 88.235 -148.405 88.565 -148.075 ;
        RECT 88.235 -149.765 88.565 -149.435 ;
        RECT 88.235 -151.125 88.565 -150.795 ;
        RECT 88.235 -152.485 88.565 -152.155 ;
        RECT 88.235 -153.845 88.565 -153.515 ;
        RECT 88.235 -155.205 88.565 -154.875 ;
        RECT 88.235 -156.565 88.565 -156.235 ;
        RECT 88.235 -157.925 88.565 -157.595 ;
        RECT 88.235 -160.17 88.565 -159.04 ;
        RECT 88.24 -160.285 88.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.71 -94.075 89.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 127.225 89.925 128.355 ;
        RECT 89.595 124.955 89.925 125.285 ;
        RECT 89.595 123.595 89.925 123.925 ;
        RECT 89.6 123.595 89.92 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 -1.525 89.925 -1.195 ;
        RECT 89.595 -2.885 89.925 -2.555 ;
        RECT 89.6 -3.56 89.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 127.225 91.285 128.355 ;
        RECT 90.955 124.955 91.285 125.285 ;
        RECT 90.955 123.595 91.285 123.925 ;
        RECT 90.96 123.595 91.28 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 -1.525 91.285 -1.195 ;
        RECT 90.955 -2.885 91.285 -2.555 ;
        RECT 90.96 -3.56 91.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 127.225 92.645 128.355 ;
        RECT 92.315 124.955 92.645 125.285 ;
        RECT 92.315 123.595 92.645 123.925 ;
        RECT 92.32 123.595 92.64 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -1.525 92.645 -1.195 ;
        RECT 92.315 -2.885 92.645 -2.555 ;
        RECT 92.32 -3.56 92.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -91.285 92.645 -90.955 ;
        RECT 92.315 -92.645 92.645 -92.315 ;
        RECT 92.315 -94.005 92.645 -93.675 ;
        RECT 92.315 -95.365 92.645 -95.035 ;
        RECT 92.315 -96.725 92.645 -96.395 ;
        RECT 92.315 -98.085 92.645 -97.755 ;
        RECT 92.315 -99.445 92.645 -99.115 ;
        RECT 92.315 -100.805 92.645 -100.475 ;
        RECT 92.315 -102.165 92.645 -101.835 ;
        RECT 92.315 -103.525 92.645 -103.195 ;
        RECT 92.315 -104.885 92.645 -104.555 ;
        RECT 92.315 -106.245 92.645 -105.915 ;
        RECT 92.315 -107.605 92.645 -107.275 ;
        RECT 92.315 -108.965 92.645 -108.635 ;
        RECT 92.315 -110.325 92.645 -109.995 ;
        RECT 92.315 -111.685 92.645 -111.355 ;
        RECT 92.315 -113.045 92.645 -112.715 ;
        RECT 92.315 -114.405 92.645 -114.075 ;
        RECT 92.315 -115.765 92.645 -115.435 ;
        RECT 92.315 -117.125 92.645 -116.795 ;
        RECT 92.315 -118.485 92.645 -118.155 ;
        RECT 92.315 -119.845 92.645 -119.515 ;
        RECT 92.315 -121.205 92.645 -120.875 ;
        RECT 92.315 -122.565 92.645 -122.235 ;
        RECT 92.315 -123.925 92.645 -123.595 ;
        RECT 92.315 -125.285 92.645 -124.955 ;
        RECT 92.315 -126.645 92.645 -126.315 ;
        RECT 92.315 -128.005 92.645 -127.675 ;
        RECT 92.315 -129.365 92.645 -129.035 ;
        RECT 92.315 -130.725 92.645 -130.395 ;
        RECT 92.315 -132.085 92.645 -131.755 ;
        RECT 92.315 -133.445 92.645 -133.115 ;
        RECT 92.315 -134.805 92.645 -134.475 ;
        RECT 92.315 -136.165 92.645 -135.835 ;
        RECT 92.315 -137.525 92.645 -137.195 ;
        RECT 92.315 -138.885 92.645 -138.555 ;
        RECT 92.315 -140.245 92.645 -139.915 ;
        RECT 92.315 -141.605 92.645 -141.275 ;
        RECT 92.315 -142.965 92.645 -142.635 ;
        RECT 92.315 -144.325 92.645 -143.995 ;
        RECT 92.315 -145.685 92.645 -145.355 ;
        RECT 92.315 -147.045 92.645 -146.715 ;
        RECT 92.315 -148.405 92.645 -148.075 ;
        RECT 92.315 -149.765 92.645 -149.435 ;
        RECT 92.315 -151.125 92.645 -150.795 ;
        RECT 92.315 -152.485 92.645 -152.155 ;
        RECT 92.315 -153.845 92.645 -153.515 ;
        RECT 92.315 -155.205 92.645 -154.875 ;
        RECT 92.315 -156.565 92.645 -156.235 ;
        RECT 92.315 -157.925 92.645 -157.595 ;
        RECT 92.315 -160.17 92.645 -159.04 ;
        RECT 92.32 -160.285 92.64 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 127.225 94.005 128.355 ;
        RECT 93.675 124.955 94.005 125.285 ;
        RECT 93.675 123.595 94.005 123.925 ;
        RECT 93.68 123.595 94 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 -95.365 94.005 -95.035 ;
        RECT 93.675 -96.725 94.005 -96.395 ;
        RECT 93.675 -98.085 94.005 -97.755 ;
        RECT 93.675 -99.445 94.005 -99.115 ;
        RECT 93.675 -100.805 94.005 -100.475 ;
        RECT 93.675 -102.165 94.005 -101.835 ;
        RECT 93.675 -103.525 94.005 -103.195 ;
        RECT 93.675 -104.885 94.005 -104.555 ;
        RECT 93.675 -106.245 94.005 -105.915 ;
        RECT 93.675 -107.605 94.005 -107.275 ;
        RECT 93.675 -108.965 94.005 -108.635 ;
        RECT 93.675 -110.325 94.005 -109.995 ;
        RECT 93.675 -111.685 94.005 -111.355 ;
        RECT 93.675 -113.045 94.005 -112.715 ;
        RECT 93.675 -114.405 94.005 -114.075 ;
        RECT 93.675 -115.765 94.005 -115.435 ;
        RECT 93.675 -117.125 94.005 -116.795 ;
        RECT 93.675 -118.485 94.005 -118.155 ;
        RECT 93.675 -119.845 94.005 -119.515 ;
        RECT 93.675 -121.205 94.005 -120.875 ;
        RECT 93.675 -122.565 94.005 -122.235 ;
        RECT 93.675 -123.925 94.005 -123.595 ;
        RECT 93.675 -125.285 94.005 -124.955 ;
        RECT 93.675 -126.645 94.005 -126.315 ;
        RECT 93.675 -128.005 94.005 -127.675 ;
        RECT 93.675 -129.365 94.005 -129.035 ;
        RECT 93.675 -130.725 94.005 -130.395 ;
        RECT 93.675 -132.085 94.005 -131.755 ;
        RECT 93.675 -133.445 94.005 -133.115 ;
        RECT 93.675 -134.805 94.005 -134.475 ;
        RECT 93.675 -136.165 94.005 -135.835 ;
        RECT 93.675 -137.525 94.005 -137.195 ;
        RECT 93.675 -138.885 94.005 -138.555 ;
        RECT 93.675 -140.245 94.005 -139.915 ;
        RECT 93.675 -141.605 94.005 -141.275 ;
        RECT 93.675 -142.965 94.005 -142.635 ;
        RECT 93.675 -144.325 94.005 -143.995 ;
        RECT 93.675 -145.685 94.005 -145.355 ;
        RECT 93.675 -147.045 94.005 -146.715 ;
        RECT 93.675 -148.405 94.005 -148.075 ;
        RECT 93.675 -149.765 94.005 -149.435 ;
        RECT 93.675 -151.125 94.005 -150.795 ;
        RECT 93.675 -152.485 94.005 -152.155 ;
        RECT 93.675 -153.845 94.005 -153.515 ;
        RECT 93.675 -155.205 94.005 -154.875 ;
        RECT 93.675 -156.565 94.005 -156.235 ;
        RECT 93.675 -157.925 94.005 -157.595 ;
        RECT 93.675 -160.17 94.005 -159.04 ;
        RECT 93.68 -160.285 94 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.81 -94.075 95.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 127.225 95.365 128.355 ;
        RECT 95.035 124.955 95.365 125.285 ;
        RECT 95.035 123.595 95.365 123.925 ;
        RECT 95.04 123.595 95.36 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 127.225 96.725 128.355 ;
        RECT 96.395 124.955 96.725 125.285 ;
        RECT 96.395 123.595 96.725 123.925 ;
        RECT 96.4 123.595 96.72 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -1.525 96.725 -1.195 ;
        RECT 96.395 -2.885 96.725 -2.555 ;
        RECT 96.4 -3.56 96.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -91.285 96.725 -90.955 ;
        RECT 96.395 -92.645 96.725 -92.315 ;
        RECT 96.395 -94.005 96.725 -93.675 ;
        RECT 96.395 -95.365 96.725 -95.035 ;
        RECT 96.395 -96.725 96.725 -96.395 ;
        RECT 96.395 -98.085 96.725 -97.755 ;
        RECT 96.395 -99.445 96.725 -99.115 ;
        RECT 96.395 -100.805 96.725 -100.475 ;
        RECT 96.395 -102.165 96.725 -101.835 ;
        RECT 96.395 -103.525 96.725 -103.195 ;
        RECT 96.395 -104.885 96.725 -104.555 ;
        RECT 96.395 -106.245 96.725 -105.915 ;
        RECT 96.395 -107.605 96.725 -107.275 ;
        RECT 96.395 -108.965 96.725 -108.635 ;
        RECT 96.395 -110.325 96.725 -109.995 ;
        RECT 96.395 -111.685 96.725 -111.355 ;
        RECT 96.395 -113.045 96.725 -112.715 ;
        RECT 96.395 -114.405 96.725 -114.075 ;
        RECT 96.395 -115.765 96.725 -115.435 ;
        RECT 96.395 -117.125 96.725 -116.795 ;
        RECT 96.395 -118.485 96.725 -118.155 ;
        RECT 96.395 -119.845 96.725 -119.515 ;
        RECT 96.395 -121.205 96.725 -120.875 ;
        RECT 96.395 -122.565 96.725 -122.235 ;
        RECT 96.395 -123.925 96.725 -123.595 ;
        RECT 96.395 -125.285 96.725 -124.955 ;
        RECT 96.395 -126.645 96.725 -126.315 ;
        RECT 96.395 -128.005 96.725 -127.675 ;
        RECT 96.395 -129.365 96.725 -129.035 ;
        RECT 96.395 -130.725 96.725 -130.395 ;
        RECT 96.395 -132.085 96.725 -131.755 ;
        RECT 96.395 -133.445 96.725 -133.115 ;
        RECT 96.395 -134.805 96.725 -134.475 ;
        RECT 96.395 -136.165 96.725 -135.835 ;
        RECT 96.395 -137.525 96.725 -137.195 ;
        RECT 96.395 -138.885 96.725 -138.555 ;
        RECT 96.395 -140.245 96.725 -139.915 ;
        RECT 96.395 -141.605 96.725 -141.275 ;
        RECT 96.395 -142.965 96.725 -142.635 ;
        RECT 96.395 -144.325 96.725 -143.995 ;
        RECT 96.395 -145.685 96.725 -145.355 ;
        RECT 96.395 -147.045 96.725 -146.715 ;
        RECT 96.395 -148.405 96.725 -148.075 ;
        RECT 96.395 -149.765 96.725 -149.435 ;
        RECT 96.395 -151.125 96.725 -150.795 ;
        RECT 96.395 -152.485 96.725 -152.155 ;
        RECT 96.395 -153.845 96.725 -153.515 ;
        RECT 96.395 -155.205 96.725 -154.875 ;
        RECT 96.395 -156.565 96.725 -156.235 ;
        RECT 96.395 -157.925 96.725 -157.595 ;
        RECT 96.395 -160.17 96.725 -159.04 ;
        RECT 96.4 -160.285 96.72 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 127.225 98.085 128.355 ;
        RECT 97.755 124.955 98.085 125.285 ;
        RECT 97.755 123.595 98.085 123.925 ;
        RECT 97.76 123.595 98.08 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 -1.525 98.085 -1.195 ;
        RECT 97.755 -2.885 98.085 -2.555 ;
        RECT 97.76 -3.56 98.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 127.225 99.445 128.355 ;
        RECT 99.115 124.955 99.445 125.285 ;
        RECT 99.115 123.595 99.445 123.925 ;
        RECT 99.12 123.595 99.44 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -1.525 99.445 -1.195 ;
        RECT 99.115 -2.885 99.445 -2.555 ;
        RECT 99.12 -3.56 99.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -91.285 99.445 -90.955 ;
        RECT 99.115 -92.645 99.445 -92.315 ;
        RECT 99.115 -94.005 99.445 -93.675 ;
        RECT 99.115 -95.365 99.445 -95.035 ;
        RECT 99.115 -96.725 99.445 -96.395 ;
        RECT 99.115 -98.085 99.445 -97.755 ;
        RECT 99.115 -99.445 99.445 -99.115 ;
        RECT 99.115 -100.805 99.445 -100.475 ;
        RECT 99.115 -102.165 99.445 -101.835 ;
        RECT 99.115 -103.525 99.445 -103.195 ;
        RECT 99.115 -104.885 99.445 -104.555 ;
        RECT 99.115 -106.245 99.445 -105.915 ;
        RECT 99.115 -107.605 99.445 -107.275 ;
        RECT 99.115 -108.965 99.445 -108.635 ;
        RECT 99.115 -110.325 99.445 -109.995 ;
        RECT 99.115 -111.685 99.445 -111.355 ;
        RECT 99.115 -113.045 99.445 -112.715 ;
        RECT 99.115 -114.405 99.445 -114.075 ;
        RECT 99.115 -115.765 99.445 -115.435 ;
        RECT 99.115 -117.125 99.445 -116.795 ;
        RECT 99.115 -118.485 99.445 -118.155 ;
        RECT 99.115 -119.845 99.445 -119.515 ;
        RECT 99.115 -121.205 99.445 -120.875 ;
        RECT 99.115 -122.565 99.445 -122.235 ;
        RECT 99.115 -123.925 99.445 -123.595 ;
        RECT 99.115 -125.285 99.445 -124.955 ;
        RECT 99.115 -126.645 99.445 -126.315 ;
        RECT 99.115 -128.005 99.445 -127.675 ;
        RECT 99.115 -129.365 99.445 -129.035 ;
        RECT 99.115 -130.725 99.445 -130.395 ;
        RECT 99.115 -132.085 99.445 -131.755 ;
        RECT 99.115 -133.445 99.445 -133.115 ;
        RECT 99.115 -134.805 99.445 -134.475 ;
        RECT 99.115 -136.165 99.445 -135.835 ;
        RECT 99.115 -137.525 99.445 -137.195 ;
        RECT 99.115 -138.885 99.445 -138.555 ;
        RECT 99.115 -140.245 99.445 -139.915 ;
        RECT 99.115 -141.605 99.445 -141.275 ;
        RECT 99.115 -142.965 99.445 -142.635 ;
        RECT 99.115 -144.325 99.445 -143.995 ;
        RECT 99.115 -145.685 99.445 -145.355 ;
        RECT 99.115 -147.045 99.445 -146.715 ;
        RECT 99.115 -148.405 99.445 -148.075 ;
        RECT 99.115 -149.765 99.445 -149.435 ;
        RECT 99.115 -151.125 99.445 -150.795 ;
        RECT 99.115 -152.485 99.445 -152.155 ;
        RECT 99.115 -153.845 99.445 -153.515 ;
        RECT 99.115 -155.205 99.445 -154.875 ;
        RECT 99.115 -156.565 99.445 -156.235 ;
        RECT 99.115 -157.925 99.445 -157.595 ;
        RECT 99.115 -160.17 99.445 -159.04 ;
        RECT 99.12 -160.285 99.44 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 127.225 100.805 128.355 ;
        RECT 100.475 124.955 100.805 125.285 ;
        RECT 100.475 123.595 100.805 123.925 ;
        RECT 100.48 123.595 100.8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 -95.365 100.805 -95.035 ;
        RECT 100.475 -96.725 100.805 -96.395 ;
        RECT 100.475 -98.085 100.805 -97.755 ;
        RECT 100.475 -99.445 100.805 -99.115 ;
        RECT 100.475 -100.805 100.805 -100.475 ;
        RECT 100.475 -102.165 100.805 -101.835 ;
        RECT 100.475 -103.525 100.805 -103.195 ;
        RECT 100.475 -104.885 100.805 -104.555 ;
        RECT 100.475 -106.245 100.805 -105.915 ;
        RECT 100.475 -107.605 100.805 -107.275 ;
        RECT 100.475 -108.965 100.805 -108.635 ;
        RECT 100.475 -110.325 100.805 -109.995 ;
        RECT 100.475 -111.685 100.805 -111.355 ;
        RECT 100.475 -113.045 100.805 -112.715 ;
        RECT 100.475 -114.405 100.805 -114.075 ;
        RECT 100.475 -115.765 100.805 -115.435 ;
        RECT 100.475 -117.125 100.805 -116.795 ;
        RECT 100.475 -118.485 100.805 -118.155 ;
        RECT 100.475 -119.845 100.805 -119.515 ;
        RECT 100.475 -121.205 100.805 -120.875 ;
        RECT 100.475 -122.565 100.805 -122.235 ;
        RECT 100.475 -123.925 100.805 -123.595 ;
        RECT 100.475 -125.285 100.805 -124.955 ;
        RECT 100.475 -126.645 100.805 -126.315 ;
        RECT 100.475 -128.005 100.805 -127.675 ;
        RECT 100.475 -129.365 100.805 -129.035 ;
        RECT 100.475 -130.725 100.805 -130.395 ;
        RECT 100.475 -132.085 100.805 -131.755 ;
        RECT 100.475 -133.445 100.805 -133.115 ;
        RECT 100.475 -134.805 100.805 -134.475 ;
        RECT 100.475 -136.165 100.805 -135.835 ;
        RECT 100.475 -137.525 100.805 -137.195 ;
        RECT 100.475 -138.885 100.805 -138.555 ;
        RECT 100.475 -140.245 100.805 -139.915 ;
        RECT 100.475 -141.605 100.805 -141.275 ;
        RECT 100.475 -142.965 100.805 -142.635 ;
        RECT 100.475 -144.325 100.805 -143.995 ;
        RECT 100.475 -145.685 100.805 -145.355 ;
        RECT 100.475 -147.045 100.805 -146.715 ;
        RECT 100.475 -148.405 100.805 -148.075 ;
        RECT 100.475 -149.765 100.805 -149.435 ;
        RECT 100.475 -151.125 100.805 -150.795 ;
        RECT 100.475 -152.485 100.805 -152.155 ;
        RECT 100.475 -153.845 100.805 -153.515 ;
        RECT 100.475 -155.205 100.805 -154.875 ;
        RECT 100.475 -156.565 100.805 -156.235 ;
        RECT 100.475 -157.925 100.805 -157.595 ;
        RECT 100.475 -160.17 100.805 -159.04 ;
        RECT 100.48 -160.285 100.8 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.91 -94.075 101.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 127.225 102.165 128.355 ;
        RECT 101.835 124.955 102.165 125.285 ;
        RECT 101.835 123.595 102.165 123.925 ;
        RECT 101.84 123.595 102.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 -1.525 102.165 -1.195 ;
        RECT 101.835 -2.885 102.165 -2.555 ;
        RECT 101.84 -3.56 102.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 127.225 103.525 128.355 ;
        RECT 103.195 124.955 103.525 125.285 ;
        RECT 103.195 123.595 103.525 123.925 ;
        RECT 103.2 123.595 103.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 -1.525 103.525 -1.195 ;
        RECT 103.195 -2.885 103.525 -2.555 ;
        RECT 103.2 -3.56 103.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 127.225 104.885 128.355 ;
        RECT 104.555 124.955 104.885 125.285 ;
        RECT 104.555 123.595 104.885 123.925 ;
        RECT 104.56 123.595 104.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 -1.525 104.885 -1.195 ;
        RECT 104.555 -2.885 104.885 -2.555 ;
        RECT 104.56 -3.56 104.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 127.225 106.245 128.355 ;
        RECT 105.915 124.955 106.245 125.285 ;
        RECT 105.915 123.595 106.245 123.925 ;
        RECT 105.92 123.595 106.24 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 -95.365 106.245 -95.035 ;
        RECT 105.915 -96.725 106.245 -96.395 ;
        RECT 105.915 -98.085 106.245 -97.755 ;
        RECT 105.915 -99.445 106.245 -99.115 ;
        RECT 105.915 -100.805 106.245 -100.475 ;
        RECT 105.915 -102.165 106.245 -101.835 ;
        RECT 105.915 -103.525 106.245 -103.195 ;
        RECT 105.915 -104.885 106.245 -104.555 ;
        RECT 105.915 -106.245 106.245 -105.915 ;
        RECT 105.915 -107.605 106.245 -107.275 ;
        RECT 105.915 -108.965 106.245 -108.635 ;
        RECT 105.915 -110.325 106.245 -109.995 ;
        RECT 105.915 -111.685 106.245 -111.355 ;
        RECT 105.915 -113.045 106.245 -112.715 ;
        RECT 105.915 -114.405 106.245 -114.075 ;
        RECT 105.915 -115.765 106.245 -115.435 ;
        RECT 105.915 -117.125 106.245 -116.795 ;
        RECT 105.915 -118.485 106.245 -118.155 ;
        RECT 105.915 -119.845 106.245 -119.515 ;
        RECT 105.915 -121.205 106.245 -120.875 ;
        RECT 105.915 -122.565 106.245 -122.235 ;
        RECT 105.915 -123.925 106.245 -123.595 ;
        RECT 105.915 -125.285 106.245 -124.955 ;
        RECT 105.915 -126.645 106.245 -126.315 ;
        RECT 105.915 -128.005 106.245 -127.675 ;
        RECT 105.915 -129.365 106.245 -129.035 ;
        RECT 105.915 -130.725 106.245 -130.395 ;
        RECT 105.915 -132.085 106.245 -131.755 ;
        RECT 105.915 -133.445 106.245 -133.115 ;
        RECT 105.915 -134.805 106.245 -134.475 ;
        RECT 105.915 -136.165 106.245 -135.835 ;
        RECT 105.915 -137.525 106.245 -137.195 ;
        RECT 105.915 -138.885 106.245 -138.555 ;
        RECT 105.915 -140.245 106.245 -139.915 ;
        RECT 105.915 -141.605 106.245 -141.275 ;
        RECT 105.915 -142.965 106.245 -142.635 ;
        RECT 105.915 -144.325 106.245 -143.995 ;
        RECT 105.915 -145.685 106.245 -145.355 ;
        RECT 105.915 -147.045 106.245 -146.715 ;
        RECT 105.915 -148.405 106.245 -148.075 ;
        RECT 105.915 -149.765 106.245 -149.435 ;
        RECT 105.915 -151.125 106.245 -150.795 ;
        RECT 105.915 -152.485 106.245 -152.155 ;
        RECT 105.915 -153.845 106.245 -153.515 ;
        RECT 105.915 -155.205 106.245 -154.875 ;
        RECT 105.915 -156.565 106.245 -156.235 ;
        RECT 105.915 -157.925 106.245 -157.595 ;
        RECT 105.915 -160.17 106.245 -159.04 ;
        RECT 105.92 -160.285 106.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.01 -94.075 107.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 127.225 107.605 128.355 ;
        RECT 107.275 124.955 107.605 125.285 ;
        RECT 107.275 123.595 107.605 123.925 ;
        RECT 107.28 123.595 107.6 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 127.225 108.965 128.355 ;
        RECT 108.635 124.955 108.965 125.285 ;
        RECT 108.635 123.595 108.965 123.925 ;
        RECT 108.64 123.595 108.96 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 -1.525 108.965 -1.195 ;
        RECT 108.635 -2.885 108.965 -2.555 ;
        RECT 108.64 -3.56 108.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 127.225 110.325 128.355 ;
        RECT 109.995 124.955 110.325 125.285 ;
        RECT 109.995 123.595 110.325 123.925 ;
        RECT 110 123.595 110.32 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 -1.525 110.325 -1.195 ;
        RECT 109.995 -2.885 110.325 -2.555 ;
        RECT 110 -3.56 110.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 127.225 111.685 128.355 ;
        RECT 111.355 124.955 111.685 125.285 ;
        RECT 111.355 123.595 111.685 123.925 ;
        RECT 111.36 123.595 111.68 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 -1.525 111.685 -1.195 ;
        RECT 111.355 -2.885 111.685 -2.555 ;
        RECT 111.36 -3.56 111.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 -91.285 111.685 -90.955 ;
        RECT 111.355 -92.645 111.685 -92.315 ;
        RECT 111.355 -94.005 111.685 -93.675 ;
        RECT 111.355 -95.365 111.685 -95.035 ;
        RECT 111.355 -96.725 111.685 -96.395 ;
        RECT 111.355 -98.085 111.685 -97.755 ;
        RECT 111.355 -99.445 111.685 -99.115 ;
        RECT 111.355 -100.805 111.685 -100.475 ;
        RECT 111.355 -102.165 111.685 -101.835 ;
        RECT 111.355 -103.525 111.685 -103.195 ;
        RECT 111.355 -104.885 111.685 -104.555 ;
        RECT 111.355 -106.245 111.685 -105.915 ;
        RECT 111.355 -107.605 111.685 -107.275 ;
        RECT 111.355 -108.965 111.685 -108.635 ;
        RECT 111.355 -110.325 111.685 -109.995 ;
        RECT 111.355 -111.685 111.685 -111.355 ;
        RECT 111.355 -113.045 111.685 -112.715 ;
        RECT 111.355 -114.405 111.685 -114.075 ;
        RECT 111.355 -115.765 111.685 -115.435 ;
        RECT 111.355 -117.125 111.685 -116.795 ;
        RECT 111.355 -118.485 111.685 -118.155 ;
        RECT 111.355 -119.845 111.685 -119.515 ;
        RECT 111.355 -121.205 111.685 -120.875 ;
        RECT 111.355 -122.565 111.685 -122.235 ;
        RECT 111.355 -123.925 111.685 -123.595 ;
        RECT 111.355 -125.285 111.685 -124.955 ;
        RECT 111.355 -126.645 111.685 -126.315 ;
        RECT 111.355 -128.005 111.685 -127.675 ;
        RECT 111.355 -129.365 111.685 -129.035 ;
        RECT 111.355 -130.725 111.685 -130.395 ;
        RECT 111.355 -132.085 111.685 -131.755 ;
        RECT 111.355 -133.445 111.685 -133.115 ;
        RECT 111.355 -134.805 111.685 -134.475 ;
        RECT 111.355 -136.165 111.685 -135.835 ;
        RECT 111.355 -137.525 111.685 -137.195 ;
        RECT 111.355 -138.885 111.685 -138.555 ;
        RECT 111.355 -140.245 111.685 -139.915 ;
        RECT 111.355 -141.605 111.685 -141.275 ;
        RECT 111.355 -142.965 111.685 -142.635 ;
        RECT 111.355 -144.325 111.685 -143.995 ;
        RECT 111.355 -145.685 111.685 -145.355 ;
        RECT 111.355 -147.045 111.685 -146.715 ;
        RECT 111.355 -148.405 111.685 -148.075 ;
        RECT 111.355 -149.765 111.685 -149.435 ;
        RECT 111.355 -151.125 111.685 -150.795 ;
        RECT 111.355 -152.485 111.685 -152.155 ;
        RECT 111.355 -153.845 111.685 -153.515 ;
        RECT 111.355 -155.205 111.685 -154.875 ;
        RECT 111.355 -156.565 111.685 -156.235 ;
        RECT 111.355 -157.925 111.685 -157.595 ;
        RECT 111.355 -160.17 111.685 -159.04 ;
        RECT 111.36 -160.285 111.68 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 127.225 113.045 128.355 ;
        RECT 112.715 124.955 113.045 125.285 ;
        RECT 112.715 123.595 113.045 123.925 ;
        RECT 112.72 123.595 113.04 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 -126.645 113.045 -126.315 ;
        RECT 112.715 -128.005 113.045 -127.675 ;
        RECT 112.715 -129.365 113.045 -129.035 ;
        RECT 112.715 -130.725 113.045 -130.395 ;
        RECT 112.715 -132.085 113.045 -131.755 ;
        RECT 112.715 -133.445 113.045 -133.115 ;
        RECT 112.715 -134.805 113.045 -134.475 ;
        RECT 112.715 -136.165 113.045 -135.835 ;
        RECT 112.715 -137.525 113.045 -137.195 ;
        RECT 112.715 -138.885 113.045 -138.555 ;
        RECT 112.715 -140.245 113.045 -139.915 ;
        RECT 112.715 -141.605 113.045 -141.275 ;
        RECT 112.715 -142.965 113.045 -142.635 ;
        RECT 112.715 -144.325 113.045 -143.995 ;
        RECT 112.715 -145.685 113.045 -145.355 ;
        RECT 112.715 -147.045 113.045 -146.715 ;
        RECT 112.715 -148.405 113.045 -148.075 ;
        RECT 112.715 -149.765 113.045 -149.435 ;
        RECT 112.715 -151.125 113.045 -150.795 ;
        RECT 112.715 -152.485 113.045 -152.155 ;
        RECT 112.715 -153.845 113.045 -153.515 ;
        RECT 112.715 -155.205 113.045 -154.875 ;
        RECT 112.715 -156.565 113.045 -156.235 ;
        RECT 112.715 -157.925 113.045 -157.595 ;
        RECT 112.715 -160.17 113.045 -159.04 ;
        RECT 112.72 -160.285 113.04 -95.035 ;
        RECT 112.715 -95.365 113.045 -95.035 ;
        RECT 112.715 -96.725 113.045 -96.395 ;
        RECT 112.715 -98.085 113.045 -97.755 ;
        RECT 112.715 -99.445 113.045 -99.115 ;
        RECT 112.715 -100.805 113.045 -100.475 ;
        RECT 112.715 -102.165 113.045 -101.835 ;
        RECT 112.715 -103.525 113.045 -103.195 ;
        RECT 112.715 -104.885 113.045 -104.555 ;
        RECT 112.715 -106.245 113.045 -105.915 ;
        RECT 112.715 -107.605 113.045 -107.275 ;
        RECT 112.715 -108.965 113.045 -108.635 ;
        RECT 112.715 -110.325 113.045 -109.995 ;
        RECT 112.715 -111.685 113.045 -111.355 ;
        RECT 112.715 -113.045 113.045 -112.715 ;
        RECT 112.715 -114.405 113.045 -114.075 ;
        RECT 112.715 -115.765 113.045 -115.435 ;
        RECT 112.715 -117.125 113.045 -116.795 ;
        RECT 112.715 -118.485 113.045 -118.155 ;
        RECT 112.715 -119.845 113.045 -119.515 ;
        RECT 112.715 -121.205 113.045 -120.875 ;
        RECT 112.715 -122.565 113.045 -122.235 ;
        RECT 112.715 -123.925 113.045 -123.595 ;
        RECT 112.715 -125.285 113.045 -124.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 -91.285 26.005 -90.955 ;
        RECT 25.675 -92.645 26.005 -92.315 ;
        RECT 25.675 -94.005 26.005 -93.675 ;
        RECT 25.675 -95.365 26.005 -95.035 ;
        RECT 25.675 -96.725 26.005 -96.395 ;
        RECT 25.675 -98.085 26.005 -97.755 ;
        RECT 25.675 -99.445 26.005 -99.115 ;
        RECT 25.675 -100.805 26.005 -100.475 ;
        RECT 25.675 -102.165 26.005 -101.835 ;
        RECT 25.675 -103.525 26.005 -103.195 ;
        RECT 25.675 -104.885 26.005 -104.555 ;
        RECT 25.675 -106.245 26.005 -105.915 ;
        RECT 25.675 -107.605 26.005 -107.275 ;
        RECT 25.675 -108.965 26.005 -108.635 ;
        RECT 25.675 -110.325 26.005 -109.995 ;
        RECT 25.675 -111.685 26.005 -111.355 ;
        RECT 25.675 -113.045 26.005 -112.715 ;
        RECT 25.675 -114.405 26.005 -114.075 ;
        RECT 25.675 -115.765 26.005 -115.435 ;
        RECT 25.675 -117.125 26.005 -116.795 ;
        RECT 25.675 -118.485 26.005 -118.155 ;
        RECT 25.675 -119.845 26.005 -119.515 ;
        RECT 25.675 -121.205 26.005 -120.875 ;
        RECT 25.675 -122.565 26.005 -122.235 ;
        RECT 25.675 -123.925 26.005 -123.595 ;
        RECT 25.675 -125.285 26.005 -124.955 ;
        RECT 25.675 -126.645 26.005 -126.315 ;
        RECT 25.675 -128.005 26.005 -127.675 ;
        RECT 25.675 -129.365 26.005 -129.035 ;
        RECT 25.675 -130.725 26.005 -130.395 ;
        RECT 25.675 -132.085 26.005 -131.755 ;
        RECT 25.675 -133.445 26.005 -133.115 ;
        RECT 25.675 -134.805 26.005 -134.475 ;
        RECT 25.675 -136.165 26.005 -135.835 ;
        RECT 25.675 -137.525 26.005 -137.195 ;
        RECT 25.675 -138.885 26.005 -138.555 ;
        RECT 25.675 -140.245 26.005 -139.915 ;
        RECT 25.675 -141.605 26.005 -141.275 ;
        RECT 25.675 -142.965 26.005 -142.635 ;
        RECT 25.675 -144.325 26.005 -143.995 ;
        RECT 25.675 -145.685 26.005 -145.355 ;
        RECT 25.675 -147.045 26.005 -146.715 ;
        RECT 25.675 -148.405 26.005 -148.075 ;
        RECT 25.675 -149.765 26.005 -149.435 ;
        RECT 25.675 -151.125 26.005 -150.795 ;
        RECT 25.675 -152.485 26.005 -152.155 ;
        RECT 25.675 -153.845 26.005 -153.515 ;
        RECT 25.675 -155.205 26.005 -154.875 ;
        RECT 25.675 -156.565 26.005 -156.235 ;
        RECT 25.675 -157.925 26.005 -157.595 ;
        RECT 25.675 -160.17 26.005 -159.04 ;
        RECT 25.68 -160.285 26 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 127.225 27.365 128.355 ;
        RECT 27.035 124.955 27.365 125.285 ;
        RECT 27.035 123.595 27.365 123.925 ;
        RECT 27.04 123.595 27.36 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 -95.365 27.365 -95.035 ;
        RECT 27.035 -96.725 27.365 -96.395 ;
        RECT 27.035 -98.085 27.365 -97.755 ;
        RECT 27.035 -99.445 27.365 -99.115 ;
        RECT 27.035 -100.805 27.365 -100.475 ;
        RECT 27.035 -102.165 27.365 -101.835 ;
        RECT 27.035 -103.525 27.365 -103.195 ;
        RECT 27.035 -104.885 27.365 -104.555 ;
        RECT 27.035 -106.245 27.365 -105.915 ;
        RECT 27.035 -107.605 27.365 -107.275 ;
        RECT 27.035 -108.965 27.365 -108.635 ;
        RECT 27.035 -110.325 27.365 -109.995 ;
        RECT 27.035 -111.685 27.365 -111.355 ;
        RECT 27.035 -113.045 27.365 -112.715 ;
        RECT 27.035 -114.405 27.365 -114.075 ;
        RECT 27.035 -115.765 27.365 -115.435 ;
        RECT 27.035 -117.125 27.365 -116.795 ;
        RECT 27.035 -118.485 27.365 -118.155 ;
        RECT 27.035 -119.845 27.365 -119.515 ;
        RECT 27.035 -121.205 27.365 -120.875 ;
        RECT 27.035 -122.565 27.365 -122.235 ;
        RECT 27.035 -123.925 27.365 -123.595 ;
        RECT 27.035 -125.285 27.365 -124.955 ;
        RECT 27.035 -126.645 27.365 -126.315 ;
        RECT 27.035 -128.005 27.365 -127.675 ;
        RECT 27.035 -129.365 27.365 -129.035 ;
        RECT 27.035 -130.725 27.365 -130.395 ;
        RECT 27.035 -132.085 27.365 -131.755 ;
        RECT 27.035 -133.445 27.365 -133.115 ;
        RECT 27.035 -134.805 27.365 -134.475 ;
        RECT 27.035 -136.165 27.365 -135.835 ;
        RECT 27.035 -137.525 27.365 -137.195 ;
        RECT 27.035 -138.885 27.365 -138.555 ;
        RECT 27.035 -140.245 27.365 -139.915 ;
        RECT 27.035 -141.605 27.365 -141.275 ;
        RECT 27.035 -142.965 27.365 -142.635 ;
        RECT 27.035 -144.325 27.365 -143.995 ;
        RECT 27.035 -145.685 27.365 -145.355 ;
        RECT 27.035 -147.045 27.365 -146.715 ;
        RECT 27.035 -148.405 27.365 -148.075 ;
        RECT 27.035 -149.765 27.365 -149.435 ;
        RECT 27.035 -151.125 27.365 -150.795 ;
        RECT 27.035 -152.485 27.365 -152.155 ;
        RECT 27.035 -153.845 27.365 -153.515 ;
        RECT 27.035 -155.205 27.365 -154.875 ;
        RECT 27.035 -156.565 27.365 -156.235 ;
        RECT 27.035 -157.925 27.365 -157.595 ;
        RECT 27.035 -160.17 27.365 -159.04 ;
        RECT 27.04 -160.285 27.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.71 -94.075 28.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 127.225 28.725 128.355 ;
        RECT 28.395 124.955 28.725 125.285 ;
        RECT 28.395 123.595 28.725 123.925 ;
        RECT 28.4 123.595 28.72 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -1.525 28.725 -1.195 ;
        RECT 28.395 -2.885 28.725 -2.555 ;
        RECT 28.4 -3.56 28.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 127.225 30.085 128.355 ;
        RECT 29.755 124.955 30.085 125.285 ;
        RECT 29.755 123.595 30.085 123.925 ;
        RECT 29.76 123.595 30.08 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -1.525 30.085 -1.195 ;
        RECT 29.755 -2.885 30.085 -2.555 ;
        RECT 29.76 -3.56 30.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 127.225 31.445 128.355 ;
        RECT 31.115 124.955 31.445 125.285 ;
        RECT 31.115 123.595 31.445 123.925 ;
        RECT 31.12 123.595 31.44 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -1.525 31.445 -1.195 ;
        RECT 31.115 -2.885 31.445 -2.555 ;
        RECT 31.12 -3.56 31.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -91.285 31.445 -90.955 ;
        RECT 31.115 -92.645 31.445 -92.315 ;
        RECT 31.115 -94.005 31.445 -93.675 ;
        RECT 31.115 -95.365 31.445 -95.035 ;
        RECT 31.115 -96.725 31.445 -96.395 ;
        RECT 31.115 -98.085 31.445 -97.755 ;
        RECT 31.115 -99.445 31.445 -99.115 ;
        RECT 31.115 -100.805 31.445 -100.475 ;
        RECT 31.115 -102.165 31.445 -101.835 ;
        RECT 31.115 -103.525 31.445 -103.195 ;
        RECT 31.115 -104.885 31.445 -104.555 ;
        RECT 31.115 -106.245 31.445 -105.915 ;
        RECT 31.115 -107.605 31.445 -107.275 ;
        RECT 31.115 -108.965 31.445 -108.635 ;
        RECT 31.115 -110.325 31.445 -109.995 ;
        RECT 31.115 -111.685 31.445 -111.355 ;
        RECT 31.115 -113.045 31.445 -112.715 ;
        RECT 31.115 -114.405 31.445 -114.075 ;
        RECT 31.115 -115.765 31.445 -115.435 ;
        RECT 31.115 -117.125 31.445 -116.795 ;
        RECT 31.115 -118.485 31.445 -118.155 ;
        RECT 31.115 -119.845 31.445 -119.515 ;
        RECT 31.115 -121.205 31.445 -120.875 ;
        RECT 31.115 -122.565 31.445 -122.235 ;
        RECT 31.115 -123.925 31.445 -123.595 ;
        RECT 31.115 -125.285 31.445 -124.955 ;
        RECT 31.115 -126.645 31.445 -126.315 ;
        RECT 31.115 -128.005 31.445 -127.675 ;
        RECT 31.115 -129.365 31.445 -129.035 ;
        RECT 31.115 -130.725 31.445 -130.395 ;
        RECT 31.115 -132.085 31.445 -131.755 ;
        RECT 31.115 -133.445 31.445 -133.115 ;
        RECT 31.115 -134.805 31.445 -134.475 ;
        RECT 31.115 -136.165 31.445 -135.835 ;
        RECT 31.115 -137.525 31.445 -137.195 ;
        RECT 31.115 -138.885 31.445 -138.555 ;
        RECT 31.115 -140.245 31.445 -139.915 ;
        RECT 31.115 -141.605 31.445 -141.275 ;
        RECT 31.115 -142.965 31.445 -142.635 ;
        RECT 31.115 -144.325 31.445 -143.995 ;
        RECT 31.115 -145.685 31.445 -145.355 ;
        RECT 31.115 -147.045 31.445 -146.715 ;
        RECT 31.115 -148.405 31.445 -148.075 ;
        RECT 31.115 -149.765 31.445 -149.435 ;
        RECT 31.115 -151.125 31.445 -150.795 ;
        RECT 31.115 -152.485 31.445 -152.155 ;
        RECT 31.115 -153.845 31.445 -153.515 ;
        RECT 31.115 -155.205 31.445 -154.875 ;
        RECT 31.115 -156.565 31.445 -156.235 ;
        RECT 31.115 -157.925 31.445 -157.595 ;
        RECT 31.115 -160.17 31.445 -159.04 ;
        RECT 31.12 -160.285 31.44 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 127.225 32.805 128.355 ;
        RECT 32.475 124.955 32.805 125.285 ;
        RECT 32.475 123.595 32.805 123.925 ;
        RECT 32.48 123.595 32.8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -1.525 32.805 -1.195 ;
        RECT 32.475 -2.885 32.805 -2.555 ;
        RECT 32.48 -3.56 32.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -91.285 32.805 -90.955 ;
        RECT 32.475 -92.645 32.805 -92.315 ;
        RECT 32.475 -94.005 32.805 -93.675 ;
        RECT 32.475 -95.365 32.805 -95.035 ;
        RECT 32.475 -96.725 32.805 -96.395 ;
        RECT 32.475 -98.085 32.805 -97.755 ;
        RECT 32.475 -99.445 32.805 -99.115 ;
        RECT 32.475 -100.805 32.805 -100.475 ;
        RECT 32.475 -102.165 32.805 -101.835 ;
        RECT 32.475 -103.525 32.805 -103.195 ;
        RECT 32.475 -104.885 32.805 -104.555 ;
        RECT 32.475 -106.245 32.805 -105.915 ;
        RECT 32.475 -107.605 32.805 -107.275 ;
        RECT 32.475 -108.965 32.805 -108.635 ;
        RECT 32.475 -110.325 32.805 -109.995 ;
        RECT 32.475 -111.685 32.805 -111.355 ;
        RECT 32.475 -113.045 32.805 -112.715 ;
        RECT 32.475 -114.405 32.805 -114.075 ;
        RECT 32.475 -115.765 32.805 -115.435 ;
        RECT 32.475 -117.125 32.805 -116.795 ;
        RECT 32.475 -118.485 32.805 -118.155 ;
        RECT 32.475 -119.845 32.805 -119.515 ;
        RECT 32.475 -121.205 32.805 -120.875 ;
        RECT 32.475 -122.565 32.805 -122.235 ;
        RECT 32.475 -123.925 32.805 -123.595 ;
        RECT 32.475 -125.285 32.805 -124.955 ;
        RECT 32.475 -126.645 32.805 -126.315 ;
        RECT 32.475 -128.005 32.805 -127.675 ;
        RECT 32.475 -129.365 32.805 -129.035 ;
        RECT 32.475 -130.725 32.805 -130.395 ;
        RECT 32.475 -132.085 32.805 -131.755 ;
        RECT 32.475 -133.445 32.805 -133.115 ;
        RECT 32.475 -134.805 32.805 -134.475 ;
        RECT 32.475 -136.165 32.805 -135.835 ;
        RECT 32.475 -137.525 32.805 -137.195 ;
        RECT 32.475 -138.885 32.805 -138.555 ;
        RECT 32.475 -140.245 32.805 -139.915 ;
        RECT 32.475 -141.605 32.805 -141.275 ;
        RECT 32.475 -142.965 32.805 -142.635 ;
        RECT 32.475 -144.325 32.805 -143.995 ;
        RECT 32.475 -145.685 32.805 -145.355 ;
        RECT 32.475 -147.045 32.805 -146.715 ;
        RECT 32.475 -148.405 32.805 -148.075 ;
        RECT 32.475 -149.765 32.805 -149.435 ;
        RECT 32.475 -151.125 32.805 -150.795 ;
        RECT 32.475 -152.485 32.805 -152.155 ;
        RECT 32.475 -153.845 32.805 -153.515 ;
        RECT 32.475 -155.205 32.805 -154.875 ;
        RECT 32.475 -156.565 32.805 -156.235 ;
        RECT 32.475 -157.925 32.805 -157.595 ;
        RECT 32.475 -160.17 32.805 -159.04 ;
        RECT 32.48 -160.285 32.8 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.81 -94.075 34.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 127.225 34.165 128.355 ;
        RECT 33.835 124.955 34.165 125.285 ;
        RECT 33.835 123.595 34.165 123.925 ;
        RECT 33.84 123.595 34.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 127.225 35.525 128.355 ;
        RECT 35.195 124.955 35.525 125.285 ;
        RECT 35.195 123.595 35.525 123.925 ;
        RECT 35.2 123.595 35.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 -1.525 35.525 -1.195 ;
        RECT 35.195 -2.885 35.525 -2.555 ;
        RECT 35.2 -3.56 35.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 127.225 36.885 128.355 ;
        RECT 36.555 124.955 36.885 125.285 ;
        RECT 36.555 123.595 36.885 123.925 ;
        RECT 36.56 123.595 36.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 -1.525 36.885 -1.195 ;
        RECT 36.555 -2.885 36.885 -2.555 ;
        RECT 36.56 -3.56 36.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 127.225 38.245 128.355 ;
        RECT 37.915 124.955 38.245 125.285 ;
        RECT 37.915 123.595 38.245 123.925 ;
        RECT 37.92 123.595 38.24 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 -1.525 38.245 -1.195 ;
        RECT 37.915 -2.885 38.245 -2.555 ;
        RECT 37.92 -3.56 38.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 -91.285 38.245 -90.955 ;
        RECT 37.915 -92.645 38.245 -92.315 ;
        RECT 37.915 -94.005 38.245 -93.675 ;
        RECT 37.915 -95.365 38.245 -95.035 ;
        RECT 37.915 -96.725 38.245 -96.395 ;
        RECT 37.915 -98.085 38.245 -97.755 ;
        RECT 37.915 -99.445 38.245 -99.115 ;
        RECT 37.915 -100.805 38.245 -100.475 ;
        RECT 37.915 -102.165 38.245 -101.835 ;
        RECT 37.915 -103.525 38.245 -103.195 ;
        RECT 37.915 -104.885 38.245 -104.555 ;
        RECT 37.915 -106.245 38.245 -105.915 ;
        RECT 37.915 -107.605 38.245 -107.275 ;
        RECT 37.915 -108.965 38.245 -108.635 ;
        RECT 37.915 -110.325 38.245 -109.995 ;
        RECT 37.915 -111.685 38.245 -111.355 ;
        RECT 37.915 -113.045 38.245 -112.715 ;
        RECT 37.915 -114.405 38.245 -114.075 ;
        RECT 37.915 -115.765 38.245 -115.435 ;
        RECT 37.915 -117.125 38.245 -116.795 ;
        RECT 37.915 -118.485 38.245 -118.155 ;
        RECT 37.915 -119.845 38.245 -119.515 ;
        RECT 37.915 -121.205 38.245 -120.875 ;
        RECT 37.915 -122.565 38.245 -122.235 ;
        RECT 37.915 -123.925 38.245 -123.595 ;
        RECT 37.915 -125.285 38.245 -124.955 ;
        RECT 37.915 -126.645 38.245 -126.315 ;
        RECT 37.915 -128.005 38.245 -127.675 ;
        RECT 37.915 -129.365 38.245 -129.035 ;
        RECT 37.915 -130.725 38.245 -130.395 ;
        RECT 37.915 -132.085 38.245 -131.755 ;
        RECT 37.915 -133.445 38.245 -133.115 ;
        RECT 37.915 -134.805 38.245 -134.475 ;
        RECT 37.915 -136.165 38.245 -135.835 ;
        RECT 37.915 -137.525 38.245 -137.195 ;
        RECT 37.915 -138.885 38.245 -138.555 ;
        RECT 37.915 -140.245 38.245 -139.915 ;
        RECT 37.915 -141.605 38.245 -141.275 ;
        RECT 37.915 -142.965 38.245 -142.635 ;
        RECT 37.915 -144.325 38.245 -143.995 ;
        RECT 37.915 -145.685 38.245 -145.355 ;
        RECT 37.915 -147.045 38.245 -146.715 ;
        RECT 37.915 -148.405 38.245 -148.075 ;
        RECT 37.915 -149.765 38.245 -149.435 ;
        RECT 37.915 -151.125 38.245 -150.795 ;
        RECT 37.915 -152.485 38.245 -152.155 ;
        RECT 37.915 -153.845 38.245 -153.515 ;
        RECT 37.915 -155.205 38.245 -154.875 ;
        RECT 37.915 -156.565 38.245 -156.235 ;
        RECT 37.915 -157.925 38.245 -157.595 ;
        RECT 37.915 -160.17 38.245 -159.04 ;
        RECT 37.92 -160.285 38.24 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 127.225 39.605 128.355 ;
        RECT 39.275 124.955 39.605 125.285 ;
        RECT 39.275 123.595 39.605 123.925 ;
        RECT 39.28 123.595 39.6 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 -95.365 39.605 -95.035 ;
        RECT 39.275 -96.725 39.605 -96.395 ;
        RECT 39.275 -98.085 39.605 -97.755 ;
        RECT 39.275 -99.445 39.605 -99.115 ;
        RECT 39.275 -100.805 39.605 -100.475 ;
        RECT 39.275 -102.165 39.605 -101.835 ;
        RECT 39.275 -103.525 39.605 -103.195 ;
        RECT 39.275 -104.885 39.605 -104.555 ;
        RECT 39.275 -106.245 39.605 -105.915 ;
        RECT 39.275 -107.605 39.605 -107.275 ;
        RECT 39.275 -108.965 39.605 -108.635 ;
        RECT 39.275 -110.325 39.605 -109.995 ;
        RECT 39.275 -111.685 39.605 -111.355 ;
        RECT 39.275 -113.045 39.605 -112.715 ;
        RECT 39.275 -114.405 39.605 -114.075 ;
        RECT 39.275 -115.765 39.605 -115.435 ;
        RECT 39.275 -117.125 39.605 -116.795 ;
        RECT 39.275 -118.485 39.605 -118.155 ;
        RECT 39.275 -119.845 39.605 -119.515 ;
        RECT 39.275 -121.205 39.605 -120.875 ;
        RECT 39.275 -122.565 39.605 -122.235 ;
        RECT 39.275 -123.925 39.605 -123.595 ;
        RECT 39.275 -125.285 39.605 -124.955 ;
        RECT 39.275 -126.645 39.605 -126.315 ;
        RECT 39.275 -128.005 39.605 -127.675 ;
        RECT 39.275 -129.365 39.605 -129.035 ;
        RECT 39.275 -130.725 39.605 -130.395 ;
        RECT 39.275 -132.085 39.605 -131.755 ;
        RECT 39.275 -133.445 39.605 -133.115 ;
        RECT 39.275 -134.805 39.605 -134.475 ;
        RECT 39.275 -136.165 39.605 -135.835 ;
        RECT 39.275 -137.525 39.605 -137.195 ;
        RECT 39.275 -138.885 39.605 -138.555 ;
        RECT 39.275 -140.245 39.605 -139.915 ;
        RECT 39.275 -141.605 39.605 -141.275 ;
        RECT 39.275 -142.965 39.605 -142.635 ;
        RECT 39.275 -144.325 39.605 -143.995 ;
        RECT 39.275 -145.685 39.605 -145.355 ;
        RECT 39.275 -147.045 39.605 -146.715 ;
        RECT 39.275 -148.405 39.605 -148.075 ;
        RECT 39.275 -149.765 39.605 -149.435 ;
        RECT 39.275 -151.125 39.605 -150.795 ;
        RECT 39.275 -152.485 39.605 -152.155 ;
        RECT 39.275 -153.845 39.605 -153.515 ;
        RECT 39.275 -155.205 39.605 -154.875 ;
        RECT 39.275 -156.565 39.605 -156.235 ;
        RECT 39.275 -157.925 39.605 -157.595 ;
        RECT 39.275 -160.17 39.605 -159.04 ;
        RECT 39.28 -160.285 39.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.91 -94.075 40.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 127.225 40.965 128.355 ;
        RECT 40.635 124.955 40.965 125.285 ;
        RECT 40.635 123.595 40.965 123.925 ;
        RECT 40.64 123.595 40.96 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 -1.525 40.965 -1.195 ;
        RECT 40.635 -2.885 40.965 -2.555 ;
        RECT 40.64 -3.56 40.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 127.225 42.325 128.355 ;
        RECT 41.995 124.955 42.325 125.285 ;
        RECT 41.995 123.595 42.325 123.925 ;
        RECT 42 123.595 42.32 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 -1.525 42.325 -1.195 ;
        RECT 41.995 -2.885 42.325 -2.555 ;
        RECT 42 -3.56 42.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 127.225 43.685 128.355 ;
        RECT 43.355 124.955 43.685 125.285 ;
        RECT 43.355 123.595 43.685 123.925 ;
        RECT 43.36 123.595 43.68 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -1.525 43.685 -1.195 ;
        RECT 43.355 -2.885 43.685 -2.555 ;
        RECT 43.36 -3.56 43.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -91.285 43.685 -90.955 ;
        RECT 43.355 -92.645 43.685 -92.315 ;
        RECT 43.355 -94.005 43.685 -93.675 ;
        RECT 43.355 -95.365 43.685 -95.035 ;
        RECT 43.355 -96.725 43.685 -96.395 ;
        RECT 43.355 -98.085 43.685 -97.755 ;
        RECT 43.355 -99.445 43.685 -99.115 ;
        RECT 43.355 -100.805 43.685 -100.475 ;
        RECT 43.355 -102.165 43.685 -101.835 ;
        RECT 43.355 -103.525 43.685 -103.195 ;
        RECT 43.355 -104.885 43.685 -104.555 ;
        RECT 43.355 -106.245 43.685 -105.915 ;
        RECT 43.355 -107.605 43.685 -107.275 ;
        RECT 43.355 -108.965 43.685 -108.635 ;
        RECT 43.355 -110.325 43.685 -109.995 ;
        RECT 43.355 -111.685 43.685 -111.355 ;
        RECT 43.355 -113.045 43.685 -112.715 ;
        RECT 43.355 -114.405 43.685 -114.075 ;
        RECT 43.355 -115.765 43.685 -115.435 ;
        RECT 43.355 -117.125 43.685 -116.795 ;
        RECT 43.355 -118.485 43.685 -118.155 ;
        RECT 43.355 -119.845 43.685 -119.515 ;
        RECT 43.355 -121.205 43.685 -120.875 ;
        RECT 43.355 -122.565 43.685 -122.235 ;
        RECT 43.355 -123.925 43.685 -123.595 ;
        RECT 43.355 -125.285 43.685 -124.955 ;
        RECT 43.355 -126.645 43.685 -126.315 ;
        RECT 43.355 -128.005 43.685 -127.675 ;
        RECT 43.355 -129.365 43.685 -129.035 ;
        RECT 43.355 -130.725 43.685 -130.395 ;
        RECT 43.355 -132.085 43.685 -131.755 ;
        RECT 43.355 -133.445 43.685 -133.115 ;
        RECT 43.355 -134.805 43.685 -134.475 ;
        RECT 43.355 -136.165 43.685 -135.835 ;
        RECT 43.355 -137.525 43.685 -137.195 ;
        RECT 43.355 -138.885 43.685 -138.555 ;
        RECT 43.355 -140.245 43.685 -139.915 ;
        RECT 43.355 -141.605 43.685 -141.275 ;
        RECT 43.355 -142.965 43.685 -142.635 ;
        RECT 43.355 -144.325 43.685 -143.995 ;
        RECT 43.355 -145.685 43.685 -145.355 ;
        RECT 43.355 -147.045 43.685 -146.715 ;
        RECT 43.355 -148.405 43.685 -148.075 ;
        RECT 43.355 -149.765 43.685 -149.435 ;
        RECT 43.355 -151.125 43.685 -150.795 ;
        RECT 43.355 -152.485 43.685 -152.155 ;
        RECT 43.355 -153.845 43.685 -153.515 ;
        RECT 43.355 -155.205 43.685 -154.875 ;
        RECT 43.355 -156.565 43.685 -156.235 ;
        RECT 43.355 -157.925 43.685 -157.595 ;
        RECT 43.355 -160.17 43.685 -159.04 ;
        RECT 43.36 -160.285 43.68 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 127.225 45.045 128.355 ;
        RECT 44.715 124.955 45.045 125.285 ;
        RECT 44.715 123.595 45.045 123.925 ;
        RECT 44.72 123.595 45.04 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 -95.365 45.045 -95.035 ;
        RECT 44.715 -96.725 45.045 -96.395 ;
        RECT 44.715 -98.085 45.045 -97.755 ;
        RECT 44.715 -99.445 45.045 -99.115 ;
        RECT 44.715 -100.805 45.045 -100.475 ;
        RECT 44.715 -102.165 45.045 -101.835 ;
        RECT 44.715 -103.525 45.045 -103.195 ;
        RECT 44.715 -104.885 45.045 -104.555 ;
        RECT 44.715 -106.245 45.045 -105.915 ;
        RECT 44.715 -107.605 45.045 -107.275 ;
        RECT 44.715 -108.965 45.045 -108.635 ;
        RECT 44.715 -110.325 45.045 -109.995 ;
        RECT 44.715 -111.685 45.045 -111.355 ;
        RECT 44.715 -113.045 45.045 -112.715 ;
        RECT 44.715 -114.405 45.045 -114.075 ;
        RECT 44.715 -115.765 45.045 -115.435 ;
        RECT 44.715 -117.125 45.045 -116.795 ;
        RECT 44.715 -118.485 45.045 -118.155 ;
        RECT 44.715 -119.845 45.045 -119.515 ;
        RECT 44.715 -121.205 45.045 -120.875 ;
        RECT 44.715 -122.565 45.045 -122.235 ;
        RECT 44.715 -123.925 45.045 -123.595 ;
        RECT 44.715 -125.285 45.045 -124.955 ;
        RECT 44.715 -126.645 45.045 -126.315 ;
        RECT 44.715 -128.005 45.045 -127.675 ;
        RECT 44.715 -129.365 45.045 -129.035 ;
        RECT 44.715 -130.725 45.045 -130.395 ;
        RECT 44.715 -132.085 45.045 -131.755 ;
        RECT 44.715 -133.445 45.045 -133.115 ;
        RECT 44.715 -134.805 45.045 -134.475 ;
        RECT 44.715 -136.165 45.045 -135.835 ;
        RECT 44.715 -137.525 45.045 -137.195 ;
        RECT 44.715 -138.885 45.045 -138.555 ;
        RECT 44.715 -140.245 45.045 -139.915 ;
        RECT 44.715 -141.605 45.045 -141.275 ;
        RECT 44.715 -142.965 45.045 -142.635 ;
        RECT 44.715 -144.325 45.045 -143.995 ;
        RECT 44.715 -145.685 45.045 -145.355 ;
        RECT 44.715 -147.045 45.045 -146.715 ;
        RECT 44.715 -148.405 45.045 -148.075 ;
        RECT 44.715 -149.765 45.045 -149.435 ;
        RECT 44.715 -151.125 45.045 -150.795 ;
        RECT 44.715 -152.485 45.045 -152.155 ;
        RECT 44.715 -153.845 45.045 -153.515 ;
        RECT 44.715 -155.205 45.045 -154.875 ;
        RECT 44.715 -156.565 45.045 -156.235 ;
        RECT 44.715 -157.925 45.045 -157.595 ;
        RECT 44.715 -160.17 45.045 -159.04 ;
        RECT 44.72 -160.285 45.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.01 -94.075 46.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 127.225 46.405 128.355 ;
        RECT 46.075 124.955 46.405 125.285 ;
        RECT 46.075 123.595 46.405 123.925 ;
        RECT 46.08 123.595 46.4 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 127.225 47.765 128.355 ;
        RECT 47.435 124.955 47.765 125.285 ;
        RECT 47.435 123.595 47.765 123.925 ;
        RECT 47.44 123.595 47.76 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 -1.525 47.765 -1.195 ;
        RECT 47.435 -2.885 47.765 -2.555 ;
        RECT 47.44 -3.56 47.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 127.225 49.125 128.355 ;
        RECT 48.795 124.955 49.125 125.285 ;
        RECT 48.795 123.595 49.125 123.925 ;
        RECT 48.8 123.595 49.12 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 -1.525 49.125 -1.195 ;
        RECT 48.795 -2.885 49.125 -2.555 ;
        RECT 48.8 -3.56 49.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 127.225 50.485 128.355 ;
        RECT 50.155 124.955 50.485 125.285 ;
        RECT 50.155 123.595 50.485 123.925 ;
        RECT 50.16 123.595 50.48 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -1.525 50.485 -1.195 ;
        RECT 50.155 -2.885 50.485 -2.555 ;
        RECT 50.16 -3.56 50.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -91.285 50.485 -90.955 ;
        RECT 50.155 -92.645 50.485 -92.315 ;
        RECT 50.155 -94.005 50.485 -93.675 ;
        RECT 50.155 -95.365 50.485 -95.035 ;
        RECT 50.155 -96.725 50.485 -96.395 ;
        RECT 50.155 -98.085 50.485 -97.755 ;
        RECT 50.155 -99.445 50.485 -99.115 ;
        RECT 50.155 -100.805 50.485 -100.475 ;
        RECT 50.155 -102.165 50.485 -101.835 ;
        RECT 50.155 -103.525 50.485 -103.195 ;
        RECT 50.155 -104.885 50.485 -104.555 ;
        RECT 50.155 -106.245 50.485 -105.915 ;
        RECT 50.155 -107.605 50.485 -107.275 ;
        RECT 50.155 -108.965 50.485 -108.635 ;
        RECT 50.155 -110.325 50.485 -109.995 ;
        RECT 50.155 -111.685 50.485 -111.355 ;
        RECT 50.155 -113.045 50.485 -112.715 ;
        RECT 50.155 -114.405 50.485 -114.075 ;
        RECT 50.155 -115.765 50.485 -115.435 ;
        RECT 50.155 -117.125 50.485 -116.795 ;
        RECT 50.155 -118.485 50.485 -118.155 ;
        RECT 50.155 -119.845 50.485 -119.515 ;
        RECT 50.155 -121.205 50.485 -120.875 ;
        RECT 50.155 -122.565 50.485 -122.235 ;
        RECT 50.155 -123.925 50.485 -123.595 ;
        RECT 50.155 -125.285 50.485 -124.955 ;
        RECT 50.155 -126.645 50.485 -126.315 ;
        RECT 50.155 -128.005 50.485 -127.675 ;
        RECT 50.155 -129.365 50.485 -129.035 ;
        RECT 50.155 -130.725 50.485 -130.395 ;
        RECT 50.155 -132.085 50.485 -131.755 ;
        RECT 50.155 -133.445 50.485 -133.115 ;
        RECT 50.155 -134.805 50.485 -134.475 ;
        RECT 50.155 -136.165 50.485 -135.835 ;
        RECT 50.155 -137.525 50.485 -137.195 ;
        RECT 50.155 -138.885 50.485 -138.555 ;
        RECT 50.155 -140.245 50.485 -139.915 ;
        RECT 50.155 -141.605 50.485 -141.275 ;
        RECT 50.155 -142.965 50.485 -142.635 ;
        RECT 50.155 -144.325 50.485 -143.995 ;
        RECT 50.155 -145.685 50.485 -145.355 ;
        RECT 50.155 -147.045 50.485 -146.715 ;
        RECT 50.155 -148.405 50.485 -148.075 ;
        RECT 50.155 -149.765 50.485 -149.435 ;
        RECT 50.155 -151.125 50.485 -150.795 ;
        RECT 50.155 -152.485 50.485 -152.155 ;
        RECT 50.155 -153.845 50.485 -153.515 ;
        RECT 50.155 -155.205 50.485 -154.875 ;
        RECT 50.155 -156.565 50.485 -156.235 ;
        RECT 50.155 -157.925 50.485 -157.595 ;
        RECT 50.155 -160.17 50.485 -159.04 ;
        RECT 50.16 -160.285 50.48 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 127.225 51.845 128.355 ;
        RECT 51.515 124.955 51.845 125.285 ;
        RECT 51.515 123.595 51.845 123.925 ;
        RECT 51.52 123.595 51.84 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 -95.365 51.845 -95.035 ;
        RECT 51.515 -96.725 51.845 -96.395 ;
        RECT 51.515 -98.085 51.845 -97.755 ;
        RECT 51.515 -99.445 51.845 -99.115 ;
        RECT 51.515 -100.805 51.845 -100.475 ;
        RECT 51.515 -102.165 51.845 -101.835 ;
        RECT 51.515 -103.525 51.845 -103.195 ;
        RECT 51.515 -104.885 51.845 -104.555 ;
        RECT 51.515 -106.245 51.845 -105.915 ;
        RECT 51.515 -107.605 51.845 -107.275 ;
        RECT 51.515 -108.965 51.845 -108.635 ;
        RECT 51.515 -110.325 51.845 -109.995 ;
        RECT 51.515 -111.685 51.845 -111.355 ;
        RECT 51.515 -113.045 51.845 -112.715 ;
        RECT 51.515 -114.405 51.845 -114.075 ;
        RECT 51.515 -115.765 51.845 -115.435 ;
        RECT 51.515 -117.125 51.845 -116.795 ;
        RECT 51.515 -118.485 51.845 -118.155 ;
        RECT 51.515 -119.845 51.845 -119.515 ;
        RECT 51.515 -121.205 51.845 -120.875 ;
        RECT 51.515 -122.565 51.845 -122.235 ;
        RECT 51.515 -123.925 51.845 -123.595 ;
        RECT 51.515 -125.285 51.845 -124.955 ;
        RECT 51.515 -126.645 51.845 -126.315 ;
        RECT 51.515 -128.005 51.845 -127.675 ;
        RECT 51.515 -129.365 51.845 -129.035 ;
        RECT 51.515 -130.725 51.845 -130.395 ;
        RECT 51.515 -132.085 51.845 -131.755 ;
        RECT 51.515 -133.445 51.845 -133.115 ;
        RECT 51.515 -134.805 51.845 -134.475 ;
        RECT 51.515 -136.165 51.845 -135.835 ;
        RECT 51.515 -137.525 51.845 -137.195 ;
        RECT 51.515 -138.885 51.845 -138.555 ;
        RECT 51.515 -140.245 51.845 -139.915 ;
        RECT 51.515 -141.605 51.845 -141.275 ;
        RECT 51.515 -142.965 51.845 -142.635 ;
        RECT 51.515 -144.325 51.845 -143.995 ;
        RECT 51.515 -145.685 51.845 -145.355 ;
        RECT 51.515 -147.045 51.845 -146.715 ;
        RECT 51.515 -148.405 51.845 -148.075 ;
        RECT 51.515 -149.765 51.845 -149.435 ;
        RECT 51.515 -151.125 51.845 -150.795 ;
        RECT 51.515 -152.485 51.845 -152.155 ;
        RECT 51.515 -153.845 51.845 -153.515 ;
        RECT 51.515 -155.205 51.845 -154.875 ;
        RECT 51.515 -156.565 51.845 -156.235 ;
        RECT 51.515 -157.925 51.845 -157.595 ;
        RECT 51.515 -160.17 51.845 -159.04 ;
        RECT 51.52 -160.285 51.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.11 -94.075 52.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 127.225 53.205 128.355 ;
        RECT 52.875 124.955 53.205 125.285 ;
        RECT 52.875 123.595 53.205 123.925 ;
        RECT 52.88 123.595 53.2 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 -1.525 53.205 -1.195 ;
        RECT 52.875 -2.885 53.205 -2.555 ;
        RECT 52.88 -3.56 53.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 127.225 54.565 128.355 ;
        RECT 54.235 124.955 54.565 125.285 ;
        RECT 54.235 123.595 54.565 123.925 ;
        RECT 54.24 123.595 54.56 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 -1.525 54.565 -1.195 ;
        RECT 54.235 -2.885 54.565 -2.555 ;
        RECT 54.24 -3.56 54.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 127.225 55.925 128.355 ;
        RECT 55.595 124.955 55.925 125.285 ;
        RECT 55.595 123.595 55.925 123.925 ;
        RECT 55.6 123.595 55.92 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 -1.525 55.925 -1.195 ;
        RECT 55.595 -2.885 55.925 -2.555 ;
        RECT 55.6 -3.56 55.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 127.225 57.285 128.355 ;
        RECT 56.955 124.955 57.285 125.285 ;
        RECT 56.955 123.595 57.285 123.925 ;
        RECT 56.96 123.595 57.28 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 -95.365 57.285 -95.035 ;
        RECT 56.955 -96.725 57.285 -96.395 ;
        RECT 56.955 -98.085 57.285 -97.755 ;
        RECT 56.955 -99.445 57.285 -99.115 ;
        RECT 56.955 -100.805 57.285 -100.475 ;
        RECT 56.955 -102.165 57.285 -101.835 ;
        RECT 56.955 -103.525 57.285 -103.195 ;
        RECT 56.955 -104.885 57.285 -104.555 ;
        RECT 56.955 -106.245 57.285 -105.915 ;
        RECT 56.955 -107.605 57.285 -107.275 ;
        RECT 56.955 -108.965 57.285 -108.635 ;
        RECT 56.955 -110.325 57.285 -109.995 ;
        RECT 56.955 -111.685 57.285 -111.355 ;
        RECT 56.955 -113.045 57.285 -112.715 ;
        RECT 56.955 -114.405 57.285 -114.075 ;
        RECT 56.955 -115.765 57.285 -115.435 ;
        RECT 56.955 -117.125 57.285 -116.795 ;
        RECT 56.955 -118.485 57.285 -118.155 ;
        RECT 56.955 -119.845 57.285 -119.515 ;
        RECT 56.955 -121.205 57.285 -120.875 ;
        RECT 56.955 -122.565 57.285 -122.235 ;
        RECT 56.955 -123.925 57.285 -123.595 ;
        RECT 56.955 -125.285 57.285 -124.955 ;
        RECT 56.955 -126.645 57.285 -126.315 ;
        RECT 56.955 -128.005 57.285 -127.675 ;
        RECT 56.955 -129.365 57.285 -129.035 ;
        RECT 56.955 -130.725 57.285 -130.395 ;
        RECT 56.955 -132.085 57.285 -131.755 ;
        RECT 56.955 -133.445 57.285 -133.115 ;
        RECT 56.955 -134.805 57.285 -134.475 ;
        RECT 56.955 -136.165 57.285 -135.835 ;
        RECT 56.955 -137.525 57.285 -137.195 ;
        RECT 56.955 -138.885 57.285 -138.555 ;
        RECT 56.955 -140.245 57.285 -139.915 ;
        RECT 56.955 -141.605 57.285 -141.275 ;
        RECT 56.955 -142.965 57.285 -142.635 ;
        RECT 56.955 -144.325 57.285 -143.995 ;
        RECT 56.955 -145.685 57.285 -145.355 ;
        RECT 56.955 -147.045 57.285 -146.715 ;
        RECT 56.955 -148.405 57.285 -148.075 ;
        RECT 56.955 -149.765 57.285 -149.435 ;
        RECT 56.955 -151.125 57.285 -150.795 ;
        RECT 56.955 -152.485 57.285 -152.155 ;
        RECT 56.955 -153.845 57.285 -153.515 ;
        RECT 56.955 -155.205 57.285 -154.875 ;
        RECT 56.955 -156.565 57.285 -156.235 ;
        RECT 56.955 -157.925 57.285 -157.595 ;
        RECT 56.955 -160.17 57.285 -159.04 ;
        RECT 56.96 -160.285 57.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.21 -94.075 58.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.315 127.225 58.645 128.355 ;
        RECT 58.315 124.955 58.645 125.285 ;
        RECT 58.315 123.595 58.645 123.925 ;
        RECT 58.32 123.595 58.64 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 127.225 60.005 128.355 ;
        RECT 59.675 124.955 60.005 125.285 ;
        RECT 59.675 123.595 60.005 123.925 ;
        RECT 59.68 123.595 60 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 -1.525 60.005 -1.195 ;
        RECT 59.675 -2.885 60.005 -2.555 ;
        RECT 59.68 -3.56 60 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 -91.285 60.005 -90.955 ;
        RECT 59.675 -92.645 60.005 -92.315 ;
        RECT 59.675 -94.005 60.005 -93.675 ;
        RECT 59.675 -95.365 60.005 -95.035 ;
        RECT 59.675 -96.725 60.005 -96.395 ;
        RECT 59.675 -98.085 60.005 -97.755 ;
        RECT 59.675 -99.445 60.005 -99.115 ;
        RECT 59.675 -100.805 60.005 -100.475 ;
        RECT 59.675 -102.165 60.005 -101.835 ;
        RECT 59.675 -103.525 60.005 -103.195 ;
        RECT 59.675 -104.885 60.005 -104.555 ;
        RECT 59.675 -106.245 60.005 -105.915 ;
        RECT 59.675 -107.605 60.005 -107.275 ;
        RECT 59.675 -108.965 60.005 -108.635 ;
        RECT 59.675 -110.325 60.005 -109.995 ;
        RECT 59.675 -111.685 60.005 -111.355 ;
        RECT 59.675 -113.045 60.005 -112.715 ;
        RECT 59.675 -114.405 60.005 -114.075 ;
        RECT 59.675 -115.765 60.005 -115.435 ;
        RECT 59.675 -117.125 60.005 -116.795 ;
        RECT 59.675 -118.485 60.005 -118.155 ;
        RECT 59.675 -119.845 60.005 -119.515 ;
        RECT 59.675 -121.205 60.005 -120.875 ;
        RECT 59.675 -122.565 60.005 -122.235 ;
        RECT 59.675 -123.925 60.005 -123.595 ;
        RECT 59.675 -125.285 60.005 -124.955 ;
        RECT 59.675 -126.645 60.005 -126.315 ;
        RECT 59.675 -128.005 60.005 -127.675 ;
        RECT 59.675 -129.365 60.005 -129.035 ;
        RECT 59.675 -130.725 60.005 -130.395 ;
        RECT 59.675 -132.085 60.005 -131.755 ;
        RECT 59.675 -133.445 60.005 -133.115 ;
        RECT 59.675 -134.805 60.005 -134.475 ;
        RECT 59.675 -136.165 60.005 -135.835 ;
        RECT 59.675 -137.525 60.005 -137.195 ;
        RECT 59.675 -138.885 60.005 -138.555 ;
        RECT 59.675 -140.245 60.005 -139.915 ;
        RECT 59.675 -141.605 60.005 -141.275 ;
        RECT 59.675 -142.965 60.005 -142.635 ;
        RECT 59.675 -144.325 60.005 -143.995 ;
        RECT 59.675 -145.685 60.005 -145.355 ;
        RECT 59.675 -147.045 60.005 -146.715 ;
        RECT 59.675 -148.405 60.005 -148.075 ;
        RECT 59.675 -149.765 60.005 -149.435 ;
        RECT 59.675 -151.125 60.005 -150.795 ;
        RECT 59.675 -152.485 60.005 -152.155 ;
        RECT 59.675 -153.845 60.005 -153.515 ;
        RECT 59.675 -155.205 60.005 -154.875 ;
        RECT 59.675 -156.565 60.005 -156.235 ;
        RECT 59.675 -157.925 60.005 -157.595 ;
        RECT 59.675 -160.17 60.005 -159.04 ;
        RECT 59.68 -160.285 60 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 127.225 61.365 128.355 ;
        RECT 61.035 124.955 61.365 125.285 ;
        RECT 61.035 123.595 61.365 123.925 ;
        RECT 61.04 123.595 61.36 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 -1.525 61.365 -1.195 ;
        RECT 61.035 -2.885 61.365 -2.555 ;
        RECT 61.04 -3.56 61.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 127.225 62.725 128.355 ;
        RECT 62.395 124.955 62.725 125.285 ;
        RECT 62.395 123.595 62.725 123.925 ;
        RECT 62.4 123.595 62.72 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -1.525 62.725 -1.195 ;
        RECT 62.395 -2.885 62.725 -2.555 ;
        RECT 62.4 -3.56 62.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -91.285 62.725 -90.955 ;
        RECT 62.395 -92.645 62.725 -92.315 ;
        RECT 62.395 -94.005 62.725 -93.675 ;
        RECT 62.395 -95.365 62.725 -95.035 ;
        RECT 62.395 -96.725 62.725 -96.395 ;
        RECT 62.395 -98.085 62.725 -97.755 ;
        RECT 62.395 -99.445 62.725 -99.115 ;
        RECT 62.395 -100.805 62.725 -100.475 ;
        RECT 62.395 -102.165 62.725 -101.835 ;
        RECT 62.395 -103.525 62.725 -103.195 ;
        RECT 62.395 -104.885 62.725 -104.555 ;
        RECT 62.395 -106.245 62.725 -105.915 ;
        RECT 62.395 -107.605 62.725 -107.275 ;
        RECT 62.395 -108.965 62.725 -108.635 ;
        RECT 62.395 -110.325 62.725 -109.995 ;
        RECT 62.395 -111.685 62.725 -111.355 ;
        RECT 62.395 -113.045 62.725 -112.715 ;
        RECT 62.395 -114.405 62.725 -114.075 ;
        RECT 62.395 -115.765 62.725 -115.435 ;
        RECT 62.395 -117.125 62.725 -116.795 ;
        RECT 62.395 -118.485 62.725 -118.155 ;
        RECT 62.395 -119.845 62.725 -119.515 ;
        RECT 62.395 -121.205 62.725 -120.875 ;
        RECT 62.395 -122.565 62.725 -122.235 ;
        RECT 62.395 -123.925 62.725 -123.595 ;
        RECT 62.395 -125.285 62.725 -124.955 ;
        RECT 62.395 -126.645 62.725 -126.315 ;
        RECT 62.395 -128.005 62.725 -127.675 ;
        RECT 62.395 -129.365 62.725 -129.035 ;
        RECT 62.395 -130.725 62.725 -130.395 ;
        RECT 62.395 -132.085 62.725 -131.755 ;
        RECT 62.395 -133.445 62.725 -133.115 ;
        RECT 62.395 -134.805 62.725 -134.475 ;
        RECT 62.395 -136.165 62.725 -135.835 ;
        RECT 62.395 -137.525 62.725 -137.195 ;
        RECT 62.395 -138.885 62.725 -138.555 ;
        RECT 62.395 -140.245 62.725 -139.915 ;
        RECT 62.395 -141.605 62.725 -141.275 ;
        RECT 62.395 -142.965 62.725 -142.635 ;
        RECT 62.395 -144.325 62.725 -143.995 ;
        RECT 62.395 -145.685 62.725 -145.355 ;
        RECT 62.395 -147.045 62.725 -146.715 ;
        RECT 62.395 -148.405 62.725 -148.075 ;
        RECT 62.395 -149.765 62.725 -149.435 ;
        RECT 62.395 -151.125 62.725 -150.795 ;
        RECT 62.395 -152.485 62.725 -152.155 ;
        RECT 62.395 -153.845 62.725 -153.515 ;
        RECT 62.395 -155.205 62.725 -154.875 ;
        RECT 62.395 -156.565 62.725 -156.235 ;
        RECT 62.395 -157.925 62.725 -157.595 ;
        RECT 62.395 -160.17 62.725 -159.04 ;
        RECT 62.4 -160.285 62.72 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 127.225 64.085 128.355 ;
        RECT 63.755 124.955 64.085 125.285 ;
        RECT 63.755 123.595 64.085 123.925 ;
        RECT 63.76 123.595 64.08 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 -95.365 64.085 -95.035 ;
        RECT 63.755 -96.725 64.085 -96.395 ;
        RECT 63.755 -98.085 64.085 -97.755 ;
        RECT 63.755 -99.445 64.085 -99.115 ;
        RECT 63.755 -100.805 64.085 -100.475 ;
        RECT 63.755 -102.165 64.085 -101.835 ;
        RECT 63.755 -103.525 64.085 -103.195 ;
        RECT 63.755 -104.885 64.085 -104.555 ;
        RECT 63.755 -106.245 64.085 -105.915 ;
        RECT 63.755 -107.605 64.085 -107.275 ;
        RECT 63.755 -108.965 64.085 -108.635 ;
        RECT 63.755 -110.325 64.085 -109.995 ;
        RECT 63.755 -111.685 64.085 -111.355 ;
        RECT 63.755 -113.045 64.085 -112.715 ;
        RECT 63.755 -114.405 64.085 -114.075 ;
        RECT 63.755 -115.765 64.085 -115.435 ;
        RECT 63.755 -117.125 64.085 -116.795 ;
        RECT 63.755 -118.485 64.085 -118.155 ;
        RECT 63.755 -119.845 64.085 -119.515 ;
        RECT 63.755 -121.205 64.085 -120.875 ;
        RECT 63.755 -122.565 64.085 -122.235 ;
        RECT 63.755 -123.925 64.085 -123.595 ;
        RECT 63.755 -125.285 64.085 -124.955 ;
        RECT 63.755 -126.645 64.085 -126.315 ;
        RECT 63.755 -128.005 64.085 -127.675 ;
        RECT 63.755 -129.365 64.085 -129.035 ;
        RECT 63.755 -130.725 64.085 -130.395 ;
        RECT 63.755 -132.085 64.085 -131.755 ;
        RECT 63.755 -133.445 64.085 -133.115 ;
        RECT 63.755 -134.805 64.085 -134.475 ;
        RECT 63.755 -136.165 64.085 -135.835 ;
        RECT 63.755 -137.525 64.085 -137.195 ;
        RECT 63.755 -138.885 64.085 -138.555 ;
        RECT 63.755 -140.245 64.085 -139.915 ;
        RECT 63.755 -141.605 64.085 -141.275 ;
        RECT 63.755 -142.965 64.085 -142.635 ;
        RECT 63.755 -144.325 64.085 -143.995 ;
        RECT 63.755 -145.685 64.085 -145.355 ;
        RECT 63.755 -147.045 64.085 -146.715 ;
        RECT 63.755 -148.405 64.085 -148.075 ;
        RECT 63.755 -149.765 64.085 -149.435 ;
        RECT 63.755 -151.125 64.085 -150.795 ;
        RECT 63.755 -152.485 64.085 -152.155 ;
        RECT 63.755 -153.845 64.085 -153.515 ;
        RECT 63.755 -155.205 64.085 -154.875 ;
        RECT 63.755 -156.565 64.085 -156.235 ;
        RECT 63.755 -157.925 64.085 -157.595 ;
        RECT 63.755 -160.17 64.085 -159.04 ;
        RECT 63.76 -160.285 64.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.31 -94.075 64.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 127.225 65.445 128.355 ;
        RECT 65.115 124.955 65.445 125.285 ;
        RECT 65.115 123.595 65.445 123.925 ;
        RECT 65.12 123.595 65.44 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 -1.525 65.445 -1.195 ;
        RECT 65.115 -2.885 65.445 -2.555 ;
        RECT 65.12 -3.56 65.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 127.225 66.805 128.355 ;
        RECT 66.475 124.955 66.805 125.285 ;
        RECT 66.475 123.595 66.805 123.925 ;
        RECT 66.48 123.595 66.8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 -1.525 66.805 -1.195 ;
        RECT 66.475 -2.885 66.805 -2.555 ;
        RECT 66.48 -3.56 66.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 127.225 68.165 128.355 ;
        RECT 67.835 124.955 68.165 125.285 ;
        RECT 67.835 123.595 68.165 123.925 ;
        RECT 67.84 123.595 68.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 -1.525 68.165 -1.195 ;
        RECT 67.835 -2.885 68.165 -2.555 ;
        RECT 67.84 -3.56 68.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 -91.285 68.165 -90.955 ;
        RECT 67.835 -92.645 68.165 -92.315 ;
        RECT 67.835 -94.005 68.165 -93.675 ;
        RECT 67.835 -95.365 68.165 -95.035 ;
        RECT 67.835 -96.725 68.165 -96.395 ;
        RECT 67.835 -98.085 68.165 -97.755 ;
        RECT 67.835 -99.445 68.165 -99.115 ;
        RECT 67.835 -100.805 68.165 -100.475 ;
        RECT 67.835 -102.165 68.165 -101.835 ;
        RECT 67.835 -103.525 68.165 -103.195 ;
        RECT 67.835 -104.885 68.165 -104.555 ;
        RECT 67.835 -106.245 68.165 -105.915 ;
        RECT 67.835 -107.605 68.165 -107.275 ;
        RECT 67.835 -108.965 68.165 -108.635 ;
        RECT 67.835 -110.325 68.165 -109.995 ;
        RECT 67.835 -111.685 68.165 -111.355 ;
        RECT 67.835 -113.045 68.165 -112.715 ;
        RECT 67.835 -114.405 68.165 -114.075 ;
        RECT 67.835 -115.765 68.165 -115.435 ;
        RECT 67.835 -117.125 68.165 -116.795 ;
        RECT 67.835 -118.485 68.165 -118.155 ;
        RECT 67.835 -119.845 68.165 -119.515 ;
        RECT 67.835 -121.205 68.165 -120.875 ;
        RECT 67.835 -122.565 68.165 -122.235 ;
        RECT 67.835 -123.925 68.165 -123.595 ;
        RECT 67.835 -125.285 68.165 -124.955 ;
        RECT 67.835 -126.645 68.165 -126.315 ;
        RECT 67.835 -128.005 68.165 -127.675 ;
        RECT 67.835 -129.365 68.165 -129.035 ;
        RECT 67.835 -130.725 68.165 -130.395 ;
        RECT 67.835 -132.085 68.165 -131.755 ;
        RECT 67.835 -133.445 68.165 -133.115 ;
        RECT 67.835 -134.805 68.165 -134.475 ;
        RECT 67.835 -136.165 68.165 -135.835 ;
        RECT 67.835 -137.525 68.165 -137.195 ;
        RECT 67.835 -138.885 68.165 -138.555 ;
        RECT 67.835 -140.245 68.165 -139.915 ;
        RECT 67.835 -141.605 68.165 -141.275 ;
        RECT 67.835 -142.965 68.165 -142.635 ;
        RECT 67.835 -144.325 68.165 -143.995 ;
        RECT 67.835 -145.685 68.165 -145.355 ;
        RECT 67.835 -147.045 68.165 -146.715 ;
        RECT 67.835 -148.405 68.165 -148.075 ;
        RECT 67.835 -149.765 68.165 -149.435 ;
        RECT 67.835 -151.125 68.165 -150.795 ;
        RECT 67.835 -152.485 68.165 -152.155 ;
        RECT 67.835 -153.845 68.165 -153.515 ;
        RECT 67.835 -155.205 68.165 -154.875 ;
        RECT 67.835 -156.565 68.165 -156.235 ;
        RECT 67.835 -157.925 68.165 -157.595 ;
        RECT 67.835 -160.17 68.165 -159.04 ;
        RECT 67.84 -160.285 68.16 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 127.225 69.525 128.355 ;
        RECT 69.195 124.955 69.525 125.285 ;
        RECT 69.195 123.595 69.525 123.925 ;
        RECT 69.2 123.595 69.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 -114.405 69.525 -114.075 ;
        RECT 69.195 -115.765 69.525 -115.435 ;
        RECT 69.195 -117.125 69.525 -116.795 ;
        RECT 69.195 -118.485 69.525 -118.155 ;
        RECT 69.195 -119.845 69.525 -119.515 ;
        RECT 69.195 -121.205 69.525 -120.875 ;
        RECT 69.195 -122.565 69.525 -122.235 ;
        RECT 69.195 -123.925 69.525 -123.595 ;
        RECT 69.195 -125.285 69.525 -124.955 ;
        RECT 69.195 -126.645 69.525 -126.315 ;
        RECT 69.195 -128.005 69.525 -127.675 ;
        RECT 69.195 -129.365 69.525 -129.035 ;
        RECT 69.195 -130.725 69.525 -130.395 ;
        RECT 69.195 -132.085 69.525 -131.755 ;
        RECT 69.195 -133.445 69.525 -133.115 ;
        RECT 69.195 -134.805 69.525 -134.475 ;
        RECT 69.195 -136.165 69.525 -135.835 ;
        RECT 69.195 -137.525 69.525 -137.195 ;
        RECT 69.195 -138.885 69.525 -138.555 ;
        RECT 69.195 -140.245 69.525 -139.915 ;
        RECT 69.195 -141.605 69.525 -141.275 ;
        RECT 69.195 -142.965 69.525 -142.635 ;
        RECT 69.195 -144.325 69.525 -143.995 ;
        RECT 69.195 -145.685 69.525 -145.355 ;
        RECT 69.195 -147.045 69.525 -146.715 ;
        RECT 69.195 -148.405 69.525 -148.075 ;
        RECT 69.195 -149.765 69.525 -149.435 ;
        RECT 69.195 -151.125 69.525 -150.795 ;
        RECT 69.195 -152.485 69.525 -152.155 ;
        RECT 69.195 -153.845 69.525 -153.515 ;
        RECT 69.195 -155.205 69.525 -154.875 ;
        RECT 69.195 -156.565 69.525 -156.235 ;
        RECT 69.195 -157.925 69.525 -157.595 ;
        RECT 69.195 -160.17 69.525 -159.04 ;
        RECT 69.2 -160.285 69.52 -95.035 ;
        RECT 69.195 -95.365 69.525 -95.035 ;
        RECT 69.195 -96.725 69.525 -96.395 ;
        RECT 69.195 -98.085 69.525 -97.755 ;
        RECT 69.195 -99.445 69.525 -99.115 ;
        RECT 69.195 -100.805 69.525 -100.475 ;
        RECT 69.195 -102.165 69.525 -101.835 ;
        RECT 69.195 -103.525 69.525 -103.195 ;
        RECT 69.195 -104.885 69.525 -104.555 ;
        RECT 69.195 -106.245 69.525 -105.915 ;
        RECT 69.195 -107.605 69.525 -107.275 ;
        RECT 69.195 -108.965 69.525 -108.635 ;
        RECT 69.195 -110.325 69.525 -109.995 ;
        RECT 69.195 -111.685 69.525 -111.355 ;
        RECT 69.195 -113.045 69.525 -112.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 127.225 -1.195 128.355 ;
        RECT -1.525 124.955 -1.195 125.285 ;
        RECT -1.525 123.595 -1.195 123.925 ;
        RECT -1.525 122.215 -1.195 122.545 ;
        RECT -1.525 120.165 -1.195 120.495 ;
        RECT -1.525 118.235 -1.195 118.565 ;
        RECT -1.525 116.395 -1.195 116.725 ;
        RECT -1.525 114.905 -1.195 115.235 ;
        RECT -1.525 113.235 -1.195 113.565 ;
        RECT -1.525 111.745 -1.195 112.075 ;
        RECT -1.525 110.075 -1.195 110.405 ;
        RECT -1.525 108.585 -1.195 108.915 ;
        RECT -1.525 106.915 -1.195 107.245 ;
        RECT -1.525 105.425 -1.195 105.755 ;
        RECT -1.525 104.015 -1.195 104.345 ;
        RECT -1.525 102.175 -1.195 102.505 ;
        RECT -1.525 100.685 -1.195 101.015 ;
        RECT -1.525 99.015 -1.195 99.345 ;
        RECT -1.525 97.525 -1.195 97.855 ;
        RECT -1.525 95.855 -1.195 96.185 ;
        RECT -1.525 94.365 -1.195 94.695 ;
        RECT -1.525 92.695 -1.195 93.025 ;
        RECT -1.525 91.205 -1.195 91.535 ;
        RECT -1.525 89.795 -1.195 90.125 ;
        RECT -1.525 87.955 -1.195 88.285 ;
        RECT -1.525 86.465 -1.195 86.795 ;
        RECT -1.525 84.795 -1.195 85.125 ;
        RECT -1.525 83.305 -1.195 83.635 ;
        RECT -1.525 81.635 -1.195 81.965 ;
        RECT -1.525 80.145 -1.195 80.475 ;
        RECT -1.525 78.475 -1.195 78.805 ;
        RECT -1.525 76.985 -1.195 77.315 ;
        RECT -1.525 75.575 -1.195 75.905 ;
        RECT -1.525 73.735 -1.195 74.065 ;
        RECT -1.525 72.245 -1.195 72.575 ;
        RECT -1.525 70.575 -1.195 70.905 ;
        RECT -1.525 69.085 -1.195 69.415 ;
        RECT -1.525 67.415 -1.195 67.745 ;
        RECT -1.525 65.925 -1.195 66.255 ;
        RECT -1.525 64.255 -1.195 64.585 ;
        RECT -1.525 62.765 -1.195 63.095 ;
        RECT -1.525 61.355 -1.195 61.685 ;
        RECT -1.525 59.515 -1.195 59.845 ;
        RECT -1.525 58.025 -1.195 58.355 ;
        RECT -1.525 56.355 -1.195 56.685 ;
        RECT -1.525 54.865 -1.195 55.195 ;
        RECT -1.525 53.195 -1.195 53.525 ;
        RECT -1.525 51.705 -1.195 52.035 ;
        RECT -1.525 50.035 -1.195 50.365 ;
        RECT -1.525 48.545 -1.195 48.875 ;
        RECT -1.525 47.135 -1.195 47.465 ;
        RECT -1.525 45.295 -1.195 45.625 ;
        RECT -1.525 43.805 -1.195 44.135 ;
        RECT -1.525 42.135 -1.195 42.465 ;
        RECT -1.525 40.645 -1.195 40.975 ;
        RECT -1.525 38.975 -1.195 39.305 ;
        RECT -1.525 37.485 -1.195 37.815 ;
        RECT -1.525 35.815 -1.195 36.145 ;
        RECT -1.525 34.325 -1.195 34.655 ;
        RECT -1.525 32.915 -1.195 33.245 ;
        RECT -1.525 31.075 -1.195 31.405 ;
        RECT -1.525 29.585 -1.195 29.915 ;
        RECT -1.525 27.915 -1.195 28.245 ;
        RECT -1.525 26.425 -1.195 26.755 ;
        RECT -1.525 24.755 -1.195 25.085 ;
        RECT -1.525 23.265 -1.195 23.595 ;
        RECT -1.525 21.595 -1.195 21.925 ;
        RECT -1.525 20.105 -1.195 20.435 ;
        RECT -1.525 18.695 -1.195 19.025 ;
        RECT -1.525 16.855 -1.195 17.185 ;
        RECT -1.525 15.365 -1.195 15.695 ;
        RECT -1.525 13.695 -1.195 14.025 ;
        RECT -1.525 12.205 -1.195 12.535 ;
        RECT -1.525 10.535 -1.195 10.865 ;
        RECT -1.525 9.045 -1.195 9.375 ;
        RECT -1.525 7.375 -1.195 7.705 ;
        RECT -1.525 5.885 -1.195 6.215 ;
        RECT -1.525 4.475 -1.195 4.805 ;
        RECT -1.525 2.115 -1.195 2.445 ;
        RECT -1.525 0.06 -1.195 0.39 ;
        RECT -1.525 -1.525 -1.195 -1.195 ;
        RECT -1.525 -2.885 -1.195 -2.555 ;
        RECT -1.525 -4.245 -1.195 -3.915 ;
        RECT -1.525 -5.605 -1.195 -5.275 ;
        RECT -1.525 -6.965 -1.195 -6.635 ;
        RECT -1.525 -8.325 -1.195 -7.995 ;
        RECT -1.525 -9.685 -1.195 -9.355 ;
        RECT -1.525 -12.405 -1.195 -12.075 ;
        RECT -1.525 -13.765 -1.195 -13.435 ;
        RECT -1.525 -15.125 -1.195 -14.795 ;
        RECT -1.525 -16.485 -1.195 -16.155 ;
        RECT -1.525 -17.845 -1.195 -17.515 ;
        RECT -1.525 -21.925 -1.195 -21.595 ;
        RECT -1.525 -23.285 -1.195 -22.955 ;
        RECT -1.525 -24.645 -1.195 -24.315 ;
        RECT -1.525 -26.005 -1.195 -25.675 ;
        RECT -1.525 -27.365 -1.195 -27.035 ;
        RECT -1.525 -28.725 -1.195 -28.395 ;
        RECT -1.525 -30.085 -1.195 -29.755 ;
        RECT -1.525 -31.445 -1.195 -31.115 ;
        RECT -1.525 -34.165 -1.195 -33.835 ;
        RECT -1.525 -35.525 -1.195 -35.195 ;
        RECT -1.525 -36.885 -1.195 -36.555 ;
        RECT -1.525 -38.245 -1.195 -37.915 ;
        RECT -1.525 -40.965 -1.195 -40.635 ;
        RECT -1.525 -42.325 -1.195 -41.995 ;
        RECT -1.525 -43.685 -1.195 -43.355 ;
        RECT -1.525 -45.045 -1.195 -44.715 ;
        RECT -1.525 -49.125 -1.195 -48.795 ;
        RECT -1.525 -50.485 -1.195 -50.155 ;
        RECT -1.525 -51.845 -1.195 -51.515 ;
        RECT -1.525 -53.205 -1.195 -52.875 ;
        RECT -1.525 -54.565 -1.195 -54.235 ;
        RECT -1.525 -55.925 -1.195 -55.595 ;
        RECT -1.525 -57.285 -1.195 -56.955 ;
        RECT -1.525 -58.645 -1.195 -58.315 ;
        RECT -1.525 -60.005 -1.195 -59.675 ;
        RECT -1.525 -61.365 -1.195 -61.035 ;
        RECT -1.525 -62.725 -1.195 -62.395 ;
        RECT -1.525 -64.085 -1.195 -63.755 ;
        RECT -1.525 -65.445 -1.195 -65.115 ;
        RECT -1.525 -66.805 -1.195 -66.475 ;
        RECT -1.525 -68.165 -1.195 -67.835 ;
        RECT -1.525 -69.525 -1.195 -69.195 ;
        RECT -1.525 -70.885 -1.195 -70.555 ;
        RECT -1.525 -72.245 -1.195 -71.915 ;
        RECT -1.525 -73.605 -1.195 -73.275 ;
        RECT -1.525 -74.965 -1.195 -74.635 ;
        RECT -1.525 -76.325 -1.195 -75.995 ;
        RECT -1.525 -77.685 -1.195 -77.355 ;
        RECT -1.525 -79.045 -1.195 -78.715 ;
        RECT -1.525 -80.405 -1.195 -80.075 ;
        RECT -1.525 -81.765 -1.195 -81.435 ;
        RECT -1.525 -83.125 -1.195 -82.795 ;
        RECT -1.525 -84.485 -1.195 -84.155 ;
        RECT -1.525 -85.845 -1.195 -85.515 ;
        RECT -1.525 -87.205 -1.195 -86.875 ;
        RECT -1.525 -88.565 -1.195 -88.235 ;
        RECT -1.525 -89.925 -1.195 -89.595 ;
        RECT -1.525 -91.285 -1.195 -90.955 ;
        RECT -1.525 -92.645 -1.195 -92.315 ;
        RECT -1.525 -94.005 -1.195 -93.675 ;
        RECT -1.525 -95.365 -1.195 -95.035 ;
        RECT -1.525 -96.725 -1.195 -96.395 ;
        RECT -1.525 -98.085 -1.195 -97.755 ;
        RECT -1.525 -99.445 -1.195 -99.115 ;
        RECT -1.525 -100.805 -1.195 -100.475 ;
        RECT -1.525 -102.165 -1.195 -101.835 ;
        RECT -1.525 -103.525 -1.195 -103.195 ;
        RECT -1.525 -104.885 -1.195 -104.555 ;
        RECT -1.525 -106.245 -1.195 -105.915 ;
        RECT -1.525 -107.605 -1.195 -107.275 ;
        RECT -1.525 -108.965 -1.195 -108.635 ;
        RECT -1.525 -110.325 -1.195 -109.995 ;
        RECT -1.525 -111.685 -1.195 -111.355 ;
        RECT -1.525 -113.045 -1.195 -112.715 ;
        RECT -1.525 -114.405 -1.195 -114.075 ;
        RECT -1.525 -115.765 -1.195 -115.435 ;
        RECT -1.525 -117.125 -1.195 -116.795 ;
        RECT -1.525 -118.485 -1.195 -118.155 ;
        RECT -1.525 -119.845 -1.195 -119.515 ;
        RECT -1.525 -121.205 -1.195 -120.875 ;
        RECT -1.525 -122.565 -1.195 -122.235 ;
        RECT -1.525 -123.925 -1.195 -123.595 ;
        RECT -1.525 -125.285 -1.195 -124.955 ;
        RECT -1.525 -126.645 -1.195 -126.315 ;
        RECT -1.525 -128.005 -1.195 -127.675 ;
        RECT -1.525 -129.365 -1.195 -129.035 ;
        RECT -1.525 -130.725 -1.195 -130.395 ;
        RECT -1.525 -132.085 -1.195 -131.755 ;
        RECT -1.525 -133.445 -1.195 -133.115 ;
        RECT -1.525 -134.805 -1.195 -134.475 ;
        RECT -1.525 -136.165 -1.195 -135.835 ;
        RECT -1.525 -137.525 -1.195 -137.195 ;
        RECT -1.525 -138.885 -1.195 -138.555 ;
        RECT -1.525 -140.245 -1.195 -139.915 ;
        RECT -1.525 -141.605 -1.195 -141.275 ;
        RECT -1.525 -142.965 -1.195 -142.635 ;
        RECT -1.525 -144.325 -1.195 -143.995 ;
        RECT -1.525 -145.685 -1.195 -145.355 ;
        RECT -1.525 -147.045 -1.195 -146.715 ;
        RECT -1.525 -148.405 -1.195 -148.075 ;
        RECT -1.525 -149.765 -1.195 -149.435 ;
        RECT -1.525 -151.125 -1.195 -150.795 ;
        RECT -1.525 -152.485 -1.195 -152.155 ;
        RECT -1.525 -153.845 -1.195 -153.515 ;
        RECT -1.525 -155.205 -1.195 -154.875 ;
        RECT -1.525 -156.565 -1.195 -156.235 ;
        RECT -1.525 -157.925 -1.195 -157.595 ;
        RECT -1.525 -160.17 -1.195 -159.04 ;
        RECT -1.52 -160.285 -1.2 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 127.225 0.165 128.355 ;
        RECT -0.165 124.955 0.165 125.285 ;
        RECT -0.165 123.595 0.165 123.925 ;
        RECT -0.16 123.595 0.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -1.525 0.165 -1.195 ;
        RECT -0.165 -2.885 0.165 -2.555 ;
        RECT -0.16 -3.56 0.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -91.285 0.165 -90.955 ;
        RECT -0.165 -92.645 0.165 -92.315 ;
        RECT -0.165 -94.005 0.165 -93.675 ;
        RECT -0.165 -95.365 0.165 -95.035 ;
        RECT -0.165 -96.725 0.165 -96.395 ;
        RECT -0.165 -98.085 0.165 -97.755 ;
        RECT -0.165 -99.445 0.165 -99.115 ;
        RECT -0.165 -100.805 0.165 -100.475 ;
        RECT -0.165 -102.165 0.165 -101.835 ;
        RECT -0.165 -103.525 0.165 -103.195 ;
        RECT -0.165 -104.885 0.165 -104.555 ;
        RECT -0.165 -106.245 0.165 -105.915 ;
        RECT -0.165 -107.605 0.165 -107.275 ;
        RECT -0.165 -108.965 0.165 -108.635 ;
        RECT -0.165 -110.325 0.165 -109.995 ;
        RECT -0.165 -111.685 0.165 -111.355 ;
        RECT -0.165 -113.045 0.165 -112.715 ;
        RECT -0.165 -114.405 0.165 -114.075 ;
        RECT -0.165 -115.765 0.165 -115.435 ;
        RECT -0.165 -117.125 0.165 -116.795 ;
        RECT -0.165 -118.485 0.165 -118.155 ;
        RECT -0.165 -119.845 0.165 -119.515 ;
        RECT -0.165 -121.205 0.165 -120.875 ;
        RECT -0.165 -122.565 0.165 -122.235 ;
        RECT -0.165 -123.925 0.165 -123.595 ;
        RECT -0.165 -125.285 0.165 -124.955 ;
        RECT -0.165 -126.645 0.165 -126.315 ;
        RECT -0.165 -128.005 0.165 -127.675 ;
        RECT -0.165 -129.365 0.165 -129.035 ;
        RECT -0.165 -130.725 0.165 -130.395 ;
        RECT -0.165 -132.085 0.165 -131.755 ;
        RECT -0.165 -133.445 0.165 -133.115 ;
        RECT -0.165 -134.805 0.165 -134.475 ;
        RECT -0.165 -136.165 0.165 -135.835 ;
        RECT -0.165 -137.525 0.165 -137.195 ;
        RECT -0.165 -138.885 0.165 -138.555 ;
        RECT -0.165 -140.245 0.165 -139.915 ;
        RECT -0.165 -141.605 0.165 -141.275 ;
        RECT -0.165 -142.965 0.165 -142.635 ;
        RECT -0.165 -144.325 0.165 -143.995 ;
        RECT -0.165 -145.685 0.165 -145.355 ;
        RECT -0.165 -147.045 0.165 -146.715 ;
        RECT -0.165 -148.405 0.165 -148.075 ;
        RECT -0.165 -149.765 0.165 -149.435 ;
        RECT -0.165 -151.125 0.165 -150.795 ;
        RECT -0.165 -152.485 0.165 -152.155 ;
        RECT -0.165 -153.845 0.165 -153.515 ;
        RECT -0.165 -155.205 0.165 -154.875 ;
        RECT -0.165 -156.565 0.165 -156.235 ;
        RECT -0.165 -157.925 0.165 -157.595 ;
        RECT -0.165 -160.17 0.165 -159.04 ;
        RECT -0.16 -160.285 0.16 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 127.225 1.525 128.355 ;
        RECT 1.195 124.955 1.525 125.285 ;
        RECT 1.195 123.595 1.525 123.925 ;
        RECT 1.2 123.595 1.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -1.525 1.525 -1.195 ;
        RECT 1.195 -2.885 1.525 -2.555 ;
        RECT 1.2 -3.56 1.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -91.285 1.525 -90.955 ;
        RECT 1.195 -92.645 1.525 -92.315 ;
        RECT 1.195 -94.005 1.525 -93.675 ;
        RECT 1.195 -95.365 1.525 -95.035 ;
        RECT 1.195 -96.725 1.525 -96.395 ;
        RECT 1.195 -98.085 1.525 -97.755 ;
        RECT 1.195 -99.445 1.525 -99.115 ;
        RECT 1.195 -100.805 1.525 -100.475 ;
        RECT 1.195 -102.165 1.525 -101.835 ;
        RECT 1.195 -103.525 1.525 -103.195 ;
        RECT 1.195 -104.885 1.525 -104.555 ;
        RECT 1.195 -106.245 1.525 -105.915 ;
        RECT 1.195 -107.605 1.525 -107.275 ;
        RECT 1.195 -108.965 1.525 -108.635 ;
        RECT 1.195 -110.325 1.525 -109.995 ;
        RECT 1.195 -111.685 1.525 -111.355 ;
        RECT 1.195 -113.045 1.525 -112.715 ;
        RECT 1.195 -114.405 1.525 -114.075 ;
        RECT 1.195 -115.765 1.525 -115.435 ;
        RECT 1.195 -117.125 1.525 -116.795 ;
        RECT 1.195 -118.485 1.525 -118.155 ;
        RECT 1.195 -119.845 1.525 -119.515 ;
        RECT 1.195 -121.205 1.525 -120.875 ;
        RECT 1.195 -122.565 1.525 -122.235 ;
        RECT 1.195 -123.925 1.525 -123.595 ;
        RECT 1.195 -125.285 1.525 -124.955 ;
        RECT 1.195 -126.645 1.525 -126.315 ;
        RECT 1.195 -128.005 1.525 -127.675 ;
        RECT 1.195 -129.365 1.525 -129.035 ;
        RECT 1.195 -130.725 1.525 -130.395 ;
        RECT 1.195 -132.085 1.525 -131.755 ;
        RECT 1.195 -133.445 1.525 -133.115 ;
        RECT 1.195 -134.805 1.525 -134.475 ;
        RECT 1.195 -136.165 1.525 -135.835 ;
        RECT 1.195 -137.525 1.525 -137.195 ;
        RECT 1.195 -138.885 1.525 -138.555 ;
        RECT 1.195 -140.245 1.525 -139.915 ;
        RECT 1.195 -141.605 1.525 -141.275 ;
        RECT 1.195 -142.965 1.525 -142.635 ;
        RECT 1.195 -144.325 1.525 -143.995 ;
        RECT 1.195 -145.685 1.525 -145.355 ;
        RECT 1.195 -147.045 1.525 -146.715 ;
        RECT 1.195 -148.405 1.525 -148.075 ;
        RECT 1.195 -149.765 1.525 -149.435 ;
        RECT 1.195 -151.125 1.525 -150.795 ;
        RECT 1.195 -152.485 1.525 -152.155 ;
        RECT 1.195 -153.845 1.525 -153.515 ;
        RECT 1.195 -155.205 1.525 -154.875 ;
        RECT 1.195 -156.565 1.525 -156.235 ;
        RECT 1.195 -157.925 1.525 -157.595 ;
        RECT 1.195 -160.17 1.525 -159.04 ;
        RECT 1.2 -160.285 1.52 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 127.225 2.885 128.355 ;
        RECT 2.555 124.955 2.885 125.285 ;
        RECT 2.555 123.595 2.885 123.925 ;
        RECT 2.56 123.595 2.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 -95.365 2.885 -95.035 ;
        RECT 2.555 -96.725 2.885 -96.395 ;
        RECT 2.555 -98.085 2.885 -97.755 ;
        RECT 2.555 -99.445 2.885 -99.115 ;
        RECT 2.555 -100.805 2.885 -100.475 ;
        RECT 2.555 -102.165 2.885 -101.835 ;
        RECT 2.555 -103.525 2.885 -103.195 ;
        RECT 2.555 -104.885 2.885 -104.555 ;
        RECT 2.555 -106.245 2.885 -105.915 ;
        RECT 2.555 -107.605 2.885 -107.275 ;
        RECT 2.555 -108.965 2.885 -108.635 ;
        RECT 2.555 -110.325 2.885 -109.995 ;
        RECT 2.555 -111.685 2.885 -111.355 ;
        RECT 2.555 -113.045 2.885 -112.715 ;
        RECT 2.555 -114.405 2.885 -114.075 ;
        RECT 2.555 -115.765 2.885 -115.435 ;
        RECT 2.555 -117.125 2.885 -116.795 ;
        RECT 2.555 -118.485 2.885 -118.155 ;
        RECT 2.555 -119.845 2.885 -119.515 ;
        RECT 2.555 -121.205 2.885 -120.875 ;
        RECT 2.555 -122.565 2.885 -122.235 ;
        RECT 2.555 -123.925 2.885 -123.595 ;
        RECT 2.555 -125.285 2.885 -124.955 ;
        RECT 2.555 -126.645 2.885 -126.315 ;
        RECT 2.555 -128.005 2.885 -127.675 ;
        RECT 2.555 -129.365 2.885 -129.035 ;
        RECT 2.555 -130.725 2.885 -130.395 ;
        RECT 2.555 -132.085 2.885 -131.755 ;
        RECT 2.555 -133.445 2.885 -133.115 ;
        RECT 2.555 -134.805 2.885 -134.475 ;
        RECT 2.555 -136.165 2.885 -135.835 ;
        RECT 2.555 -137.525 2.885 -137.195 ;
        RECT 2.555 -138.885 2.885 -138.555 ;
        RECT 2.555 -140.245 2.885 -139.915 ;
        RECT 2.555 -141.605 2.885 -141.275 ;
        RECT 2.555 -142.965 2.885 -142.635 ;
        RECT 2.555 -144.325 2.885 -143.995 ;
        RECT 2.555 -145.685 2.885 -145.355 ;
        RECT 2.555 -147.045 2.885 -146.715 ;
        RECT 2.555 -148.405 2.885 -148.075 ;
        RECT 2.555 -149.765 2.885 -149.435 ;
        RECT 2.555 -151.125 2.885 -150.795 ;
        RECT 2.555 -152.485 2.885 -152.155 ;
        RECT 2.555 -153.845 2.885 -153.515 ;
        RECT 2.555 -155.205 2.885 -154.875 ;
        RECT 2.555 -156.565 2.885 -156.235 ;
        RECT 2.555 -157.925 2.885 -157.595 ;
        RECT 2.555 -160.17 2.885 -159.04 ;
        RECT 2.56 -160.285 2.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.31 -94.075 3.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 127.225 4.245 128.355 ;
        RECT 3.915 124.955 4.245 125.285 ;
        RECT 3.915 123.595 4.245 123.925 ;
        RECT 3.92 123.595 4.24 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 127.225 5.605 128.355 ;
        RECT 5.275 124.955 5.605 125.285 ;
        RECT 5.275 123.595 5.605 123.925 ;
        RECT 5.28 123.595 5.6 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 -1.525 5.605 -1.195 ;
        RECT 5.275 -2.885 5.605 -2.555 ;
        RECT 5.28 -3.56 5.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 127.225 6.965 128.355 ;
        RECT 6.635 124.955 6.965 125.285 ;
        RECT 6.635 123.595 6.965 123.925 ;
        RECT 6.64 123.595 6.96 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 -1.525 6.965 -1.195 ;
        RECT 6.635 -2.885 6.965 -2.555 ;
        RECT 6.64 -3.56 6.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 127.225 8.325 128.355 ;
        RECT 7.995 124.955 8.325 125.285 ;
        RECT 7.995 123.595 8.325 123.925 ;
        RECT 8 123.595 8.32 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -1.525 8.325 -1.195 ;
        RECT 7.995 -2.885 8.325 -2.555 ;
        RECT 8 -3.56 8.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -91.285 8.325 -90.955 ;
        RECT 7.995 -92.645 8.325 -92.315 ;
        RECT 7.995 -94.005 8.325 -93.675 ;
        RECT 7.995 -95.365 8.325 -95.035 ;
        RECT 7.995 -96.725 8.325 -96.395 ;
        RECT 7.995 -98.085 8.325 -97.755 ;
        RECT 7.995 -99.445 8.325 -99.115 ;
        RECT 7.995 -100.805 8.325 -100.475 ;
        RECT 7.995 -102.165 8.325 -101.835 ;
        RECT 7.995 -103.525 8.325 -103.195 ;
        RECT 7.995 -104.885 8.325 -104.555 ;
        RECT 7.995 -106.245 8.325 -105.915 ;
        RECT 7.995 -107.605 8.325 -107.275 ;
        RECT 7.995 -108.965 8.325 -108.635 ;
        RECT 7.995 -110.325 8.325 -109.995 ;
        RECT 7.995 -111.685 8.325 -111.355 ;
        RECT 7.995 -113.045 8.325 -112.715 ;
        RECT 7.995 -114.405 8.325 -114.075 ;
        RECT 7.995 -115.765 8.325 -115.435 ;
        RECT 7.995 -117.125 8.325 -116.795 ;
        RECT 7.995 -118.485 8.325 -118.155 ;
        RECT 7.995 -119.845 8.325 -119.515 ;
        RECT 7.995 -121.205 8.325 -120.875 ;
        RECT 7.995 -122.565 8.325 -122.235 ;
        RECT 7.995 -123.925 8.325 -123.595 ;
        RECT 7.995 -125.285 8.325 -124.955 ;
        RECT 7.995 -126.645 8.325 -126.315 ;
        RECT 7.995 -128.005 8.325 -127.675 ;
        RECT 7.995 -129.365 8.325 -129.035 ;
        RECT 7.995 -130.725 8.325 -130.395 ;
        RECT 7.995 -132.085 8.325 -131.755 ;
        RECT 7.995 -133.445 8.325 -133.115 ;
        RECT 7.995 -134.805 8.325 -134.475 ;
        RECT 7.995 -136.165 8.325 -135.835 ;
        RECT 7.995 -137.525 8.325 -137.195 ;
        RECT 7.995 -138.885 8.325 -138.555 ;
        RECT 7.995 -140.245 8.325 -139.915 ;
        RECT 7.995 -141.605 8.325 -141.275 ;
        RECT 7.995 -142.965 8.325 -142.635 ;
        RECT 7.995 -144.325 8.325 -143.995 ;
        RECT 7.995 -145.685 8.325 -145.355 ;
        RECT 7.995 -147.045 8.325 -146.715 ;
        RECT 7.995 -148.405 8.325 -148.075 ;
        RECT 7.995 -149.765 8.325 -149.435 ;
        RECT 7.995 -151.125 8.325 -150.795 ;
        RECT 7.995 -152.485 8.325 -152.155 ;
        RECT 7.995 -153.845 8.325 -153.515 ;
        RECT 7.995 -155.205 8.325 -154.875 ;
        RECT 7.995 -156.565 8.325 -156.235 ;
        RECT 7.995 -157.925 8.325 -157.595 ;
        RECT 7.995 -160.17 8.325 -159.04 ;
        RECT 8 -160.285 8.32 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 127.225 9.685 128.355 ;
        RECT 9.355 124.955 9.685 125.285 ;
        RECT 9.355 123.595 9.685 123.925 ;
        RECT 9.36 123.595 9.68 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 -95.365 9.685 -95.035 ;
        RECT 9.355 -96.725 9.685 -96.395 ;
        RECT 9.355 -98.085 9.685 -97.755 ;
        RECT 9.355 -99.445 9.685 -99.115 ;
        RECT 9.355 -100.805 9.685 -100.475 ;
        RECT 9.355 -102.165 9.685 -101.835 ;
        RECT 9.355 -103.525 9.685 -103.195 ;
        RECT 9.355 -104.885 9.685 -104.555 ;
        RECT 9.355 -106.245 9.685 -105.915 ;
        RECT 9.355 -107.605 9.685 -107.275 ;
        RECT 9.355 -108.965 9.685 -108.635 ;
        RECT 9.355 -110.325 9.685 -109.995 ;
        RECT 9.355 -111.685 9.685 -111.355 ;
        RECT 9.355 -113.045 9.685 -112.715 ;
        RECT 9.355 -114.405 9.685 -114.075 ;
        RECT 9.355 -115.765 9.685 -115.435 ;
        RECT 9.355 -117.125 9.685 -116.795 ;
        RECT 9.355 -118.485 9.685 -118.155 ;
        RECT 9.355 -119.845 9.685 -119.515 ;
        RECT 9.355 -121.205 9.685 -120.875 ;
        RECT 9.355 -122.565 9.685 -122.235 ;
        RECT 9.355 -123.925 9.685 -123.595 ;
        RECT 9.355 -125.285 9.685 -124.955 ;
        RECT 9.355 -126.645 9.685 -126.315 ;
        RECT 9.355 -128.005 9.685 -127.675 ;
        RECT 9.355 -129.365 9.685 -129.035 ;
        RECT 9.355 -130.725 9.685 -130.395 ;
        RECT 9.355 -132.085 9.685 -131.755 ;
        RECT 9.355 -133.445 9.685 -133.115 ;
        RECT 9.355 -134.805 9.685 -134.475 ;
        RECT 9.355 -136.165 9.685 -135.835 ;
        RECT 9.355 -137.525 9.685 -137.195 ;
        RECT 9.355 -138.885 9.685 -138.555 ;
        RECT 9.355 -140.245 9.685 -139.915 ;
        RECT 9.355 -141.605 9.685 -141.275 ;
        RECT 9.355 -142.965 9.685 -142.635 ;
        RECT 9.355 -144.325 9.685 -143.995 ;
        RECT 9.355 -145.685 9.685 -145.355 ;
        RECT 9.355 -147.045 9.685 -146.715 ;
        RECT 9.355 -148.405 9.685 -148.075 ;
        RECT 9.355 -149.765 9.685 -149.435 ;
        RECT 9.355 -151.125 9.685 -150.795 ;
        RECT 9.355 -152.485 9.685 -152.155 ;
        RECT 9.355 -153.845 9.685 -153.515 ;
        RECT 9.355 -155.205 9.685 -154.875 ;
        RECT 9.355 -156.565 9.685 -156.235 ;
        RECT 9.355 -157.925 9.685 -157.595 ;
        RECT 9.355 -160.17 9.685 -159.04 ;
        RECT 9.36 -160.285 9.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.41 -94.075 9.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 127.225 11.045 128.355 ;
        RECT 10.715 124.955 11.045 125.285 ;
        RECT 10.715 123.595 11.045 123.925 ;
        RECT 10.72 123.595 11.04 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -1.525 11.045 -1.195 ;
        RECT 10.715 -2.885 11.045 -2.555 ;
        RECT 10.72 -3.56 11.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 127.225 12.405 128.355 ;
        RECT 12.075 124.955 12.405 125.285 ;
        RECT 12.075 123.595 12.405 123.925 ;
        RECT 12.08 123.595 12.4 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 -1.525 12.405 -1.195 ;
        RECT 12.075 -2.885 12.405 -2.555 ;
        RECT 12.08 -3.56 12.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 127.225 13.765 128.355 ;
        RECT 13.435 124.955 13.765 125.285 ;
        RECT 13.435 123.595 13.765 123.925 ;
        RECT 13.44 123.595 13.76 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -1.525 13.765 -1.195 ;
        RECT 13.435 -2.885 13.765 -2.555 ;
        RECT 13.44 -3.56 13.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -91.285 13.765 -90.955 ;
        RECT 13.435 -92.645 13.765 -92.315 ;
        RECT 13.435 -94.005 13.765 -93.675 ;
        RECT 13.435 -95.365 13.765 -95.035 ;
        RECT 13.435 -96.725 13.765 -96.395 ;
        RECT 13.435 -98.085 13.765 -97.755 ;
        RECT 13.435 -99.445 13.765 -99.115 ;
        RECT 13.435 -100.805 13.765 -100.475 ;
        RECT 13.435 -102.165 13.765 -101.835 ;
        RECT 13.435 -103.525 13.765 -103.195 ;
        RECT 13.435 -104.885 13.765 -104.555 ;
        RECT 13.435 -106.245 13.765 -105.915 ;
        RECT 13.435 -107.605 13.765 -107.275 ;
        RECT 13.435 -108.965 13.765 -108.635 ;
        RECT 13.435 -110.325 13.765 -109.995 ;
        RECT 13.435 -111.685 13.765 -111.355 ;
        RECT 13.435 -113.045 13.765 -112.715 ;
        RECT 13.435 -114.405 13.765 -114.075 ;
        RECT 13.435 -115.765 13.765 -115.435 ;
        RECT 13.435 -117.125 13.765 -116.795 ;
        RECT 13.435 -118.485 13.765 -118.155 ;
        RECT 13.435 -119.845 13.765 -119.515 ;
        RECT 13.435 -121.205 13.765 -120.875 ;
        RECT 13.435 -122.565 13.765 -122.235 ;
        RECT 13.435 -123.925 13.765 -123.595 ;
        RECT 13.435 -125.285 13.765 -124.955 ;
        RECT 13.435 -126.645 13.765 -126.315 ;
        RECT 13.435 -128.005 13.765 -127.675 ;
        RECT 13.435 -129.365 13.765 -129.035 ;
        RECT 13.435 -130.725 13.765 -130.395 ;
        RECT 13.435 -132.085 13.765 -131.755 ;
        RECT 13.435 -133.445 13.765 -133.115 ;
        RECT 13.435 -134.805 13.765 -134.475 ;
        RECT 13.435 -136.165 13.765 -135.835 ;
        RECT 13.435 -137.525 13.765 -137.195 ;
        RECT 13.435 -138.885 13.765 -138.555 ;
        RECT 13.435 -140.245 13.765 -139.915 ;
        RECT 13.435 -141.605 13.765 -141.275 ;
        RECT 13.435 -142.965 13.765 -142.635 ;
        RECT 13.435 -144.325 13.765 -143.995 ;
        RECT 13.435 -145.685 13.765 -145.355 ;
        RECT 13.435 -147.045 13.765 -146.715 ;
        RECT 13.435 -148.405 13.765 -148.075 ;
        RECT 13.435 -149.765 13.765 -149.435 ;
        RECT 13.435 -151.125 13.765 -150.795 ;
        RECT 13.435 -152.485 13.765 -152.155 ;
        RECT 13.435 -153.845 13.765 -153.515 ;
        RECT 13.435 -155.205 13.765 -154.875 ;
        RECT 13.435 -156.565 13.765 -156.235 ;
        RECT 13.435 -157.925 13.765 -157.595 ;
        RECT 13.435 -160.17 13.765 -159.04 ;
        RECT 13.44 -160.285 13.76 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 127.225 15.125 128.355 ;
        RECT 14.795 124.955 15.125 125.285 ;
        RECT 14.795 123.595 15.125 123.925 ;
        RECT 14.8 123.595 15.12 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 -95.365 15.125 -95.035 ;
        RECT 14.795 -96.725 15.125 -96.395 ;
        RECT 14.795 -98.085 15.125 -97.755 ;
        RECT 14.795 -99.445 15.125 -99.115 ;
        RECT 14.795 -100.805 15.125 -100.475 ;
        RECT 14.795 -102.165 15.125 -101.835 ;
        RECT 14.795 -103.525 15.125 -103.195 ;
        RECT 14.795 -104.885 15.125 -104.555 ;
        RECT 14.795 -106.245 15.125 -105.915 ;
        RECT 14.795 -107.605 15.125 -107.275 ;
        RECT 14.795 -108.965 15.125 -108.635 ;
        RECT 14.795 -110.325 15.125 -109.995 ;
        RECT 14.795 -111.685 15.125 -111.355 ;
        RECT 14.795 -113.045 15.125 -112.715 ;
        RECT 14.795 -114.405 15.125 -114.075 ;
        RECT 14.795 -115.765 15.125 -115.435 ;
        RECT 14.795 -117.125 15.125 -116.795 ;
        RECT 14.795 -118.485 15.125 -118.155 ;
        RECT 14.795 -119.845 15.125 -119.515 ;
        RECT 14.795 -121.205 15.125 -120.875 ;
        RECT 14.795 -122.565 15.125 -122.235 ;
        RECT 14.795 -123.925 15.125 -123.595 ;
        RECT 14.795 -125.285 15.125 -124.955 ;
        RECT 14.795 -126.645 15.125 -126.315 ;
        RECT 14.795 -128.005 15.125 -127.675 ;
        RECT 14.795 -129.365 15.125 -129.035 ;
        RECT 14.795 -130.725 15.125 -130.395 ;
        RECT 14.795 -132.085 15.125 -131.755 ;
        RECT 14.795 -133.445 15.125 -133.115 ;
        RECT 14.795 -134.805 15.125 -134.475 ;
        RECT 14.795 -136.165 15.125 -135.835 ;
        RECT 14.795 -137.525 15.125 -137.195 ;
        RECT 14.795 -138.885 15.125 -138.555 ;
        RECT 14.795 -140.245 15.125 -139.915 ;
        RECT 14.795 -141.605 15.125 -141.275 ;
        RECT 14.795 -142.965 15.125 -142.635 ;
        RECT 14.795 -144.325 15.125 -143.995 ;
        RECT 14.795 -145.685 15.125 -145.355 ;
        RECT 14.795 -147.045 15.125 -146.715 ;
        RECT 14.795 -148.405 15.125 -148.075 ;
        RECT 14.795 -149.765 15.125 -149.435 ;
        RECT 14.795 -151.125 15.125 -150.795 ;
        RECT 14.795 -152.485 15.125 -152.155 ;
        RECT 14.795 -153.845 15.125 -153.515 ;
        RECT 14.795 -155.205 15.125 -154.875 ;
        RECT 14.795 -156.565 15.125 -156.235 ;
        RECT 14.795 -157.925 15.125 -157.595 ;
        RECT 14.795 -160.17 15.125 -159.04 ;
        RECT 14.8 -160.285 15.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.51 -94.075 15.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 127.225 16.485 128.355 ;
        RECT 16.155 124.955 16.485 125.285 ;
        RECT 16.155 123.595 16.485 123.925 ;
        RECT 16.16 123.595 16.48 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 127.225 17.845 128.355 ;
        RECT 17.515 124.955 17.845 125.285 ;
        RECT 17.515 123.595 17.845 123.925 ;
        RECT 17.52 123.595 17.84 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -1.525 17.845 -1.195 ;
        RECT 17.515 -2.885 17.845 -2.555 ;
        RECT 17.52 -3.56 17.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 127.225 19.205 128.355 ;
        RECT 18.875 124.955 19.205 125.285 ;
        RECT 18.875 123.595 19.205 123.925 ;
        RECT 18.88 123.595 19.2 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -1.525 19.205 -1.195 ;
        RECT 18.875 -2.885 19.205 -2.555 ;
        RECT 18.88 -3.56 19.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -91.285 19.205 -90.955 ;
        RECT 18.875 -92.645 19.205 -92.315 ;
        RECT 18.875 -94.005 19.205 -93.675 ;
        RECT 18.875 -95.365 19.205 -95.035 ;
        RECT 18.875 -96.725 19.205 -96.395 ;
        RECT 18.875 -98.085 19.205 -97.755 ;
        RECT 18.875 -99.445 19.205 -99.115 ;
        RECT 18.875 -100.805 19.205 -100.475 ;
        RECT 18.875 -102.165 19.205 -101.835 ;
        RECT 18.875 -103.525 19.205 -103.195 ;
        RECT 18.875 -104.885 19.205 -104.555 ;
        RECT 18.875 -106.245 19.205 -105.915 ;
        RECT 18.875 -107.605 19.205 -107.275 ;
        RECT 18.875 -108.965 19.205 -108.635 ;
        RECT 18.875 -110.325 19.205 -109.995 ;
        RECT 18.875 -111.685 19.205 -111.355 ;
        RECT 18.875 -113.045 19.205 -112.715 ;
        RECT 18.875 -114.405 19.205 -114.075 ;
        RECT 18.875 -115.765 19.205 -115.435 ;
        RECT 18.875 -117.125 19.205 -116.795 ;
        RECT 18.875 -118.485 19.205 -118.155 ;
        RECT 18.875 -119.845 19.205 -119.515 ;
        RECT 18.875 -121.205 19.205 -120.875 ;
        RECT 18.875 -122.565 19.205 -122.235 ;
        RECT 18.875 -123.925 19.205 -123.595 ;
        RECT 18.875 -125.285 19.205 -124.955 ;
        RECT 18.875 -126.645 19.205 -126.315 ;
        RECT 18.875 -128.005 19.205 -127.675 ;
        RECT 18.875 -129.365 19.205 -129.035 ;
        RECT 18.875 -130.725 19.205 -130.395 ;
        RECT 18.875 -132.085 19.205 -131.755 ;
        RECT 18.875 -133.445 19.205 -133.115 ;
        RECT 18.875 -134.805 19.205 -134.475 ;
        RECT 18.875 -136.165 19.205 -135.835 ;
        RECT 18.875 -137.525 19.205 -137.195 ;
        RECT 18.875 -138.885 19.205 -138.555 ;
        RECT 18.875 -140.245 19.205 -139.915 ;
        RECT 18.875 -141.605 19.205 -141.275 ;
        RECT 18.875 -142.965 19.205 -142.635 ;
        RECT 18.875 -144.325 19.205 -143.995 ;
        RECT 18.875 -145.685 19.205 -145.355 ;
        RECT 18.875 -147.045 19.205 -146.715 ;
        RECT 18.875 -148.405 19.205 -148.075 ;
        RECT 18.875 -149.765 19.205 -149.435 ;
        RECT 18.875 -151.125 19.205 -150.795 ;
        RECT 18.875 -152.485 19.205 -152.155 ;
        RECT 18.875 -153.845 19.205 -153.515 ;
        RECT 18.875 -155.205 19.205 -154.875 ;
        RECT 18.875 -156.565 19.205 -156.235 ;
        RECT 18.875 -157.925 19.205 -157.595 ;
        RECT 18.875 -160.17 19.205 -159.04 ;
        RECT 18.88 -160.285 19.2 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 127.225 20.565 128.355 ;
        RECT 20.235 124.955 20.565 125.285 ;
        RECT 20.235 123.595 20.565 123.925 ;
        RECT 20.24 123.595 20.56 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -1.525 20.565 -1.195 ;
        RECT 20.235 -2.885 20.565 -2.555 ;
        RECT 20.24 -3.56 20.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -91.285 20.565 -90.955 ;
        RECT 20.235 -92.645 20.565 -92.315 ;
        RECT 20.235 -94.005 20.565 -93.675 ;
        RECT 20.235 -95.365 20.565 -95.035 ;
        RECT 20.235 -96.725 20.565 -96.395 ;
        RECT 20.235 -98.085 20.565 -97.755 ;
        RECT 20.235 -99.445 20.565 -99.115 ;
        RECT 20.235 -100.805 20.565 -100.475 ;
        RECT 20.235 -102.165 20.565 -101.835 ;
        RECT 20.235 -103.525 20.565 -103.195 ;
        RECT 20.235 -104.885 20.565 -104.555 ;
        RECT 20.235 -106.245 20.565 -105.915 ;
        RECT 20.235 -107.605 20.565 -107.275 ;
        RECT 20.235 -108.965 20.565 -108.635 ;
        RECT 20.235 -110.325 20.565 -109.995 ;
        RECT 20.235 -111.685 20.565 -111.355 ;
        RECT 20.235 -113.045 20.565 -112.715 ;
        RECT 20.235 -114.405 20.565 -114.075 ;
        RECT 20.235 -115.765 20.565 -115.435 ;
        RECT 20.235 -117.125 20.565 -116.795 ;
        RECT 20.235 -118.485 20.565 -118.155 ;
        RECT 20.235 -119.845 20.565 -119.515 ;
        RECT 20.235 -121.205 20.565 -120.875 ;
        RECT 20.235 -122.565 20.565 -122.235 ;
        RECT 20.235 -123.925 20.565 -123.595 ;
        RECT 20.235 -125.285 20.565 -124.955 ;
        RECT 20.235 -126.645 20.565 -126.315 ;
        RECT 20.235 -128.005 20.565 -127.675 ;
        RECT 20.235 -129.365 20.565 -129.035 ;
        RECT 20.235 -130.725 20.565 -130.395 ;
        RECT 20.235 -132.085 20.565 -131.755 ;
        RECT 20.235 -133.445 20.565 -133.115 ;
        RECT 20.235 -134.805 20.565 -134.475 ;
        RECT 20.235 -136.165 20.565 -135.835 ;
        RECT 20.235 -137.525 20.565 -137.195 ;
        RECT 20.235 -138.885 20.565 -138.555 ;
        RECT 20.235 -140.245 20.565 -139.915 ;
        RECT 20.235 -141.605 20.565 -141.275 ;
        RECT 20.235 -142.965 20.565 -142.635 ;
        RECT 20.235 -144.325 20.565 -143.995 ;
        RECT 20.235 -145.685 20.565 -145.355 ;
        RECT 20.235 -147.045 20.565 -146.715 ;
        RECT 20.235 -148.405 20.565 -148.075 ;
        RECT 20.235 -149.765 20.565 -149.435 ;
        RECT 20.235 -151.125 20.565 -150.795 ;
        RECT 20.235 -152.485 20.565 -152.155 ;
        RECT 20.235 -153.845 20.565 -153.515 ;
        RECT 20.235 -155.205 20.565 -154.875 ;
        RECT 20.235 -156.565 20.565 -156.235 ;
        RECT 20.235 -157.925 20.565 -157.595 ;
        RECT 20.235 -160.17 20.565 -159.04 ;
        RECT 20.24 -160.285 20.56 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 127.225 21.925 128.355 ;
        RECT 21.595 124.955 21.925 125.285 ;
        RECT 21.595 123.595 21.925 123.925 ;
        RECT 21.6 123.595 21.92 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 -95.365 21.925 -95.035 ;
        RECT 21.595 -96.725 21.925 -96.395 ;
        RECT 21.595 -98.085 21.925 -97.755 ;
        RECT 21.595 -99.445 21.925 -99.115 ;
        RECT 21.595 -100.805 21.925 -100.475 ;
        RECT 21.595 -102.165 21.925 -101.835 ;
        RECT 21.595 -103.525 21.925 -103.195 ;
        RECT 21.595 -104.885 21.925 -104.555 ;
        RECT 21.595 -106.245 21.925 -105.915 ;
        RECT 21.595 -107.605 21.925 -107.275 ;
        RECT 21.595 -108.965 21.925 -108.635 ;
        RECT 21.595 -110.325 21.925 -109.995 ;
        RECT 21.595 -111.685 21.925 -111.355 ;
        RECT 21.595 -113.045 21.925 -112.715 ;
        RECT 21.595 -114.405 21.925 -114.075 ;
        RECT 21.595 -115.765 21.925 -115.435 ;
        RECT 21.595 -117.125 21.925 -116.795 ;
        RECT 21.595 -118.485 21.925 -118.155 ;
        RECT 21.595 -119.845 21.925 -119.515 ;
        RECT 21.595 -121.205 21.925 -120.875 ;
        RECT 21.595 -122.565 21.925 -122.235 ;
        RECT 21.595 -123.925 21.925 -123.595 ;
        RECT 21.595 -125.285 21.925 -124.955 ;
        RECT 21.595 -126.645 21.925 -126.315 ;
        RECT 21.595 -128.005 21.925 -127.675 ;
        RECT 21.595 -129.365 21.925 -129.035 ;
        RECT 21.595 -130.725 21.925 -130.395 ;
        RECT 21.595 -132.085 21.925 -131.755 ;
        RECT 21.595 -133.445 21.925 -133.115 ;
        RECT 21.595 -134.805 21.925 -134.475 ;
        RECT 21.595 -136.165 21.925 -135.835 ;
        RECT 21.595 -137.525 21.925 -137.195 ;
        RECT 21.595 -138.885 21.925 -138.555 ;
        RECT 21.595 -140.245 21.925 -139.915 ;
        RECT 21.595 -141.605 21.925 -141.275 ;
        RECT 21.595 -142.965 21.925 -142.635 ;
        RECT 21.595 -144.325 21.925 -143.995 ;
        RECT 21.595 -145.685 21.925 -145.355 ;
        RECT 21.595 -147.045 21.925 -146.715 ;
        RECT 21.595 -148.405 21.925 -148.075 ;
        RECT 21.595 -149.765 21.925 -149.435 ;
        RECT 21.595 -151.125 21.925 -150.795 ;
        RECT 21.595 -152.485 21.925 -152.155 ;
        RECT 21.595 -153.845 21.925 -153.515 ;
        RECT 21.595 -155.205 21.925 -154.875 ;
        RECT 21.595 -156.565 21.925 -156.235 ;
        RECT 21.595 -157.925 21.925 -157.595 ;
        RECT 21.595 -160.17 21.925 -159.04 ;
        RECT 21.6 -160.285 21.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.61 -94.075 21.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 127.225 23.285 128.355 ;
        RECT 22.955 124.955 23.285 125.285 ;
        RECT 22.955 123.595 23.285 123.925 ;
        RECT 22.96 123.595 23.28 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 -1.525 23.285 -1.195 ;
        RECT 22.955 -2.885 23.285 -2.555 ;
        RECT 22.96 -3.56 23.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 127.225 24.645 128.355 ;
        RECT 24.315 124.955 24.645 125.285 ;
        RECT 24.315 123.595 24.645 123.925 ;
        RECT 24.32 123.595 24.64 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 -1.525 24.645 -1.195 ;
        RECT 24.315 -2.885 24.645 -2.555 ;
        RECT 24.32 -3.56 24.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 127.225 26.005 128.355 ;
        RECT 25.675 124.955 26.005 125.285 ;
        RECT 25.675 123.595 26.005 123.925 ;
        RECT 25.68 123.595 26 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.68 -3.56 26 -0.52 ;
        RECT 25.675 -1.525 26.005 -1.195 ;
        RECT 25.675 -2.885 26.005 -2.555 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 -24.645 -12.075 -24.315 ;
        RECT -12.405 -26.005 -12.075 -25.675 ;
        RECT -12.405 -27.365 -12.075 -27.035 ;
        RECT -12.405 -28.725 -12.075 -28.395 ;
        RECT -12.405 -30.085 -12.075 -29.755 ;
        RECT -12.405 -34.165 -12.075 -33.835 ;
        RECT -12.405 -35.39 -12.075 -35.06 ;
        RECT -12.405 -38.245 -12.075 -37.915 ;
        RECT -12.405 -40.23 -12.075 -39.9 ;
        RECT -12.405 -40.965 -12.075 -40.635 ;
        RECT -12.405 -49.125 -12.075 -48.795 ;
        RECT -12.405 -50.485 -12.075 -50.155 ;
        RECT -12.405 -51.845 -12.075 -51.515 ;
        RECT -12.405 -54.565 -12.075 -54.235 ;
        RECT -12.405 -56.27 -12.075 -55.94 ;
        RECT -12.405 -57.285 -12.075 -56.955 ;
        RECT -12.405 -58.645 -12.075 -58.315 ;
        RECT -12.405 -61.365 -12.075 -61.035 ;
        RECT -12.405 -62.725 -12.075 -62.395 ;
        RECT -12.405 -64.085 -12.075 -63.755 ;
        RECT -12.405 -64.81 -12.075 -64.48 ;
        RECT -12.405 -66.805 -12.075 -66.475 ;
        RECT -12.405 -69.525 -12.075 -69.195 ;
        RECT -12.405 -70.885 -12.075 -70.555 ;
        RECT -12.405 -72.245 -12.075 -71.915 ;
        RECT -12.405 -73.605 -12.075 -73.275 ;
        RECT -12.405 -76.325 -12.075 -75.995 ;
        RECT -12.405 -77.685 -12.075 -77.355 ;
        RECT -12.405 -78.45 -12.075 -78.12 ;
        RECT -12.405 -80.405 -12.075 -80.075 ;
        RECT -12.405 -81.765 -12.075 -81.435 ;
        RECT -12.405 -84.485 -12.075 -84.155 ;
        RECT -12.405 -85.845 -12.075 -85.515 ;
        RECT -12.405 -86.99 -12.075 -86.66 ;
        RECT -12.405 -92.645 -12.075 -92.315 ;
        RECT -12.405 -94.005 -12.075 -93.675 ;
        RECT -12.405 -95.365 -12.075 -95.035 ;
        RECT -12.405 -96.725 -12.075 -96.395 ;
        RECT -12.405 -98.085 -12.075 -97.755 ;
        RECT -12.405 -99.445 -12.075 -99.115 ;
        RECT -12.405 -108.965 -12.075 -108.635 ;
        RECT -12.405 -113.045 -12.075 -112.715 ;
        RECT -12.405 -115.765 -12.075 -115.435 ;
        RECT -12.405 -118.485 -12.075 -118.155 ;
        RECT -12.405 -119.845 -12.075 -119.515 ;
        RECT -12.405 -121.205 -12.075 -120.875 ;
        RECT -12.405 -125.285 -12.075 -124.955 ;
        RECT -12.405 -126.645 -12.075 -126.315 ;
        RECT -12.405 -128.005 -12.075 -127.675 ;
        RECT -12.405 -129.365 -12.075 -129.035 ;
        RECT -12.405 -132.085 -12.075 -131.755 ;
        RECT -12.405 -133.445 -12.075 -133.115 ;
        RECT -12.405 -134.805 -12.075 -134.475 ;
        RECT -12.405 -136.165 -12.075 -135.835 ;
        RECT -12.405 -138.885 -12.075 -138.555 ;
        RECT -12.405 -140.245 -12.075 -139.915 ;
        RECT -12.405 -141.605 -12.075 -141.275 ;
        RECT -12.405 -142.965 -12.075 -142.635 ;
        RECT -12.405 -144.325 -12.075 -143.995 ;
        RECT -12.405 -145.685 -12.075 -145.355 ;
        RECT -12.405 -149.765 -12.075 -149.435 ;
        RECT -12.405 -152.485 -12.075 -152.155 ;
        RECT -12.405 -153.845 -12.075 -153.515 ;
        RECT -12.405 -155.285 -12.075 -154.955 ;
        RECT -12.405 -156.565 -12.075 -156.235 ;
        RECT -12.405 -157.925 -12.075 -157.595 ;
        RECT -12.405 -160.17 -12.075 -159.04 ;
        RECT -12.4 -160.285 -12.08 -23.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 127.225 -10.715 128.355 ;
        RECT -11.045 124.955 -10.715 125.285 ;
        RECT -11.045 123.595 -10.715 123.925 ;
        RECT -11.045 122.235 -10.715 122.565 ;
        RECT -11.045 120.875 -10.715 121.205 ;
        RECT -11.045 119.515 -10.715 119.845 ;
        RECT -11.045 118.155 -10.715 118.485 ;
        RECT -11.045 116.795 -10.715 117.125 ;
        RECT -11.045 115.435 -10.715 115.765 ;
        RECT -11.045 114.075 -10.715 114.405 ;
        RECT -11.045 112.715 -10.715 113.045 ;
        RECT -11.045 111.355 -10.715 111.685 ;
        RECT -11.045 109.995 -10.715 110.325 ;
        RECT -11.045 108.635 -10.715 108.965 ;
        RECT -11.045 107.275 -10.715 107.605 ;
        RECT -11.045 105.915 -10.715 106.245 ;
        RECT -11.045 104.555 -10.715 104.885 ;
        RECT -11.045 103.195 -10.715 103.525 ;
        RECT -11.045 101.835 -10.715 102.165 ;
        RECT -11.045 100.475 -10.715 100.805 ;
        RECT -11.045 99.115 -10.715 99.445 ;
        RECT -11.045 97.755 -10.715 98.085 ;
        RECT -11.045 96.395 -10.715 96.725 ;
        RECT -11.045 95.035 -10.715 95.365 ;
        RECT -11.045 93.675 -10.715 94.005 ;
        RECT -11.045 92.315 -10.715 92.645 ;
        RECT -11.045 90.955 -10.715 91.285 ;
        RECT -11.045 89.595 -10.715 89.925 ;
        RECT -11.045 88.235 -10.715 88.565 ;
        RECT -11.045 86.875 -10.715 87.205 ;
        RECT -11.045 85.515 -10.715 85.845 ;
        RECT -11.045 84.155 -10.715 84.485 ;
        RECT -11.045 82.795 -10.715 83.125 ;
        RECT -11.045 81.435 -10.715 81.765 ;
        RECT -11.045 80.075 -10.715 80.405 ;
        RECT -11.045 78.715 -10.715 79.045 ;
        RECT -11.045 77.355 -10.715 77.685 ;
        RECT -11.045 75.995 -10.715 76.325 ;
        RECT -11.045 74.635 -10.715 74.965 ;
        RECT -11.045 73.275 -10.715 73.605 ;
        RECT -11.045 71.915 -10.715 72.245 ;
        RECT -11.045 70.555 -10.715 70.885 ;
        RECT -11.045 69.195 -10.715 69.525 ;
        RECT -11.045 67.835 -10.715 68.165 ;
        RECT -11.045 66.475 -10.715 66.805 ;
        RECT -11.045 65.115 -10.715 65.445 ;
        RECT -11.045 63.755 -10.715 64.085 ;
        RECT -11.045 62.395 -10.715 62.725 ;
        RECT -11.045 61.035 -10.715 61.365 ;
        RECT -11.045 59.675 -10.715 60.005 ;
        RECT -11.045 58.315 -10.715 58.645 ;
        RECT -11.045 56.955 -10.715 57.285 ;
        RECT -11.045 55.595 -10.715 55.925 ;
        RECT -11.045 54.235 -10.715 54.565 ;
        RECT -11.045 52.875 -10.715 53.205 ;
        RECT -11.045 51.515 -10.715 51.845 ;
        RECT -11.045 50.155 -10.715 50.485 ;
        RECT -11.045 48.795 -10.715 49.125 ;
        RECT -11.045 47.435 -10.715 47.765 ;
        RECT -11.045 46.075 -10.715 46.405 ;
        RECT -11.045 44.715 -10.715 45.045 ;
        RECT -11.045 43.355 -10.715 43.685 ;
        RECT -11.045 41.995 -10.715 42.325 ;
        RECT -11.045 40.635 -10.715 40.965 ;
        RECT -11.045 39.275 -10.715 39.605 ;
        RECT -11.045 37.915 -10.715 38.245 ;
        RECT -11.045 36.555 -10.715 36.885 ;
        RECT -11.045 35.195 -10.715 35.525 ;
        RECT -11.045 33.835 -10.715 34.165 ;
        RECT -11.045 32.475 -10.715 32.805 ;
        RECT -11.045 31.115 -10.715 31.445 ;
        RECT -11.045 29.755 -10.715 30.085 ;
        RECT -11.045 28.395 -10.715 28.725 ;
        RECT -11.045 27.035 -10.715 27.365 ;
        RECT -11.045 25.675 -10.715 26.005 ;
        RECT -11.045 24.315 -10.715 24.645 ;
        RECT -11.045 22.955 -10.715 23.285 ;
        RECT -11.045 21.595 -10.715 21.925 ;
        RECT -11.045 20.235 -10.715 20.565 ;
        RECT -11.045 18.875 -10.715 19.205 ;
        RECT -11.045 17.515 -10.715 17.845 ;
        RECT -11.045 16.155 -10.715 16.485 ;
        RECT -11.045 14.795 -10.715 15.125 ;
        RECT -11.045 13.435 -10.715 13.765 ;
        RECT -11.045 12.075 -10.715 12.405 ;
        RECT -11.045 10.715 -10.715 11.045 ;
        RECT -11.045 9.355 -10.715 9.685 ;
        RECT -11.045 7.995 -10.715 8.325 ;
        RECT -11.045 6.635 -10.715 6.965 ;
        RECT -11.045 5.275 -10.715 5.605 ;
        RECT -11.045 3.915 -10.715 4.245 ;
        RECT -11.045 2.555 -10.715 2.885 ;
        RECT -11.045 1.195 -10.715 1.525 ;
        RECT -11.045 -0.165 -10.715 0.165 ;
        RECT -11.045 -1.525 -10.715 -1.195 ;
        RECT -11.045 -2.885 -10.715 -2.555 ;
        RECT -11.045 -4.245 -10.715 -3.915 ;
        RECT -11.045 -5.605 -10.715 -5.275 ;
        RECT -11.045 -6.965 -10.715 -6.635 ;
        RECT -11.045 -9.685 -10.715 -9.355 ;
        RECT -11.04 -10.36 -10.72 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 -106.245 -10.715 -105.915 ;
        RECT -11.045 -108.965 -10.715 -108.635 ;
        RECT -11.045 -110.325 -10.715 -109.995 ;
        RECT -11.045 -113.045 -10.715 -112.715 ;
        RECT -11.045 -114.405 -10.715 -114.075 ;
        RECT -11.045 -115.765 -10.715 -115.435 ;
        RECT -11.045 -117.125 -10.715 -116.795 ;
        RECT -11.045 -118.485 -10.715 -118.155 ;
        RECT -11.045 -119.845 -10.715 -119.515 ;
        RECT -11.045 -121.205 -10.715 -120.875 ;
        RECT -11.045 -125.285 -10.715 -124.955 ;
        RECT -11.045 -126.645 -10.715 -126.315 ;
        RECT -11.045 -128.005 -10.715 -127.675 ;
        RECT -11.045 -129.365 -10.715 -129.035 ;
        RECT -11.045 -130.725 -10.715 -130.395 ;
        RECT -11.045 -132.085 -10.715 -131.755 ;
        RECT -11.045 -133.445 -10.715 -133.115 ;
        RECT -11.045 -134.805 -10.715 -134.475 ;
        RECT -11.045 -136.165 -10.715 -135.835 ;
        RECT -11.045 -138.885 -10.715 -138.555 ;
        RECT -11.045 -140.245 -10.715 -139.915 ;
        RECT -11.045 -141.605 -10.715 -141.275 ;
        RECT -11.045 -142.965 -10.715 -142.635 ;
        RECT -11.045 -144.325 -10.715 -143.995 ;
        RECT -11.045 -145.685 -10.715 -145.355 ;
        RECT -11.045 -149.765 -10.715 -149.435 ;
        RECT -11.045 -153.845 -10.715 -153.515 ;
        RECT -11.045 -155.285 -10.715 -154.955 ;
        RECT -11.045 -156.565 -10.715 -156.235 ;
        RECT -11.045 -157.925 -10.715 -157.595 ;
        RECT -11.045 -160.17 -10.715 -159.04 ;
        RECT -11.04 -160.285 -10.72 -101.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.685 127.225 -9.355 128.355 ;
        RECT -9.685 124.955 -9.355 125.285 ;
        RECT -9.685 123.595 -9.355 123.925 ;
        RECT -9.685 122.235 -9.355 122.565 ;
        RECT -9.685 120.875 -9.355 121.205 ;
        RECT -9.685 119.515 -9.355 119.845 ;
        RECT -9.685 118.155 -9.355 118.485 ;
        RECT -9.685 114.075 -9.355 114.405 ;
        RECT -9.685 104.555 -9.355 104.885 ;
        RECT -9.685 103.195 -9.355 103.525 ;
        RECT -9.685 96.395 -9.355 96.725 ;
        RECT -9.685 93.675 -9.355 94.005 ;
        RECT -9.685 89.595 -9.355 89.925 ;
        RECT -9.685 85.515 -9.355 85.845 ;
        RECT -9.685 82.795 -9.355 83.125 ;
        RECT -9.685 75.995 -9.355 76.325 ;
        RECT -9.685 74.635 -9.355 74.965 ;
        RECT -9.685 65.115 -9.355 65.445 ;
        RECT -9.685 61.035 -9.355 61.365 ;
        RECT -9.685 56.955 -9.355 57.285 ;
        RECT -9.685 54.235 -9.355 54.565 ;
        RECT -9.685 47.435 -9.355 47.765 ;
        RECT -9.685 46.075 -9.355 46.405 ;
        RECT -9.685 43.355 -9.355 43.685 ;
        RECT -9.685 36.555 -9.355 36.885 ;
        RECT -9.685 33.835 -9.355 34.165 ;
        RECT -9.685 32.475 -9.355 32.805 ;
        RECT -9.685 28.395 -9.355 28.725 ;
        RECT -9.685 25.675 -9.355 26.005 ;
        RECT -9.685 18.875 -9.355 19.205 ;
        RECT -9.685 17.515 -9.355 17.845 ;
        RECT -9.685 14.795 -9.355 15.125 ;
        RECT -9.685 7.995 -9.355 8.325 ;
        RECT -9.685 5.275 -9.355 5.605 ;
        RECT -9.685 3.915 -9.355 4.245 ;
        RECT -9.685 2.555 -9.355 2.885 ;
        RECT -9.685 1.195 -9.355 1.525 ;
        RECT -9.685 -0.165 -9.355 0.165 ;
        RECT -9.685 -1.525 -9.355 -1.195 ;
        RECT -9.685 -2.885 -9.355 -2.555 ;
        RECT -9.685 -4.245 -9.355 -3.915 ;
        RECT -9.685 -5.605 -9.355 -5.275 ;
        RECT -9.685 -6.965 -9.355 -6.635 ;
        RECT -9.685 -9.685 -9.355 -9.355 ;
        RECT -9.685 -15.125 -9.355 -14.795 ;
        RECT -9.685 -16.485 -9.355 -16.155 ;
        RECT -9.685 -23.285 -9.355 -22.955 ;
        RECT -9.685 -24.645 -9.355 -24.315 ;
        RECT -9.685 -26.005 -9.355 -25.675 ;
        RECT -9.685 -27.365 -9.355 -27.035 ;
        RECT -9.685 -28.725 -9.355 -28.395 ;
        RECT -9.685 -30.085 -9.355 -29.755 ;
        RECT -9.685 -34.165 -9.355 -33.835 ;
        RECT -9.685 -38.245 -9.355 -37.915 ;
        RECT -9.685 -40.965 -9.355 -40.635 ;
        RECT -9.685 -49.125 -9.355 -48.795 ;
        RECT -9.685 -50.485 -9.355 -50.155 ;
        RECT -9.685 -51.845 -9.355 -51.515 ;
        RECT -9.685 -54.565 -9.355 -54.235 ;
        RECT -9.685 -57.285 -9.355 -56.955 ;
        RECT -9.685 -58.645 -9.355 -58.315 ;
        RECT -9.685 -61.365 -9.355 -61.035 ;
        RECT -9.685 -62.725 -9.355 -62.395 ;
        RECT -9.685 -64.085 -9.355 -63.755 ;
        RECT -9.685 -66.805 -9.355 -66.475 ;
        RECT -9.685 -69.525 -9.355 -69.195 ;
        RECT -9.685 -70.885 -9.355 -70.555 ;
        RECT -9.685 -72.245 -9.355 -71.915 ;
        RECT -9.685 -73.605 -9.355 -73.275 ;
        RECT -9.685 -76.325 -9.355 -75.995 ;
        RECT -9.685 -77.685 -9.355 -77.355 ;
        RECT -9.685 -80.405 -9.355 -80.075 ;
        RECT -9.685 -81.765 -9.355 -81.435 ;
        RECT -9.685 -84.485 -9.355 -84.155 ;
        RECT -9.685 -85.845 -9.355 -85.515 ;
        RECT -9.685 -92.645 -9.355 -92.315 ;
        RECT -9.685 -94.005 -9.355 -93.675 ;
        RECT -9.685 -95.365 -9.355 -95.035 ;
        RECT -9.685 -96.725 -9.355 -96.395 ;
        RECT -9.685 -98.085 -9.355 -97.755 ;
        RECT -9.685 -99.445 -9.355 -99.115 ;
        RECT -9.685 -100.805 -9.355 -100.475 ;
        RECT -9.685 -102.165 -9.355 -101.835 ;
        RECT -9.685 -103.525 -9.355 -103.195 ;
        RECT -9.685 -106.245 -9.355 -105.915 ;
        RECT -9.685 -107.605 -9.355 -107.275 ;
        RECT -9.685 -108.965 -9.355 -108.635 ;
        RECT -9.685 -110.325 -9.355 -109.995 ;
        RECT -9.685 -113.045 -9.355 -112.715 ;
        RECT -9.685 -114.405 -9.355 -114.075 ;
        RECT -9.685 -115.765 -9.355 -115.435 ;
        RECT -9.685 -117.125 -9.355 -116.795 ;
        RECT -9.685 -118.485 -9.355 -118.155 ;
        RECT -9.685 -119.845 -9.355 -119.515 ;
        RECT -9.685 -121.205 -9.355 -120.875 ;
        RECT -9.685 -122.565 -9.355 -122.235 ;
        RECT -9.685 -123.925 -9.355 -123.595 ;
        RECT -9.685 -125.285 -9.355 -124.955 ;
        RECT -9.685 -126.645 -9.355 -126.315 ;
        RECT -9.685 -128.005 -9.355 -127.675 ;
        RECT -9.685 -129.365 -9.355 -129.035 ;
        RECT -9.685 -130.725 -9.355 -130.395 ;
        RECT -9.685 -132.085 -9.355 -131.755 ;
        RECT -9.685 -133.445 -9.355 -133.115 ;
        RECT -9.685 -134.805 -9.355 -134.475 ;
        RECT -9.685 -136.165 -9.355 -135.835 ;
        RECT -9.68 -136.84 -9.36 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 127.225 -7.995 128.355 ;
        RECT -8.325 124.955 -7.995 125.285 ;
        RECT -8.325 123.595 -7.995 123.925 ;
        RECT -8.325 122.235 -7.995 122.565 ;
        RECT -8.325 120.875 -7.995 121.205 ;
        RECT -8.325 119.515 -7.995 119.845 ;
        RECT -8.325 118.155 -7.995 118.485 ;
        RECT -8.325 114.075 -7.995 114.405 ;
        RECT -8.325 104.555 -7.995 104.885 ;
        RECT -8.325 103.195 -7.995 103.525 ;
        RECT -8.325 96.395 -7.995 96.725 ;
        RECT -8.325 93.675 -7.995 94.005 ;
        RECT -8.325 89.595 -7.995 89.925 ;
        RECT -8.325 85.515 -7.995 85.845 ;
        RECT -8.325 82.795 -7.995 83.125 ;
        RECT -8.325 75.995 -7.995 76.325 ;
        RECT -8.325 74.635 -7.995 74.965 ;
        RECT -8.325 65.115 -7.995 65.445 ;
        RECT -8.325 61.035 -7.995 61.365 ;
        RECT -8.325 56.955 -7.995 57.285 ;
        RECT -8.325 54.235 -7.995 54.565 ;
        RECT -8.325 47.435 -7.995 47.765 ;
        RECT -8.325 46.075 -7.995 46.405 ;
        RECT -8.325 43.355 -7.995 43.685 ;
        RECT -8.325 36.555 -7.995 36.885 ;
        RECT -8.325 33.835 -7.995 34.165 ;
        RECT -8.325 32.475 -7.995 32.805 ;
        RECT -8.325 28.395 -7.995 28.725 ;
        RECT -8.325 25.675 -7.995 26.005 ;
        RECT -8.325 18.875 -7.995 19.205 ;
        RECT -8.325 17.515 -7.995 17.845 ;
        RECT -8.325 14.795 -7.995 15.125 ;
        RECT -8.325 7.995 -7.995 8.325 ;
        RECT -8.325 5.275 -7.995 5.605 ;
        RECT -8.325 3.915 -7.995 4.245 ;
        RECT -8.325 2.555 -7.995 2.885 ;
        RECT -8.325 1.195 -7.995 1.525 ;
        RECT -8.325 -0.165 -7.995 0.165 ;
        RECT -8.325 -1.525 -7.995 -1.195 ;
        RECT -8.325 -2.885 -7.995 -2.555 ;
        RECT -8.325 -4.245 -7.995 -3.915 ;
        RECT -8.325 -5.605 -7.995 -5.275 ;
        RECT -8.325 -6.965 -7.995 -6.635 ;
        RECT -8.325 -8.325 -7.995 -7.995 ;
        RECT -8.325 -9.685 -7.995 -9.355 ;
        RECT -8.325 -12.405 -7.995 -12.075 ;
        RECT -8.325 -13.765 -7.995 -13.435 ;
        RECT -8.325 -15.125 -7.995 -14.795 ;
        RECT -8.325 -16.485 -7.995 -16.155 ;
        RECT -8.325 -17.845 -7.995 -17.515 ;
        RECT -8.325 -21.925 -7.995 -21.595 ;
        RECT -8.325 -23.285 -7.995 -22.955 ;
        RECT -8.325 -24.645 -7.995 -24.315 ;
        RECT -8.325 -26.005 -7.995 -25.675 ;
        RECT -8.325 -27.365 -7.995 -27.035 ;
        RECT -8.325 -28.725 -7.995 -28.395 ;
        RECT -8.325 -30.085 -7.995 -29.755 ;
        RECT -8.325 -31.445 -7.995 -31.115 ;
        RECT -8.325 -34.165 -7.995 -33.835 ;
        RECT -8.325 -35.525 -7.995 -35.195 ;
        RECT -8.325 -36.885 -7.995 -36.555 ;
        RECT -8.325 -38.245 -7.995 -37.915 ;
        RECT -8.32 -38.92 -8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 -100.805 -7.995 -100.475 ;
        RECT -8.325 -102.165 -7.995 -101.835 ;
        RECT -8.325 -103.525 -7.995 -103.195 ;
        RECT -8.325 -104.885 -7.995 -104.555 ;
        RECT -8.325 -106.245 -7.995 -105.915 ;
        RECT -8.325 -107.605 -7.995 -107.275 ;
        RECT -8.325 -108.965 -7.995 -108.635 ;
        RECT -8.325 -110.325 -7.995 -109.995 ;
        RECT -8.325 -111.685 -7.995 -111.355 ;
        RECT -8.325 -113.045 -7.995 -112.715 ;
        RECT -8.325 -114.405 -7.995 -114.075 ;
        RECT -8.325 -115.765 -7.995 -115.435 ;
        RECT -8.325 -117.125 -7.995 -116.795 ;
        RECT -8.325 -118.485 -7.995 -118.155 ;
        RECT -8.325 -119.845 -7.995 -119.515 ;
        RECT -8.325 -121.205 -7.995 -120.875 ;
        RECT -8.325 -122.565 -7.995 -122.235 ;
        RECT -8.325 -123.925 -7.995 -123.595 ;
        RECT -8.325 -125.285 -7.995 -124.955 ;
        RECT -8.325 -126.645 -7.995 -126.315 ;
        RECT -8.325 -128.005 -7.995 -127.675 ;
        RECT -8.325 -129.365 -7.995 -129.035 ;
        RECT -8.325 -130.725 -7.995 -130.395 ;
        RECT -8.325 -132.085 -7.995 -131.755 ;
        RECT -8.325 -133.445 -7.995 -133.115 ;
        RECT -8.325 -134.805 -7.995 -134.475 ;
        RECT -8.325 -136.165 -7.995 -135.835 ;
        RECT -8.325 -137.525 -7.995 -137.195 ;
        RECT -8.325 -138.885 -7.995 -138.555 ;
        RECT -8.325 -140.245 -7.995 -139.915 ;
        RECT -8.325 -141.605 -7.995 -141.275 ;
        RECT -8.325 -142.965 -7.995 -142.635 ;
        RECT -8.325 -144.325 -7.995 -143.995 ;
        RECT -8.325 -145.685 -7.995 -145.355 ;
        RECT -8.325 -147.045 -7.995 -146.715 ;
        RECT -8.325 -148.405 -7.995 -148.075 ;
        RECT -8.325 -149.765 -7.995 -149.435 ;
        RECT -8.325 -151.125 -7.995 -150.795 ;
        RECT -8.325 -152.485 -7.995 -152.155 ;
        RECT -8.325 -153.845 -7.995 -153.515 ;
        RECT -8.325 -155.205 -7.995 -154.875 ;
        RECT -8.325 -156.565 -7.995 -156.235 ;
        RECT -8.325 -157.925 -7.995 -157.595 ;
        RECT -8.325 -160.17 -7.995 -159.04 ;
        RECT -8.32 -160.285 -8 -100.475 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.965 127.225 -6.635 128.355 ;
        RECT -6.965 124.955 -6.635 125.285 ;
        RECT -6.965 123.595 -6.635 123.925 ;
        RECT -6.965 122.235 -6.635 122.565 ;
        RECT -6.965 120.875 -6.635 121.205 ;
        RECT -6.965 119.515 -6.635 119.845 ;
        RECT -6.965 118.155 -6.635 118.485 ;
        RECT -6.965 114.075 -6.635 114.405 ;
        RECT -6.965 104.555 -6.635 104.885 ;
        RECT -6.965 103.195 -6.635 103.525 ;
        RECT -6.965 96.395 -6.635 96.725 ;
        RECT -6.965 93.675 -6.635 94.005 ;
        RECT -6.965 89.595 -6.635 89.925 ;
        RECT -6.965 85.515 -6.635 85.845 ;
        RECT -6.965 82.795 -6.635 83.125 ;
        RECT -6.965 75.995 -6.635 76.325 ;
        RECT -6.965 74.635 -6.635 74.965 ;
        RECT -6.965 65.115 -6.635 65.445 ;
        RECT -6.965 61.035 -6.635 61.365 ;
        RECT -6.965 56.955 -6.635 57.285 ;
        RECT -6.965 54.235 -6.635 54.565 ;
        RECT -6.965 47.435 -6.635 47.765 ;
        RECT -6.965 46.075 -6.635 46.405 ;
        RECT -6.965 43.355 -6.635 43.685 ;
        RECT -6.965 36.555 -6.635 36.885 ;
        RECT -6.965 33.835 -6.635 34.165 ;
        RECT -6.965 32.475 -6.635 32.805 ;
        RECT -6.965 28.395 -6.635 28.725 ;
        RECT -6.965 25.675 -6.635 26.005 ;
        RECT -6.965 18.875 -6.635 19.205 ;
        RECT -6.965 17.515 -6.635 17.845 ;
        RECT -6.965 14.795 -6.635 15.125 ;
        RECT -6.965 7.995 -6.635 8.325 ;
        RECT -6.965 5.275 -6.635 5.605 ;
        RECT -6.965 3.915 -6.635 4.245 ;
        RECT -6.965 2.555 -6.635 2.885 ;
        RECT -6.965 1.195 -6.635 1.525 ;
        RECT -6.965 -0.165 -6.635 0.165 ;
        RECT -6.965 -1.525 -6.635 -1.195 ;
        RECT -6.965 -2.885 -6.635 -2.555 ;
        RECT -6.965 -4.245 -6.635 -3.915 ;
        RECT -6.965 -5.605 -6.635 -5.275 ;
        RECT -6.965 -6.965 -6.635 -6.635 ;
        RECT -6.965 -8.325 -6.635 -7.995 ;
        RECT -6.965 -9.685 -6.635 -9.355 ;
        RECT -6.965 -12.405 -6.635 -12.075 ;
        RECT -6.965 -13.765 -6.635 -13.435 ;
        RECT -6.965 -15.125 -6.635 -14.795 ;
        RECT -6.965 -16.485 -6.635 -16.155 ;
        RECT -6.965 -17.845 -6.635 -17.515 ;
        RECT -6.965 -21.925 -6.635 -21.595 ;
        RECT -6.965 -23.285 -6.635 -22.955 ;
        RECT -6.965 -24.645 -6.635 -24.315 ;
        RECT -6.965 -26.005 -6.635 -25.675 ;
        RECT -6.965 -27.365 -6.635 -27.035 ;
        RECT -6.965 -28.725 -6.635 -28.395 ;
        RECT -6.965 -30.085 -6.635 -29.755 ;
        RECT -6.965 -31.445 -6.635 -31.115 ;
        RECT -6.965 -34.165 -6.635 -33.835 ;
        RECT -6.965 -35.525 -6.635 -35.195 ;
        RECT -6.965 -36.885 -6.635 -36.555 ;
        RECT -6.965 -38.245 -6.635 -37.915 ;
        RECT -6.965 -40.965 -6.635 -40.635 ;
        RECT -6.965 -42.325 -6.635 -41.995 ;
        RECT -6.965 -43.685 -6.635 -43.355 ;
        RECT -6.965 -45.045 -6.635 -44.715 ;
        RECT -6.965 -49.125 -6.635 -48.795 ;
        RECT -6.965 -50.485 -6.635 -50.155 ;
        RECT -6.965 -51.845 -6.635 -51.515 ;
        RECT -6.965 -53.205 -6.635 -52.875 ;
        RECT -6.965 -54.565 -6.635 -54.235 ;
        RECT -6.965 -55.925 -6.635 -55.595 ;
        RECT -6.965 -57.285 -6.635 -56.955 ;
        RECT -6.965 -58.645 -6.635 -58.315 ;
        RECT -6.965 -60.005 -6.635 -59.675 ;
        RECT -6.965 -61.365 -6.635 -61.035 ;
        RECT -6.965 -62.725 -6.635 -62.395 ;
        RECT -6.965 -64.085 -6.635 -63.755 ;
        RECT -6.965 -65.445 -6.635 -65.115 ;
        RECT -6.965 -66.805 -6.635 -66.475 ;
        RECT -6.965 -68.165 -6.635 -67.835 ;
        RECT -6.965 -69.525 -6.635 -69.195 ;
        RECT -6.965 -70.885 -6.635 -70.555 ;
        RECT -6.965 -72.245 -6.635 -71.915 ;
        RECT -6.965 -73.605 -6.635 -73.275 ;
        RECT -6.965 -74.965 -6.635 -74.635 ;
        RECT -6.965 -76.325 -6.635 -75.995 ;
        RECT -6.965 -77.685 -6.635 -77.355 ;
        RECT -6.965 -79.045 -6.635 -78.715 ;
        RECT -6.965 -80.405 -6.635 -80.075 ;
        RECT -6.965 -81.765 -6.635 -81.435 ;
        RECT -6.965 -83.125 -6.635 -82.795 ;
        RECT -6.965 -84.485 -6.635 -84.155 ;
        RECT -6.965 -85.845 -6.635 -85.515 ;
        RECT -6.965 -87.205 -6.635 -86.875 ;
        RECT -6.965 -88.565 -6.635 -88.235 ;
        RECT -6.965 -89.925 -6.635 -89.595 ;
        RECT -6.965 -91.285 -6.635 -90.955 ;
        RECT -6.965 -92.645 -6.635 -92.315 ;
        RECT -6.965 -94.005 -6.635 -93.675 ;
        RECT -6.965 -95.365 -6.635 -95.035 ;
        RECT -6.965 -96.725 -6.635 -96.395 ;
        RECT -6.965 -98.085 -6.635 -97.755 ;
        RECT -6.965 -99.445 -6.635 -99.115 ;
        RECT -6.965 -100.805 -6.635 -100.475 ;
        RECT -6.965 -102.165 -6.635 -101.835 ;
        RECT -6.965 -103.525 -6.635 -103.195 ;
        RECT -6.965 -104.885 -6.635 -104.555 ;
        RECT -6.965 -106.245 -6.635 -105.915 ;
        RECT -6.965 -107.605 -6.635 -107.275 ;
        RECT -6.965 -108.965 -6.635 -108.635 ;
        RECT -6.965 -110.325 -6.635 -109.995 ;
        RECT -6.965 -111.685 -6.635 -111.355 ;
        RECT -6.965 -113.045 -6.635 -112.715 ;
        RECT -6.965 -114.405 -6.635 -114.075 ;
        RECT -6.965 -115.765 -6.635 -115.435 ;
        RECT -6.965 -117.125 -6.635 -116.795 ;
        RECT -6.965 -118.485 -6.635 -118.155 ;
        RECT -6.965 -119.845 -6.635 -119.515 ;
        RECT -6.965 -121.205 -6.635 -120.875 ;
        RECT -6.965 -122.565 -6.635 -122.235 ;
        RECT -6.965 -123.925 -6.635 -123.595 ;
        RECT -6.965 -125.285 -6.635 -124.955 ;
        RECT -6.965 -126.645 -6.635 -126.315 ;
        RECT -6.965 -128.005 -6.635 -127.675 ;
        RECT -6.965 -129.365 -6.635 -129.035 ;
        RECT -6.965 -130.725 -6.635 -130.395 ;
        RECT -6.965 -132.085 -6.635 -131.755 ;
        RECT -6.965 -133.445 -6.635 -133.115 ;
        RECT -6.965 -134.805 -6.635 -134.475 ;
        RECT -6.965 -136.165 -6.635 -135.835 ;
        RECT -6.965 -137.525 -6.635 -137.195 ;
        RECT -6.965 -138.885 -6.635 -138.555 ;
        RECT -6.965 -140.245 -6.635 -139.915 ;
        RECT -6.965 -141.605 -6.635 -141.275 ;
        RECT -6.965 -142.965 -6.635 -142.635 ;
        RECT -6.965 -144.325 -6.635 -143.995 ;
        RECT -6.965 -145.685 -6.635 -145.355 ;
        RECT -6.965 -147.045 -6.635 -146.715 ;
        RECT -6.965 -148.405 -6.635 -148.075 ;
        RECT -6.965 -149.765 -6.635 -149.435 ;
        RECT -6.965 -151.125 -6.635 -150.795 ;
        RECT -6.965 -152.485 -6.635 -152.155 ;
        RECT -6.965 -153.845 -6.635 -153.515 ;
        RECT -6.965 -155.205 -6.635 -154.875 ;
        RECT -6.965 -156.565 -6.635 -156.235 ;
        RECT -6.965 -157.925 -6.635 -157.595 ;
        RECT -6.965 -160.17 -6.635 -159.04 ;
        RECT -6.96 -160.285 -6.64 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.605 127.225 -5.275 128.355 ;
        RECT -5.605 124.955 -5.275 125.285 ;
        RECT -5.605 123.595 -5.275 123.925 ;
        RECT -5.605 122.215 -5.275 122.545 ;
        RECT -5.605 120.165 -5.275 120.495 ;
        RECT -5.605 118.235 -5.275 118.565 ;
        RECT -5.605 116.395 -5.275 116.725 ;
        RECT -5.605 114.905 -5.275 115.235 ;
        RECT -5.605 113.235 -5.275 113.565 ;
        RECT -5.605 111.745 -5.275 112.075 ;
        RECT -5.605 110.075 -5.275 110.405 ;
        RECT -5.605 108.585 -5.275 108.915 ;
        RECT -5.605 106.915 -5.275 107.245 ;
        RECT -5.605 105.425 -5.275 105.755 ;
        RECT -5.605 104.015 -5.275 104.345 ;
        RECT -5.605 102.175 -5.275 102.505 ;
        RECT -5.605 100.685 -5.275 101.015 ;
        RECT -5.605 99.015 -5.275 99.345 ;
        RECT -5.605 97.525 -5.275 97.855 ;
        RECT -5.605 95.855 -5.275 96.185 ;
        RECT -5.605 94.365 -5.275 94.695 ;
        RECT -5.605 92.695 -5.275 93.025 ;
        RECT -5.605 91.205 -5.275 91.535 ;
        RECT -5.605 89.795 -5.275 90.125 ;
        RECT -5.605 87.955 -5.275 88.285 ;
        RECT -5.605 86.465 -5.275 86.795 ;
        RECT -5.605 84.795 -5.275 85.125 ;
        RECT -5.605 83.305 -5.275 83.635 ;
        RECT -5.605 81.635 -5.275 81.965 ;
        RECT -5.605 80.145 -5.275 80.475 ;
        RECT -5.605 78.475 -5.275 78.805 ;
        RECT -5.605 76.985 -5.275 77.315 ;
        RECT -5.605 75.575 -5.275 75.905 ;
        RECT -5.605 73.735 -5.275 74.065 ;
        RECT -5.605 72.245 -5.275 72.575 ;
        RECT -5.605 70.575 -5.275 70.905 ;
        RECT -5.605 69.085 -5.275 69.415 ;
        RECT -5.605 67.415 -5.275 67.745 ;
        RECT -5.605 65.925 -5.275 66.255 ;
        RECT -5.605 64.255 -5.275 64.585 ;
        RECT -5.605 62.765 -5.275 63.095 ;
        RECT -5.605 61.355 -5.275 61.685 ;
        RECT -5.605 59.515 -5.275 59.845 ;
        RECT -5.605 58.025 -5.275 58.355 ;
        RECT -5.605 56.355 -5.275 56.685 ;
        RECT -5.605 54.865 -5.275 55.195 ;
        RECT -5.605 53.195 -5.275 53.525 ;
        RECT -5.605 51.705 -5.275 52.035 ;
        RECT -5.605 50.035 -5.275 50.365 ;
        RECT -5.605 48.545 -5.275 48.875 ;
        RECT -5.605 47.135 -5.275 47.465 ;
        RECT -5.605 45.295 -5.275 45.625 ;
        RECT -5.605 43.805 -5.275 44.135 ;
        RECT -5.605 42.135 -5.275 42.465 ;
        RECT -5.605 40.645 -5.275 40.975 ;
        RECT -5.605 38.975 -5.275 39.305 ;
        RECT -5.605 37.485 -5.275 37.815 ;
        RECT -5.605 35.815 -5.275 36.145 ;
        RECT -5.605 34.325 -5.275 34.655 ;
        RECT -5.605 32.915 -5.275 33.245 ;
        RECT -5.605 31.075 -5.275 31.405 ;
        RECT -5.605 29.585 -5.275 29.915 ;
        RECT -5.605 27.915 -5.275 28.245 ;
        RECT -5.605 26.425 -5.275 26.755 ;
        RECT -5.605 24.755 -5.275 25.085 ;
        RECT -5.605 23.265 -5.275 23.595 ;
        RECT -5.605 21.595 -5.275 21.925 ;
        RECT -5.605 20.105 -5.275 20.435 ;
        RECT -5.605 18.695 -5.275 19.025 ;
        RECT -5.605 16.855 -5.275 17.185 ;
        RECT -5.605 15.365 -5.275 15.695 ;
        RECT -5.605 13.695 -5.275 14.025 ;
        RECT -5.605 12.205 -5.275 12.535 ;
        RECT -5.605 10.535 -5.275 10.865 ;
        RECT -5.605 9.045 -5.275 9.375 ;
        RECT -5.605 7.375 -5.275 7.705 ;
        RECT -5.605 5.885 -5.275 6.215 ;
        RECT -5.605 4.475 -5.275 4.805 ;
        RECT -5.605 2.115 -5.275 2.445 ;
        RECT -5.605 0.06 -5.275 0.39 ;
        RECT -5.605 -1.525 -5.275 -1.195 ;
        RECT -5.605 -2.885 -5.275 -2.555 ;
        RECT -5.605 -4.245 -5.275 -3.915 ;
        RECT -5.605 -5.605 -5.275 -5.275 ;
        RECT -5.605 -6.965 -5.275 -6.635 ;
        RECT -5.605 -8.325 -5.275 -7.995 ;
        RECT -5.605 -9.685 -5.275 -9.355 ;
        RECT -5.605 -12.405 -5.275 -12.075 ;
        RECT -5.605 -13.765 -5.275 -13.435 ;
        RECT -5.605 -15.125 -5.275 -14.795 ;
        RECT -5.605 -16.485 -5.275 -16.155 ;
        RECT -5.605 -17.845 -5.275 -17.515 ;
        RECT -5.605 -21.925 -5.275 -21.595 ;
        RECT -5.605 -23.285 -5.275 -22.955 ;
        RECT -5.605 -24.645 -5.275 -24.315 ;
        RECT -5.605 -26.005 -5.275 -25.675 ;
        RECT -5.605 -27.365 -5.275 -27.035 ;
        RECT -5.605 -28.725 -5.275 -28.395 ;
        RECT -5.605 -30.085 -5.275 -29.755 ;
        RECT -5.605 -31.445 -5.275 -31.115 ;
        RECT -5.605 -34.165 -5.275 -33.835 ;
        RECT -5.605 -35.525 -5.275 -35.195 ;
        RECT -5.605 -36.885 -5.275 -36.555 ;
        RECT -5.605 -38.245 -5.275 -37.915 ;
        RECT -5.605 -40.965 -5.275 -40.635 ;
        RECT -5.605 -42.325 -5.275 -41.995 ;
        RECT -5.605 -43.685 -5.275 -43.355 ;
        RECT -5.605 -45.045 -5.275 -44.715 ;
        RECT -5.605 -49.125 -5.275 -48.795 ;
        RECT -5.605 -50.485 -5.275 -50.155 ;
        RECT -5.605 -51.845 -5.275 -51.515 ;
        RECT -5.605 -53.205 -5.275 -52.875 ;
        RECT -5.605 -54.565 -5.275 -54.235 ;
        RECT -5.605 -55.925 -5.275 -55.595 ;
        RECT -5.605 -57.285 -5.275 -56.955 ;
        RECT -5.605 -58.645 -5.275 -58.315 ;
        RECT -5.605 -60.005 -5.275 -59.675 ;
        RECT -5.605 -61.365 -5.275 -61.035 ;
        RECT -5.605 -62.725 -5.275 -62.395 ;
        RECT -5.605 -64.085 -5.275 -63.755 ;
        RECT -5.605 -65.445 -5.275 -65.115 ;
        RECT -5.605 -66.805 -5.275 -66.475 ;
        RECT -5.605 -68.165 -5.275 -67.835 ;
        RECT -5.605 -69.525 -5.275 -69.195 ;
        RECT -5.605 -70.885 -5.275 -70.555 ;
        RECT -5.605 -72.245 -5.275 -71.915 ;
        RECT -5.605 -73.605 -5.275 -73.275 ;
        RECT -5.605 -74.965 -5.275 -74.635 ;
        RECT -5.605 -76.325 -5.275 -75.995 ;
        RECT -5.605 -77.685 -5.275 -77.355 ;
        RECT -5.605 -79.045 -5.275 -78.715 ;
        RECT -5.605 -80.405 -5.275 -80.075 ;
        RECT -5.605 -81.765 -5.275 -81.435 ;
        RECT -5.605 -83.125 -5.275 -82.795 ;
        RECT -5.605 -84.485 -5.275 -84.155 ;
        RECT -5.605 -85.845 -5.275 -85.515 ;
        RECT -5.605 -87.205 -5.275 -86.875 ;
        RECT -5.605 -88.565 -5.275 -88.235 ;
        RECT -5.605 -89.925 -5.275 -89.595 ;
        RECT -5.605 -91.285 -5.275 -90.955 ;
        RECT -5.605 -92.645 -5.275 -92.315 ;
        RECT -5.605 -94.005 -5.275 -93.675 ;
        RECT -5.605 -95.365 -5.275 -95.035 ;
        RECT -5.605 -96.725 -5.275 -96.395 ;
        RECT -5.605 -98.085 -5.275 -97.755 ;
        RECT -5.605 -99.445 -5.275 -99.115 ;
        RECT -5.605 -100.805 -5.275 -100.475 ;
        RECT -5.605 -102.165 -5.275 -101.835 ;
        RECT -5.605 -103.525 -5.275 -103.195 ;
        RECT -5.605 -104.885 -5.275 -104.555 ;
        RECT -5.605 -106.245 -5.275 -105.915 ;
        RECT -5.605 -107.605 -5.275 -107.275 ;
        RECT -5.605 -108.965 -5.275 -108.635 ;
        RECT -5.605 -110.325 -5.275 -109.995 ;
        RECT -5.605 -111.685 -5.275 -111.355 ;
        RECT -5.605 -113.045 -5.275 -112.715 ;
        RECT -5.605 -114.405 -5.275 -114.075 ;
        RECT -5.605 -115.765 -5.275 -115.435 ;
        RECT -5.605 -117.125 -5.275 -116.795 ;
        RECT -5.605 -118.485 -5.275 -118.155 ;
        RECT -5.605 -119.845 -5.275 -119.515 ;
        RECT -5.605 -121.205 -5.275 -120.875 ;
        RECT -5.605 -122.565 -5.275 -122.235 ;
        RECT -5.605 -123.925 -5.275 -123.595 ;
        RECT -5.605 -125.285 -5.275 -124.955 ;
        RECT -5.605 -126.645 -5.275 -126.315 ;
        RECT -5.605 -128.005 -5.275 -127.675 ;
        RECT -5.605 -129.365 -5.275 -129.035 ;
        RECT -5.605 -130.725 -5.275 -130.395 ;
        RECT -5.605 -132.085 -5.275 -131.755 ;
        RECT -5.605 -133.445 -5.275 -133.115 ;
        RECT -5.605 -134.805 -5.275 -134.475 ;
        RECT -5.605 -136.165 -5.275 -135.835 ;
        RECT -5.605 -137.525 -5.275 -137.195 ;
        RECT -5.605 -138.885 -5.275 -138.555 ;
        RECT -5.605 -140.245 -5.275 -139.915 ;
        RECT -5.605 -141.605 -5.275 -141.275 ;
        RECT -5.605 -142.965 -5.275 -142.635 ;
        RECT -5.605 -144.325 -5.275 -143.995 ;
        RECT -5.605 -145.685 -5.275 -145.355 ;
        RECT -5.605 -147.045 -5.275 -146.715 ;
        RECT -5.605 -148.405 -5.275 -148.075 ;
        RECT -5.605 -149.765 -5.275 -149.435 ;
        RECT -5.605 -151.125 -5.275 -150.795 ;
        RECT -5.605 -152.485 -5.275 -152.155 ;
        RECT -5.605 -153.845 -5.275 -153.515 ;
        RECT -5.605 -155.205 -5.275 -154.875 ;
        RECT -5.605 -156.565 -5.275 -156.235 ;
        RECT -5.605 -157.925 -5.275 -157.595 ;
        RECT -5.605 -160.17 -5.275 -159.04 ;
        RECT -5.6 -160.285 -5.28 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.245 127.225 -3.915 128.355 ;
        RECT -4.245 124.955 -3.915 125.285 ;
        RECT -4.245 123.595 -3.915 123.925 ;
        RECT -4.245 122.215 -3.915 122.545 ;
        RECT -4.245 120.165 -3.915 120.495 ;
        RECT -4.245 118.235 -3.915 118.565 ;
        RECT -4.245 116.395 -3.915 116.725 ;
        RECT -4.245 114.905 -3.915 115.235 ;
        RECT -4.245 113.235 -3.915 113.565 ;
        RECT -4.245 111.745 -3.915 112.075 ;
        RECT -4.245 110.075 -3.915 110.405 ;
        RECT -4.245 108.585 -3.915 108.915 ;
        RECT -4.245 106.915 -3.915 107.245 ;
        RECT -4.245 105.425 -3.915 105.755 ;
        RECT -4.245 104.015 -3.915 104.345 ;
        RECT -4.245 102.175 -3.915 102.505 ;
        RECT -4.245 100.685 -3.915 101.015 ;
        RECT -4.245 99.015 -3.915 99.345 ;
        RECT -4.245 97.525 -3.915 97.855 ;
        RECT -4.245 95.855 -3.915 96.185 ;
        RECT -4.245 94.365 -3.915 94.695 ;
        RECT -4.245 92.695 -3.915 93.025 ;
        RECT -4.245 91.205 -3.915 91.535 ;
        RECT -4.245 89.795 -3.915 90.125 ;
        RECT -4.245 87.955 -3.915 88.285 ;
        RECT -4.245 86.465 -3.915 86.795 ;
        RECT -4.245 84.795 -3.915 85.125 ;
        RECT -4.245 83.305 -3.915 83.635 ;
        RECT -4.245 81.635 -3.915 81.965 ;
        RECT -4.245 80.145 -3.915 80.475 ;
        RECT -4.245 78.475 -3.915 78.805 ;
        RECT -4.245 76.985 -3.915 77.315 ;
        RECT -4.245 75.575 -3.915 75.905 ;
        RECT -4.245 73.735 -3.915 74.065 ;
        RECT -4.245 72.245 -3.915 72.575 ;
        RECT -4.245 70.575 -3.915 70.905 ;
        RECT -4.245 69.085 -3.915 69.415 ;
        RECT -4.245 67.415 -3.915 67.745 ;
        RECT -4.245 65.925 -3.915 66.255 ;
        RECT -4.245 64.255 -3.915 64.585 ;
        RECT -4.245 62.765 -3.915 63.095 ;
        RECT -4.245 61.355 -3.915 61.685 ;
        RECT -4.245 59.515 -3.915 59.845 ;
        RECT -4.245 58.025 -3.915 58.355 ;
        RECT -4.245 56.355 -3.915 56.685 ;
        RECT -4.245 54.865 -3.915 55.195 ;
        RECT -4.245 53.195 -3.915 53.525 ;
        RECT -4.245 51.705 -3.915 52.035 ;
        RECT -4.245 50.035 -3.915 50.365 ;
        RECT -4.245 48.545 -3.915 48.875 ;
        RECT -4.245 47.135 -3.915 47.465 ;
        RECT -4.245 45.295 -3.915 45.625 ;
        RECT -4.245 43.805 -3.915 44.135 ;
        RECT -4.245 42.135 -3.915 42.465 ;
        RECT -4.245 40.645 -3.915 40.975 ;
        RECT -4.245 38.975 -3.915 39.305 ;
        RECT -4.245 37.485 -3.915 37.815 ;
        RECT -4.245 35.815 -3.915 36.145 ;
        RECT -4.245 34.325 -3.915 34.655 ;
        RECT -4.245 32.915 -3.915 33.245 ;
        RECT -4.245 31.075 -3.915 31.405 ;
        RECT -4.245 29.585 -3.915 29.915 ;
        RECT -4.245 27.915 -3.915 28.245 ;
        RECT -4.245 26.425 -3.915 26.755 ;
        RECT -4.245 24.755 -3.915 25.085 ;
        RECT -4.245 23.265 -3.915 23.595 ;
        RECT -4.245 21.595 -3.915 21.925 ;
        RECT -4.245 20.105 -3.915 20.435 ;
        RECT -4.245 18.695 -3.915 19.025 ;
        RECT -4.245 16.855 -3.915 17.185 ;
        RECT -4.245 15.365 -3.915 15.695 ;
        RECT -4.245 13.695 -3.915 14.025 ;
        RECT -4.245 12.205 -3.915 12.535 ;
        RECT -4.245 10.535 -3.915 10.865 ;
        RECT -4.245 9.045 -3.915 9.375 ;
        RECT -4.245 7.375 -3.915 7.705 ;
        RECT -4.245 5.885 -3.915 6.215 ;
        RECT -4.245 4.475 -3.915 4.805 ;
        RECT -4.245 2.115 -3.915 2.445 ;
        RECT -4.245 0.06 -3.915 0.39 ;
        RECT -4.245 -1.525 -3.915 -1.195 ;
        RECT -4.245 -2.885 -3.915 -2.555 ;
        RECT -4.245 -4.245 -3.915 -3.915 ;
        RECT -4.245 -5.605 -3.915 -5.275 ;
        RECT -4.245 -6.965 -3.915 -6.635 ;
        RECT -4.245 -8.325 -3.915 -7.995 ;
        RECT -4.245 -9.685 -3.915 -9.355 ;
        RECT -4.245 -12.405 -3.915 -12.075 ;
        RECT -4.245 -13.765 -3.915 -13.435 ;
        RECT -4.245 -15.125 -3.915 -14.795 ;
        RECT -4.245 -16.485 -3.915 -16.155 ;
        RECT -4.245 -17.845 -3.915 -17.515 ;
        RECT -4.245 -21.925 -3.915 -21.595 ;
        RECT -4.245 -23.285 -3.915 -22.955 ;
        RECT -4.245 -24.645 -3.915 -24.315 ;
        RECT -4.245 -26.005 -3.915 -25.675 ;
        RECT -4.245 -27.365 -3.915 -27.035 ;
        RECT -4.245 -28.725 -3.915 -28.395 ;
        RECT -4.245 -30.085 -3.915 -29.755 ;
        RECT -4.245 -31.445 -3.915 -31.115 ;
        RECT -4.245 -34.165 -3.915 -33.835 ;
        RECT -4.245 -35.525 -3.915 -35.195 ;
        RECT -4.245 -36.885 -3.915 -36.555 ;
        RECT -4.245 -38.245 -3.915 -37.915 ;
        RECT -4.245 -40.965 -3.915 -40.635 ;
        RECT -4.245 -42.325 -3.915 -41.995 ;
        RECT -4.245 -43.685 -3.915 -43.355 ;
        RECT -4.245 -45.045 -3.915 -44.715 ;
        RECT -4.245 -49.125 -3.915 -48.795 ;
        RECT -4.245 -50.485 -3.915 -50.155 ;
        RECT -4.245 -51.845 -3.915 -51.515 ;
        RECT -4.245 -53.205 -3.915 -52.875 ;
        RECT -4.245 -54.565 -3.915 -54.235 ;
        RECT -4.245 -55.925 -3.915 -55.595 ;
        RECT -4.245 -57.285 -3.915 -56.955 ;
        RECT -4.245 -58.645 -3.915 -58.315 ;
        RECT -4.245 -60.005 -3.915 -59.675 ;
        RECT -4.245 -61.365 -3.915 -61.035 ;
        RECT -4.245 -62.725 -3.915 -62.395 ;
        RECT -4.245 -64.085 -3.915 -63.755 ;
        RECT -4.245 -65.445 -3.915 -65.115 ;
        RECT -4.245 -66.805 -3.915 -66.475 ;
        RECT -4.245 -68.165 -3.915 -67.835 ;
        RECT -4.245 -69.525 -3.915 -69.195 ;
        RECT -4.245 -70.885 -3.915 -70.555 ;
        RECT -4.245 -72.245 -3.915 -71.915 ;
        RECT -4.245 -73.605 -3.915 -73.275 ;
        RECT -4.245 -74.965 -3.915 -74.635 ;
        RECT -4.245 -76.325 -3.915 -75.995 ;
        RECT -4.245 -77.685 -3.915 -77.355 ;
        RECT -4.245 -79.045 -3.915 -78.715 ;
        RECT -4.245 -80.405 -3.915 -80.075 ;
        RECT -4.245 -81.765 -3.915 -81.435 ;
        RECT -4.245 -83.125 -3.915 -82.795 ;
        RECT -4.245 -84.485 -3.915 -84.155 ;
        RECT -4.245 -85.845 -3.915 -85.515 ;
        RECT -4.245 -87.205 -3.915 -86.875 ;
        RECT -4.245 -88.565 -3.915 -88.235 ;
        RECT -4.245 -89.925 -3.915 -89.595 ;
        RECT -4.245 -91.285 -3.915 -90.955 ;
        RECT -4.245 -92.645 -3.915 -92.315 ;
        RECT -4.245 -94.005 -3.915 -93.675 ;
        RECT -4.245 -95.365 -3.915 -95.035 ;
        RECT -4.245 -96.725 -3.915 -96.395 ;
        RECT -4.245 -98.085 -3.915 -97.755 ;
        RECT -4.245 -99.445 -3.915 -99.115 ;
        RECT -4.245 -100.805 -3.915 -100.475 ;
        RECT -4.245 -102.165 -3.915 -101.835 ;
        RECT -4.245 -103.525 -3.915 -103.195 ;
        RECT -4.245 -104.885 -3.915 -104.555 ;
        RECT -4.245 -106.245 -3.915 -105.915 ;
        RECT -4.245 -107.605 -3.915 -107.275 ;
        RECT -4.245 -108.965 -3.915 -108.635 ;
        RECT -4.245 -110.325 -3.915 -109.995 ;
        RECT -4.245 -111.685 -3.915 -111.355 ;
        RECT -4.245 -113.045 -3.915 -112.715 ;
        RECT -4.245 -114.405 -3.915 -114.075 ;
        RECT -4.245 -115.765 -3.915 -115.435 ;
        RECT -4.245 -117.125 -3.915 -116.795 ;
        RECT -4.245 -118.485 -3.915 -118.155 ;
        RECT -4.245 -119.845 -3.915 -119.515 ;
        RECT -4.245 -121.205 -3.915 -120.875 ;
        RECT -4.245 -122.565 -3.915 -122.235 ;
        RECT -4.245 -123.925 -3.915 -123.595 ;
        RECT -4.245 -125.285 -3.915 -124.955 ;
        RECT -4.245 -126.645 -3.915 -126.315 ;
        RECT -4.245 -128.005 -3.915 -127.675 ;
        RECT -4.245 -129.365 -3.915 -129.035 ;
        RECT -4.245 -130.725 -3.915 -130.395 ;
        RECT -4.245 -132.085 -3.915 -131.755 ;
        RECT -4.245 -133.445 -3.915 -133.115 ;
        RECT -4.245 -134.805 -3.915 -134.475 ;
        RECT -4.245 -136.165 -3.915 -135.835 ;
        RECT -4.245 -137.525 -3.915 -137.195 ;
        RECT -4.245 -138.885 -3.915 -138.555 ;
        RECT -4.245 -140.245 -3.915 -139.915 ;
        RECT -4.245 -141.605 -3.915 -141.275 ;
        RECT -4.245 -142.965 -3.915 -142.635 ;
        RECT -4.245 -144.325 -3.915 -143.995 ;
        RECT -4.245 -145.685 -3.915 -145.355 ;
        RECT -4.245 -147.045 -3.915 -146.715 ;
        RECT -4.245 -148.405 -3.915 -148.075 ;
        RECT -4.245 -149.765 -3.915 -149.435 ;
        RECT -4.245 -151.125 -3.915 -150.795 ;
        RECT -4.245 -152.485 -3.915 -152.155 ;
        RECT -4.245 -153.845 -3.915 -153.515 ;
        RECT -4.245 -155.205 -3.915 -154.875 ;
        RECT -4.245 -156.565 -3.915 -156.235 ;
        RECT -4.245 -157.925 -3.915 -157.595 ;
        RECT -4.245 -160.17 -3.915 -159.04 ;
        RECT -4.24 -160.285 -3.92 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.885 -142.965 -2.555 -142.635 ;
        RECT -2.885 -144.325 -2.555 -143.995 ;
        RECT -2.885 -145.685 -2.555 -145.355 ;
        RECT -2.885 -147.045 -2.555 -146.715 ;
        RECT -2.885 -148.405 -2.555 -148.075 ;
        RECT -2.885 -149.765 -2.555 -149.435 ;
        RECT -2.885 -151.125 -2.555 -150.795 ;
        RECT -2.885 -152.485 -2.555 -152.155 ;
        RECT -2.885 -153.845 -2.555 -153.515 ;
        RECT -2.885 -155.205 -2.555 -154.875 ;
        RECT -2.885 -156.565 -2.555 -156.235 ;
        RECT -2.885 -157.925 -2.555 -157.595 ;
        RECT -2.885 -160.17 -2.555 -159.04 ;
        RECT -2.88 -160.285 -2.56 128.47 ;
        RECT -2.885 127.225 -2.555 128.355 ;
        RECT -2.885 124.955 -2.555 125.285 ;
        RECT -2.885 123.595 -2.555 123.925 ;
        RECT -2.885 122.215 -2.555 122.545 ;
        RECT -2.885 120.165 -2.555 120.495 ;
        RECT -2.885 118.235 -2.555 118.565 ;
        RECT -2.885 116.395 -2.555 116.725 ;
        RECT -2.885 114.905 -2.555 115.235 ;
        RECT -2.885 113.235 -2.555 113.565 ;
        RECT -2.885 111.745 -2.555 112.075 ;
        RECT -2.885 110.075 -2.555 110.405 ;
        RECT -2.885 108.585 -2.555 108.915 ;
        RECT -2.885 106.915 -2.555 107.245 ;
        RECT -2.885 105.425 -2.555 105.755 ;
        RECT -2.885 104.015 -2.555 104.345 ;
        RECT -2.885 102.175 -2.555 102.505 ;
        RECT -2.885 100.685 -2.555 101.015 ;
        RECT -2.885 99.015 -2.555 99.345 ;
        RECT -2.885 97.525 -2.555 97.855 ;
        RECT -2.885 95.855 -2.555 96.185 ;
        RECT -2.885 94.365 -2.555 94.695 ;
        RECT -2.885 92.695 -2.555 93.025 ;
        RECT -2.885 91.205 -2.555 91.535 ;
        RECT -2.885 89.795 -2.555 90.125 ;
        RECT -2.885 87.955 -2.555 88.285 ;
        RECT -2.885 86.465 -2.555 86.795 ;
        RECT -2.885 84.795 -2.555 85.125 ;
        RECT -2.885 83.305 -2.555 83.635 ;
        RECT -2.885 81.635 -2.555 81.965 ;
        RECT -2.885 80.145 -2.555 80.475 ;
        RECT -2.885 78.475 -2.555 78.805 ;
        RECT -2.885 76.985 -2.555 77.315 ;
        RECT -2.885 75.575 -2.555 75.905 ;
        RECT -2.885 73.735 -2.555 74.065 ;
        RECT -2.885 72.245 -2.555 72.575 ;
        RECT -2.885 70.575 -2.555 70.905 ;
        RECT -2.885 69.085 -2.555 69.415 ;
        RECT -2.885 67.415 -2.555 67.745 ;
        RECT -2.885 65.925 -2.555 66.255 ;
        RECT -2.885 64.255 -2.555 64.585 ;
        RECT -2.885 62.765 -2.555 63.095 ;
        RECT -2.885 61.355 -2.555 61.685 ;
        RECT -2.885 59.515 -2.555 59.845 ;
        RECT -2.885 58.025 -2.555 58.355 ;
        RECT -2.885 56.355 -2.555 56.685 ;
        RECT -2.885 54.865 -2.555 55.195 ;
        RECT -2.885 53.195 -2.555 53.525 ;
        RECT -2.885 51.705 -2.555 52.035 ;
        RECT -2.885 50.035 -2.555 50.365 ;
        RECT -2.885 48.545 -2.555 48.875 ;
        RECT -2.885 47.135 -2.555 47.465 ;
        RECT -2.885 45.295 -2.555 45.625 ;
        RECT -2.885 43.805 -2.555 44.135 ;
        RECT -2.885 42.135 -2.555 42.465 ;
        RECT -2.885 40.645 -2.555 40.975 ;
        RECT -2.885 38.975 -2.555 39.305 ;
        RECT -2.885 37.485 -2.555 37.815 ;
        RECT -2.885 35.815 -2.555 36.145 ;
        RECT -2.885 34.325 -2.555 34.655 ;
        RECT -2.885 32.915 -2.555 33.245 ;
        RECT -2.885 31.075 -2.555 31.405 ;
        RECT -2.885 29.585 -2.555 29.915 ;
        RECT -2.885 27.915 -2.555 28.245 ;
        RECT -2.885 26.425 -2.555 26.755 ;
        RECT -2.885 24.755 -2.555 25.085 ;
        RECT -2.885 23.265 -2.555 23.595 ;
        RECT -2.885 21.595 -2.555 21.925 ;
        RECT -2.885 20.105 -2.555 20.435 ;
        RECT -2.885 18.695 -2.555 19.025 ;
        RECT -2.885 16.855 -2.555 17.185 ;
        RECT -2.885 15.365 -2.555 15.695 ;
        RECT -2.885 13.695 -2.555 14.025 ;
        RECT -2.885 12.205 -2.555 12.535 ;
        RECT -2.885 10.535 -2.555 10.865 ;
        RECT -2.885 9.045 -2.555 9.375 ;
        RECT -2.885 7.375 -2.555 7.705 ;
        RECT -2.885 5.885 -2.555 6.215 ;
        RECT -2.885 4.475 -2.555 4.805 ;
        RECT -2.885 2.115 -2.555 2.445 ;
        RECT -2.885 0.06 -2.555 0.39 ;
        RECT -2.885 -1.525 -2.555 -1.195 ;
        RECT -2.885 -2.885 -2.555 -2.555 ;
        RECT -2.885 -4.245 -2.555 -3.915 ;
        RECT -2.885 -5.605 -2.555 -5.275 ;
        RECT -2.885 -6.965 -2.555 -6.635 ;
        RECT -2.885 -8.325 -2.555 -7.995 ;
        RECT -2.885 -9.685 -2.555 -9.355 ;
        RECT -2.885 -12.405 -2.555 -12.075 ;
        RECT -2.885 -13.765 -2.555 -13.435 ;
        RECT -2.885 -15.125 -2.555 -14.795 ;
        RECT -2.885 -16.485 -2.555 -16.155 ;
        RECT -2.885 -17.845 -2.555 -17.515 ;
        RECT -2.885 -21.925 -2.555 -21.595 ;
        RECT -2.885 -23.285 -2.555 -22.955 ;
        RECT -2.885 -24.645 -2.555 -24.315 ;
        RECT -2.885 -26.005 -2.555 -25.675 ;
        RECT -2.885 -27.365 -2.555 -27.035 ;
        RECT -2.885 -28.725 -2.555 -28.395 ;
        RECT -2.885 -30.085 -2.555 -29.755 ;
        RECT -2.885 -31.445 -2.555 -31.115 ;
        RECT -2.885 -34.165 -2.555 -33.835 ;
        RECT -2.885 -35.525 -2.555 -35.195 ;
        RECT -2.885 -36.885 -2.555 -36.555 ;
        RECT -2.885 -38.245 -2.555 -37.915 ;
        RECT -2.885 -40.965 -2.555 -40.635 ;
        RECT -2.885 -42.325 -2.555 -41.995 ;
        RECT -2.885 -43.685 -2.555 -43.355 ;
        RECT -2.885 -45.045 -2.555 -44.715 ;
        RECT -2.885 -49.125 -2.555 -48.795 ;
        RECT -2.885 -50.485 -2.555 -50.155 ;
        RECT -2.885 -51.845 -2.555 -51.515 ;
        RECT -2.885 -53.205 -2.555 -52.875 ;
        RECT -2.885 -54.565 -2.555 -54.235 ;
        RECT -2.885 -55.925 -2.555 -55.595 ;
        RECT -2.885 -57.285 -2.555 -56.955 ;
        RECT -2.885 -58.645 -2.555 -58.315 ;
        RECT -2.885 -60.005 -2.555 -59.675 ;
        RECT -2.885 -61.365 -2.555 -61.035 ;
        RECT -2.885 -62.725 -2.555 -62.395 ;
        RECT -2.885 -64.085 -2.555 -63.755 ;
        RECT -2.885 -65.445 -2.555 -65.115 ;
        RECT -2.885 -66.805 -2.555 -66.475 ;
        RECT -2.885 -68.165 -2.555 -67.835 ;
        RECT -2.885 -69.525 -2.555 -69.195 ;
        RECT -2.885 -70.885 -2.555 -70.555 ;
        RECT -2.885 -72.245 -2.555 -71.915 ;
        RECT -2.885 -73.605 -2.555 -73.275 ;
        RECT -2.885 -74.965 -2.555 -74.635 ;
        RECT -2.885 -76.325 -2.555 -75.995 ;
        RECT -2.885 -77.685 -2.555 -77.355 ;
        RECT -2.885 -79.045 -2.555 -78.715 ;
        RECT -2.885 -80.405 -2.555 -80.075 ;
        RECT -2.885 -81.765 -2.555 -81.435 ;
        RECT -2.885 -83.125 -2.555 -82.795 ;
        RECT -2.885 -84.485 -2.555 -84.155 ;
        RECT -2.885 -85.845 -2.555 -85.515 ;
        RECT -2.885 -87.205 -2.555 -86.875 ;
        RECT -2.885 -88.565 -2.555 -88.235 ;
        RECT -2.885 -89.925 -2.555 -89.595 ;
        RECT -2.885 -91.285 -2.555 -90.955 ;
        RECT -2.885 -92.645 -2.555 -92.315 ;
        RECT -2.885 -94.005 -2.555 -93.675 ;
        RECT -2.885 -95.365 -2.555 -95.035 ;
        RECT -2.885 -96.725 -2.555 -96.395 ;
        RECT -2.885 -98.085 -2.555 -97.755 ;
        RECT -2.885 -99.445 -2.555 -99.115 ;
        RECT -2.885 -100.805 -2.555 -100.475 ;
        RECT -2.885 -102.165 -2.555 -101.835 ;
        RECT -2.885 -103.525 -2.555 -103.195 ;
        RECT -2.885 -104.885 -2.555 -104.555 ;
        RECT -2.885 -106.245 -2.555 -105.915 ;
        RECT -2.885 -107.605 -2.555 -107.275 ;
        RECT -2.885 -108.965 -2.555 -108.635 ;
        RECT -2.885 -110.325 -2.555 -109.995 ;
        RECT -2.885 -111.685 -2.555 -111.355 ;
        RECT -2.885 -113.045 -2.555 -112.715 ;
        RECT -2.885 -114.405 -2.555 -114.075 ;
        RECT -2.885 -115.765 -2.555 -115.435 ;
        RECT -2.885 -117.125 -2.555 -116.795 ;
        RECT -2.885 -118.485 -2.555 -118.155 ;
        RECT -2.885 -119.845 -2.555 -119.515 ;
        RECT -2.885 -121.205 -2.555 -120.875 ;
        RECT -2.885 -122.565 -2.555 -122.235 ;
        RECT -2.885 -123.925 -2.555 -123.595 ;
        RECT -2.885 -125.285 -2.555 -124.955 ;
        RECT -2.885 -126.645 -2.555 -126.315 ;
        RECT -2.885 -128.005 -2.555 -127.675 ;
        RECT -2.885 -129.365 -2.555 -129.035 ;
        RECT -2.885 -130.725 -2.555 -130.395 ;
        RECT -2.885 -132.085 -2.555 -131.755 ;
        RECT -2.885 -133.445 -2.555 -133.115 ;
        RECT -2.885 -134.805 -2.555 -134.475 ;
        RECT -2.885 -136.165 -2.555 -135.835 ;
        RECT -2.885 -137.525 -2.555 -137.195 ;
        RECT -2.885 -138.885 -2.555 -138.555 ;
        RECT -2.885 -140.245 -2.555 -139.915 ;
        RECT -2.885 -141.605 -2.555 -141.275 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 127.225 -20.235 128.355 ;
        RECT -20.565 124.955 -20.235 125.285 ;
        RECT -20.565 123.595 -20.235 123.925 ;
        RECT -20.565 122.235 -20.235 122.565 ;
        RECT -20.565 120.875 -20.235 121.205 ;
        RECT -20.565 119.515 -20.235 119.845 ;
        RECT -20.565 118.155 -20.235 118.485 ;
        RECT -20.565 116.795 -20.235 117.125 ;
        RECT -20.565 115.435 -20.235 115.765 ;
        RECT -20.565 114.075 -20.235 114.405 ;
        RECT -20.565 112.715 -20.235 113.045 ;
        RECT -20.565 111.355 -20.235 111.685 ;
        RECT -20.565 109.995 -20.235 110.325 ;
        RECT -20.565 108.635 -20.235 108.965 ;
        RECT -20.565 107.275 -20.235 107.605 ;
        RECT -20.565 105.915 -20.235 106.245 ;
        RECT -20.565 104.555 -20.235 104.885 ;
        RECT -20.565 103.195 -20.235 103.525 ;
        RECT -20.565 101.835 -20.235 102.165 ;
        RECT -20.565 100.475 -20.235 100.805 ;
        RECT -20.565 99.115 -20.235 99.445 ;
        RECT -20.565 97.755 -20.235 98.085 ;
        RECT -20.565 96.395 -20.235 96.725 ;
        RECT -20.565 95.035 -20.235 95.365 ;
        RECT -20.565 93.675 -20.235 94.005 ;
        RECT -20.565 92.315 -20.235 92.645 ;
        RECT -20.565 90.955 -20.235 91.285 ;
        RECT -20.565 89.595 -20.235 89.925 ;
        RECT -20.565 88.235 -20.235 88.565 ;
        RECT -20.565 86.875 -20.235 87.205 ;
        RECT -20.565 85.515 -20.235 85.845 ;
        RECT -20.565 84.155 -20.235 84.485 ;
        RECT -20.565 82.795 -20.235 83.125 ;
        RECT -20.565 81.435 -20.235 81.765 ;
        RECT -20.565 80.075 -20.235 80.405 ;
        RECT -20.565 78.715 -20.235 79.045 ;
        RECT -20.565 77.355 -20.235 77.685 ;
        RECT -20.565 75.995 -20.235 76.325 ;
        RECT -20.565 74.635 -20.235 74.965 ;
        RECT -20.565 73.275 -20.235 73.605 ;
        RECT -20.565 71.915 -20.235 72.245 ;
        RECT -20.565 70.555 -20.235 70.885 ;
        RECT -20.565 69.195 -20.235 69.525 ;
        RECT -20.565 67.835 -20.235 68.165 ;
        RECT -20.565 66.475 -20.235 66.805 ;
        RECT -20.565 65.115 -20.235 65.445 ;
        RECT -20.565 63.755 -20.235 64.085 ;
        RECT -20.565 62.395 -20.235 62.725 ;
        RECT -20.565 61.035 -20.235 61.365 ;
        RECT -20.565 59.675 -20.235 60.005 ;
        RECT -20.565 58.315 -20.235 58.645 ;
        RECT -20.565 56.955 -20.235 57.285 ;
        RECT -20.565 55.595 -20.235 55.925 ;
        RECT -20.565 54.235 -20.235 54.565 ;
        RECT -20.565 52.875 -20.235 53.205 ;
        RECT -20.565 51.515 -20.235 51.845 ;
        RECT -20.565 50.155 -20.235 50.485 ;
        RECT -20.565 48.795 -20.235 49.125 ;
        RECT -20.565 47.435 -20.235 47.765 ;
        RECT -20.565 46.075 -20.235 46.405 ;
        RECT -20.565 44.715 -20.235 45.045 ;
        RECT -20.565 43.355 -20.235 43.685 ;
        RECT -20.565 41.995 -20.235 42.325 ;
        RECT -20.565 40.635 -20.235 40.965 ;
        RECT -20.565 39.275 -20.235 39.605 ;
        RECT -20.565 37.915 -20.235 38.245 ;
        RECT -20.565 36.555 -20.235 36.885 ;
        RECT -20.565 35.195 -20.235 35.525 ;
        RECT -20.565 33.835 -20.235 34.165 ;
        RECT -20.565 32.475 -20.235 32.805 ;
        RECT -20.565 31.115 -20.235 31.445 ;
        RECT -20.565 29.755 -20.235 30.085 ;
        RECT -20.565 28.395 -20.235 28.725 ;
        RECT -20.565 27.035 -20.235 27.365 ;
        RECT -20.565 25.675 -20.235 26.005 ;
        RECT -20.565 24.315 -20.235 24.645 ;
        RECT -20.565 22.955 -20.235 23.285 ;
        RECT -20.565 21.595 -20.235 21.925 ;
        RECT -20.565 20.235 -20.235 20.565 ;
        RECT -20.565 18.875 -20.235 19.205 ;
        RECT -20.565 17.515 -20.235 17.845 ;
        RECT -20.565 16.155 -20.235 16.485 ;
        RECT -20.565 14.795 -20.235 15.125 ;
        RECT -20.565 13.435 -20.235 13.765 ;
        RECT -20.565 12.075 -20.235 12.405 ;
        RECT -20.565 10.715 -20.235 11.045 ;
        RECT -20.565 9.355 -20.235 9.685 ;
        RECT -20.565 7.995 -20.235 8.325 ;
        RECT -20.565 6.635 -20.235 6.965 ;
        RECT -20.565 5.275 -20.235 5.605 ;
        RECT -20.565 3.915 -20.235 4.245 ;
        RECT -20.565 2.555 -20.235 2.885 ;
        RECT -20.565 1.195 -20.235 1.525 ;
        RECT -20.565 -0.165 -20.235 0.165 ;
        RECT -20.565 -1.525 -20.235 -1.195 ;
        RECT -20.565 -2.885 -20.235 -2.555 ;
        RECT -20.565 -6.965 -20.235 -6.635 ;
        RECT -20.565 -12.41 -20.235 -12.08 ;
        RECT -20.565 -15.125 -20.235 -14.795 ;
        RECT -20.565 -16.485 -20.235 -16.155 ;
        RECT -20.565 -17.25 -20.235 -16.92 ;
        RECT -20.565 -19.205 -20.235 -18.875 ;
        RECT -20.56 -20.56 -20.24 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -27.365 -20.235 -27.035 ;
        RECT -20.565 -28.725 -20.235 -28.395 ;
        RECT -20.565 -30.085 -20.235 -29.755 ;
        RECT -20.565 -32.805 -20.235 -32.475 ;
        RECT -20.565 -34.165 -20.235 -33.835 ;
        RECT -20.565 -35.39 -20.235 -35.06 ;
        RECT -20.565 -38.245 -20.235 -37.915 ;
        RECT -20.565 -40.23 -20.235 -39.9 ;
        RECT -20.565 -40.965 -20.235 -40.635 ;
        RECT -20.56 -43.68 -20.24 -26.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -50.485 -20.235 -50.155 ;
        RECT -20.565 -51.845 -20.235 -51.515 ;
        RECT -20.565 -54.565 -20.235 -54.235 ;
        RECT -20.565 -57.285 -20.235 -56.955 ;
        RECT -20.565 -58.645 -20.235 -58.315 ;
        RECT -20.565 -61.365 -20.235 -61.035 ;
        RECT -20.565 -62.725 -20.235 -62.395 ;
        RECT -20.565 -64.085 -20.235 -63.755 ;
        RECT -20.565 -66.805 -20.235 -66.475 ;
        RECT -20.56 -67.48 -20.24 -49.48 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -103.525 -20.235 -103.195 ;
        RECT -20.565 -104.885 -20.235 -104.555 ;
        RECT -20.565 -106.245 -20.235 -105.915 ;
        RECT -20.565 -107.605 -20.235 -107.275 ;
        RECT -20.565 -114.405 -20.235 -114.075 ;
        RECT -20.565 -118.485 -20.235 -118.155 ;
        RECT -20.565 -122.565 -20.235 -122.235 ;
        RECT -20.565 -125.285 -20.235 -124.955 ;
        RECT -20.565 -126.645 -20.235 -126.315 ;
        RECT -20.565 -128.005 -20.235 -127.675 ;
        RECT -20.565 -130.725 -20.235 -130.395 ;
        RECT -20.565 -132.085 -20.235 -131.755 ;
        RECT -20.565 -137.525 -20.235 -137.195 ;
        RECT -20.565 -138.885 -20.235 -138.555 ;
        RECT -20.565 -140.245 -20.235 -139.915 ;
        RECT -20.565 -141.605 -20.235 -141.275 ;
        RECT -20.565 -142.965 -20.235 -142.635 ;
        RECT -20.565 -144.325 -20.235 -143.995 ;
        RECT -20.565 -145.685 -20.235 -145.355 ;
        RECT -20.565 -147.045 -20.235 -146.715 ;
        RECT -20.565 -149.765 -20.235 -149.435 ;
        RECT -20.565 -152.485 -20.235 -152.155 ;
        RECT -20.565 -153.845 -20.235 -153.515 ;
        RECT -20.565 -155.285 -20.235 -154.955 ;
        RECT -20.565 -156.565 -20.235 -156.235 ;
        RECT -20.565 -157.925 -20.235 -157.595 ;
        RECT -20.565 -160.17 -20.235 -159.04 ;
        RECT -20.56 -160.285 -20.24 -99.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 127.225 -18.875 128.355 ;
        RECT -19.205 124.955 -18.875 125.285 ;
        RECT -19.205 123.595 -18.875 123.925 ;
        RECT -19.205 122.235 -18.875 122.565 ;
        RECT -19.205 120.875 -18.875 121.205 ;
        RECT -19.205 119.515 -18.875 119.845 ;
        RECT -19.205 118.155 -18.875 118.485 ;
        RECT -19.205 116.795 -18.875 117.125 ;
        RECT -19.205 115.435 -18.875 115.765 ;
        RECT -19.205 114.075 -18.875 114.405 ;
        RECT -19.205 112.715 -18.875 113.045 ;
        RECT -19.205 111.355 -18.875 111.685 ;
        RECT -19.205 109.995 -18.875 110.325 ;
        RECT -19.205 108.635 -18.875 108.965 ;
        RECT -19.205 107.275 -18.875 107.605 ;
        RECT -19.205 105.915 -18.875 106.245 ;
        RECT -19.205 104.555 -18.875 104.885 ;
        RECT -19.205 103.195 -18.875 103.525 ;
        RECT -19.205 101.835 -18.875 102.165 ;
        RECT -19.205 100.475 -18.875 100.805 ;
        RECT -19.205 99.115 -18.875 99.445 ;
        RECT -19.205 97.755 -18.875 98.085 ;
        RECT -19.205 96.395 -18.875 96.725 ;
        RECT -19.205 95.035 -18.875 95.365 ;
        RECT -19.205 93.675 -18.875 94.005 ;
        RECT -19.205 92.315 -18.875 92.645 ;
        RECT -19.205 90.955 -18.875 91.285 ;
        RECT -19.205 89.595 -18.875 89.925 ;
        RECT -19.205 88.235 -18.875 88.565 ;
        RECT -19.205 86.875 -18.875 87.205 ;
        RECT -19.205 85.515 -18.875 85.845 ;
        RECT -19.205 84.155 -18.875 84.485 ;
        RECT -19.205 82.795 -18.875 83.125 ;
        RECT -19.205 81.435 -18.875 81.765 ;
        RECT -19.205 80.075 -18.875 80.405 ;
        RECT -19.205 78.715 -18.875 79.045 ;
        RECT -19.205 77.355 -18.875 77.685 ;
        RECT -19.205 75.995 -18.875 76.325 ;
        RECT -19.205 74.635 -18.875 74.965 ;
        RECT -19.205 73.275 -18.875 73.605 ;
        RECT -19.205 71.915 -18.875 72.245 ;
        RECT -19.205 70.555 -18.875 70.885 ;
        RECT -19.205 69.195 -18.875 69.525 ;
        RECT -19.205 67.835 -18.875 68.165 ;
        RECT -19.205 66.475 -18.875 66.805 ;
        RECT -19.205 65.115 -18.875 65.445 ;
        RECT -19.205 63.755 -18.875 64.085 ;
        RECT -19.205 62.395 -18.875 62.725 ;
        RECT -19.205 61.035 -18.875 61.365 ;
        RECT -19.205 59.675 -18.875 60.005 ;
        RECT -19.205 58.315 -18.875 58.645 ;
        RECT -19.205 56.955 -18.875 57.285 ;
        RECT -19.205 55.595 -18.875 55.925 ;
        RECT -19.205 54.235 -18.875 54.565 ;
        RECT -19.205 52.875 -18.875 53.205 ;
        RECT -19.205 51.515 -18.875 51.845 ;
        RECT -19.205 50.155 -18.875 50.485 ;
        RECT -19.205 48.795 -18.875 49.125 ;
        RECT -19.205 47.435 -18.875 47.765 ;
        RECT -19.205 46.075 -18.875 46.405 ;
        RECT -19.205 44.715 -18.875 45.045 ;
        RECT -19.205 43.355 -18.875 43.685 ;
        RECT -19.205 41.995 -18.875 42.325 ;
        RECT -19.205 40.635 -18.875 40.965 ;
        RECT -19.205 39.275 -18.875 39.605 ;
        RECT -19.205 37.915 -18.875 38.245 ;
        RECT -19.205 36.555 -18.875 36.885 ;
        RECT -19.205 35.195 -18.875 35.525 ;
        RECT -19.205 33.835 -18.875 34.165 ;
        RECT -19.205 32.475 -18.875 32.805 ;
        RECT -19.205 31.115 -18.875 31.445 ;
        RECT -19.205 29.755 -18.875 30.085 ;
        RECT -19.205 28.395 -18.875 28.725 ;
        RECT -19.205 27.035 -18.875 27.365 ;
        RECT -19.205 25.675 -18.875 26.005 ;
        RECT -19.205 24.315 -18.875 24.645 ;
        RECT -19.205 22.955 -18.875 23.285 ;
        RECT -19.205 21.595 -18.875 21.925 ;
        RECT -19.205 20.235 -18.875 20.565 ;
        RECT -19.205 18.875 -18.875 19.205 ;
        RECT -19.205 17.515 -18.875 17.845 ;
        RECT -19.205 16.155 -18.875 16.485 ;
        RECT -19.205 14.795 -18.875 15.125 ;
        RECT -19.205 13.435 -18.875 13.765 ;
        RECT -19.205 12.075 -18.875 12.405 ;
        RECT -19.205 10.715 -18.875 11.045 ;
        RECT -19.205 9.355 -18.875 9.685 ;
        RECT -19.205 7.995 -18.875 8.325 ;
        RECT -19.205 6.635 -18.875 6.965 ;
        RECT -19.205 5.275 -18.875 5.605 ;
        RECT -19.205 3.915 -18.875 4.245 ;
        RECT -19.205 2.555 -18.875 2.885 ;
        RECT -19.205 1.195 -18.875 1.525 ;
        RECT -19.205 -0.165 -18.875 0.165 ;
        RECT -19.205 -1.525 -18.875 -1.195 ;
        RECT -19.205 -2.885 -18.875 -2.555 ;
        RECT -19.205 -6.965 -18.875 -6.635 ;
        RECT -19.205 -12.41 -18.875 -12.08 ;
        RECT -19.205 -15.125 -18.875 -14.795 ;
        RECT -19.205 -16.485 -18.875 -16.155 ;
        RECT -19.205 -17.25 -18.875 -16.92 ;
        RECT -19.205 -19.205 -18.875 -18.875 ;
        RECT -19.2 -19.88 -18.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -27.365 -18.875 -27.035 ;
        RECT -19.205 -28.725 -18.875 -28.395 ;
        RECT -19.205 -30.085 -18.875 -29.755 ;
        RECT -19.205 -32.805 -18.875 -32.475 ;
        RECT -19.205 -34.165 -18.875 -33.835 ;
        RECT -19.205 -35.39 -18.875 -35.06 ;
        RECT -19.205 -38.245 -18.875 -37.915 ;
        RECT -19.205 -40.23 -18.875 -39.9 ;
        RECT -19.205 -40.965 -18.875 -40.635 ;
        RECT -19.2 -43 -18.88 -25 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -49.125 -18.875 -48.795 ;
        RECT -19.205 -50.485 -18.875 -50.155 ;
        RECT -19.205 -51.845 -18.875 -51.515 ;
        RECT -19.205 -54.565 -18.875 -54.235 ;
        RECT -19.205 -56.27 -18.875 -55.94 ;
        RECT -19.205 -57.285 -18.875 -56.955 ;
        RECT -19.205 -58.645 -18.875 -58.315 ;
        RECT -19.205 -61.365 -18.875 -61.035 ;
        RECT -19.205 -62.725 -18.875 -62.395 ;
        RECT -19.205 -64.085 -18.875 -63.755 ;
        RECT -19.205 -64.81 -18.875 -64.48 ;
        RECT -19.205 -66.805 -18.875 -66.475 ;
        RECT -19.205 -69.525 -18.875 -69.195 ;
        RECT -19.205 -70.885 -18.875 -70.555 ;
        RECT -19.205 -72.245 -18.875 -71.915 ;
        RECT -19.205 -73.605 -18.875 -73.275 ;
        RECT -19.205 -76.325 -18.875 -75.995 ;
        RECT -19.205 -77.685 -18.875 -77.355 ;
        RECT -19.205 -78.45 -18.875 -78.12 ;
        RECT -19.205 -80.405 -18.875 -80.075 ;
        RECT -19.205 -81.765 -18.875 -81.435 ;
        RECT -19.205 -84.485 -18.875 -84.155 ;
        RECT -19.205 -85.845 -18.875 -85.515 ;
        RECT -19.205 -86.99 -18.875 -86.66 ;
        RECT -19.205 -88.565 -18.875 -88.235 ;
        RECT -19.205 -94.005 -18.875 -93.675 ;
        RECT -19.205 -95.365 -18.875 -95.035 ;
        RECT -19.205 -96.725 -18.875 -96.395 ;
        RECT -19.205 -98.085 -18.875 -97.755 ;
        RECT -19.205 -103.525 -18.875 -103.195 ;
        RECT -19.205 -104.885 -18.875 -104.555 ;
        RECT -19.205 -106.245 -18.875 -105.915 ;
        RECT -19.205 -114.405 -18.875 -114.075 ;
        RECT -19.205 -118.485 -18.875 -118.155 ;
        RECT -19.205 -122.565 -18.875 -122.235 ;
        RECT -19.205 -123.925 -18.875 -123.595 ;
        RECT -19.205 -125.285 -18.875 -124.955 ;
        RECT -19.205 -128.005 -18.875 -127.675 ;
        RECT -19.205 -130.725 -18.875 -130.395 ;
        RECT -19.205 -132.085 -18.875 -131.755 ;
        RECT -19.205 -137.525 -18.875 -137.195 ;
        RECT -19.205 -138.885 -18.875 -138.555 ;
        RECT -19.205 -140.245 -18.875 -139.915 ;
        RECT -19.205 -141.605 -18.875 -141.275 ;
        RECT -19.205 -142.965 -18.875 -142.635 ;
        RECT -19.205 -144.325 -18.875 -143.995 ;
        RECT -19.205 -145.685 -18.875 -145.355 ;
        RECT -19.205 -147.045 -18.875 -146.715 ;
        RECT -19.205 -149.765 -18.875 -149.435 ;
        RECT -19.205 -152.485 -18.875 -152.155 ;
        RECT -19.205 -153.845 -18.875 -153.515 ;
        RECT -19.205 -155.285 -18.875 -154.955 ;
        RECT -19.205 -156.565 -18.875 -156.235 ;
        RECT -19.205 -157.925 -18.875 -157.595 ;
        RECT -19.205 -160.17 -18.875 -159.04 ;
        RECT -19.2 -160.285 -18.88 -48.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 127.225 -17.515 128.355 ;
        RECT -17.845 124.955 -17.515 125.285 ;
        RECT -17.845 123.595 -17.515 123.925 ;
        RECT -17.845 122.235 -17.515 122.565 ;
        RECT -17.845 120.875 -17.515 121.205 ;
        RECT -17.845 119.515 -17.515 119.845 ;
        RECT -17.845 118.155 -17.515 118.485 ;
        RECT -17.845 116.795 -17.515 117.125 ;
        RECT -17.845 115.435 -17.515 115.765 ;
        RECT -17.845 114.075 -17.515 114.405 ;
        RECT -17.845 112.715 -17.515 113.045 ;
        RECT -17.845 111.355 -17.515 111.685 ;
        RECT -17.845 109.995 -17.515 110.325 ;
        RECT -17.845 108.635 -17.515 108.965 ;
        RECT -17.845 107.275 -17.515 107.605 ;
        RECT -17.845 105.915 -17.515 106.245 ;
        RECT -17.845 104.555 -17.515 104.885 ;
        RECT -17.845 103.195 -17.515 103.525 ;
        RECT -17.845 101.835 -17.515 102.165 ;
        RECT -17.845 100.475 -17.515 100.805 ;
        RECT -17.845 99.115 -17.515 99.445 ;
        RECT -17.845 97.755 -17.515 98.085 ;
        RECT -17.845 96.395 -17.515 96.725 ;
        RECT -17.845 95.035 -17.515 95.365 ;
        RECT -17.845 93.675 -17.515 94.005 ;
        RECT -17.845 92.315 -17.515 92.645 ;
        RECT -17.845 90.955 -17.515 91.285 ;
        RECT -17.845 89.595 -17.515 89.925 ;
        RECT -17.845 88.235 -17.515 88.565 ;
        RECT -17.845 86.875 -17.515 87.205 ;
        RECT -17.845 85.515 -17.515 85.845 ;
        RECT -17.845 84.155 -17.515 84.485 ;
        RECT -17.845 82.795 -17.515 83.125 ;
        RECT -17.845 81.435 -17.515 81.765 ;
        RECT -17.845 80.075 -17.515 80.405 ;
        RECT -17.845 78.715 -17.515 79.045 ;
        RECT -17.845 77.355 -17.515 77.685 ;
        RECT -17.845 75.995 -17.515 76.325 ;
        RECT -17.845 74.635 -17.515 74.965 ;
        RECT -17.845 73.275 -17.515 73.605 ;
        RECT -17.845 71.915 -17.515 72.245 ;
        RECT -17.845 70.555 -17.515 70.885 ;
        RECT -17.845 69.195 -17.515 69.525 ;
        RECT -17.845 67.835 -17.515 68.165 ;
        RECT -17.845 66.475 -17.515 66.805 ;
        RECT -17.845 65.115 -17.515 65.445 ;
        RECT -17.845 63.755 -17.515 64.085 ;
        RECT -17.845 62.395 -17.515 62.725 ;
        RECT -17.845 61.035 -17.515 61.365 ;
        RECT -17.845 59.675 -17.515 60.005 ;
        RECT -17.845 58.315 -17.515 58.645 ;
        RECT -17.845 56.955 -17.515 57.285 ;
        RECT -17.845 55.595 -17.515 55.925 ;
        RECT -17.845 54.235 -17.515 54.565 ;
        RECT -17.845 52.875 -17.515 53.205 ;
        RECT -17.845 51.515 -17.515 51.845 ;
        RECT -17.845 50.155 -17.515 50.485 ;
        RECT -17.845 48.795 -17.515 49.125 ;
        RECT -17.845 47.435 -17.515 47.765 ;
        RECT -17.845 46.075 -17.515 46.405 ;
        RECT -17.845 44.715 -17.515 45.045 ;
        RECT -17.845 43.355 -17.515 43.685 ;
        RECT -17.845 41.995 -17.515 42.325 ;
        RECT -17.845 40.635 -17.515 40.965 ;
        RECT -17.845 39.275 -17.515 39.605 ;
        RECT -17.845 37.915 -17.515 38.245 ;
        RECT -17.845 36.555 -17.515 36.885 ;
        RECT -17.845 35.195 -17.515 35.525 ;
        RECT -17.845 33.835 -17.515 34.165 ;
        RECT -17.845 32.475 -17.515 32.805 ;
        RECT -17.845 31.115 -17.515 31.445 ;
        RECT -17.845 29.755 -17.515 30.085 ;
        RECT -17.845 28.395 -17.515 28.725 ;
        RECT -17.845 27.035 -17.515 27.365 ;
        RECT -17.845 25.675 -17.515 26.005 ;
        RECT -17.845 24.315 -17.515 24.645 ;
        RECT -17.845 22.955 -17.515 23.285 ;
        RECT -17.845 21.595 -17.515 21.925 ;
        RECT -17.845 20.235 -17.515 20.565 ;
        RECT -17.845 18.875 -17.515 19.205 ;
        RECT -17.845 17.515 -17.515 17.845 ;
        RECT -17.845 16.155 -17.515 16.485 ;
        RECT -17.845 14.795 -17.515 15.125 ;
        RECT -17.845 13.435 -17.515 13.765 ;
        RECT -17.845 12.075 -17.515 12.405 ;
        RECT -17.845 10.715 -17.515 11.045 ;
        RECT -17.845 9.355 -17.515 9.685 ;
        RECT -17.845 7.995 -17.515 8.325 ;
        RECT -17.845 6.635 -17.515 6.965 ;
        RECT -17.845 5.275 -17.515 5.605 ;
        RECT -17.845 3.915 -17.515 4.245 ;
        RECT -17.845 2.555 -17.515 2.885 ;
        RECT -17.845 1.195 -17.515 1.525 ;
        RECT -17.845 -0.165 -17.515 0.165 ;
        RECT -17.845 -1.525 -17.515 -1.195 ;
        RECT -17.845 -2.885 -17.515 -2.555 ;
        RECT -17.845 -6.965 -17.515 -6.635 ;
        RECT -17.845 -12.41 -17.515 -12.08 ;
        RECT -17.845 -15.125 -17.515 -14.795 ;
        RECT -17.845 -16.485 -17.515 -16.155 ;
        RECT -17.845 -17.25 -17.515 -16.92 ;
        RECT -17.845 -19.205 -17.515 -18.875 ;
        RECT -17.84 -19.205 -17.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 -24.645 -17.515 -24.315 ;
        RECT -17.845 -27.365 -17.515 -27.035 ;
        RECT -17.845 -28.725 -17.515 -28.395 ;
        RECT -17.845 -30.085 -17.515 -29.755 ;
        RECT -17.845 -32.805 -17.515 -32.475 ;
        RECT -17.845 -34.165 -17.515 -33.835 ;
        RECT -17.845 -35.39 -17.515 -35.06 ;
        RECT -17.845 -38.245 -17.515 -37.915 ;
        RECT -17.845 -40.23 -17.515 -39.9 ;
        RECT -17.845 -40.965 -17.515 -40.635 ;
        RECT -17.84 -41.64 -17.52 -23.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 -47.765 -17.515 -47.435 ;
        RECT -17.845 -49.125 -17.515 -48.795 ;
        RECT -17.845 -50.485 -17.515 -50.155 ;
        RECT -17.845 -51.845 -17.515 -51.515 ;
        RECT -17.845 -54.565 -17.515 -54.235 ;
        RECT -17.845 -56.27 -17.515 -55.94 ;
        RECT -17.845 -57.285 -17.515 -56.955 ;
        RECT -17.845 -58.645 -17.515 -58.315 ;
        RECT -17.845 -61.365 -17.515 -61.035 ;
        RECT -17.845 -62.725 -17.515 -62.395 ;
        RECT -17.845 -64.085 -17.515 -63.755 ;
        RECT -17.845 -64.81 -17.515 -64.48 ;
        RECT -17.845 -66.805 -17.515 -66.475 ;
        RECT -17.845 -69.525 -17.515 -69.195 ;
        RECT -17.845 -70.885 -17.515 -70.555 ;
        RECT -17.845 -72.245 -17.515 -71.915 ;
        RECT -17.845 -73.605 -17.515 -73.275 ;
        RECT -17.845 -76.325 -17.515 -75.995 ;
        RECT -17.845 -77.685 -17.515 -77.355 ;
        RECT -17.845 -78.45 -17.515 -78.12 ;
        RECT -17.845 -80.405 -17.515 -80.075 ;
        RECT -17.845 -81.765 -17.515 -81.435 ;
        RECT -17.845 -84.485 -17.515 -84.155 ;
        RECT -17.845 -85.845 -17.515 -85.515 ;
        RECT -17.845 -86.99 -17.515 -86.66 ;
        RECT -17.845 -88.565 -17.515 -88.235 ;
        RECT -17.845 -94.005 -17.515 -93.675 ;
        RECT -17.845 -95.365 -17.515 -95.035 ;
        RECT -17.845 -96.725 -17.515 -96.395 ;
        RECT -17.845 -106.245 -17.515 -105.915 ;
        RECT -17.845 -118.485 -17.515 -118.155 ;
        RECT -17.845 -123.925 -17.515 -123.595 ;
        RECT -17.845 -125.285 -17.515 -124.955 ;
        RECT -17.845 -130.725 -17.515 -130.395 ;
        RECT -17.845 -132.085 -17.515 -131.755 ;
        RECT -17.845 -136.165 -17.515 -135.835 ;
        RECT -17.845 -137.525 -17.515 -137.195 ;
        RECT -17.845 -138.885 -17.515 -138.555 ;
        RECT -17.845 -140.245 -17.515 -139.915 ;
        RECT -17.845 -141.605 -17.515 -141.275 ;
        RECT -17.845 -142.965 -17.515 -142.635 ;
        RECT -17.845 -144.325 -17.515 -143.995 ;
        RECT -17.845 -145.685 -17.515 -145.355 ;
        RECT -17.845 -147.045 -17.515 -146.715 ;
        RECT -17.845 -149.765 -17.515 -149.435 ;
        RECT -17.845 -152.485 -17.515 -152.155 ;
        RECT -17.845 -153.845 -17.515 -153.515 ;
        RECT -17.845 -155.285 -17.515 -154.955 ;
        RECT -17.845 -156.565 -17.515 -156.235 ;
        RECT -17.845 -157.925 -17.515 -157.595 ;
        RECT -17.845 -160.17 -17.515 -159.04 ;
        RECT -17.84 -160.285 -17.52 -46.76 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 127.225 -16.155 128.355 ;
        RECT -16.485 124.955 -16.155 125.285 ;
        RECT -16.485 123.595 -16.155 123.925 ;
        RECT -16.485 122.235 -16.155 122.565 ;
        RECT -16.485 120.875 -16.155 121.205 ;
        RECT -16.485 119.515 -16.155 119.845 ;
        RECT -16.485 118.155 -16.155 118.485 ;
        RECT -16.485 116.795 -16.155 117.125 ;
        RECT -16.485 115.435 -16.155 115.765 ;
        RECT -16.485 114.075 -16.155 114.405 ;
        RECT -16.485 112.715 -16.155 113.045 ;
        RECT -16.485 111.355 -16.155 111.685 ;
        RECT -16.485 109.995 -16.155 110.325 ;
        RECT -16.485 108.635 -16.155 108.965 ;
        RECT -16.485 107.275 -16.155 107.605 ;
        RECT -16.485 105.915 -16.155 106.245 ;
        RECT -16.485 104.555 -16.155 104.885 ;
        RECT -16.485 103.195 -16.155 103.525 ;
        RECT -16.485 101.835 -16.155 102.165 ;
        RECT -16.485 100.475 -16.155 100.805 ;
        RECT -16.485 99.115 -16.155 99.445 ;
        RECT -16.485 97.755 -16.155 98.085 ;
        RECT -16.485 96.395 -16.155 96.725 ;
        RECT -16.485 95.035 -16.155 95.365 ;
        RECT -16.485 93.675 -16.155 94.005 ;
        RECT -16.485 92.315 -16.155 92.645 ;
        RECT -16.485 90.955 -16.155 91.285 ;
        RECT -16.485 89.595 -16.155 89.925 ;
        RECT -16.485 88.235 -16.155 88.565 ;
        RECT -16.485 86.875 -16.155 87.205 ;
        RECT -16.485 85.515 -16.155 85.845 ;
        RECT -16.485 84.155 -16.155 84.485 ;
        RECT -16.485 82.795 -16.155 83.125 ;
        RECT -16.485 81.435 -16.155 81.765 ;
        RECT -16.485 80.075 -16.155 80.405 ;
        RECT -16.485 78.715 -16.155 79.045 ;
        RECT -16.485 77.355 -16.155 77.685 ;
        RECT -16.485 75.995 -16.155 76.325 ;
        RECT -16.485 74.635 -16.155 74.965 ;
        RECT -16.485 73.275 -16.155 73.605 ;
        RECT -16.485 71.915 -16.155 72.245 ;
        RECT -16.485 70.555 -16.155 70.885 ;
        RECT -16.485 69.195 -16.155 69.525 ;
        RECT -16.485 67.835 -16.155 68.165 ;
        RECT -16.485 66.475 -16.155 66.805 ;
        RECT -16.485 65.115 -16.155 65.445 ;
        RECT -16.485 63.755 -16.155 64.085 ;
        RECT -16.485 62.395 -16.155 62.725 ;
        RECT -16.485 61.035 -16.155 61.365 ;
        RECT -16.485 59.675 -16.155 60.005 ;
        RECT -16.485 58.315 -16.155 58.645 ;
        RECT -16.485 56.955 -16.155 57.285 ;
        RECT -16.485 55.595 -16.155 55.925 ;
        RECT -16.485 54.235 -16.155 54.565 ;
        RECT -16.485 52.875 -16.155 53.205 ;
        RECT -16.485 51.515 -16.155 51.845 ;
        RECT -16.485 50.155 -16.155 50.485 ;
        RECT -16.485 48.795 -16.155 49.125 ;
        RECT -16.485 47.435 -16.155 47.765 ;
        RECT -16.485 46.075 -16.155 46.405 ;
        RECT -16.485 44.715 -16.155 45.045 ;
        RECT -16.485 43.355 -16.155 43.685 ;
        RECT -16.485 41.995 -16.155 42.325 ;
        RECT -16.485 40.635 -16.155 40.965 ;
        RECT -16.485 39.275 -16.155 39.605 ;
        RECT -16.485 37.915 -16.155 38.245 ;
        RECT -16.485 36.555 -16.155 36.885 ;
        RECT -16.485 35.195 -16.155 35.525 ;
        RECT -16.485 33.835 -16.155 34.165 ;
        RECT -16.485 32.475 -16.155 32.805 ;
        RECT -16.485 31.115 -16.155 31.445 ;
        RECT -16.485 29.755 -16.155 30.085 ;
        RECT -16.485 28.395 -16.155 28.725 ;
        RECT -16.485 27.035 -16.155 27.365 ;
        RECT -16.485 25.675 -16.155 26.005 ;
        RECT -16.485 24.315 -16.155 24.645 ;
        RECT -16.485 22.955 -16.155 23.285 ;
        RECT -16.485 21.595 -16.155 21.925 ;
        RECT -16.485 20.235 -16.155 20.565 ;
        RECT -16.485 18.875 -16.155 19.205 ;
        RECT -16.485 17.515 -16.155 17.845 ;
        RECT -16.485 16.155 -16.155 16.485 ;
        RECT -16.485 14.795 -16.155 15.125 ;
        RECT -16.485 13.435 -16.155 13.765 ;
        RECT -16.485 12.075 -16.155 12.405 ;
        RECT -16.485 10.715 -16.155 11.045 ;
        RECT -16.485 9.355 -16.155 9.685 ;
        RECT -16.485 7.995 -16.155 8.325 ;
        RECT -16.485 6.635 -16.155 6.965 ;
        RECT -16.485 5.275 -16.155 5.605 ;
        RECT -16.485 3.915 -16.155 4.245 ;
        RECT -16.485 2.555 -16.155 2.885 ;
        RECT -16.485 1.195 -16.155 1.525 ;
        RECT -16.485 -0.165 -16.155 0.165 ;
        RECT -16.485 -1.525 -16.155 -1.195 ;
        RECT -16.485 -2.885 -16.155 -2.555 ;
        RECT -16.485 -4.245 -16.155 -3.915 ;
        RECT -16.485 -6.965 -16.155 -6.635 ;
        RECT -16.48 -9 -16.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -24.645 -16.155 -24.315 ;
        RECT -16.485 -26.005 -16.155 -25.675 ;
        RECT -16.485 -27.365 -16.155 -27.035 ;
        RECT -16.485 -28.725 -16.155 -28.395 ;
        RECT -16.485 -30.085 -16.155 -29.755 ;
        RECT -16.48 -32.12 -16.16 -23.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -100.805 -16.155 -100.475 ;
        RECT -16.485 -106.245 -16.155 -105.915 ;
        RECT -16.485 -118.485 -16.155 -118.155 ;
        RECT -16.485 -123.925 -16.155 -123.595 ;
        RECT -16.485 -125.285 -16.155 -124.955 ;
        RECT -16.485 -130.725 -16.155 -130.395 ;
        RECT -16.485 -136.165 -16.155 -135.835 ;
        RECT -16.485 -137.525 -16.155 -137.195 ;
        RECT -16.485 -138.885 -16.155 -138.555 ;
        RECT -16.485 -140.245 -16.155 -139.915 ;
        RECT -16.485 -141.605 -16.155 -141.275 ;
        RECT -16.485 -142.965 -16.155 -142.635 ;
        RECT -16.485 -144.325 -16.155 -143.995 ;
        RECT -16.485 -145.685 -16.155 -145.355 ;
        RECT -16.485 -147.045 -16.155 -146.715 ;
        RECT -16.485 -149.765 -16.155 -149.435 ;
        RECT -16.485 -153.845 -16.155 -153.515 ;
        RECT -16.485 -155.285 -16.155 -154.955 ;
        RECT -16.485 -156.565 -16.155 -156.235 ;
        RECT -16.485 -157.925 -16.155 -157.595 ;
        RECT -16.485 -160.17 -16.155 -159.04 ;
        RECT -16.48 -160.285 -16.16 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 127.225 -14.795 128.355 ;
        RECT -15.125 124.955 -14.795 125.285 ;
        RECT -15.125 123.595 -14.795 123.925 ;
        RECT -15.125 122.235 -14.795 122.565 ;
        RECT -15.125 120.875 -14.795 121.205 ;
        RECT -15.125 119.515 -14.795 119.845 ;
        RECT -15.125 118.155 -14.795 118.485 ;
        RECT -15.125 116.795 -14.795 117.125 ;
        RECT -15.125 115.435 -14.795 115.765 ;
        RECT -15.125 114.075 -14.795 114.405 ;
        RECT -15.125 112.715 -14.795 113.045 ;
        RECT -15.125 111.355 -14.795 111.685 ;
        RECT -15.125 109.995 -14.795 110.325 ;
        RECT -15.125 108.635 -14.795 108.965 ;
        RECT -15.125 107.275 -14.795 107.605 ;
        RECT -15.125 105.915 -14.795 106.245 ;
        RECT -15.125 104.555 -14.795 104.885 ;
        RECT -15.125 103.195 -14.795 103.525 ;
        RECT -15.125 101.835 -14.795 102.165 ;
        RECT -15.125 100.475 -14.795 100.805 ;
        RECT -15.125 99.115 -14.795 99.445 ;
        RECT -15.125 97.755 -14.795 98.085 ;
        RECT -15.125 96.395 -14.795 96.725 ;
        RECT -15.125 95.035 -14.795 95.365 ;
        RECT -15.125 93.675 -14.795 94.005 ;
        RECT -15.125 92.315 -14.795 92.645 ;
        RECT -15.125 90.955 -14.795 91.285 ;
        RECT -15.125 89.595 -14.795 89.925 ;
        RECT -15.125 88.235 -14.795 88.565 ;
        RECT -15.125 86.875 -14.795 87.205 ;
        RECT -15.125 85.515 -14.795 85.845 ;
        RECT -15.125 84.155 -14.795 84.485 ;
        RECT -15.125 82.795 -14.795 83.125 ;
        RECT -15.125 81.435 -14.795 81.765 ;
        RECT -15.125 80.075 -14.795 80.405 ;
        RECT -15.125 78.715 -14.795 79.045 ;
        RECT -15.125 77.355 -14.795 77.685 ;
        RECT -15.125 75.995 -14.795 76.325 ;
        RECT -15.125 74.635 -14.795 74.965 ;
        RECT -15.125 73.275 -14.795 73.605 ;
        RECT -15.125 71.915 -14.795 72.245 ;
        RECT -15.125 70.555 -14.795 70.885 ;
        RECT -15.125 69.195 -14.795 69.525 ;
        RECT -15.125 67.835 -14.795 68.165 ;
        RECT -15.125 66.475 -14.795 66.805 ;
        RECT -15.125 65.115 -14.795 65.445 ;
        RECT -15.125 63.755 -14.795 64.085 ;
        RECT -15.125 62.395 -14.795 62.725 ;
        RECT -15.125 61.035 -14.795 61.365 ;
        RECT -15.125 59.675 -14.795 60.005 ;
        RECT -15.125 58.315 -14.795 58.645 ;
        RECT -15.125 56.955 -14.795 57.285 ;
        RECT -15.125 55.595 -14.795 55.925 ;
        RECT -15.125 54.235 -14.795 54.565 ;
        RECT -15.125 52.875 -14.795 53.205 ;
        RECT -15.125 51.515 -14.795 51.845 ;
        RECT -15.125 50.155 -14.795 50.485 ;
        RECT -15.125 48.795 -14.795 49.125 ;
        RECT -15.125 47.435 -14.795 47.765 ;
        RECT -15.125 46.075 -14.795 46.405 ;
        RECT -15.125 44.715 -14.795 45.045 ;
        RECT -15.125 43.355 -14.795 43.685 ;
        RECT -15.125 41.995 -14.795 42.325 ;
        RECT -15.125 40.635 -14.795 40.965 ;
        RECT -15.125 39.275 -14.795 39.605 ;
        RECT -15.125 37.915 -14.795 38.245 ;
        RECT -15.125 36.555 -14.795 36.885 ;
        RECT -15.125 35.195 -14.795 35.525 ;
        RECT -15.125 33.835 -14.795 34.165 ;
        RECT -15.125 32.475 -14.795 32.805 ;
        RECT -15.125 31.115 -14.795 31.445 ;
        RECT -15.125 29.755 -14.795 30.085 ;
        RECT -15.125 28.395 -14.795 28.725 ;
        RECT -15.125 27.035 -14.795 27.365 ;
        RECT -15.125 25.675 -14.795 26.005 ;
        RECT -15.125 24.315 -14.795 24.645 ;
        RECT -15.125 22.955 -14.795 23.285 ;
        RECT -15.125 21.595 -14.795 21.925 ;
        RECT -15.125 20.235 -14.795 20.565 ;
        RECT -15.125 18.875 -14.795 19.205 ;
        RECT -15.125 17.515 -14.795 17.845 ;
        RECT -15.125 16.155 -14.795 16.485 ;
        RECT -15.125 14.795 -14.795 15.125 ;
        RECT -15.125 13.435 -14.795 13.765 ;
        RECT -15.125 12.075 -14.795 12.405 ;
        RECT -15.125 10.715 -14.795 11.045 ;
        RECT -15.125 9.355 -14.795 9.685 ;
        RECT -15.125 7.995 -14.795 8.325 ;
        RECT -15.125 6.635 -14.795 6.965 ;
        RECT -15.125 5.275 -14.795 5.605 ;
        RECT -15.125 3.915 -14.795 4.245 ;
        RECT -15.125 2.555 -14.795 2.885 ;
        RECT -15.125 1.195 -14.795 1.525 ;
        RECT -15.125 -0.165 -14.795 0.165 ;
        RECT -15.125 -1.525 -14.795 -1.195 ;
        RECT -15.125 -2.885 -14.795 -2.555 ;
        RECT -15.125 -4.245 -14.795 -3.915 ;
        RECT -15.125 -6.965 -14.795 -6.635 ;
        RECT -15.125 -9.685 -14.795 -9.355 ;
        RECT -15.125 -12.41 -14.795 -12.08 ;
        RECT -15.125 -15.125 -14.795 -14.795 ;
        RECT -15.125 -16.485 -14.795 -16.155 ;
        RECT -15.125 -17.25 -14.795 -16.92 ;
        RECT -15.125 -19.205 -14.795 -18.875 ;
        RECT -15.125 -24.645 -14.795 -24.315 ;
        RECT -15.125 -26.005 -14.795 -25.675 ;
        RECT -15.125 -27.365 -14.795 -27.035 ;
        RECT -15.125 -28.725 -14.795 -28.395 ;
        RECT -15.125 -30.085 -14.795 -29.755 ;
        RECT -15.125 -34.165 -14.795 -33.835 ;
        RECT -15.125 -35.39 -14.795 -35.06 ;
        RECT -15.125 -38.245 -14.795 -37.915 ;
        RECT -15.125 -40.23 -14.795 -39.9 ;
        RECT -15.125 -40.965 -14.795 -40.635 ;
        RECT -15.125 -47.765 -14.795 -47.435 ;
        RECT -15.125 -49.125 -14.795 -48.795 ;
        RECT -15.125 -50.485 -14.795 -50.155 ;
        RECT -15.125 -51.845 -14.795 -51.515 ;
        RECT -15.125 -54.565 -14.795 -54.235 ;
        RECT -15.125 -56.27 -14.795 -55.94 ;
        RECT -15.125 -57.285 -14.795 -56.955 ;
        RECT -15.125 -58.645 -14.795 -58.315 ;
        RECT -15.125 -61.365 -14.795 -61.035 ;
        RECT -15.125 -62.725 -14.795 -62.395 ;
        RECT -15.125 -64.085 -14.795 -63.755 ;
        RECT -15.125 -64.81 -14.795 -64.48 ;
        RECT -15.125 -66.805 -14.795 -66.475 ;
        RECT -15.125 -69.525 -14.795 -69.195 ;
        RECT -15.125 -70.885 -14.795 -70.555 ;
        RECT -15.125 -72.245 -14.795 -71.915 ;
        RECT -15.125 -73.605 -14.795 -73.275 ;
        RECT -15.125 -76.325 -14.795 -75.995 ;
        RECT -15.125 -77.685 -14.795 -77.355 ;
        RECT -15.125 -78.45 -14.795 -78.12 ;
        RECT -15.125 -80.405 -14.795 -80.075 ;
        RECT -15.125 -81.765 -14.795 -81.435 ;
        RECT -15.125 -84.485 -14.795 -84.155 ;
        RECT -15.125 -85.845 -14.795 -85.515 ;
        RECT -15.125 -86.99 -14.795 -86.66 ;
        RECT -15.12 -89.92 -14.8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 127.225 -13.435 128.355 ;
        RECT -13.765 124.955 -13.435 125.285 ;
        RECT -13.765 123.595 -13.435 123.925 ;
        RECT -13.765 122.235 -13.435 122.565 ;
        RECT -13.765 120.875 -13.435 121.205 ;
        RECT -13.765 119.515 -13.435 119.845 ;
        RECT -13.765 118.155 -13.435 118.485 ;
        RECT -13.765 116.795 -13.435 117.125 ;
        RECT -13.765 115.435 -13.435 115.765 ;
        RECT -13.765 114.075 -13.435 114.405 ;
        RECT -13.765 112.715 -13.435 113.045 ;
        RECT -13.765 111.355 -13.435 111.685 ;
        RECT -13.765 109.995 -13.435 110.325 ;
        RECT -13.765 108.635 -13.435 108.965 ;
        RECT -13.765 107.275 -13.435 107.605 ;
        RECT -13.765 105.915 -13.435 106.245 ;
        RECT -13.765 104.555 -13.435 104.885 ;
        RECT -13.765 103.195 -13.435 103.525 ;
        RECT -13.765 101.835 -13.435 102.165 ;
        RECT -13.765 100.475 -13.435 100.805 ;
        RECT -13.765 99.115 -13.435 99.445 ;
        RECT -13.765 97.755 -13.435 98.085 ;
        RECT -13.765 96.395 -13.435 96.725 ;
        RECT -13.765 95.035 -13.435 95.365 ;
        RECT -13.765 93.675 -13.435 94.005 ;
        RECT -13.765 92.315 -13.435 92.645 ;
        RECT -13.765 90.955 -13.435 91.285 ;
        RECT -13.765 89.595 -13.435 89.925 ;
        RECT -13.765 88.235 -13.435 88.565 ;
        RECT -13.765 86.875 -13.435 87.205 ;
        RECT -13.765 85.515 -13.435 85.845 ;
        RECT -13.765 84.155 -13.435 84.485 ;
        RECT -13.765 82.795 -13.435 83.125 ;
        RECT -13.765 81.435 -13.435 81.765 ;
        RECT -13.765 80.075 -13.435 80.405 ;
        RECT -13.765 78.715 -13.435 79.045 ;
        RECT -13.765 77.355 -13.435 77.685 ;
        RECT -13.765 75.995 -13.435 76.325 ;
        RECT -13.765 74.635 -13.435 74.965 ;
        RECT -13.765 73.275 -13.435 73.605 ;
        RECT -13.765 71.915 -13.435 72.245 ;
        RECT -13.765 70.555 -13.435 70.885 ;
        RECT -13.765 69.195 -13.435 69.525 ;
        RECT -13.765 67.835 -13.435 68.165 ;
        RECT -13.765 66.475 -13.435 66.805 ;
        RECT -13.765 65.115 -13.435 65.445 ;
        RECT -13.765 63.755 -13.435 64.085 ;
        RECT -13.765 62.395 -13.435 62.725 ;
        RECT -13.765 61.035 -13.435 61.365 ;
        RECT -13.765 59.675 -13.435 60.005 ;
        RECT -13.765 58.315 -13.435 58.645 ;
        RECT -13.765 56.955 -13.435 57.285 ;
        RECT -13.765 55.595 -13.435 55.925 ;
        RECT -13.765 54.235 -13.435 54.565 ;
        RECT -13.765 52.875 -13.435 53.205 ;
        RECT -13.765 51.515 -13.435 51.845 ;
        RECT -13.765 50.155 -13.435 50.485 ;
        RECT -13.765 48.795 -13.435 49.125 ;
        RECT -13.765 47.435 -13.435 47.765 ;
        RECT -13.765 46.075 -13.435 46.405 ;
        RECT -13.765 44.715 -13.435 45.045 ;
        RECT -13.765 43.355 -13.435 43.685 ;
        RECT -13.765 41.995 -13.435 42.325 ;
        RECT -13.765 40.635 -13.435 40.965 ;
        RECT -13.765 39.275 -13.435 39.605 ;
        RECT -13.765 37.915 -13.435 38.245 ;
        RECT -13.765 36.555 -13.435 36.885 ;
        RECT -13.765 35.195 -13.435 35.525 ;
        RECT -13.765 33.835 -13.435 34.165 ;
        RECT -13.765 32.475 -13.435 32.805 ;
        RECT -13.765 31.115 -13.435 31.445 ;
        RECT -13.765 29.755 -13.435 30.085 ;
        RECT -13.765 28.395 -13.435 28.725 ;
        RECT -13.765 27.035 -13.435 27.365 ;
        RECT -13.765 25.675 -13.435 26.005 ;
        RECT -13.765 24.315 -13.435 24.645 ;
        RECT -13.765 22.955 -13.435 23.285 ;
        RECT -13.765 21.595 -13.435 21.925 ;
        RECT -13.765 20.235 -13.435 20.565 ;
        RECT -13.765 18.875 -13.435 19.205 ;
        RECT -13.765 17.515 -13.435 17.845 ;
        RECT -13.765 16.155 -13.435 16.485 ;
        RECT -13.765 14.795 -13.435 15.125 ;
        RECT -13.765 13.435 -13.435 13.765 ;
        RECT -13.765 12.075 -13.435 12.405 ;
        RECT -13.765 10.715 -13.435 11.045 ;
        RECT -13.765 9.355 -13.435 9.685 ;
        RECT -13.765 7.995 -13.435 8.325 ;
        RECT -13.765 6.635 -13.435 6.965 ;
        RECT -13.765 5.275 -13.435 5.605 ;
        RECT -13.765 3.915 -13.435 4.245 ;
        RECT -13.765 2.555 -13.435 2.885 ;
        RECT -13.765 1.195 -13.435 1.525 ;
        RECT -13.765 -0.165 -13.435 0.165 ;
        RECT -13.765 -1.525 -13.435 -1.195 ;
        RECT -13.765 -2.885 -13.435 -2.555 ;
        RECT -13.765 -4.245 -13.435 -3.915 ;
        RECT -13.765 -6.965 -13.435 -6.635 ;
        RECT -13.765 -9.685 -13.435 -9.355 ;
        RECT -13.765 -12.41 -13.435 -12.08 ;
        RECT -13.765 -15.125 -13.435 -14.795 ;
        RECT -13.765 -16.485 -13.435 -16.155 ;
        RECT -13.765 -17.25 -13.435 -16.92 ;
        RECT -13.765 -19.205 -13.435 -18.875 ;
        RECT -13.765 -24.645 -13.435 -24.315 ;
        RECT -13.765 -26.005 -13.435 -25.675 ;
        RECT -13.765 -27.365 -13.435 -27.035 ;
        RECT -13.765 -28.725 -13.435 -28.395 ;
        RECT -13.765 -30.085 -13.435 -29.755 ;
        RECT -13.765 -34.165 -13.435 -33.835 ;
        RECT -13.765 -35.39 -13.435 -35.06 ;
        RECT -13.765 -38.245 -13.435 -37.915 ;
        RECT -13.765 -40.23 -13.435 -39.9 ;
        RECT -13.765 -40.965 -13.435 -40.635 ;
        RECT -13.765 -47.765 -13.435 -47.435 ;
        RECT -13.765 -49.125 -13.435 -48.795 ;
        RECT -13.765 -50.485 -13.435 -50.155 ;
        RECT -13.765 -51.845 -13.435 -51.515 ;
        RECT -13.765 -54.565 -13.435 -54.235 ;
        RECT -13.765 -56.27 -13.435 -55.94 ;
        RECT -13.765 -57.285 -13.435 -56.955 ;
        RECT -13.765 -58.645 -13.435 -58.315 ;
        RECT -13.765 -61.365 -13.435 -61.035 ;
        RECT -13.765 -62.725 -13.435 -62.395 ;
        RECT -13.765 -64.085 -13.435 -63.755 ;
        RECT -13.765 -64.81 -13.435 -64.48 ;
        RECT -13.765 -66.805 -13.435 -66.475 ;
        RECT -13.765 -69.525 -13.435 -69.195 ;
        RECT -13.765 -70.885 -13.435 -70.555 ;
        RECT -13.765 -72.245 -13.435 -71.915 ;
        RECT -13.765 -73.605 -13.435 -73.275 ;
        RECT -13.765 -76.325 -13.435 -75.995 ;
        RECT -13.765 -77.685 -13.435 -77.355 ;
        RECT -13.765 -78.45 -13.435 -78.12 ;
        RECT -13.765 -80.405 -13.435 -80.075 ;
        RECT -13.765 -81.765 -13.435 -81.435 ;
        RECT -13.765 -84.485 -13.435 -84.155 ;
        RECT -13.765 -85.845 -13.435 -85.515 ;
        RECT -13.765 -86.99 -13.435 -86.66 ;
        RECT -13.76 -88.56 -13.44 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 -92.645 -13.435 -92.315 ;
        RECT -13.765 -94.005 -13.435 -93.675 ;
        RECT -13.765 -95.365 -13.435 -95.035 ;
        RECT -13.765 -96.725 -13.435 -96.395 ;
        RECT -13.765 -98.085 -13.435 -97.755 ;
        RECT -13.765 -99.445 -13.435 -99.115 ;
        RECT -13.765 -100.805 -13.435 -100.475 ;
        RECT -13.765 -108.965 -13.435 -108.635 ;
        RECT -13.765 -113.045 -13.435 -112.715 ;
        RECT -13.765 -115.765 -13.435 -115.435 ;
        RECT -13.765 -118.485 -13.435 -118.155 ;
        RECT -13.765 -121.205 -13.435 -120.875 ;
        RECT -13.765 -125.285 -13.435 -124.955 ;
        RECT -13.765 -126.645 -13.435 -126.315 ;
        RECT -13.765 -129.365 -13.435 -129.035 ;
        RECT -13.765 -133.445 -13.435 -133.115 ;
        RECT -13.765 -136.165 -13.435 -135.835 ;
        RECT -13.765 -137.525 -13.435 -137.195 ;
        RECT -13.765 -138.885 -13.435 -138.555 ;
        RECT -13.765 -140.245 -13.435 -139.915 ;
        RECT -13.765 -141.605 -13.435 -141.275 ;
        RECT -13.765 -142.965 -13.435 -142.635 ;
        RECT -13.765 -144.325 -13.435 -143.995 ;
        RECT -13.765 -145.685 -13.435 -145.355 ;
        RECT -13.765 -149.765 -13.435 -149.435 ;
        RECT -13.765 -152.485 -13.435 -152.155 ;
        RECT -13.765 -153.845 -13.435 -153.515 ;
        RECT -13.765 -155.285 -13.435 -154.955 ;
        RECT -13.765 -156.565 -13.435 -156.235 ;
        RECT -13.765 -157.925 -13.435 -157.595 ;
        RECT -13.765 -160.17 -13.435 -159.04 ;
        RECT -13.76 -160.285 -13.44 -92.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 73.275 -12.075 73.605 ;
        RECT -12.405 71.915 -12.075 72.245 ;
        RECT -12.405 70.555 -12.075 70.885 ;
        RECT -12.405 69.195 -12.075 69.525 ;
        RECT -12.405 67.835 -12.075 68.165 ;
        RECT -12.405 66.475 -12.075 66.805 ;
        RECT -12.405 65.115 -12.075 65.445 ;
        RECT -12.405 63.755 -12.075 64.085 ;
        RECT -12.405 62.395 -12.075 62.725 ;
        RECT -12.405 61.035 -12.075 61.365 ;
        RECT -12.405 59.675 -12.075 60.005 ;
        RECT -12.405 58.315 -12.075 58.645 ;
        RECT -12.405 56.955 -12.075 57.285 ;
        RECT -12.405 55.595 -12.075 55.925 ;
        RECT -12.405 54.235 -12.075 54.565 ;
        RECT -12.405 52.875 -12.075 53.205 ;
        RECT -12.405 51.515 -12.075 51.845 ;
        RECT -12.405 50.155 -12.075 50.485 ;
        RECT -12.405 48.795 -12.075 49.125 ;
        RECT -12.405 47.435 -12.075 47.765 ;
        RECT -12.405 46.075 -12.075 46.405 ;
        RECT -12.405 44.715 -12.075 45.045 ;
        RECT -12.405 43.355 -12.075 43.685 ;
        RECT -12.405 41.995 -12.075 42.325 ;
        RECT -12.405 40.635 -12.075 40.965 ;
        RECT -12.405 39.275 -12.075 39.605 ;
        RECT -12.405 37.915 -12.075 38.245 ;
        RECT -12.405 36.555 -12.075 36.885 ;
        RECT -12.405 35.195 -12.075 35.525 ;
        RECT -12.405 33.835 -12.075 34.165 ;
        RECT -12.405 32.475 -12.075 32.805 ;
        RECT -12.405 31.115 -12.075 31.445 ;
        RECT -12.405 29.755 -12.075 30.085 ;
        RECT -12.405 28.395 -12.075 28.725 ;
        RECT -12.405 27.035 -12.075 27.365 ;
        RECT -12.405 25.675 -12.075 26.005 ;
        RECT -12.405 24.315 -12.075 24.645 ;
        RECT -12.405 22.955 -12.075 23.285 ;
        RECT -12.405 21.595 -12.075 21.925 ;
        RECT -12.405 20.235 -12.075 20.565 ;
        RECT -12.405 18.875 -12.075 19.205 ;
        RECT -12.405 17.515 -12.075 17.845 ;
        RECT -12.405 16.155 -12.075 16.485 ;
        RECT -12.405 14.795 -12.075 15.125 ;
        RECT -12.405 13.435 -12.075 13.765 ;
        RECT -12.405 12.075 -12.075 12.405 ;
        RECT -12.405 10.715 -12.075 11.045 ;
        RECT -12.405 9.355 -12.075 9.685 ;
        RECT -12.405 7.995 -12.075 8.325 ;
        RECT -12.405 6.635 -12.075 6.965 ;
        RECT -12.405 5.275 -12.075 5.605 ;
        RECT -12.405 3.915 -12.075 4.245 ;
        RECT -12.405 2.555 -12.075 2.885 ;
        RECT -12.405 1.195 -12.075 1.525 ;
        RECT -12.405 -0.165 -12.075 0.165 ;
        RECT -12.405 -1.525 -12.075 -1.195 ;
        RECT -12.405 -2.885 -12.075 -2.555 ;
        RECT -12.405 -4.245 -12.075 -3.915 ;
        RECT -12.405 -6.965 -12.075 -6.635 ;
        RECT -12.405 -9.685 -12.075 -9.355 ;
        RECT -12.4 -9.685 -12.08 128.47 ;
        RECT -12.405 127.225 -12.075 128.355 ;
        RECT -12.405 124.955 -12.075 125.285 ;
        RECT -12.405 123.595 -12.075 123.925 ;
        RECT -12.405 122.235 -12.075 122.565 ;
        RECT -12.405 120.875 -12.075 121.205 ;
        RECT -12.405 119.515 -12.075 119.845 ;
        RECT -12.405 118.155 -12.075 118.485 ;
        RECT -12.405 116.795 -12.075 117.125 ;
        RECT -12.405 115.435 -12.075 115.765 ;
        RECT -12.405 114.075 -12.075 114.405 ;
        RECT -12.405 112.715 -12.075 113.045 ;
        RECT -12.405 111.355 -12.075 111.685 ;
        RECT -12.405 109.995 -12.075 110.325 ;
        RECT -12.405 108.635 -12.075 108.965 ;
        RECT -12.405 107.275 -12.075 107.605 ;
        RECT -12.405 105.915 -12.075 106.245 ;
        RECT -12.405 104.555 -12.075 104.885 ;
        RECT -12.405 103.195 -12.075 103.525 ;
        RECT -12.405 101.835 -12.075 102.165 ;
        RECT -12.405 100.475 -12.075 100.805 ;
        RECT -12.405 99.115 -12.075 99.445 ;
        RECT -12.405 97.755 -12.075 98.085 ;
        RECT -12.405 96.395 -12.075 96.725 ;
        RECT -12.405 95.035 -12.075 95.365 ;
        RECT -12.405 93.675 -12.075 94.005 ;
        RECT -12.405 92.315 -12.075 92.645 ;
        RECT -12.405 90.955 -12.075 91.285 ;
        RECT -12.405 89.595 -12.075 89.925 ;
        RECT -12.405 88.235 -12.075 88.565 ;
        RECT -12.405 86.875 -12.075 87.205 ;
        RECT -12.405 85.515 -12.075 85.845 ;
        RECT -12.405 84.155 -12.075 84.485 ;
        RECT -12.405 82.795 -12.075 83.125 ;
        RECT -12.405 81.435 -12.075 81.765 ;
        RECT -12.405 80.075 -12.075 80.405 ;
        RECT -12.405 78.715 -12.075 79.045 ;
        RECT -12.405 77.355 -12.075 77.685 ;
        RECT -12.405 75.995 -12.075 76.325 ;
        RECT -12.405 74.635 -12.075 74.965 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 127.225 -28.395 128.355 ;
        RECT -28.725 124.955 -28.395 125.285 ;
        RECT -28.725 123.595 -28.395 123.925 ;
        RECT -28.725 122.235 -28.395 122.565 ;
        RECT -28.725 120.875 -28.395 121.205 ;
        RECT -28.725 119.515 -28.395 119.845 ;
        RECT -28.725 118.155 -28.395 118.485 ;
        RECT -28.725 116.795 -28.395 117.125 ;
        RECT -28.725 115.435 -28.395 115.765 ;
        RECT -28.725 114.075 -28.395 114.405 ;
        RECT -28.725 112.715 -28.395 113.045 ;
        RECT -28.725 111.355 -28.395 111.685 ;
        RECT -28.725 109.995 -28.395 110.325 ;
        RECT -28.725 108.635 -28.395 108.965 ;
        RECT -28.725 107.275 -28.395 107.605 ;
        RECT -28.725 105.915 -28.395 106.245 ;
        RECT -28.725 104.555 -28.395 104.885 ;
        RECT -28.725 103.195 -28.395 103.525 ;
        RECT -28.725 101.835 -28.395 102.165 ;
        RECT -28.725 100.475 -28.395 100.805 ;
        RECT -28.725 99.115 -28.395 99.445 ;
        RECT -28.725 97.755 -28.395 98.085 ;
        RECT -28.725 96.395 -28.395 96.725 ;
        RECT -28.725 95.035 -28.395 95.365 ;
        RECT -28.725 93.675 -28.395 94.005 ;
        RECT -28.725 92.315 -28.395 92.645 ;
        RECT -28.725 90.955 -28.395 91.285 ;
        RECT -28.725 89.595 -28.395 89.925 ;
        RECT -28.725 88.235 -28.395 88.565 ;
        RECT -28.725 86.875 -28.395 87.205 ;
        RECT -28.725 85.515 -28.395 85.845 ;
        RECT -28.725 84.155 -28.395 84.485 ;
        RECT -28.725 82.795 -28.395 83.125 ;
        RECT -28.725 81.435 -28.395 81.765 ;
        RECT -28.725 80.075 -28.395 80.405 ;
        RECT -28.725 78.715 -28.395 79.045 ;
        RECT -28.725 77.355 -28.395 77.685 ;
        RECT -28.725 75.995 -28.395 76.325 ;
        RECT -28.725 74.635 -28.395 74.965 ;
        RECT -28.725 73.275 -28.395 73.605 ;
        RECT -28.725 71.915 -28.395 72.245 ;
        RECT -28.725 70.555 -28.395 70.885 ;
        RECT -28.725 69.195 -28.395 69.525 ;
        RECT -28.725 67.835 -28.395 68.165 ;
        RECT -28.725 66.475 -28.395 66.805 ;
        RECT -28.725 65.115 -28.395 65.445 ;
        RECT -28.725 63.755 -28.395 64.085 ;
        RECT -28.725 62.395 -28.395 62.725 ;
        RECT -28.725 61.035 -28.395 61.365 ;
        RECT -28.725 59.675 -28.395 60.005 ;
        RECT -28.725 58.315 -28.395 58.645 ;
        RECT -28.725 56.955 -28.395 57.285 ;
        RECT -28.725 55.595 -28.395 55.925 ;
        RECT -28.725 54.235 -28.395 54.565 ;
        RECT -28.725 52.875 -28.395 53.205 ;
        RECT -28.725 51.515 -28.395 51.845 ;
        RECT -28.725 50.155 -28.395 50.485 ;
        RECT -28.725 48.795 -28.395 49.125 ;
        RECT -28.725 47.435 -28.395 47.765 ;
        RECT -28.725 46.075 -28.395 46.405 ;
        RECT -28.725 44.715 -28.395 45.045 ;
        RECT -28.725 43.355 -28.395 43.685 ;
        RECT -28.725 41.995 -28.395 42.325 ;
        RECT -28.725 40.635 -28.395 40.965 ;
        RECT -28.725 39.275 -28.395 39.605 ;
        RECT -28.725 37.915 -28.395 38.245 ;
        RECT -28.725 36.555 -28.395 36.885 ;
        RECT -28.725 35.195 -28.395 35.525 ;
        RECT -28.725 33.835 -28.395 34.165 ;
        RECT -28.725 32.475 -28.395 32.805 ;
        RECT -28.725 31.115 -28.395 31.445 ;
        RECT -28.725 29.755 -28.395 30.085 ;
        RECT -28.725 28.395 -28.395 28.725 ;
        RECT -28.725 27.035 -28.395 27.365 ;
        RECT -28.725 25.675 -28.395 26.005 ;
        RECT -28.725 24.315 -28.395 24.645 ;
        RECT -28.725 22.955 -28.395 23.285 ;
        RECT -28.725 21.595 -28.395 21.925 ;
        RECT -28.725 20.235 -28.395 20.565 ;
        RECT -28.725 18.875 -28.395 19.205 ;
        RECT -28.725 17.515 -28.395 17.845 ;
        RECT -28.725 16.155 -28.395 16.485 ;
        RECT -28.725 14.795 -28.395 15.125 ;
        RECT -28.725 13.435 -28.395 13.765 ;
        RECT -28.725 12.075 -28.395 12.405 ;
        RECT -28.725 10.715 -28.395 11.045 ;
        RECT -28.725 9.355 -28.395 9.685 ;
        RECT -28.725 7.995 -28.395 8.325 ;
        RECT -28.725 6.635 -28.395 6.965 ;
        RECT -28.725 5.275 -28.395 5.605 ;
        RECT -28.725 3.915 -28.395 4.245 ;
        RECT -28.725 2.555 -28.395 2.885 ;
        RECT -28.725 1.195 -28.395 1.525 ;
        RECT -28.725 -0.165 -28.395 0.165 ;
        RECT -28.725 -12.41 -28.395 -12.08 ;
        RECT -28.725 -15.125 -28.395 -14.795 ;
        RECT -28.725 -16.485 -28.395 -16.155 ;
        RECT -28.725 -17.25 -28.395 -16.92 ;
        RECT -28.725 -19.205 -28.395 -18.875 ;
        RECT -28.725 -28.725 -28.395 -28.395 ;
        RECT -28.725 -30.085 -28.395 -29.755 ;
        RECT -28.725 -32.805 -28.395 -32.475 ;
        RECT -28.725 -34.165 -28.395 -33.835 ;
        RECT -28.725 -35.39 -28.395 -35.06 ;
        RECT -28.725 -38.245 -28.395 -37.915 ;
        RECT -28.725 -40.23 -28.395 -39.9 ;
        RECT -28.725 -40.965 -28.395 -40.635 ;
        RECT -28.725 -50.485 -28.395 -50.155 ;
        RECT -28.725 -51.845 -28.395 -51.515 ;
        RECT -28.725 -53.205 -28.395 -52.875 ;
        RECT -28.725 -54.565 -28.395 -54.235 ;
        RECT -28.725 -55.925 -28.395 -55.595 ;
        RECT -28.725 -57.285 -28.395 -56.955 ;
        RECT -28.725 -58.645 -28.395 -58.315 ;
        RECT -28.725 -60.005 -28.395 -59.675 ;
        RECT -28.725 -61.365 -28.395 -61.035 ;
        RECT -28.725 -62.725 -28.395 -62.395 ;
        RECT -28.725 -64.085 -28.395 -63.755 ;
        RECT -28.725 -65.445 -28.395 -65.115 ;
        RECT -28.725 -66.805 -28.395 -66.475 ;
        RECT -28.725 -68.165 -28.395 -67.835 ;
        RECT -28.725 -69.525 -28.395 -69.195 ;
        RECT -28.725 -72.245 -28.395 -71.915 ;
        RECT -28.725 -73.605 -28.395 -73.275 ;
        RECT -28.725 -74.965 -28.395 -74.635 ;
        RECT -28.725 -76.325 -28.395 -75.995 ;
        RECT -28.725 -78.29 -28.395 -77.96 ;
        RECT -28.725 -79.045 -28.395 -78.715 ;
        RECT -28.725 -81.765 -28.395 -81.435 ;
        RECT -28.725 -83.125 -28.395 -82.795 ;
        RECT -28.725 -84.485 -28.395 -84.155 ;
        RECT -28.725 -86.43 -28.395 -86.1 ;
        RECT -28.725 -87.205 -28.395 -86.875 ;
        RECT -28.725 -88.565 -28.395 -88.235 ;
        RECT -28.725 -89.925 -28.395 -89.595 ;
        RECT -28.72 -91.28 -28.4 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 -153.845 -28.395 -153.515 ;
        RECT -28.725 -156.565 -28.395 -156.235 ;
        RECT -28.725 -157.925 -28.395 -157.595 ;
        RECT -28.725 -160.17 -28.395 -159.04 ;
        RECT -28.72 -160.285 -28.4 -152.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.365 127.225 -27.035 128.355 ;
        RECT -27.365 124.955 -27.035 125.285 ;
        RECT -27.365 123.595 -27.035 123.925 ;
        RECT -27.365 122.235 -27.035 122.565 ;
        RECT -27.365 120.875 -27.035 121.205 ;
        RECT -27.365 119.515 -27.035 119.845 ;
        RECT -27.365 118.155 -27.035 118.485 ;
        RECT -27.365 116.795 -27.035 117.125 ;
        RECT -27.365 115.435 -27.035 115.765 ;
        RECT -27.365 114.075 -27.035 114.405 ;
        RECT -27.365 112.715 -27.035 113.045 ;
        RECT -27.365 111.355 -27.035 111.685 ;
        RECT -27.365 109.995 -27.035 110.325 ;
        RECT -27.365 108.635 -27.035 108.965 ;
        RECT -27.365 107.275 -27.035 107.605 ;
        RECT -27.365 105.915 -27.035 106.245 ;
        RECT -27.365 104.555 -27.035 104.885 ;
        RECT -27.365 103.195 -27.035 103.525 ;
        RECT -27.365 101.835 -27.035 102.165 ;
        RECT -27.365 100.475 -27.035 100.805 ;
        RECT -27.365 99.115 -27.035 99.445 ;
        RECT -27.365 97.755 -27.035 98.085 ;
        RECT -27.365 96.395 -27.035 96.725 ;
        RECT -27.365 95.035 -27.035 95.365 ;
        RECT -27.365 93.675 -27.035 94.005 ;
        RECT -27.365 92.315 -27.035 92.645 ;
        RECT -27.365 90.955 -27.035 91.285 ;
        RECT -27.365 89.595 -27.035 89.925 ;
        RECT -27.365 88.235 -27.035 88.565 ;
        RECT -27.365 86.875 -27.035 87.205 ;
        RECT -27.365 85.515 -27.035 85.845 ;
        RECT -27.365 84.155 -27.035 84.485 ;
        RECT -27.365 82.795 -27.035 83.125 ;
        RECT -27.365 81.435 -27.035 81.765 ;
        RECT -27.365 80.075 -27.035 80.405 ;
        RECT -27.365 78.715 -27.035 79.045 ;
        RECT -27.365 77.355 -27.035 77.685 ;
        RECT -27.365 75.995 -27.035 76.325 ;
        RECT -27.365 74.635 -27.035 74.965 ;
        RECT -27.365 73.275 -27.035 73.605 ;
        RECT -27.365 71.915 -27.035 72.245 ;
        RECT -27.365 70.555 -27.035 70.885 ;
        RECT -27.365 69.195 -27.035 69.525 ;
        RECT -27.365 67.835 -27.035 68.165 ;
        RECT -27.365 66.475 -27.035 66.805 ;
        RECT -27.365 65.115 -27.035 65.445 ;
        RECT -27.365 63.755 -27.035 64.085 ;
        RECT -27.365 62.395 -27.035 62.725 ;
        RECT -27.365 61.035 -27.035 61.365 ;
        RECT -27.365 59.675 -27.035 60.005 ;
        RECT -27.365 58.315 -27.035 58.645 ;
        RECT -27.365 56.955 -27.035 57.285 ;
        RECT -27.365 55.595 -27.035 55.925 ;
        RECT -27.365 54.235 -27.035 54.565 ;
        RECT -27.365 52.875 -27.035 53.205 ;
        RECT -27.365 51.515 -27.035 51.845 ;
        RECT -27.365 50.155 -27.035 50.485 ;
        RECT -27.365 48.795 -27.035 49.125 ;
        RECT -27.365 47.435 -27.035 47.765 ;
        RECT -27.365 46.075 -27.035 46.405 ;
        RECT -27.365 44.715 -27.035 45.045 ;
        RECT -27.365 43.355 -27.035 43.685 ;
        RECT -27.365 41.995 -27.035 42.325 ;
        RECT -27.365 40.635 -27.035 40.965 ;
        RECT -27.365 39.275 -27.035 39.605 ;
        RECT -27.365 37.915 -27.035 38.245 ;
        RECT -27.365 36.555 -27.035 36.885 ;
        RECT -27.365 35.195 -27.035 35.525 ;
        RECT -27.365 33.835 -27.035 34.165 ;
        RECT -27.365 32.475 -27.035 32.805 ;
        RECT -27.365 31.115 -27.035 31.445 ;
        RECT -27.365 29.755 -27.035 30.085 ;
        RECT -27.365 28.395 -27.035 28.725 ;
        RECT -27.365 27.035 -27.035 27.365 ;
        RECT -27.365 25.675 -27.035 26.005 ;
        RECT -27.365 24.315 -27.035 24.645 ;
        RECT -27.365 22.955 -27.035 23.285 ;
        RECT -27.365 21.595 -27.035 21.925 ;
        RECT -27.365 20.235 -27.035 20.565 ;
        RECT -27.365 18.875 -27.035 19.205 ;
        RECT -27.365 17.515 -27.035 17.845 ;
        RECT -27.365 16.155 -27.035 16.485 ;
        RECT -27.365 14.795 -27.035 15.125 ;
        RECT -27.365 13.435 -27.035 13.765 ;
        RECT -27.365 12.075 -27.035 12.405 ;
        RECT -27.365 10.715 -27.035 11.045 ;
        RECT -27.365 9.355 -27.035 9.685 ;
        RECT -27.365 7.995 -27.035 8.325 ;
        RECT -27.365 6.635 -27.035 6.965 ;
        RECT -27.365 5.275 -27.035 5.605 ;
        RECT -27.365 3.915 -27.035 4.245 ;
        RECT -27.365 2.555 -27.035 2.885 ;
        RECT -27.365 1.195 -27.035 1.525 ;
        RECT -27.365 -0.165 -27.035 0.165 ;
        RECT -27.365 -12.41 -27.035 -12.08 ;
        RECT -27.365 -15.125 -27.035 -14.795 ;
        RECT -27.365 -16.485 -27.035 -16.155 ;
        RECT -27.365 -17.25 -27.035 -16.92 ;
        RECT -27.365 -19.205 -27.035 -18.875 ;
        RECT -27.365 -28.725 -27.035 -28.395 ;
        RECT -27.365 -30.085 -27.035 -29.755 ;
        RECT -27.365 -32.805 -27.035 -32.475 ;
        RECT -27.365 -34.165 -27.035 -33.835 ;
        RECT -27.365 -35.39 -27.035 -35.06 ;
        RECT -27.365 -38.245 -27.035 -37.915 ;
        RECT -27.365 -40.23 -27.035 -39.9 ;
        RECT -27.365 -40.965 -27.035 -40.635 ;
        RECT -27.365 -50.485 -27.035 -50.155 ;
        RECT -27.365 -51.845 -27.035 -51.515 ;
        RECT -27.365 -53.205 -27.035 -52.875 ;
        RECT -27.365 -54.565 -27.035 -54.235 ;
        RECT -27.365 -55.925 -27.035 -55.595 ;
        RECT -27.365 -57.285 -27.035 -56.955 ;
        RECT -27.365 -58.645 -27.035 -58.315 ;
        RECT -27.365 -60.005 -27.035 -59.675 ;
        RECT -27.365 -61.365 -27.035 -61.035 ;
        RECT -27.365 -62.725 -27.035 -62.395 ;
        RECT -27.365 -64.085 -27.035 -63.755 ;
        RECT -27.365 -65.445 -27.035 -65.115 ;
        RECT -27.365 -66.805 -27.035 -66.475 ;
        RECT -27.365 -68.165 -27.035 -67.835 ;
        RECT -27.365 -69.525 -27.035 -69.195 ;
        RECT -27.365 -72.245 -27.035 -71.915 ;
        RECT -27.365 -73.605 -27.035 -73.275 ;
        RECT -27.365 -74.965 -27.035 -74.635 ;
        RECT -27.365 -76.325 -27.035 -75.995 ;
        RECT -27.365 -78.29 -27.035 -77.96 ;
        RECT -27.365 -79.045 -27.035 -78.715 ;
        RECT -27.365 -81.765 -27.035 -81.435 ;
        RECT -27.365 -83.125 -27.035 -82.795 ;
        RECT -27.365 -84.485 -27.035 -84.155 ;
        RECT -27.365 -86.43 -27.035 -86.1 ;
        RECT -27.365 -87.205 -27.035 -86.875 ;
        RECT -27.365 -88.565 -27.035 -88.235 ;
        RECT -27.365 -89.925 -27.035 -89.595 ;
        RECT -27.365 -92.645 -27.035 -92.315 ;
        RECT -27.365 -94.005 -27.035 -93.675 ;
        RECT -27.365 -95.365 -27.035 -95.035 ;
        RECT -27.365 -96.725 -27.035 -96.395 ;
        RECT -27.365 -98.085 -27.035 -97.755 ;
        RECT -27.365 -102.165 -27.035 -101.835 ;
        RECT -27.365 -104.885 -27.035 -104.555 ;
        RECT -27.365 -106.245 -27.035 -105.915 ;
        RECT -27.365 -107.605 -27.035 -107.275 ;
        RECT -27.365 -108.965 -27.035 -108.635 ;
        RECT -27.365 -113.045 -27.035 -112.715 ;
        RECT -27.365 -114.405 -27.035 -114.075 ;
        RECT -27.365 -115.765 -27.035 -115.435 ;
        RECT -27.365 -118.485 -27.035 -118.155 ;
        RECT -27.365 -121.205 -27.035 -120.875 ;
        RECT -27.365 -122.565 -27.035 -122.235 ;
        RECT -27.365 -123.925 -27.035 -123.595 ;
        RECT -27.365 -125.285 -27.035 -124.955 ;
        RECT -27.365 -126.645 -27.035 -126.315 ;
        RECT -27.365 -128.005 -27.035 -127.675 ;
        RECT -27.365 -130.725 -27.035 -130.395 ;
        RECT -27.365 -132.085 -27.035 -131.755 ;
        RECT -27.365 -136.165 -27.035 -135.835 ;
        RECT -27.365 -137.525 -27.035 -137.195 ;
        RECT -27.365 -138.885 -27.035 -138.555 ;
        RECT -27.365 -140.245 -27.035 -139.915 ;
        RECT -27.365 -141.605 -27.035 -141.275 ;
        RECT -27.365 -142.965 -27.035 -142.635 ;
        RECT -27.365 -144.325 -27.035 -143.995 ;
        RECT -27.365 -145.685 -27.035 -145.355 ;
        RECT -27.365 -147.045 -27.035 -146.715 ;
        RECT -27.365 -149.765 -27.035 -149.435 ;
        RECT -27.36 -151.8 -27.04 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.005 127.225 -25.675 128.355 ;
        RECT -26.005 124.955 -25.675 125.285 ;
        RECT -26.005 123.595 -25.675 123.925 ;
        RECT -26.005 122.235 -25.675 122.565 ;
        RECT -26.005 120.875 -25.675 121.205 ;
        RECT -26.005 119.515 -25.675 119.845 ;
        RECT -26.005 118.155 -25.675 118.485 ;
        RECT -26.005 116.795 -25.675 117.125 ;
        RECT -26.005 115.435 -25.675 115.765 ;
        RECT -26.005 114.075 -25.675 114.405 ;
        RECT -26.005 112.715 -25.675 113.045 ;
        RECT -26.005 111.355 -25.675 111.685 ;
        RECT -26.005 109.995 -25.675 110.325 ;
        RECT -26.005 108.635 -25.675 108.965 ;
        RECT -26.005 107.275 -25.675 107.605 ;
        RECT -26.005 105.915 -25.675 106.245 ;
        RECT -26.005 104.555 -25.675 104.885 ;
        RECT -26.005 103.195 -25.675 103.525 ;
        RECT -26.005 101.835 -25.675 102.165 ;
        RECT -26.005 100.475 -25.675 100.805 ;
        RECT -26.005 99.115 -25.675 99.445 ;
        RECT -26.005 97.755 -25.675 98.085 ;
        RECT -26.005 96.395 -25.675 96.725 ;
        RECT -26.005 95.035 -25.675 95.365 ;
        RECT -26.005 93.675 -25.675 94.005 ;
        RECT -26.005 92.315 -25.675 92.645 ;
        RECT -26.005 90.955 -25.675 91.285 ;
        RECT -26.005 89.595 -25.675 89.925 ;
        RECT -26.005 88.235 -25.675 88.565 ;
        RECT -26.005 86.875 -25.675 87.205 ;
        RECT -26.005 85.515 -25.675 85.845 ;
        RECT -26.005 84.155 -25.675 84.485 ;
        RECT -26.005 82.795 -25.675 83.125 ;
        RECT -26.005 81.435 -25.675 81.765 ;
        RECT -26.005 80.075 -25.675 80.405 ;
        RECT -26.005 78.715 -25.675 79.045 ;
        RECT -26.005 77.355 -25.675 77.685 ;
        RECT -26.005 75.995 -25.675 76.325 ;
        RECT -26.005 74.635 -25.675 74.965 ;
        RECT -26.005 73.275 -25.675 73.605 ;
        RECT -26.005 71.915 -25.675 72.245 ;
        RECT -26.005 70.555 -25.675 70.885 ;
        RECT -26.005 69.195 -25.675 69.525 ;
        RECT -26.005 67.835 -25.675 68.165 ;
        RECT -26.005 66.475 -25.675 66.805 ;
        RECT -26.005 65.115 -25.675 65.445 ;
        RECT -26.005 63.755 -25.675 64.085 ;
        RECT -26.005 62.395 -25.675 62.725 ;
        RECT -26.005 61.035 -25.675 61.365 ;
        RECT -26.005 59.675 -25.675 60.005 ;
        RECT -26.005 58.315 -25.675 58.645 ;
        RECT -26.005 56.955 -25.675 57.285 ;
        RECT -26.005 55.595 -25.675 55.925 ;
        RECT -26.005 54.235 -25.675 54.565 ;
        RECT -26.005 52.875 -25.675 53.205 ;
        RECT -26.005 51.515 -25.675 51.845 ;
        RECT -26.005 50.155 -25.675 50.485 ;
        RECT -26.005 48.795 -25.675 49.125 ;
        RECT -26.005 47.435 -25.675 47.765 ;
        RECT -26.005 46.075 -25.675 46.405 ;
        RECT -26.005 44.715 -25.675 45.045 ;
        RECT -26.005 43.355 -25.675 43.685 ;
        RECT -26.005 41.995 -25.675 42.325 ;
        RECT -26.005 40.635 -25.675 40.965 ;
        RECT -26.005 39.275 -25.675 39.605 ;
        RECT -26.005 37.915 -25.675 38.245 ;
        RECT -26.005 36.555 -25.675 36.885 ;
        RECT -26.005 35.195 -25.675 35.525 ;
        RECT -26.005 33.835 -25.675 34.165 ;
        RECT -26.005 32.475 -25.675 32.805 ;
        RECT -26.005 31.115 -25.675 31.445 ;
        RECT -26.005 29.755 -25.675 30.085 ;
        RECT -26.005 28.395 -25.675 28.725 ;
        RECT -26.005 27.035 -25.675 27.365 ;
        RECT -26.005 25.675 -25.675 26.005 ;
        RECT -26.005 24.315 -25.675 24.645 ;
        RECT -26.005 22.955 -25.675 23.285 ;
        RECT -26.005 21.595 -25.675 21.925 ;
        RECT -26.005 20.235 -25.675 20.565 ;
        RECT -26.005 18.875 -25.675 19.205 ;
        RECT -26.005 17.515 -25.675 17.845 ;
        RECT -26.005 16.155 -25.675 16.485 ;
        RECT -26.005 14.795 -25.675 15.125 ;
        RECT -26.005 13.435 -25.675 13.765 ;
        RECT -26.005 12.075 -25.675 12.405 ;
        RECT -26.005 10.715 -25.675 11.045 ;
        RECT -26.005 9.355 -25.675 9.685 ;
        RECT -26.005 7.995 -25.675 8.325 ;
        RECT -26.005 6.635 -25.675 6.965 ;
        RECT -26.005 5.275 -25.675 5.605 ;
        RECT -26.005 3.915 -25.675 4.245 ;
        RECT -26.005 2.555 -25.675 2.885 ;
        RECT -26.005 1.195 -25.675 1.525 ;
        RECT -26.005 -0.165 -25.675 0.165 ;
        RECT -26.005 -1.525 -25.675 -1.195 ;
        RECT -26.005 -12.41 -25.675 -12.08 ;
        RECT -26.005 -15.125 -25.675 -14.795 ;
        RECT -26.005 -16.485 -25.675 -16.155 ;
        RECT -26.005 -17.25 -25.675 -16.92 ;
        RECT -26.005 -19.205 -25.675 -18.875 ;
        RECT -26.005 -28.725 -25.675 -28.395 ;
        RECT -26.005 -30.085 -25.675 -29.755 ;
        RECT -26.005 -32.805 -25.675 -32.475 ;
        RECT -26.005 -34.165 -25.675 -33.835 ;
        RECT -26.005 -35.39 -25.675 -35.06 ;
        RECT -26.005 -38.245 -25.675 -37.915 ;
        RECT -26.005 -40.23 -25.675 -39.9 ;
        RECT -26.005 -40.965 -25.675 -40.635 ;
        RECT -26.005 -50.485 -25.675 -50.155 ;
        RECT -26.005 -51.845 -25.675 -51.515 ;
        RECT -26.005 -53.205 -25.675 -52.875 ;
        RECT -26.005 -54.565 -25.675 -54.235 ;
        RECT -26.005 -55.925 -25.675 -55.595 ;
        RECT -26.005 -57.285 -25.675 -56.955 ;
        RECT -26.005 -58.645 -25.675 -58.315 ;
        RECT -26.005 -60.005 -25.675 -59.675 ;
        RECT -26.005 -61.365 -25.675 -61.035 ;
        RECT -26.005 -62.725 -25.675 -62.395 ;
        RECT -26.005 -64.085 -25.675 -63.755 ;
        RECT -26.005 -65.445 -25.675 -65.115 ;
        RECT -26.005 -66.805 -25.675 -66.475 ;
        RECT -26.005 -68.165 -25.675 -67.835 ;
        RECT -26.005 -69.525 -25.675 -69.195 ;
        RECT -26.005 -70.885 -25.675 -70.555 ;
        RECT -26.005 -72.245 -25.675 -71.915 ;
        RECT -26.005 -73.605 -25.675 -73.275 ;
        RECT -26.005 -74.965 -25.675 -74.635 ;
        RECT -26.005 -76.325 -25.675 -75.995 ;
        RECT -26.005 -77.685 -25.675 -77.355 ;
        RECT -26.005 -79.045 -25.675 -78.715 ;
        RECT -26.005 -80.405 -25.675 -80.075 ;
        RECT -26.005 -81.765 -25.675 -81.435 ;
        RECT -26.005 -83.125 -25.675 -82.795 ;
        RECT -26.005 -84.485 -25.675 -84.155 ;
        RECT -26.005 -85.845 -25.675 -85.515 ;
        RECT -26.005 -87.205 -25.675 -86.875 ;
        RECT -26.005 -88.565 -25.675 -88.235 ;
        RECT -26.005 -89.925 -25.675 -89.595 ;
        RECT -26.005 -91.285 -25.675 -90.955 ;
        RECT -26.005 -92.645 -25.675 -92.315 ;
        RECT -26.005 -94.005 -25.675 -93.675 ;
        RECT -26.005 -95.365 -25.675 -95.035 ;
        RECT -26.005 -96.725 -25.675 -96.395 ;
        RECT -26.005 -98.085 -25.675 -97.755 ;
        RECT -26.005 -102.165 -25.675 -101.835 ;
        RECT -26.005 -104.885 -25.675 -104.555 ;
        RECT -26.005 -106.245 -25.675 -105.915 ;
        RECT -26.005 -107.605 -25.675 -107.275 ;
        RECT -26.005 -108.965 -25.675 -108.635 ;
        RECT -26.005 -114.405 -25.675 -114.075 ;
        RECT -26.005 -115.765 -25.675 -115.435 ;
        RECT -26.005 -118.485 -25.675 -118.155 ;
        RECT -26.005 -121.205 -25.675 -120.875 ;
        RECT -26.005 -122.565 -25.675 -122.235 ;
        RECT -26.005 -125.285 -25.675 -124.955 ;
        RECT -26.005 -126.645 -25.675 -126.315 ;
        RECT -26.005 -128.005 -25.675 -127.675 ;
        RECT -26.005 -130.725 -25.675 -130.395 ;
        RECT -26.005 -132.085 -25.675 -131.755 ;
        RECT -26.005 -136.165 -25.675 -135.835 ;
        RECT -26.005 -137.525 -25.675 -137.195 ;
        RECT -26.005 -138.885 -25.675 -138.555 ;
        RECT -26.005 -140.245 -25.675 -139.915 ;
        RECT -26.005 -141.605 -25.675 -141.275 ;
        RECT -26.005 -142.965 -25.675 -142.635 ;
        RECT -26.005 -144.325 -25.675 -143.995 ;
        RECT -26.005 -145.685 -25.675 -145.355 ;
        RECT -26.005 -147.045 -25.675 -146.715 ;
        RECT -26.005 -149.765 -25.675 -149.435 ;
        RECT -26.005 -152.485 -25.675 -152.155 ;
        RECT -26.005 -153.845 -25.675 -153.515 ;
        RECT -26.005 -155.285 -25.675 -154.955 ;
        RECT -26.005 -156.565 -25.675 -156.235 ;
        RECT -26.005 -157.925 -25.675 -157.595 ;
        RECT -26.005 -160.17 -25.675 -159.04 ;
        RECT -26 -160.285 -25.68 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.645 127.225 -24.315 128.355 ;
        RECT -24.645 124.955 -24.315 125.285 ;
        RECT -24.645 123.595 -24.315 123.925 ;
        RECT -24.645 122.235 -24.315 122.565 ;
        RECT -24.645 120.875 -24.315 121.205 ;
        RECT -24.645 119.515 -24.315 119.845 ;
        RECT -24.645 118.155 -24.315 118.485 ;
        RECT -24.645 116.795 -24.315 117.125 ;
        RECT -24.645 115.435 -24.315 115.765 ;
        RECT -24.645 114.075 -24.315 114.405 ;
        RECT -24.645 112.715 -24.315 113.045 ;
        RECT -24.645 111.355 -24.315 111.685 ;
        RECT -24.645 109.995 -24.315 110.325 ;
        RECT -24.645 108.635 -24.315 108.965 ;
        RECT -24.645 107.275 -24.315 107.605 ;
        RECT -24.645 105.915 -24.315 106.245 ;
        RECT -24.645 104.555 -24.315 104.885 ;
        RECT -24.645 103.195 -24.315 103.525 ;
        RECT -24.645 101.835 -24.315 102.165 ;
        RECT -24.645 100.475 -24.315 100.805 ;
        RECT -24.645 99.115 -24.315 99.445 ;
        RECT -24.645 97.755 -24.315 98.085 ;
        RECT -24.645 96.395 -24.315 96.725 ;
        RECT -24.645 95.035 -24.315 95.365 ;
        RECT -24.645 93.675 -24.315 94.005 ;
        RECT -24.645 92.315 -24.315 92.645 ;
        RECT -24.645 90.955 -24.315 91.285 ;
        RECT -24.645 89.595 -24.315 89.925 ;
        RECT -24.645 88.235 -24.315 88.565 ;
        RECT -24.645 86.875 -24.315 87.205 ;
        RECT -24.645 85.515 -24.315 85.845 ;
        RECT -24.645 84.155 -24.315 84.485 ;
        RECT -24.645 82.795 -24.315 83.125 ;
        RECT -24.645 81.435 -24.315 81.765 ;
        RECT -24.645 80.075 -24.315 80.405 ;
        RECT -24.645 78.715 -24.315 79.045 ;
        RECT -24.645 77.355 -24.315 77.685 ;
        RECT -24.645 75.995 -24.315 76.325 ;
        RECT -24.645 74.635 -24.315 74.965 ;
        RECT -24.645 73.275 -24.315 73.605 ;
        RECT -24.645 71.915 -24.315 72.245 ;
        RECT -24.645 70.555 -24.315 70.885 ;
        RECT -24.645 69.195 -24.315 69.525 ;
        RECT -24.645 67.835 -24.315 68.165 ;
        RECT -24.645 66.475 -24.315 66.805 ;
        RECT -24.645 65.115 -24.315 65.445 ;
        RECT -24.645 63.755 -24.315 64.085 ;
        RECT -24.645 62.395 -24.315 62.725 ;
        RECT -24.645 61.035 -24.315 61.365 ;
        RECT -24.645 59.675 -24.315 60.005 ;
        RECT -24.645 58.315 -24.315 58.645 ;
        RECT -24.645 56.955 -24.315 57.285 ;
        RECT -24.645 55.595 -24.315 55.925 ;
        RECT -24.645 54.235 -24.315 54.565 ;
        RECT -24.645 52.875 -24.315 53.205 ;
        RECT -24.645 51.515 -24.315 51.845 ;
        RECT -24.645 50.155 -24.315 50.485 ;
        RECT -24.645 48.795 -24.315 49.125 ;
        RECT -24.645 47.435 -24.315 47.765 ;
        RECT -24.645 46.075 -24.315 46.405 ;
        RECT -24.645 44.715 -24.315 45.045 ;
        RECT -24.645 43.355 -24.315 43.685 ;
        RECT -24.645 41.995 -24.315 42.325 ;
        RECT -24.645 40.635 -24.315 40.965 ;
        RECT -24.645 39.275 -24.315 39.605 ;
        RECT -24.645 37.915 -24.315 38.245 ;
        RECT -24.645 36.555 -24.315 36.885 ;
        RECT -24.645 35.195 -24.315 35.525 ;
        RECT -24.645 33.835 -24.315 34.165 ;
        RECT -24.645 32.475 -24.315 32.805 ;
        RECT -24.645 31.115 -24.315 31.445 ;
        RECT -24.645 29.755 -24.315 30.085 ;
        RECT -24.645 28.395 -24.315 28.725 ;
        RECT -24.645 27.035 -24.315 27.365 ;
        RECT -24.645 25.675 -24.315 26.005 ;
        RECT -24.645 24.315 -24.315 24.645 ;
        RECT -24.645 22.955 -24.315 23.285 ;
        RECT -24.645 21.595 -24.315 21.925 ;
        RECT -24.645 20.235 -24.315 20.565 ;
        RECT -24.645 18.875 -24.315 19.205 ;
        RECT -24.645 17.515 -24.315 17.845 ;
        RECT -24.645 16.155 -24.315 16.485 ;
        RECT -24.645 14.795 -24.315 15.125 ;
        RECT -24.645 13.435 -24.315 13.765 ;
        RECT -24.645 12.075 -24.315 12.405 ;
        RECT -24.645 10.715 -24.315 11.045 ;
        RECT -24.645 9.355 -24.315 9.685 ;
        RECT -24.645 7.995 -24.315 8.325 ;
        RECT -24.645 6.635 -24.315 6.965 ;
        RECT -24.645 5.275 -24.315 5.605 ;
        RECT -24.645 3.915 -24.315 4.245 ;
        RECT -24.645 2.555 -24.315 2.885 ;
        RECT -24.645 1.195 -24.315 1.525 ;
        RECT -24.645 -0.165 -24.315 0.165 ;
        RECT -24.645 -1.525 -24.315 -1.195 ;
        RECT -24.645 -12.41 -24.315 -12.08 ;
        RECT -24.645 -15.125 -24.315 -14.795 ;
        RECT -24.645 -16.485 -24.315 -16.155 ;
        RECT -24.645 -17.25 -24.315 -16.92 ;
        RECT -24.645 -19.205 -24.315 -18.875 ;
        RECT -24.645 -28.725 -24.315 -28.395 ;
        RECT -24.645 -30.085 -24.315 -29.755 ;
        RECT -24.645 -32.805 -24.315 -32.475 ;
        RECT -24.645 -34.165 -24.315 -33.835 ;
        RECT -24.645 -35.39 -24.315 -35.06 ;
        RECT -24.645 -38.245 -24.315 -37.915 ;
        RECT -24.645 -40.23 -24.315 -39.9 ;
        RECT -24.645 -40.965 -24.315 -40.635 ;
        RECT -24.645 -50.485 -24.315 -50.155 ;
        RECT -24.645 -51.845 -24.315 -51.515 ;
        RECT -24.645 -53.205 -24.315 -52.875 ;
        RECT -24.645 -54.565 -24.315 -54.235 ;
        RECT -24.645 -55.925 -24.315 -55.595 ;
        RECT -24.645 -57.285 -24.315 -56.955 ;
        RECT -24.645 -58.645 -24.315 -58.315 ;
        RECT -24.645 -60.005 -24.315 -59.675 ;
        RECT -24.645 -61.365 -24.315 -61.035 ;
        RECT -24.645 -62.725 -24.315 -62.395 ;
        RECT -24.645 -64.085 -24.315 -63.755 ;
        RECT -24.645 -65.445 -24.315 -65.115 ;
        RECT -24.645 -66.805 -24.315 -66.475 ;
        RECT -24.645 -68.165 -24.315 -67.835 ;
        RECT -24.645 -69.525 -24.315 -69.195 ;
        RECT -24.645 -70.885 -24.315 -70.555 ;
        RECT -24.645 -72.245 -24.315 -71.915 ;
        RECT -24.645 -73.605 -24.315 -73.275 ;
        RECT -24.645 -74.965 -24.315 -74.635 ;
        RECT -24.645 -76.325 -24.315 -75.995 ;
        RECT -24.645 -77.685 -24.315 -77.355 ;
        RECT -24.645 -79.045 -24.315 -78.715 ;
        RECT -24.645 -80.405 -24.315 -80.075 ;
        RECT -24.645 -81.765 -24.315 -81.435 ;
        RECT -24.645 -83.125 -24.315 -82.795 ;
        RECT -24.645 -84.485 -24.315 -84.155 ;
        RECT -24.645 -85.845 -24.315 -85.515 ;
        RECT -24.645 -87.205 -24.315 -86.875 ;
        RECT -24.645 -88.565 -24.315 -88.235 ;
        RECT -24.645 -89.925 -24.315 -89.595 ;
        RECT -24.645 -91.285 -24.315 -90.955 ;
        RECT -24.645 -92.645 -24.315 -92.315 ;
        RECT -24.645 -94.005 -24.315 -93.675 ;
        RECT -24.645 -95.365 -24.315 -95.035 ;
        RECT -24.645 -96.725 -24.315 -96.395 ;
        RECT -24.645 -98.085 -24.315 -97.755 ;
        RECT -24.645 -102.165 -24.315 -101.835 ;
        RECT -24.645 -103.525 -24.315 -103.195 ;
        RECT -24.645 -104.885 -24.315 -104.555 ;
        RECT -24.645 -106.245 -24.315 -105.915 ;
        RECT -24.645 -107.605 -24.315 -107.275 ;
        RECT -24.645 -108.965 -24.315 -108.635 ;
        RECT -24.645 -114.405 -24.315 -114.075 ;
        RECT -24.645 -115.765 -24.315 -115.435 ;
        RECT -24.645 -118.485 -24.315 -118.155 ;
        RECT -24.645 -121.205 -24.315 -120.875 ;
        RECT -24.645 -122.565 -24.315 -122.235 ;
        RECT -24.645 -125.285 -24.315 -124.955 ;
        RECT -24.645 -126.645 -24.315 -126.315 ;
        RECT -24.645 -128.005 -24.315 -127.675 ;
        RECT -24.645 -130.725 -24.315 -130.395 ;
        RECT -24.645 -132.085 -24.315 -131.755 ;
        RECT -24.645 -136.165 -24.315 -135.835 ;
        RECT -24.645 -137.525 -24.315 -137.195 ;
        RECT -24.645 -138.885 -24.315 -138.555 ;
        RECT -24.645 -140.245 -24.315 -139.915 ;
        RECT -24.645 -141.605 -24.315 -141.275 ;
        RECT -24.645 -142.965 -24.315 -142.635 ;
        RECT -24.645 -144.325 -24.315 -143.995 ;
        RECT -24.645 -145.685 -24.315 -145.355 ;
        RECT -24.645 -147.045 -24.315 -146.715 ;
        RECT -24.645 -149.765 -24.315 -149.435 ;
        RECT -24.645 -152.485 -24.315 -152.155 ;
        RECT -24.645 -153.845 -24.315 -153.515 ;
        RECT -24.645 -155.285 -24.315 -154.955 ;
        RECT -24.645 -156.565 -24.315 -156.235 ;
        RECT -24.645 -157.925 -24.315 -157.595 ;
        RECT -24.645 -160.17 -24.315 -159.04 ;
        RECT -24.64 -160.285 -24.32 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 127.225 -22.955 128.355 ;
        RECT -23.285 124.955 -22.955 125.285 ;
        RECT -23.285 123.595 -22.955 123.925 ;
        RECT -23.285 122.235 -22.955 122.565 ;
        RECT -23.285 120.875 -22.955 121.205 ;
        RECT -23.285 119.515 -22.955 119.845 ;
        RECT -23.285 118.155 -22.955 118.485 ;
        RECT -23.285 116.795 -22.955 117.125 ;
        RECT -23.285 115.435 -22.955 115.765 ;
        RECT -23.285 114.075 -22.955 114.405 ;
        RECT -23.285 112.715 -22.955 113.045 ;
        RECT -23.285 111.355 -22.955 111.685 ;
        RECT -23.285 109.995 -22.955 110.325 ;
        RECT -23.285 108.635 -22.955 108.965 ;
        RECT -23.285 107.275 -22.955 107.605 ;
        RECT -23.285 105.915 -22.955 106.245 ;
        RECT -23.285 104.555 -22.955 104.885 ;
        RECT -23.285 103.195 -22.955 103.525 ;
        RECT -23.285 101.835 -22.955 102.165 ;
        RECT -23.285 100.475 -22.955 100.805 ;
        RECT -23.285 99.115 -22.955 99.445 ;
        RECT -23.285 97.755 -22.955 98.085 ;
        RECT -23.285 96.395 -22.955 96.725 ;
        RECT -23.285 95.035 -22.955 95.365 ;
        RECT -23.285 93.675 -22.955 94.005 ;
        RECT -23.285 92.315 -22.955 92.645 ;
        RECT -23.285 90.955 -22.955 91.285 ;
        RECT -23.285 89.595 -22.955 89.925 ;
        RECT -23.285 88.235 -22.955 88.565 ;
        RECT -23.285 86.875 -22.955 87.205 ;
        RECT -23.285 85.515 -22.955 85.845 ;
        RECT -23.285 84.155 -22.955 84.485 ;
        RECT -23.285 82.795 -22.955 83.125 ;
        RECT -23.285 81.435 -22.955 81.765 ;
        RECT -23.285 80.075 -22.955 80.405 ;
        RECT -23.285 78.715 -22.955 79.045 ;
        RECT -23.285 77.355 -22.955 77.685 ;
        RECT -23.285 75.995 -22.955 76.325 ;
        RECT -23.285 74.635 -22.955 74.965 ;
        RECT -23.285 73.275 -22.955 73.605 ;
        RECT -23.285 71.915 -22.955 72.245 ;
        RECT -23.285 70.555 -22.955 70.885 ;
        RECT -23.285 69.195 -22.955 69.525 ;
        RECT -23.285 67.835 -22.955 68.165 ;
        RECT -23.285 66.475 -22.955 66.805 ;
        RECT -23.285 65.115 -22.955 65.445 ;
        RECT -23.285 63.755 -22.955 64.085 ;
        RECT -23.285 62.395 -22.955 62.725 ;
        RECT -23.285 61.035 -22.955 61.365 ;
        RECT -23.285 59.675 -22.955 60.005 ;
        RECT -23.285 58.315 -22.955 58.645 ;
        RECT -23.285 56.955 -22.955 57.285 ;
        RECT -23.285 55.595 -22.955 55.925 ;
        RECT -23.285 54.235 -22.955 54.565 ;
        RECT -23.285 52.875 -22.955 53.205 ;
        RECT -23.285 51.515 -22.955 51.845 ;
        RECT -23.285 50.155 -22.955 50.485 ;
        RECT -23.285 48.795 -22.955 49.125 ;
        RECT -23.285 47.435 -22.955 47.765 ;
        RECT -23.285 46.075 -22.955 46.405 ;
        RECT -23.285 44.715 -22.955 45.045 ;
        RECT -23.285 43.355 -22.955 43.685 ;
        RECT -23.285 41.995 -22.955 42.325 ;
        RECT -23.285 40.635 -22.955 40.965 ;
        RECT -23.285 39.275 -22.955 39.605 ;
        RECT -23.285 37.915 -22.955 38.245 ;
        RECT -23.285 36.555 -22.955 36.885 ;
        RECT -23.285 35.195 -22.955 35.525 ;
        RECT -23.285 33.835 -22.955 34.165 ;
        RECT -23.285 32.475 -22.955 32.805 ;
        RECT -23.285 31.115 -22.955 31.445 ;
        RECT -23.285 29.755 -22.955 30.085 ;
        RECT -23.285 28.395 -22.955 28.725 ;
        RECT -23.285 27.035 -22.955 27.365 ;
        RECT -23.285 25.675 -22.955 26.005 ;
        RECT -23.285 24.315 -22.955 24.645 ;
        RECT -23.285 22.955 -22.955 23.285 ;
        RECT -23.285 21.595 -22.955 21.925 ;
        RECT -23.285 20.235 -22.955 20.565 ;
        RECT -23.285 18.875 -22.955 19.205 ;
        RECT -23.285 17.515 -22.955 17.845 ;
        RECT -23.285 16.155 -22.955 16.485 ;
        RECT -23.285 14.795 -22.955 15.125 ;
        RECT -23.285 13.435 -22.955 13.765 ;
        RECT -23.285 12.075 -22.955 12.405 ;
        RECT -23.285 10.715 -22.955 11.045 ;
        RECT -23.285 9.355 -22.955 9.685 ;
        RECT -23.285 7.995 -22.955 8.325 ;
        RECT -23.285 6.635 -22.955 6.965 ;
        RECT -23.285 5.275 -22.955 5.605 ;
        RECT -23.285 3.915 -22.955 4.245 ;
        RECT -23.285 2.555 -22.955 2.885 ;
        RECT -23.285 1.195 -22.955 1.525 ;
        RECT -23.285 -0.165 -22.955 0.165 ;
        RECT -23.285 -1.525 -22.955 -1.195 ;
        RECT -23.285 -12.41 -22.955 -12.08 ;
        RECT -23.285 -15.125 -22.955 -14.795 ;
        RECT -23.285 -16.485 -22.955 -16.155 ;
        RECT -23.285 -17.25 -22.955 -16.92 ;
        RECT -23.285 -19.205 -22.955 -18.875 ;
        RECT -23.285 -28.725 -22.955 -28.395 ;
        RECT -23.285 -30.085 -22.955 -29.755 ;
        RECT -23.285 -32.805 -22.955 -32.475 ;
        RECT -23.285 -34.165 -22.955 -33.835 ;
        RECT -23.285 -35.39 -22.955 -35.06 ;
        RECT -23.285 -38.245 -22.955 -37.915 ;
        RECT -23.285 -40.23 -22.955 -39.9 ;
        RECT -23.285 -40.965 -22.955 -40.635 ;
        RECT -23.285 -50.485 -22.955 -50.155 ;
        RECT -23.285 -51.845 -22.955 -51.515 ;
        RECT -23.285 -53.205 -22.955 -52.875 ;
        RECT -23.285 -54.565 -22.955 -54.235 ;
        RECT -23.285 -55.925 -22.955 -55.595 ;
        RECT -23.285 -57.285 -22.955 -56.955 ;
        RECT -23.285 -58.645 -22.955 -58.315 ;
        RECT -23.285 -60.005 -22.955 -59.675 ;
        RECT -23.285 -61.365 -22.955 -61.035 ;
        RECT -23.285 -62.725 -22.955 -62.395 ;
        RECT -23.285 -64.085 -22.955 -63.755 ;
        RECT -23.285 -65.445 -22.955 -65.115 ;
        RECT -23.285 -66.805 -22.955 -66.475 ;
        RECT -23.285 -68.165 -22.955 -67.835 ;
        RECT -23.285 -69.525 -22.955 -69.195 ;
        RECT -23.285 -70.885 -22.955 -70.555 ;
        RECT -23.285 -72.245 -22.955 -71.915 ;
        RECT -23.285 -73.605 -22.955 -73.275 ;
        RECT -23.285 -74.965 -22.955 -74.635 ;
        RECT -23.285 -76.325 -22.955 -75.995 ;
        RECT -23.285 -77.685 -22.955 -77.355 ;
        RECT -23.285 -79.045 -22.955 -78.715 ;
        RECT -23.285 -80.405 -22.955 -80.075 ;
        RECT -23.285 -81.765 -22.955 -81.435 ;
        RECT -23.285 -83.125 -22.955 -82.795 ;
        RECT -23.285 -84.485 -22.955 -84.155 ;
        RECT -23.285 -85.845 -22.955 -85.515 ;
        RECT -23.285 -87.205 -22.955 -86.875 ;
        RECT -23.285 -88.565 -22.955 -88.235 ;
        RECT -23.285 -89.925 -22.955 -89.595 ;
        RECT -23.285 -91.285 -22.955 -90.955 ;
        RECT -23.28 -91.96 -22.96 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 -153.845 -22.955 -153.515 ;
        RECT -23.285 -155.285 -22.955 -154.955 ;
        RECT -23.285 -156.565 -22.955 -156.235 ;
        RECT -23.285 -157.925 -22.955 -157.595 ;
        RECT -23.285 -160.17 -22.955 -159.04 ;
        RECT -23.28 -160.285 -22.96 -153.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 127.225 -21.595 128.355 ;
        RECT -21.925 124.955 -21.595 125.285 ;
        RECT -21.925 123.595 -21.595 123.925 ;
        RECT -21.925 122.235 -21.595 122.565 ;
        RECT -21.925 120.875 -21.595 121.205 ;
        RECT -21.925 119.515 -21.595 119.845 ;
        RECT -21.925 118.155 -21.595 118.485 ;
        RECT -21.925 116.795 -21.595 117.125 ;
        RECT -21.925 115.435 -21.595 115.765 ;
        RECT -21.925 114.075 -21.595 114.405 ;
        RECT -21.925 112.715 -21.595 113.045 ;
        RECT -21.925 111.355 -21.595 111.685 ;
        RECT -21.925 109.995 -21.595 110.325 ;
        RECT -21.925 108.635 -21.595 108.965 ;
        RECT -21.925 107.275 -21.595 107.605 ;
        RECT -21.925 105.915 -21.595 106.245 ;
        RECT -21.925 104.555 -21.595 104.885 ;
        RECT -21.925 103.195 -21.595 103.525 ;
        RECT -21.925 101.835 -21.595 102.165 ;
        RECT -21.925 100.475 -21.595 100.805 ;
        RECT -21.925 99.115 -21.595 99.445 ;
        RECT -21.925 97.755 -21.595 98.085 ;
        RECT -21.925 96.395 -21.595 96.725 ;
        RECT -21.925 95.035 -21.595 95.365 ;
        RECT -21.925 93.675 -21.595 94.005 ;
        RECT -21.925 92.315 -21.595 92.645 ;
        RECT -21.925 90.955 -21.595 91.285 ;
        RECT -21.925 89.595 -21.595 89.925 ;
        RECT -21.925 88.235 -21.595 88.565 ;
        RECT -21.925 86.875 -21.595 87.205 ;
        RECT -21.925 85.515 -21.595 85.845 ;
        RECT -21.925 84.155 -21.595 84.485 ;
        RECT -21.925 82.795 -21.595 83.125 ;
        RECT -21.925 81.435 -21.595 81.765 ;
        RECT -21.925 80.075 -21.595 80.405 ;
        RECT -21.925 78.715 -21.595 79.045 ;
        RECT -21.925 77.355 -21.595 77.685 ;
        RECT -21.925 75.995 -21.595 76.325 ;
        RECT -21.925 74.635 -21.595 74.965 ;
        RECT -21.925 73.275 -21.595 73.605 ;
        RECT -21.925 71.915 -21.595 72.245 ;
        RECT -21.925 70.555 -21.595 70.885 ;
        RECT -21.925 69.195 -21.595 69.525 ;
        RECT -21.925 67.835 -21.595 68.165 ;
        RECT -21.925 66.475 -21.595 66.805 ;
        RECT -21.925 65.115 -21.595 65.445 ;
        RECT -21.925 63.755 -21.595 64.085 ;
        RECT -21.925 62.395 -21.595 62.725 ;
        RECT -21.925 61.035 -21.595 61.365 ;
        RECT -21.925 59.675 -21.595 60.005 ;
        RECT -21.925 58.315 -21.595 58.645 ;
        RECT -21.925 56.955 -21.595 57.285 ;
        RECT -21.925 55.595 -21.595 55.925 ;
        RECT -21.925 54.235 -21.595 54.565 ;
        RECT -21.925 52.875 -21.595 53.205 ;
        RECT -21.925 51.515 -21.595 51.845 ;
        RECT -21.925 50.155 -21.595 50.485 ;
        RECT -21.925 48.795 -21.595 49.125 ;
        RECT -21.925 47.435 -21.595 47.765 ;
        RECT -21.925 46.075 -21.595 46.405 ;
        RECT -21.925 44.715 -21.595 45.045 ;
        RECT -21.925 43.355 -21.595 43.685 ;
        RECT -21.925 41.995 -21.595 42.325 ;
        RECT -21.925 40.635 -21.595 40.965 ;
        RECT -21.925 39.275 -21.595 39.605 ;
        RECT -21.925 37.915 -21.595 38.245 ;
        RECT -21.925 36.555 -21.595 36.885 ;
        RECT -21.925 35.195 -21.595 35.525 ;
        RECT -21.925 33.835 -21.595 34.165 ;
        RECT -21.925 32.475 -21.595 32.805 ;
        RECT -21.925 31.115 -21.595 31.445 ;
        RECT -21.925 29.755 -21.595 30.085 ;
        RECT -21.925 28.395 -21.595 28.725 ;
        RECT -21.925 27.035 -21.595 27.365 ;
        RECT -21.925 25.675 -21.595 26.005 ;
        RECT -21.925 24.315 -21.595 24.645 ;
        RECT -21.925 22.955 -21.595 23.285 ;
        RECT -21.925 21.595 -21.595 21.925 ;
        RECT -21.925 20.235 -21.595 20.565 ;
        RECT -21.925 18.875 -21.595 19.205 ;
        RECT -21.925 17.515 -21.595 17.845 ;
        RECT -21.925 16.155 -21.595 16.485 ;
        RECT -21.925 14.795 -21.595 15.125 ;
        RECT -21.925 13.435 -21.595 13.765 ;
        RECT -21.925 12.075 -21.595 12.405 ;
        RECT -21.925 10.715 -21.595 11.045 ;
        RECT -21.925 9.355 -21.595 9.685 ;
        RECT -21.925 7.995 -21.595 8.325 ;
        RECT -21.925 6.635 -21.595 6.965 ;
        RECT -21.925 5.275 -21.595 5.605 ;
        RECT -21.925 3.915 -21.595 4.245 ;
        RECT -21.925 2.555 -21.595 2.885 ;
        RECT -21.925 1.195 -21.595 1.525 ;
        RECT -21.925 -0.165 -21.595 0.165 ;
        RECT -21.925 -1.525 -21.595 -1.195 ;
        RECT -21.92 -6.28 -21.6 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 -58.645 -21.595 -58.315 ;
        RECT -21.925 -60.005 -21.595 -59.675 ;
        RECT -21.925 -61.365 -21.595 -61.035 ;
        RECT -21.925 -62.725 -21.595 -62.395 ;
        RECT -21.925 -64.085 -21.595 -63.755 ;
        RECT -21.925 -65.445 -21.595 -65.115 ;
        RECT -21.925 -66.805 -21.595 -66.475 ;
        RECT -21.925 -68.165 -21.595 -67.835 ;
        RECT -21.925 -69.525 -21.595 -69.195 ;
        RECT -21.925 -70.885 -21.595 -70.555 ;
        RECT -21.925 -72.245 -21.595 -71.915 ;
        RECT -21.925 -73.605 -21.595 -73.275 ;
        RECT -21.925 -74.965 -21.595 -74.635 ;
        RECT -21.925 -76.325 -21.595 -75.995 ;
        RECT -21.925 -77.685 -21.595 -77.355 ;
        RECT -21.925 -79.045 -21.595 -78.715 ;
        RECT -21.925 -80.405 -21.595 -80.075 ;
        RECT -21.925 -81.765 -21.595 -81.435 ;
        RECT -21.925 -83.125 -21.595 -82.795 ;
        RECT -21.925 -84.485 -21.595 -84.155 ;
        RECT -21.925 -85.845 -21.595 -85.515 ;
        RECT -21.925 -87.205 -21.595 -86.875 ;
        RECT -21.925 -88.565 -21.595 -88.235 ;
        RECT -21.925 -89.925 -21.595 -89.595 ;
        RECT -21.925 -91.285 -21.595 -90.955 ;
        RECT -21.925 -94.005 -21.595 -93.675 ;
        RECT -21.925 -95.365 -21.595 -95.035 ;
        RECT -21.925 -96.725 -21.595 -96.395 ;
        RECT -21.925 -98.085 -21.595 -97.755 ;
        RECT -21.925 -102.165 -21.595 -101.835 ;
        RECT -21.925 -103.525 -21.595 -103.195 ;
        RECT -21.925 -104.885 -21.595 -104.555 ;
        RECT -21.925 -106.245 -21.595 -105.915 ;
        RECT -21.925 -107.605 -21.595 -107.275 ;
        RECT -21.925 -114.405 -21.595 -114.075 ;
        RECT -21.925 -115.765 -21.595 -115.435 ;
        RECT -21.925 -118.485 -21.595 -118.155 ;
        RECT -21.925 -121.205 -21.595 -120.875 ;
        RECT -21.925 -122.565 -21.595 -122.235 ;
        RECT -21.925 -125.285 -21.595 -124.955 ;
        RECT -21.925 -126.645 -21.595 -126.315 ;
        RECT -21.925 -128.005 -21.595 -127.675 ;
        RECT -21.925 -130.725 -21.595 -130.395 ;
        RECT -21.925 -132.085 -21.595 -131.755 ;
        RECT -21.925 -136.165 -21.595 -135.835 ;
        RECT -21.925 -137.525 -21.595 -137.195 ;
        RECT -21.925 -138.885 -21.595 -138.555 ;
        RECT -21.925 -140.245 -21.595 -139.915 ;
        RECT -21.925 -141.605 -21.595 -141.275 ;
        RECT -21.925 -142.965 -21.595 -142.635 ;
        RECT -21.925 -144.325 -21.595 -143.995 ;
        RECT -21.925 -145.685 -21.595 -145.355 ;
        RECT -21.925 -147.045 -21.595 -146.715 ;
        RECT -21.925 -149.765 -21.595 -149.435 ;
        RECT -21.925 -153.845 -21.595 -153.515 ;
        RECT -21.925 -155.285 -21.595 -154.955 ;
        RECT -21.925 -156.565 -21.595 -156.235 ;
        RECT -21.925 -157.925 -21.595 -157.595 ;
        RECT -21.925 -160.17 -21.595 -159.04 ;
        RECT -21.92 -160.285 -21.6 -27.72 ;
        RECT -21.925 -28.725 -21.595 -28.395 ;
        RECT -21.925 -30.085 -21.595 -29.755 ;
        RECT -21.925 -32.805 -21.595 -32.475 ;
        RECT -21.925 -34.165 -21.595 -33.835 ;
        RECT -21.925 -35.39 -21.595 -35.06 ;
        RECT -21.925 -38.245 -21.595 -37.915 ;
        RECT -21.925 -40.23 -21.595 -39.9 ;
        RECT -21.925 -40.965 -21.595 -40.635 ;
        RECT -21.925 -50.485 -21.595 -50.155 ;
        RECT -21.925 -51.845 -21.595 -51.515 ;
        RECT -21.925 -53.205 -21.595 -52.875 ;
        RECT -21.925 -54.565 -21.595 -54.235 ;
        RECT -21.925 -55.925 -21.595 -55.595 ;
        RECT -21.925 -57.285 -21.595 -56.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.885 127.225 -36.555 128.355 ;
        RECT -36.885 124.955 -36.555 125.285 ;
        RECT -36.885 123.595 -36.555 123.925 ;
        RECT -36.885 122.235 -36.555 122.565 ;
        RECT -36.885 120.875 -36.555 121.205 ;
        RECT -36.885 119.515 -36.555 119.845 ;
        RECT -36.885 118.155 -36.555 118.485 ;
        RECT -36.885 116.795 -36.555 117.125 ;
        RECT -36.885 115.435 -36.555 115.765 ;
        RECT -36.885 114.075 -36.555 114.405 ;
        RECT -36.885 112.715 -36.555 113.045 ;
        RECT -36.885 111.355 -36.555 111.685 ;
        RECT -36.885 109.995 -36.555 110.325 ;
        RECT -36.885 108.635 -36.555 108.965 ;
        RECT -36.885 107.275 -36.555 107.605 ;
        RECT -36.885 105.915 -36.555 106.245 ;
        RECT -36.885 104.555 -36.555 104.885 ;
        RECT -36.885 103.195 -36.555 103.525 ;
        RECT -36.885 101.835 -36.555 102.165 ;
        RECT -36.885 100.475 -36.555 100.805 ;
        RECT -36.885 99.115 -36.555 99.445 ;
        RECT -36.885 97.755 -36.555 98.085 ;
        RECT -36.885 96.395 -36.555 96.725 ;
        RECT -36.885 95.035 -36.555 95.365 ;
        RECT -36.885 93.675 -36.555 94.005 ;
        RECT -36.885 92.315 -36.555 92.645 ;
        RECT -36.885 90.955 -36.555 91.285 ;
        RECT -36.885 89.595 -36.555 89.925 ;
        RECT -36.885 88.235 -36.555 88.565 ;
        RECT -36.885 86.875 -36.555 87.205 ;
        RECT -36.885 85.515 -36.555 85.845 ;
        RECT -36.885 84.155 -36.555 84.485 ;
        RECT -36.885 82.795 -36.555 83.125 ;
        RECT -36.885 81.435 -36.555 81.765 ;
        RECT -36.885 80.075 -36.555 80.405 ;
        RECT -36.885 78.715 -36.555 79.045 ;
        RECT -36.885 77.355 -36.555 77.685 ;
        RECT -36.885 75.995 -36.555 76.325 ;
        RECT -36.885 74.635 -36.555 74.965 ;
        RECT -36.885 73.275 -36.555 73.605 ;
        RECT -36.885 71.915 -36.555 72.245 ;
        RECT -36.885 70.555 -36.555 70.885 ;
        RECT -36.885 69.195 -36.555 69.525 ;
        RECT -36.885 67.835 -36.555 68.165 ;
        RECT -36.885 66.475 -36.555 66.805 ;
        RECT -36.885 65.115 -36.555 65.445 ;
        RECT -36.885 63.755 -36.555 64.085 ;
        RECT -36.885 62.395 -36.555 62.725 ;
        RECT -36.885 61.035 -36.555 61.365 ;
        RECT -36.885 59.675 -36.555 60.005 ;
        RECT -36.885 58.315 -36.555 58.645 ;
        RECT -36.885 56.955 -36.555 57.285 ;
        RECT -36.885 55.595 -36.555 55.925 ;
        RECT -36.885 54.235 -36.555 54.565 ;
        RECT -36.885 52.875 -36.555 53.205 ;
        RECT -36.885 51.515 -36.555 51.845 ;
        RECT -36.885 50.155 -36.555 50.485 ;
        RECT -36.885 48.795 -36.555 49.125 ;
        RECT -36.885 47.435 -36.555 47.765 ;
        RECT -36.885 46.075 -36.555 46.405 ;
        RECT -36.885 44.715 -36.555 45.045 ;
        RECT -36.885 43.355 -36.555 43.685 ;
        RECT -36.885 41.995 -36.555 42.325 ;
        RECT -36.885 40.635 -36.555 40.965 ;
        RECT -36.885 39.275 -36.555 39.605 ;
        RECT -36.885 37.915 -36.555 38.245 ;
        RECT -36.885 36.555 -36.555 36.885 ;
        RECT -36.885 35.195 -36.555 35.525 ;
        RECT -36.885 33.835 -36.555 34.165 ;
        RECT -36.885 32.475 -36.555 32.805 ;
        RECT -36.885 31.115 -36.555 31.445 ;
        RECT -36.885 29.755 -36.555 30.085 ;
        RECT -36.885 28.395 -36.555 28.725 ;
        RECT -36.885 27.035 -36.555 27.365 ;
        RECT -36.885 25.675 -36.555 26.005 ;
        RECT -36.885 24.315 -36.555 24.645 ;
        RECT -36.885 22.955 -36.555 23.285 ;
        RECT -36.885 21.595 -36.555 21.925 ;
        RECT -36.885 20.235 -36.555 20.565 ;
        RECT -36.885 18.875 -36.555 19.205 ;
        RECT -36.885 17.515 -36.555 17.845 ;
        RECT -36.885 16.155 -36.555 16.485 ;
        RECT -36.885 14.795 -36.555 15.125 ;
        RECT -36.885 13.435 -36.555 13.765 ;
        RECT -36.885 12.075 -36.555 12.405 ;
        RECT -36.885 10.715 -36.555 11.045 ;
        RECT -36.885 9.355 -36.555 9.685 ;
        RECT -36.885 7.995 -36.555 8.325 ;
        RECT -36.885 6.635 -36.555 6.965 ;
        RECT -36.885 5.275 -36.555 5.605 ;
        RECT -36.885 3.915 -36.555 4.245 ;
        RECT -36.885 2.555 -36.555 2.885 ;
        RECT -36.885 1.195 -36.555 1.525 ;
        RECT -36.885 -0.165 -36.555 0.165 ;
        RECT -36.885 -8.325 -36.555 -7.995 ;
        RECT -36.885 -12.405 -36.555 -12.075 ;
        RECT -36.885 -13.765 -36.555 -13.435 ;
        RECT -36.885 -15.125 -36.555 -14.795 ;
        RECT -36.885 -16.485 -36.555 -16.155 ;
        RECT -36.885 -17.845 -36.555 -17.515 ;
        RECT -36.885 -19.205 -36.555 -18.875 ;
        RECT -36.885 -20.565 -36.555 -20.235 ;
        RECT -36.885 -21.925 -36.555 -21.595 ;
        RECT -36.885 -28.725 -36.555 -28.395 ;
        RECT -36.885 -30.085 -36.555 -29.755 ;
        RECT -36.885 -31.445 -36.555 -31.115 ;
        RECT -36.885 -32.805 -36.555 -32.475 ;
        RECT -36.885 -34.165 -36.555 -33.835 ;
        RECT -36.885 -35.525 -36.555 -35.195 ;
        RECT -36.885 -36.885 -36.555 -36.555 ;
        RECT -36.885 -38.245 -36.555 -37.915 ;
        RECT -36.885 -39.605 -36.555 -39.275 ;
        RECT -36.885 -40.965 -36.555 -40.635 ;
        RECT -36.885 -42.325 -36.555 -41.995 ;
        RECT -36.885 -43.685 -36.555 -43.355 ;
        RECT -36.885 -45.045 -36.555 -44.715 ;
        RECT -36.885 -47.765 -36.555 -47.435 ;
        RECT -36.885 -49.125 -36.555 -48.795 ;
        RECT -36.885 -50.485 -36.555 -50.155 ;
        RECT -36.885 -51.845 -36.555 -51.515 ;
        RECT -36.885 -53.205 -36.555 -52.875 ;
        RECT -36.885 -54.565 -36.555 -54.235 ;
        RECT -36.885 -55.925 -36.555 -55.595 ;
        RECT -36.885 -57.285 -36.555 -56.955 ;
        RECT -36.885 -58.645 -36.555 -58.315 ;
        RECT -36.885 -60.005 -36.555 -59.675 ;
        RECT -36.885 -61.365 -36.555 -61.035 ;
        RECT -36.885 -62.725 -36.555 -62.395 ;
        RECT -36.885 -64.085 -36.555 -63.755 ;
        RECT -36.885 -65.445 -36.555 -65.115 ;
        RECT -36.885 -66.805 -36.555 -66.475 ;
        RECT -36.885 -68.165 -36.555 -67.835 ;
        RECT -36.885 -69.525 -36.555 -69.195 ;
        RECT -36.885 -72.245 -36.555 -71.915 ;
        RECT -36.885 -73.605 -36.555 -73.275 ;
        RECT -36.885 -74.965 -36.555 -74.635 ;
        RECT -36.885 -76.325 -36.555 -75.995 ;
        RECT -36.885 -78.29 -36.555 -77.96 ;
        RECT -36.885 -79.045 -36.555 -78.715 ;
        RECT -36.885 -81.765 -36.555 -81.435 ;
        RECT -36.885 -83.125 -36.555 -82.795 ;
        RECT -36.885 -84.485 -36.555 -84.155 ;
        RECT -36.885 -86.43 -36.555 -86.1 ;
        RECT -36.885 -87.205 -36.555 -86.875 ;
        RECT -36.885 -88.565 -36.555 -88.235 ;
        RECT -36.885 -89.925 -36.555 -89.595 ;
        RECT -36.885 -92.645 -36.555 -92.315 ;
        RECT -36.885 -94.005 -36.555 -93.675 ;
        RECT -36.885 -95.365 -36.555 -95.035 ;
        RECT -36.885 -96.725 -36.555 -96.395 ;
        RECT -36.885 -98.085 -36.555 -97.755 ;
        RECT -36.885 -102.165 -36.555 -101.835 ;
        RECT -36.885 -103.525 -36.555 -103.195 ;
        RECT -36.885 -104.885 -36.555 -104.555 ;
        RECT -36.885 -106.245 -36.555 -105.915 ;
        RECT -36.885 -107.605 -36.555 -107.275 ;
        RECT -36.885 -108.965 -36.555 -108.635 ;
        RECT -36.885 -113.045 -36.555 -112.715 ;
        RECT -36.885 -114.405 -36.555 -114.075 ;
        RECT -36.885 -115.765 -36.555 -115.435 ;
        RECT -36.885 -117.125 -36.555 -116.795 ;
        RECT -36.885 -118.485 -36.555 -118.155 ;
        RECT -36.885 -119.845 -36.555 -119.515 ;
        RECT -36.885 -121.205 -36.555 -120.875 ;
        RECT -36.885 -122.565 -36.555 -122.235 ;
        RECT -36.885 -123.925 -36.555 -123.595 ;
        RECT -36.885 -125.285 -36.555 -124.955 ;
        RECT -36.885 -126.645 -36.555 -126.315 ;
        RECT -36.885 -128.005 -36.555 -127.675 ;
        RECT -36.885 -130.725 -36.555 -130.395 ;
        RECT -36.885 -132.085 -36.555 -131.755 ;
        RECT -36.885 -136.165 -36.555 -135.835 ;
        RECT -36.885 -137.525 -36.555 -137.195 ;
        RECT -36.885 -138.885 -36.555 -138.555 ;
        RECT -36.885 -140.245 -36.555 -139.915 ;
        RECT -36.885 -141.605 -36.555 -141.275 ;
        RECT -36.885 -142.965 -36.555 -142.635 ;
        RECT -36.885 -144.325 -36.555 -143.995 ;
        RECT -36.885 -145.685 -36.555 -145.355 ;
        RECT -36.885 -147.045 -36.555 -146.715 ;
        RECT -36.885 -149.765 -36.555 -149.435 ;
        RECT -36.885 -152.485 -36.555 -152.155 ;
        RECT -36.885 -153.845 -36.555 -153.515 ;
        RECT -36.885 -155.285 -36.555 -154.955 ;
        RECT -36.885 -156.565 -36.555 -156.235 ;
        RECT -36.885 -157.925 -36.555 -157.595 ;
        RECT -36.885 -160.17 -36.555 -159.04 ;
        RECT -36.88 -160.285 -36.56 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 127.225 -35.195 128.355 ;
        RECT -35.525 124.955 -35.195 125.285 ;
        RECT -35.525 123.595 -35.195 123.925 ;
        RECT -35.525 122.235 -35.195 122.565 ;
        RECT -35.525 120.875 -35.195 121.205 ;
        RECT -35.525 119.515 -35.195 119.845 ;
        RECT -35.525 118.155 -35.195 118.485 ;
        RECT -35.525 116.795 -35.195 117.125 ;
        RECT -35.525 115.435 -35.195 115.765 ;
        RECT -35.525 114.075 -35.195 114.405 ;
        RECT -35.525 112.715 -35.195 113.045 ;
        RECT -35.525 111.355 -35.195 111.685 ;
        RECT -35.525 109.995 -35.195 110.325 ;
        RECT -35.525 108.635 -35.195 108.965 ;
        RECT -35.525 107.275 -35.195 107.605 ;
        RECT -35.525 105.915 -35.195 106.245 ;
        RECT -35.525 104.555 -35.195 104.885 ;
        RECT -35.525 103.195 -35.195 103.525 ;
        RECT -35.525 101.835 -35.195 102.165 ;
        RECT -35.525 100.475 -35.195 100.805 ;
        RECT -35.525 99.115 -35.195 99.445 ;
        RECT -35.525 97.755 -35.195 98.085 ;
        RECT -35.525 96.395 -35.195 96.725 ;
        RECT -35.525 95.035 -35.195 95.365 ;
        RECT -35.525 93.675 -35.195 94.005 ;
        RECT -35.525 92.315 -35.195 92.645 ;
        RECT -35.525 90.955 -35.195 91.285 ;
        RECT -35.525 89.595 -35.195 89.925 ;
        RECT -35.525 88.235 -35.195 88.565 ;
        RECT -35.525 86.875 -35.195 87.205 ;
        RECT -35.525 85.515 -35.195 85.845 ;
        RECT -35.525 84.155 -35.195 84.485 ;
        RECT -35.525 82.795 -35.195 83.125 ;
        RECT -35.525 81.435 -35.195 81.765 ;
        RECT -35.525 80.075 -35.195 80.405 ;
        RECT -35.525 78.715 -35.195 79.045 ;
        RECT -35.525 77.355 -35.195 77.685 ;
        RECT -35.525 75.995 -35.195 76.325 ;
        RECT -35.525 74.635 -35.195 74.965 ;
        RECT -35.525 73.275 -35.195 73.605 ;
        RECT -35.525 71.915 -35.195 72.245 ;
        RECT -35.525 70.555 -35.195 70.885 ;
        RECT -35.525 69.195 -35.195 69.525 ;
        RECT -35.525 67.835 -35.195 68.165 ;
        RECT -35.525 66.475 -35.195 66.805 ;
        RECT -35.525 65.115 -35.195 65.445 ;
        RECT -35.525 63.755 -35.195 64.085 ;
        RECT -35.525 62.395 -35.195 62.725 ;
        RECT -35.525 61.035 -35.195 61.365 ;
        RECT -35.525 59.675 -35.195 60.005 ;
        RECT -35.525 58.315 -35.195 58.645 ;
        RECT -35.525 56.955 -35.195 57.285 ;
        RECT -35.525 55.595 -35.195 55.925 ;
        RECT -35.525 54.235 -35.195 54.565 ;
        RECT -35.525 52.875 -35.195 53.205 ;
        RECT -35.525 51.515 -35.195 51.845 ;
        RECT -35.525 50.155 -35.195 50.485 ;
        RECT -35.525 48.795 -35.195 49.125 ;
        RECT -35.525 47.435 -35.195 47.765 ;
        RECT -35.525 46.075 -35.195 46.405 ;
        RECT -35.525 44.715 -35.195 45.045 ;
        RECT -35.525 43.355 -35.195 43.685 ;
        RECT -35.525 41.995 -35.195 42.325 ;
        RECT -35.525 40.635 -35.195 40.965 ;
        RECT -35.525 39.275 -35.195 39.605 ;
        RECT -35.525 37.915 -35.195 38.245 ;
        RECT -35.525 36.555 -35.195 36.885 ;
        RECT -35.525 35.195 -35.195 35.525 ;
        RECT -35.525 33.835 -35.195 34.165 ;
        RECT -35.525 32.475 -35.195 32.805 ;
        RECT -35.525 31.115 -35.195 31.445 ;
        RECT -35.525 29.755 -35.195 30.085 ;
        RECT -35.525 28.395 -35.195 28.725 ;
        RECT -35.525 27.035 -35.195 27.365 ;
        RECT -35.525 25.675 -35.195 26.005 ;
        RECT -35.525 24.315 -35.195 24.645 ;
        RECT -35.525 22.955 -35.195 23.285 ;
        RECT -35.525 21.595 -35.195 21.925 ;
        RECT -35.525 20.235 -35.195 20.565 ;
        RECT -35.525 18.875 -35.195 19.205 ;
        RECT -35.525 17.515 -35.195 17.845 ;
        RECT -35.525 16.155 -35.195 16.485 ;
        RECT -35.525 14.795 -35.195 15.125 ;
        RECT -35.525 13.435 -35.195 13.765 ;
        RECT -35.525 12.075 -35.195 12.405 ;
        RECT -35.525 10.715 -35.195 11.045 ;
        RECT -35.525 9.355 -35.195 9.685 ;
        RECT -35.525 7.995 -35.195 8.325 ;
        RECT -35.525 6.635 -35.195 6.965 ;
        RECT -35.525 5.275 -35.195 5.605 ;
        RECT -35.525 3.915 -35.195 4.245 ;
        RECT -35.525 2.555 -35.195 2.885 ;
        RECT -35.525 1.195 -35.195 1.525 ;
        RECT -35.525 -0.165 -35.195 0.165 ;
        RECT -35.525 -8.325 -35.195 -7.995 ;
        RECT -35.525 -12.405 -35.195 -12.075 ;
        RECT -35.525 -13.765 -35.195 -13.435 ;
        RECT -35.525 -15.125 -35.195 -14.795 ;
        RECT -35.525 -16.485 -35.195 -16.155 ;
        RECT -35.525 -17.845 -35.195 -17.515 ;
        RECT -35.525 -19.205 -35.195 -18.875 ;
        RECT -35.525 -20.565 -35.195 -20.235 ;
        RECT -35.525 -21.925 -35.195 -21.595 ;
        RECT -35.525 -28.725 -35.195 -28.395 ;
        RECT -35.525 -30.085 -35.195 -29.755 ;
        RECT -35.525 -31.445 -35.195 -31.115 ;
        RECT -35.525 -32.805 -35.195 -32.475 ;
        RECT -35.525 -34.165 -35.195 -33.835 ;
        RECT -35.525 -35.525 -35.195 -35.195 ;
        RECT -35.525 -36.885 -35.195 -36.555 ;
        RECT -35.525 -38.245 -35.195 -37.915 ;
        RECT -35.525 -39.605 -35.195 -39.275 ;
        RECT -35.525 -40.965 -35.195 -40.635 ;
        RECT -35.525 -42.325 -35.195 -41.995 ;
        RECT -35.525 -43.685 -35.195 -43.355 ;
        RECT -35.525 -45.045 -35.195 -44.715 ;
        RECT -35.525 -47.765 -35.195 -47.435 ;
        RECT -35.525 -49.125 -35.195 -48.795 ;
        RECT -35.525 -50.485 -35.195 -50.155 ;
        RECT -35.525 -51.845 -35.195 -51.515 ;
        RECT -35.525 -53.205 -35.195 -52.875 ;
        RECT -35.525 -54.565 -35.195 -54.235 ;
        RECT -35.525 -55.925 -35.195 -55.595 ;
        RECT -35.525 -57.285 -35.195 -56.955 ;
        RECT -35.525 -58.645 -35.195 -58.315 ;
        RECT -35.525 -60.005 -35.195 -59.675 ;
        RECT -35.525 -61.365 -35.195 -61.035 ;
        RECT -35.525 -62.725 -35.195 -62.395 ;
        RECT -35.525 -64.085 -35.195 -63.755 ;
        RECT -35.525 -65.445 -35.195 -65.115 ;
        RECT -35.525 -66.805 -35.195 -66.475 ;
        RECT -35.525 -68.165 -35.195 -67.835 ;
        RECT -35.525 -69.525 -35.195 -69.195 ;
        RECT -35.525 -72.245 -35.195 -71.915 ;
        RECT -35.525 -73.605 -35.195 -73.275 ;
        RECT -35.525 -74.965 -35.195 -74.635 ;
        RECT -35.525 -76.325 -35.195 -75.995 ;
        RECT -35.525 -78.29 -35.195 -77.96 ;
        RECT -35.525 -79.045 -35.195 -78.715 ;
        RECT -35.525 -81.765 -35.195 -81.435 ;
        RECT -35.525 -83.125 -35.195 -82.795 ;
        RECT -35.525 -84.485 -35.195 -84.155 ;
        RECT -35.525 -86.43 -35.195 -86.1 ;
        RECT -35.525 -87.205 -35.195 -86.875 ;
        RECT -35.525 -88.565 -35.195 -88.235 ;
        RECT -35.525 -89.925 -35.195 -89.595 ;
        RECT -35.52 -91.28 -35.2 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 -153.845 -35.195 -153.515 ;
        RECT -35.525 -155.285 -35.195 -154.955 ;
        RECT -35.525 -156.565 -35.195 -156.235 ;
        RECT -35.525 -157.925 -35.195 -157.595 ;
        RECT -35.525 -160.17 -35.195 -159.04 ;
        RECT -35.52 -160.285 -35.2 -152.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.165 127.225 -33.835 128.355 ;
        RECT -34.165 124.955 -33.835 125.285 ;
        RECT -34.165 123.595 -33.835 123.925 ;
        RECT -34.165 122.235 -33.835 122.565 ;
        RECT -34.165 120.875 -33.835 121.205 ;
        RECT -34.165 119.515 -33.835 119.845 ;
        RECT -34.165 118.155 -33.835 118.485 ;
        RECT -34.165 116.795 -33.835 117.125 ;
        RECT -34.165 115.435 -33.835 115.765 ;
        RECT -34.165 114.075 -33.835 114.405 ;
        RECT -34.165 112.715 -33.835 113.045 ;
        RECT -34.165 111.355 -33.835 111.685 ;
        RECT -34.165 109.995 -33.835 110.325 ;
        RECT -34.165 108.635 -33.835 108.965 ;
        RECT -34.165 107.275 -33.835 107.605 ;
        RECT -34.165 105.915 -33.835 106.245 ;
        RECT -34.165 104.555 -33.835 104.885 ;
        RECT -34.165 103.195 -33.835 103.525 ;
        RECT -34.165 101.835 -33.835 102.165 ;
        RECT -34.165 100.475 -33.835 100.805 ;
        RECT -34.165 99.115 -33.835 99.445 ;
        RECT -34.165 97.755 -33.835 98.085 ;
        RECT -34.165 96.395 -33.835 96.725 ;
        RECT -34.165 95.035 -33.835 95.365 ;
        RECT -34.165 93.675 -33.835 94.005 ;
        RECT -34.165 92.315 -33.835 92.645 ;
        RECT -34.165 90.955 -33.835 91.285 ;
        RECT -34.165 89.595 -33.835 89.925 ;
        RECT -34.165 88.235 -33.835 88.565 ;
        RECT -34.165 86.875 -33.835 87.205 ;
        RECT -34.165 85.515 -33.835 85.845 ;
        RECT -34.165 84.155 -33.835 84.485 ;
        RECT -34.165 82.795 -33.835 83.125 ;
        RECT -34.165 81.435 -33.835 81.765 ;
        RECT -34.165 80.075 -33.835 80.405 ;
        RECT -34.165 78.715 -33.835 79.045 ;
        RECT -34.165 77.355 -33.835 77.685 ;
        RECT -34.165 75.995 -33.835 76.325 ;
        RECT -34.165 74.635 -33.835 74.965 ;
        RECT -34.165 73.275 -33.835 73.605 ;
        RECT -34.165 71.915 -33.835 72.245 ;
        RECT -34.165 70.555 -33.835 70.885 ;
        RECT -34.165 69.195 -33.835 69.525 ;
        RECT -34.165 67.835 -33.835 68.165 ;
        RECT -34.165 66.475 -33.835 66.805 ;
        RECT -34.165 65.115 -33.835 65.445 ;
        RECT -34.165 63.755 -33.835 64.085 ;
        RECT -34.165 62.395 -33.835 62.725 ;
        RECT -34.165 61.035 -33.835 61.365 ;
        RECT -34.165 59.675 -33.835 60.005 ;
        RECT -34.165 58.315 -33.835 58.645 ;
        RECT -34.165 56.955 -33.835 57.285 ;
        RECT -34.165 55.595 -33.835 55.925 ;
        RECT -34.165 54.235 -33.835 54.565 ;
        RECT -34.165 52.875 -33.835 53.205 ;
        RECT -34.165 51.515 -33.835 51.845 ;
        RECT -34.165 50.155 -33.835 50.485 ;
        RECT -34.165 48.795 -33.835 49.125 ;
        RECT -34.165 47.435 -33.835 47.765 ;
        RECT -34.165 46.075 -33.835 46.405 ;
        RECT -34.165 44.715 -33.835 45.045 ;
        RECT -34.165 43.355 -33.835 43.685 ;
        RECT -34.165 41.995 -33.835 42.325 ;
        RECT -34.165 40.635 -33.835 40.965 ;
        RECT -34.165 39.275 -33.835 39.605 ;
        RECT -34.165 37.915 -33.835 38.245 ;
        RECT -34.165 36.555 -33.835 36.885 ;
        RECT -34.165 35.195 -33.835 35.525 ;
        RECT -34.165 33.835 -33.835 34.165 ;
        RECT -34.165 32.475 -33.835 32.805 ;
        RECT -34.165 31.115 -33.835 31.445 ;
        RECT -34.165 29.755 -33.835 30.085 ;
        RECT -34.165 28.395 -33.835 28.725 ;
        RECT -34.165 27.035 -33.835 27.365 ;
        RECT -34.165 25.675 -33.835 26.005 ;
        RECT -34.165 24.315 -33.835 24.645 ;
        RECT -34.165 22.955 -33.835 23.285 ;
        RECT -34.165 21.595 -33.835 21.925 ;
        RECT -34.165 20.235 -33.835 20.565 ;
        RECT -34.165 18.875 -33.835 19.205 ;
        RECT -34.165 17.515 -33.835 17.845 ;
        RECT -34.165 16.155 -33.835 16.485 ;
        RECT -34.165 14.795 -33.835 15.125 ;
        RECT -34.165 13.435 -33.835 13.765 ;
        RECT -34.165 12.075 -33.835 12.405 ;
        RECT -34.165 10.715 -33.835 11.045 ;
        RECT -34.165 9.355 -33.835 9.685 ;
        RECT -34.165 7.995 -33.835 8.325 ;
        RECT -34.165 6.635 -33.835 6.965 ;
        RECT -34.165 5.275 -33.835 5.605 ;
        RECT -34.165 3.915 -33.835 4.245 ;
        RECT -34.165 2.555 -33.835 2.885 ;
        RECT -34.165 1.195 -33.835 1.525 ;
        RECT -34.165 -0.165 -33.835 0.165 ;
        RECT -34.165 -8.325 -33.835 -7.995 ;
        RECT -34.165 -12.405 -33.835 -12.075 ;
        RECT -34.165 -13.765 -33.835 -13.435 ;
        RECT -34.165 -15.125 -33.835 -14.795 ;
        RECT -34.165 -16.485 -33.835 -16.155 ;
        RECT -34.165 -17.845 -33.835 -17.515 ;
        RECT -34.165 -19.205 -33.835 -18.875 ;
        RECT -34.165 -20.565 -33.835 -20.235 ;
        RECT -34.165 -21.925 -33.835 -21.595 ;
        RECT -34.165 -28.725 -33.835 -28.395 ;
        RECT -34.165 -30.085 -33.835 -29.755 ;
        RECT -34.165 -31.445 -33.835 -31.115 ;
        RECT -34.165 -32.805 -33.835 -32.475 ;
        RECT -34.165 -34.165 -33.835 -33.835 ;
        RECT -34.165 -35.525 -33.835 -35.195 ;
        RECT -34.165 -36.885 -33.835 -36.555 ;
        RECT -34.165 -38.245 -33.835 -37.915 ;
        RECT -34.165 -39.605 -33.835 -39.275 ;
        RECT -34.165 -40.965 -33.835 -40.635 ;
        RECT -34.165 -42.325 -33.835 -41.995 ;
        RECT -34.165 -43.685 -33.835 -43.355 ;
        RECT -34.165 -45.045 -33.835 -44.715 ;
        RECT -34.165 -49.125 -33.835 -48.795 ;
        RECT -34.165 -50.485 -33.835 -50.155 ;
        RECT -34.165 -51.845 -33.835 -51.515 ;
        RECT -34.165 -53.205 -33.835 -52.875 ;
        RECT -34.165 -54.565 -33.835 -54.235 ;
        RECT -34.165 -55.925 -33.835 -55.595 ;
        RECT -34.165 -57.285 -33.835 -56.955 ;
        RECT -34.165 -58.645 -33.835 -58.315 ;
        RECT -34.165 -60.005 -33.835 -59.675 ;
        RECT -34.165 -61.365 -33.835 -61.035 ;
        RECT -34.165 -62.725 -33.835 -62.395 ;
        RECT -34.165 -64.085 -33.835 -63.755 ;
        RECT -34.165 -65.445 -33.835 -65.115 ;
        RECT -34.165 -66.805 -33.835 -66.475 ;
        RECT -34.165 -68.165 -33.835 -67.835 ;
        RECT -34.165 -69.525 -33.835 -69.195 ;
        RECT -34.165 -72.245 -33.835 -71.915 ;
        RECT -34.165 -73.605 -33.835 -73.275 ;
        RECT -34.165 -74.965 -33.835 -74.635 ;
        RECT -34.165 -76.325 -33.835 -75.995 ;
        RECT -34.165 -78.29 -33.835 -77.96 ;
        RECT -34.165 -79.045 -33.835 -78.715 ;
        RECT -34.165 -81.765 -33.835 -81.435 ;
        RECT -34.165 -83.125 -33.835 -82.795 ;
        RECT -34.165 -84.485 -33.835 -84.155 ;
        RECT -34.165 -86.43 -33.835 -86.1 ;
        RECT -34.165 -87.205 -33.835 -86.875 ;
        RECT -34.165 -88.565 -33.835 -88.235 ;
        RECT -34.165 -89.925 -33.835 -89.595 ;
        RECT -34.16 -91.28 -33.84 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.165 -153.845 -33.835 -153.515 ;
        RECT -34.165 -155.285 -33.835 -154.955 ;
        RECT -34.165 -156.565 -33.835 -156.235 ;
        RECT -34.165 -157.925 -33.835 -157.595 ;
        RECT -34.165 -160.17 -33.835 -159.04 ;
        RECT -34.16 -160.285 -33.84 -153.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.805 127.225 -32.475 128.355 ;
        RECT -32.805 124.955 -32.475 125.285 ;
        RECT -32.805 123.595 -32.475 123.925 ;
        RECT -32.805 122.235 -32.475 122.565 ;
        RECT -32.805 120.875 -32.475 121.205 ;
        RECT -32.805 119.515 -32.475 119.845 ;
        RECT -32.805 118.155 -32.475 118.485 ;
        RECT -32.805 116.795 -32.475 117.125 ;
        RECT -32.805 115.435 -32.475 115.765 ;
        RECT -32.805 114.075 -32.475 114.405 ;
        RECT -32.805 112.715 -32.475 113.045 ;
        RECT -32.805 111.355 -32.475 111.685 ;
        RECT -32.805 109.995 -32.475 110.325 ;
        RECT -32.805 108.635 -32.475 108.965 ;
        RECT -32.805 107.275 -32.475 107.605 ;
        RECT -32.805 105.915 -32.475 106.245 ;
        RECT -32.805 104.555 -32.475 104.885 ;
        RECT -32.805 103.195 -32.475 103.525 ;
        RECT -32.805 101.835 -32.475 102.165 ;
        RECT -32.805 100.475 -32.475 100.805 ;
        RECT -32.805 99.115 -32.475 99.445 ;
        RECT -32.805 97.755 -32.475 98.085 ;
        RECT -32.805 96.395 -32.475 96.725 ;
        RECT -32.805 95.035 -32.475 95.365 ;
        RECT -32.805 93.675 -32.475 94.005 ;
        RECT -32.805 92.315 -32.475 92.645 ;
        RECT -32.805 90.955 -32.475 91.285 ;
        RECT -32.805 89.595 -32.475 89.925 ;
        RECT -32.805 88.235 -32.475 88.565 ;
        RECT -32.805 86.875 -32.475 87.205 ;
        RECT -32.805 85.515 -32.475 85.845 ;
        RECT -32.805 84.155 -32.475 84.485 ;
        RECT -32.805 82.795 -32.475 83.125 ;
        RECT -32.805 81.435 -32.475 81.765 ;
        RECT -32.805 80.075 -32.475 80.405 ;
        RECT -32.805 78.715 -32.475 79.045 ;
        RECT -32.805 77.355 -32.475 77.685 ;
        RECT -32.805 75.995 -32.475 76.325 ;
        RECT -32.805 74.635 -32.475 74.965 ;
        RECT -32.805 73.275 -32.475 73.605 ;
        RECT -32.805 71.915 -32.475 72.245 ;
        RECT -32.805 70.555 -32.475 70.885 ;
        RECT -32.805 69.195 -32.475 69.525 ;
        RECT -32.805 67.835 -32.475 68.165 ;
        RECT -32.805 66.475 -32.475 66.805 ;
        RECT -32.805 65.115 -32.475 65.445 ;
        RECT -32.805 63.755 -32.475 64.085 ;
        RECT -32.805 62.395 -32.475 62.725 ;
        RECT -32.805 61.035 -32.475 61.365 ;
        RECT -32.805 59.675 -32.475 60.005 ;
        RECT -32.805 58.315 -32.475 58.645 ;
        RECT -32.805 56.955 -32.475 57.285 ;
        RECT -32.805 55.595 -32.475 55.925 ;
        RECT -32.805 54.235 -32.475 54.565 ;
        RECT -32.805 52.875 -32.475 53.205 ;
        RECT -32.805 51.515 -32.475 51.845 ;
        RECT -32.805 50.155 -32.475 50.485 ;
        RECT -32.805 48.795 -32.475 49.125 ;
        RECT -32.805 47.435 -32.475 47.765 ;
        RECT -32.805 46.075 -32.475 46.405 ;
        RECT -32.805 44.715 -32.475 45.045 ;
        RECT -32.805 43.355 -32.475 43.685 ;
        RECT -32.805 41.995 -32.475 42.325 ;
        RECT -32.805 40.635 -32.475 40.965 ;
        RECT -32.805 39.275 -32.475 39.605 ;
        RECT -32.805 37.915 -32.475 38.245 ;
        RECT -32.805 36.555 -32.475 36.885 ;
        RECT -32.805 35.195 -32.475 35.525 ;
        RECT -32.805 33.835 -32.475 34.165 ;
        RECT -32.805 32.475 -32.475 32.805 ;
        RECT -32.805 31.115 -32.475 31.445 ;
        RECT -32.805 29.755 -32.475 30.085 ;
        RECT -32.805 28.395 -32.475 28.725 ;
        RECT -32.805 27.035 -32.475 27.365 ;
        RECT -32.805 25.675 -32.475 26.005 ;
        RECT -32.805 24.315 -32.475 24.645 ;
        RECT -32.805 22.955 -32.475 23.285 ;
        RECT -32.805 21.595 -32.475 21.925 ;
        RECT -32.805 20.235 -32.475 20.565 ;
        RECT -32.805 18.875 -32.475 19.205 ;
        RECT -32.805 17.515 -32.475 17.845 ;
        RECT -32.805 16.155 -32.475 16.485 ;
        RECT -32.805 14.795 -32.475 15.125 ;
        RECT -32.805 13.435 -32.475 13.765 ;
        RECT -32.805 12.075 -32.475 12.405 ;
        RECT -32.805 10.715 -32.475 11.045 ;
        RECT -32.805 9.355 -32.475 9.685 ;
        RECT -32.805 7.995 -32.475 8.325 ;
        RECT -32.805 6.635 -32.475 6.965 ;
        RECT -32.805 5.275 -32.475 5.605 ;
        RECT -32.805 3.915 -32.475 4.245 ;
        RECT -32.805 2.555 -32.475 2.885 ;
        RECT -32.805 1.195 -32.475 1.525 ;
        RECT -32.805 -0.165 -32.475 0.165 ;
        RECT -32.805 -8.325 -32.475 -7.995 ;
        RECT -32.805 -12.405 -32.475 -12.075 ;
        RECT -32.805 -13.765 -32.475 -13.435 ;
        RECT -32.805 -15.125 -32.475 -14.795 ;
        RECT -32.805 -16.485 -32.475 -16.155 ;
        RECT -32.805 -17.845 -32.475 -17.515 ;
        RECT -32.805 -19.205 -32.475 -18.875 ;
        RECT -32.805 -20.565 -32.475 -20.235 ;
        RECT -32.805 -21.925 -32.475 -21.595 ;
        RECT -32.805 -28.725 -32.475 -28.395 ;
        RECT -32.805 -30.085 -32.475 -29.755 ;
        RECT -32.805 -31.445 -32.475 -31.115 ;
        RECT -32.805 -32.805 -32.475 -32.475 ;
        RECT -32.805 -34.165 -32.475 -33.835 ;
        RECT -32.805 -35.525 -32.475 -35.195 ;
        RECT -32.805 -36.885 -32.475 -36.555 ;
        RECT -32.805 -38.245 -32.475 -37.915 ;
        RECT -32.805 -39.605 -32.475 -39.275 ;
        RECT -32.805 -40.965 -32.475 -40.635 ;
        RECT -32.805 -42.325 -32.475 -41.995 ;
        RECT -32.805 -43.685 -32.475 -43.355 ;
        RECT -32.805 -45.045 -32.475 -44.715 ;
        RECT -32.805 -49.125 -32.475 -48.795 ;
        RECT -32.805 -50.485 -32.475 -50.155 ;
        RECT -32.805 -51.845 -32.475 -51.515 ;
        RECT -32.805 -53.205 -32.475 -52.875 ;
        RECT -32.805 -54.565 -32.475 -54.235 ;
        RECT -32.805 -55.925 -32.475 -55.595 ;
        RECT -32.805 -57.285 -32.475 -56.955 ;
        RECT -32.805 -58.645 -32.475 -58.315 ;
        RECT -32.805 -60.005 -32.475 -59.675 ;
        RECT -32.805 -61.365 -32.475 -61.035 ;
        RECT -32.805 -62.725 -32.475 -62.395 ;
        RECT -32.805 -64.085 -32.475 -63.755 ;
        RECT -32.805 -65.445 -32.475 -65.115 ;
        RECT -32.805 -66.805 -32.475 -66.475 ;
        RECT -32.805 -68.165 -32.475 -67.835 ;
        RECT -32.805 -69.525 -32.475 -69.195 ;
        RECT -32.805 -72.245 -32.475 -71.915 ;
        RECT -32.805 -73.605 -32.475 -73.275 ;
        RECT -32.805 -74.965 -32.475 -74.635 ;
        RECT -32.805 -76.325 -32.475 -75.995 ;
        RECT -32.805 -78.29 -32.475 -77.96 ;
        RECT -32.805 -79.045 -32.475 -78.715 ;
        RECT -32.805 -81.765 -32.475 -81.435 ;
        RECT -32.805 -83.125 -32.475 -82.795 ;
        RECT -32.805 -84.485 -32.475 -84.155 ;
        RECT -32.805 -86.43 -32.475 -86.1 ;
        RECT -32.805 -87.205 -32.475 -86.875 ;
        RECT -32.805 -88.565 -32.475 -88.235 ;
        RECT -32.805 -89.925 -32.475 -89.595 ;
        RECT -32.805 -92.645 -32.475 -92.315 ;
        RECT -32.805 -94.005 -32.475 -93.675 ;
        RECT -32.805 -95.365 -32.475 -95.035 ;
        RECT -32.805 -96.725 -32.475 -96.395 ;
        RECT -32.805 -98.085 -32.475 -97.755 ;
        RECT -32.805 -102.165 -32.475 -101.835 ;
        RECT -32.805 -104.885 -32.475 -104.555 ;
        RECT -32.805 -106.245 -32.475 -105.915 ;
        RECT -32.805 -107.605 -32.475 -107.275 ;
        RECT -32.805 -108.965 -32.475 -108.635 ;
        RECT -32.805 -113.045 -32.475 -112.715 ;
        RECT -32.805 -114.405 -32.475 -114.075 ;
        RECT -32.805 -115.765 -32.475 -115.435 ;
        RECT -32.805 -117.125 -32.475 -116.795 ;
        RECT -32.805 -118.485 -32.475 -118.155 ;
        RECT -32.805 -121.205 -32.475 -120.875 ;
        RECT -32.805 -122.565 -32.475 -122.235 ;
        RECT -32.805 -123.925 -32.475 -123.595 ;
        RECT -32.805 -125.285 -32.475 -124.955 ;
        RECT -32.805 -126.645 -32.475 -126.315 ;
        RECT -32.805 -128.005 -32.475 -127.675 ;
        RECT -32.805 -130.725 -32.475 -130.395 ;
        RECT -32.805 -132.085 -32.475 -131.755 ;
        RECT -32.805 -136.165 -32.475 -135.835 ;
        RECT -32.805 -137.525 -32.475 -137.195 ;
        RECT -32.805 -138.885 -32.475 -138.555 ;
        RECT -32.805 -140.245 -32.475 -139.915 ;
        RECT -32.805 -141.605 -32.475 -141.275 ;
        RECT -32.805 -142.965 -32.475 -142.635 ;
        RECT -32.805 -144.325 -32.475 -143.995 ;
        RECT -32.805 -145.685 -32.475 -145.355 ;
        RECT -32.805 -147.045 -32.475 -146.715 ;
        RECT -32.805 -149.765 -32.475 -149.435 ;
        RECT -32.805 -152.485 -32.475 -152.155 ;
        RECT -32.805 -153.845 -32.475 -153.515 ;
        RECT -32.805 -155.285 -32.475 -154.955 ;
        RECT -32.805 -156.565 -32.475 -156.235 ;
        RECT -32.805 -157.925 -32.475 -157.595 ;
        RECT -32.805 -160.17 -32.475 -159.04 ;
        RECT -32.8 -160.285 -32.48 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.445 127.225 -31.115 128.355 ;
        RECT -31.445 124.955 -31.115 125.285 ;
        RECT -31.445 123.595 -31.115 123.925 ;
        RECT -31.445 122.235 -31.115 122.565 ;
        RECT -31.445 120.875 -31.115 121.205 ;
        RECT -31.445 119.515 -31.115 119.845 ;
        RECT -31.445 118.155 -31.115 118.485 ;
        RECT -31.445 116.795 -31.115 117.125 ;
        RECT -31.445 115.435 -31.115 115.765 ;
        RECT -31.445 114.075 -31.115 114.405 ;
        RECT -31.445 112.715 -31.115 113.045 ;
        RECT -31.445 111.355 -31.115 111.685 ;
        RECT -31.445 109.995 -31.115 110.325 ;
        RECT -31.445 108.635 -31.115 108.965 ;
        RECT -31.445 107.275 -31.115 107.605 ;
        RECT -31.445 105.915 -31.115 106.245 ;
        RECT -31.445 104.555 -31.115 104.885 ;
        RECT -31.445 103.195 -31.115 103.525 ;
        RECT -31.445 101.835 -31.115 102.165 ;
        RECT -31.445 100.475 -31.115 100.805 ;
        RECT -31.445 99.115 -31.115 99.445 ;
        RECT -31.445 97.755 -31.115 98.085 ;
        RECT -31.445 96.395 -31.115 96.725 ;
        RECT -31.445 95.035 -31.115 95.365 ;
        RECT -31.445 93.675 -31.115 94.005 ;
        RECT -31.445 92.315 -31.115 92.645 ;
        RECT -31.445 90.955 -31.115 91.285 ;
        RECT -31.445 89.595 -31.115 89.925 ;
        RECT -31.445 88.235 -31.115 88.565 ;
        RECT -31.445 86.875 -31.115 87.205 ;
        RECT -31.445 85.515 -31.115 85.845 ;
        RECT -31.445 84.155 -31.115 84.485 ;
        RECT -31.445 82.795 -31.115 83.125 ;
        RECT -31.445 81.435 -31.115 81.765 ;
        RECT -31.445 80.075 -31.115 80.405 ;
        RECT -31.445 78.715 -31.115 79.045 ;
        RECT -31.445 77.355 -31.115 77.685 ;
        RECT -31.445 75.995 -31.115 76.325 ;
        RECT -31.445 74.635 -31.115 74.965 ;
        RECT -31.445 73.275 -31.115 73.605 ;
        RECT -31.445 71.915 -31.115 72.245 ;
        RECT -31.445 70.555 -31.115 70.885 ;
        RECT -31.445 69.195 -31.115 69.525 ;
        RECT -31.445 67.835 -31.115 68.165 ;
        RECT -31.445 66.475 -31.115 66.805 ;
        RECT -31.445 65.115 -31.115 65.445 ;
        RECT -31.445 63.755 -31.115 64.085 ;
        RECT -31.445 62.395 -31.115 62.725 ;
        RECT -31.445 61.035 -31.115 61.365 ;
        RECT -31.445 59.675 -31.115 60.005 ;
        RECT -31.445 58.315 -31.115 58.645 ;
        RECT -31.445 56.955 -31.115 57.285 ;
        RECT -31.445 55.595 -31.115 55.925 ;
        RECT -31.445 54.235 -31.115 54.565 ;
        RECT -31.445 52.875 -31.115 53.205 ;
        RECT -31.445 51.515 -31.115 51.845 ;
        RECT -31.445 50.155 -31.115 50.485 ;
        RECT -31.445 48.795 -31.115 49.125 ;
        RECT -31.445 47.435 -31.115 47.765 ;
        RECT -31.445 46.075 -31.115 46.405 ;
        RECT -31.445 44.715 -31.115 45.045 ;
        RECT -31.445 43.355 -31.115 43.685 ;
        RECT -31.445 41.995 -31.115 42.325 ;
        RECT -31.445 40.635 -31.115 40.965 ;
        RECT -31.445 39.275 -31.115 39.605 ;
        RECT -31.445 37.915 -31.115 38.245 ;
        RECT -31.445 36.555 -31.115 36.885 ;
        RECT -31.445 35.195 -31.115 35.525 ;
        RECT -31.445 33.835 -31.115 34.165 ;
        RECT -31.445 32.475 -31.115 32.805 ;
        RECT -31.445 31.115 -31.115 31.445 ;
        RECT -31.445 29.755 -31.115 30.085 ;
        RECT -31.445 28.395 -31.115 28.725 ;
        RECT -31.445 27.035 -31.115 27.365 ;
        RECT -31.445 25.675 -31.115 26.005 ;
        RECT -31.445 24.315 -31.115 24.645 ;
        RECT -31.445 22.955 -31.115 23.285 ;
        RECT -31.445 21.595 -31.115 21.925 ;
        RECT -31.445 20.235 -31.115 20.565 ;
        RECT -31.445 18.875 -31.115 19.205 ;
        RECT -31.445 17.515 -31.115 17.845 ;
        RECT -31.445 16.155 -31.115 16.485 ;
        RECT -31.445 14.795 -31.115 15.125 ;
        RECT -31.445 13.435 -31.115 13.765 ;
        RECT -31.445 12.075 -31.115 12.405 ;
        RECT -31.445 10.715 -31.115 11.045 ;
        RECT -31.445 9.355 -31.115 9.685 ;
        RECT -31.445 7.995 -31.115 8.325 ;
        RECT -31.445 6.635 -31.115 6.965 ;
        RECT -31.445 5.275 -31.115 5.605 ;
        RECT -31.445 3.915 -31.115 4.245 ;
        RECT -31.445 2.555 -31.115 2.885 ;
        RECT -31.445 1.195 -31.115 1.525 ;
        RECT -31.445 -0.165 -31.115 0.165 ;
        RECT -31.445 -8.325 -31.115 -7.995 ;
        RECT -31.445 -12.405 -31.115 -12.075 ;
        RECT -31.445 -13.765 -31.115 -13.435 ;
        RECT -31.445 -15.125 -31.115 -14.795 ;
        RECT -31.445 -16.485 -31.115 -16.155 ;
        RECT -31.445 -17.845 -31.115 -17.515 ;
        RECT -31.445 -19.205 -31.115 -18.875 ;
        RECT -31.445 -20.565 -31.115 -20.235 ;
        RECT -31.445 -21.925 -31.115 -21.595 ;
        RECT -31.445 -28.725 -31.115 -28.395 ;
        RECT -31.445 -30.085 -31.115 -29.755 ;
        RECT -31.445 -31.445 -31.115 -31.115 ;
        RECT -31.445 -32.805 -31.115 -32.475 ;
        RECT -31.445 -34.165 -31.115 -33.835 ;
        RECT -31.445 -35.525 -31.115 -35.195 ;
        RECT -31.445 -36.885 -31.115 -36.555 ;
        RECT -31.445 -38.245 -31.115 -37.915 ;
        RECT -31.445 -39.605 -31.115 -39.275 ;
        RECT -31.445 -40.965 -31.115 -40.635 ;
        RECT -31.445 -42.325 -31.115 -41.995 ;
        RECT -31.445 -43.685 -31.115 -43.355 ;
        RECT -31.445 -45.045 -31.115 -44.715 ;
        RECT -31.445 -49.125 -31.115 -48.795 ;
        RECT -31.445 -50.485 -31.115 -50.155 ;
        RECT -31.445 -51.845 -31.115 -51.515 ;
        RECT -31.445 -53.205 -31.115 -52.875 ;
        RECT -31.445 -54.565 -31.115 -54.235 ;
        RECT -31.445 -55.925 -31.115 -55.595 ;
        RECT -31.445 -57.285 -31.115 -56.955 ;
        RECT -31.445 -58.645 -31.115 -58.315 ;
        RECT -31.445 -60.005 -31.115 -59.675 ;
        RECT -31.445 -61.365 -31.115 -61.035 ;
        RECT -31.445 -62.725 -31.115 -62.395 ;
        RECT -31.445 -64.085 -31.115 -63.755 ;
        RECT -31.445 -65.445 -31.115 -65.115 ;
        RECT -31.445 -66.805 -31.115 -66.475 ;
        RECT -31.445 -68.165 -31.115 -67.835 ;
        RECT -31.445 -69.525 -31.115 -69.195 ;
        RECT -31.445 -72.245 -31.115 -71.915 ;
        RECT -31.445 -73.605 -31.115 -73.275 ;
        RECT -31.445 -74.965 -31.115 -74.635 ;
        RECT -31.445 -76.325 -31.115 -75.995 ;
        RECT -31.445 -78.29 -31.115 -77.96 ;
        RECT -31.445 -79.045 -31.115 -78.715 ;
        RECT -31.445 -81.765 -31.115 -81.435 ;
        RECT -31.445 -83.125 -31.115 -82.795 ;
        RECT -31.445 -84.485 -31.115 -84.155 ;
        RECT -31.445 -86.43 -31.115 -86.1 ;
        RECT -31.445 -87.205 -31.115 -86.875 ;
        RECT -31.445 -88.565 -31.115 -88.235 ;
        RECT -31.445 -89.925 -31.115 -89.595 ;
        RECT -31.445 -92.645 -31.115 -92.315 ;
        RECT -31.445 -94.005 -31.115 -93.675 ;
        RECT -31.445 -95.365 -31.115 -95.035 ;
        RECT -31.445 -96.725 -31.115 -96.395 ;
        RECT -31.445 -98.085 -31.115 -97.755 ;
        RECT -31.445 -102.165 -31.115 -101.835 ;
        RECT -31.445 -104.885 -31.115 -104.555 ;
        RECT -31.445 -106.245 -31.115 -105.915 ;
        RECT -31.445 -107.605 -31.115 -107.275 ;
        RECT -31.445 -108.965 -31.115 -108.635 ;
        RECT -31.445 -113.045 -31.115 -112.715 ;
        RECT -31.445 -114.405 -31.115 -114.075 ;
        RECT -31.445 -115.765 -31.115 -115.435 ;
        RECT -31.445 -118.485 -31.115 -118.155 ;
        RECT -31.445 -121.205 -31.115 -120.875 ;
        RECT -31.445 -122.565 -31.115 -122.235 ;
        RECT -31.445 -123.925 -31.115 -123.595 ;
        RECT -31.445 -125.285 -31.115 -124.955 ;
        RECT -31.445 -126.645 -31.115 -126.315 ;
        RECT -31.445 -128.005 -31.115 -127.675 ;
        RECT -31.445 -130.725 -31.115 -130.395 ;
        RECT -31.445 -132.085 -31.115 -131.755 ;
        RECT -31.445 -136.165 -31.115 -135.835 ;
        RECT -31.445 -137.525 -31.115 -137.195 ;
        RECT -31.445 -138.885 -31.115 -138.555 ;
        RECT -31.445 -140.245 -31.115 -139.915 ;
        RECT -31.445 -141.605 -31.115 -141.275 ;
        RECT -31.445 -142.965 -31.115 -142.635 ;
        RECT -31.445 -144.325 -31.115 -143.995 ;
        RECT -31.445 -145.685 -31.115 -145.355 ;
        RECT -31.445 -147.045 -31.115 -146.715 ;
        RECT -31.445 -149.765 -31.115 -149.435 ;
        RECT -31.445 -152.485 -31.115 -152.155 ;
        RECT -31.445 -153.845 -31.115 -153.515 ;
        RECT -31.445 -155.285 -31.115 -154.955 ;
        RECT -31.445 -156.565 -31.115 -156.235 ;
        RECT -31.445 -157.925 -31.115 -157.595 ;
        RECT -31.445 -160.17 -31.115 -159.04 ;
        RECT -31.44 -160.285 -31.12 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 77.355 -29.755 77.685 ;
        RECT -30.085 75.995 -29.755 76.325 ;
        RECT -30.085 74.635 -29.755 74.965 ;
        RECT -30.085 73.275 -29.755 73.605 ;
        RECT -30.085 71.915 -29.755 72.245 ;
        RECT -30.085 70.555 -29.755 70.885 ;
        RECT -30.085 69.195 -29.755 69.525 ;
        RECT -30.085 67.835 -29.755 68.165 ;
        RECT -30.085 66.475 -29.755 66.805 ;
        RECT -30.085 65.115 -29.755 65.445 ;
        RECT -30.085 63.755 -29.755 64.085 ;
        RECT -30.085 62.395 -29.755 62.725 ;
        RECT -30.085 61.035 -29.755 61.365 ;
        RECT -30.085 59.675 -29.755 60.005 ;
        RECT -30.085 58.315 -29.755 58.645 ;
        RECT -30.085 56.955 -29.755 57.285 ;
        RECT -30.085 55.595 -29.755 55.925 ;
        RECT -30.085 54.235 -29.755 54.565 ;
        RECT -30.085 52.875 -29.755 53.205 ;
        RECT -30.085 51.515 -29.755 51.845 ;
        RECT -30.085 50.155 -29.755 50.485 ;
        RECT -30.085 48.795 -29.755 49.125 ;
        RECT -30.085 47.435 -29.755 47.765 ;
        RECT -30.085 46.075 -29.755 46.405 ;
        RECT -30.085 44.715 -29.755 45.045 ;
        RECT -30.085 43.355 -29.755 43.685 ;
        RECT -30.085 41.995 -29.755 42.325 ;
        RECT -30.085 40.635 -29.755 40.965 ;
        RECT -30.085 39.275 -29.755 39.605 ;
        RECT -30.085 37.915 -29.755 38.245 ;
        RECT -30.085 36.555 -29.755 36.885 ;
        RECT -30.085 35.195 -29.755 35.525 ;
        RECT -30.085 33.835 -29.755 34.165 ;
        RECT -30.085 32.475 -29.755 32.805 ;
        RECT -30.085 31.115 -29.755 31.445 ;
        RECT -30.085 29.755 -29.755 30.085 ;
        RECT -30.085 28.395 -29.755 28.725 ;
        RECT -30.085 27.035 -29.755 27.365 ;
        RECT -30.085 25.675 -29.755 26.005 ;
        RECT -30.085 24.315 -29.755 24.645 ;
        RECT -30.085 22.955 -29.755 23.285 ;
        RECT -30.085 21.595 -29.755 21.925 ;
        RECT -30.085 20.235 -29.755 20.565 ;
        RECT -30.085 18.875 -29.755 19.205 ;
        RECT -30.085 17.515 -29.755 17.845 ;
        RECT -30.085 16.155 -29.755 16.485 ;
        RECT -30.085 14.795 -29.755 15.125 ;
        RECT -30.085 13.435 -29.755 13.765 ;
        RECT -30.085 12.075 -29.755 12.405 ;
        RECT -30.085 10.715 -29.755 11.045 ;
        RECT -30.085 9.355 -29.755 9.685 ;
        RECT -30.085 7.995 -29.755 8.325 ;
        RECT -30.085 6.635 -29.755 6.965 ;
        RECT -30.085 5.275 -29.755 5.605 ;
        RECT -30.085 3.915 -29.755 4.245 ;
        RECT -30.085 2.555 -29.755 2.885 ;
        RECT -30.085 1.195 -29.755 1.525 ;
        RECT -30.085 -0.165 -29.755 0.165 ;
        RECT -30.085 -15.125 -29.755 -14.795 ;
        RECT -30.085 -16.485 -29.755 -16.155 ;
        RECT -30.085 -19.205 -29.755 -18.875 ;
        RECT -30.085 -28.725 -29.755 -28.395 ;
        RECT -30.085 -30.085 -29.755 -29.755 ;
        RECT -30.085 -32.805 -29.755 -32.475 ;
        RECT -30.085 -34.165 -29.755 -33.835 ;
        RECT -30.085 -38.245 -29.755 -37.915 ;
        RECT -30.085 -40.965 -29.755 -40.635 ;
        RECT -30.085 -50.485 -29.755 -50.155 ;
        RECT -30.085 -51.845 -29.755 -51.515 ;
        RECT -30.085 -53.205 -29.755 -52.875 ;
        RECT -30.085 -54.565 -29.755 -54.235 ;
        RECT -30.085 -55.925 -29.755 -55.595 ;
        RECT -30.085 -57.285 -29.755 -56.955 ;
        RECT -30.085 -58.645 -29.755 -58.315 ;
        RECT -30.085 -60.005 -29.755 -59.675 ;
        RECT -30.085 -61.365 -29.755 -61.035 ;
        RECT -30.085 -62.725 -29.755 -62.395 ;
        RECT -30.085 -64.085 -29.755 -63.755 ;
        RECT -30.085 -65.445 -29.755 -65.115 ;
        RECT -30.085 -66.805 -29.755 -66.475 ;
        RECT -30.085 -68.165 -29.755 -67.835 ;
        RECT -30.085 -69.525 -29.755 -69.195 ;
        RECT -30.085 -72.245 -29.755 -71.915 ;
        RECT -30.085 -73.605 -29.755 -73.275 ;
        RECT -30.085 -74.965 -29.755 -74.635 ;
        RECT -30.085 -76.325 -29.755 -75.995 ;
        RECT -30.085 -78.29 -29.755 -77.96 ;
        RECT -30.085 -79.045 -29.755 -78.715 ;
        RECT -30.085 -81.765 -29.755 -81.435 ;
        RECT -30.085 -83.125 -29.755 -82.795 ;
        RECT -30.085 -84.485 -29.755 -84.155 ;
        RECT -30.085 -86.43 -29.755 -86.1 ;
        RECT -30.085 -87.205 -29.755 -86.875 ;
        RECT -30.085 -88.565 -29.755 -88.235 ;
        RECT -30.085 -89.925 -29.755 -89.595 ;
        RECT -30.085 -92.645 -29.755 -92.315 ;
        RECT -30.085 -94.005 -29.755 -93.675 ;
        RECT -30.085 -95.365 -29.755 -95.035 ;
        RECT -30.085 -96.725 -29.755 -96.395 ;
        RECT -30.085 -98.085 -29.755 -97.755 ;
        RECT -30.085 -102.165 -29.755 -101.835 ;
        RECT -30.085 -104.885 -29.755 -104.555 ;
        RECT -30.085 -106.245 -29.755 -105.915 ;
        RECT -30.085 -107.605 -29.755 -107.275 ;
        RECT -30.085 -108.965 -29.755 -108.635 ;
        RECT -30.085 -113.045 -29.755 -112.715 ;
        RECT -30.085 -114.405 -29.755 -114.075 ;
        RECT -30.085 -115.765 -29.755 -115.435 ;
        RECT -30.085 -118.485 -29.755 -118.155 ;
        RECT -30.085 -121.205 -29.755 -120.875 ;
        RECT -30.085 -122.565 -29.755 -122.235 ;
        RECT -30.085 -123.925 -29.755 -123.595 ;
        RECT -30.085 -125.285 -29.755 -124.955 ;
        RECT -30.085 -126.645 -29.755 -126.315 ;
        RECT -30.085 -128.005 -29.755 -127.675 ;
        RECT -30.085 -130.725 -29.755 -130.395 ;
        RECT -30.085 -132.085 -29.755 -131.755 ;
        RECT -30.085 -136.165 -29.755 -135.835 ;
        RECT -30.085 -137.525 -29.755 -137.195 ;
        RECT -30.085 -138.885 -29.755 -138.555 ;
        RECT -30.085 -140.245 -29.755 -139.915 ;
        RECT -30.085 -141.605 -29.755 -141.275 ;
        RECT -30.085 -142.965 -29.755 -142.635 ;
        RECT -30.085 -144.325 -29.755 -143.995 ;
        RECT -30.085 -145.685 -29.755 -145.355 ;
        RECT -30.085 -147.045 -29.755 -146.715 ;
        RECT -30.085 -149.765 -29.755 -149.435 ;
        RECT -30.085 -152.485 -29.755 -152.155 ;
        RECT -30.085 -153.845 -29.755 -153.515 ;
        RECT -30.085 -155.285 -29.755 -154.955 ;
        RECT -30.085 -156.565 -29.755 -156.235 ;
        RECT -30.085 -157.925 -29.755 -157.595 ;
        RECT -30.085 -160.17 -29.755 -159.04 ;
        RECT -30.08 -160.285 -29.76 128.47 ;
        RECT -30.085 127.225 -29.755 128.355 ;
        RECT -30.085 124.955 -29.755 125.285 ;
        RECT -30.085 123.595 -29.755 123.925 ;
        RECT -30.085 122.235 -29.755 122.565 ;
        RECT -30.085 120.875 -29.755 121.205 ;
        RECT -30.085 119.515 -29.755 119.845 ;
        RECT -30.085 118.155 -29.755 118.485 ;
        RECT -30.085 116.795 -29.755 117.125 ;
        RECT -30.085 115.435 -29.755 115.765 ;
        RECT -30.085 114.075 -29.755 114.405 ;
        RECT -30.085 112.715 -29.755 113.045 ;
        RECT -30.085 111.355 -29.755 111.685 ;
        RECT -30.085 109.995 -29.755 110.325 ;
        RECT -30.085 108.635 -29.755 108.965 ;
        RECT -30.085 107.275 -29.755 107.605 ;
        RECT -30.085 105.915 -29.755 106.245 ;
        RECT -30.085 104.555 -29.755 104.885 ;
        RECT -30.085 103.195 -29.755 103.525 ;
        RECT -30.085 101.835 -29.755 102.165 ;
        RECT -30.085 100.475 -29.755 100.805 ;
        RECT -30.085 99.115 -29.755 99.445 ;
        RECT -30.085 97.755 -29.755 98.085 ;
        RECT -30.085 96.395 -29.755 96.725 ;
        RECT -30.085 95.035 -29.755 95.365 ;
        RECT -30.085 93.675 -29.755 94.005 ;
        RECT -30.085 92.315 -29.755 92.645 ;
        RECT -30.085 90.955 -29.755 91.285 ;
        RECT -30.085 89.595 -29.755 89.925 ;
        RECT -30.085 88.235 -29.755 88.565 ;
        RECT -30.085 86.875 -29.755 87.205 ;
        RECT -30.085 85.515 -29.755 85.845 ;
        RECT -30.085 84.155 -29.755 84.485 ;
        RECT -30.085 82.795 -29.755 83.125 ;
        RECT -30.085 81.435 -29.755 81.765 ;
        RECT -30.085 80.075 -29.755 80.405 ;
        RECT -30.085 78.715 -29.755 79.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 127.225 -43.355 128.355 ;
        RECT -43.685 124.955 -43.355 125.285 ;
        RECT -43.685 123.595 -43.355 123.925 ;
        RECT -43.685 122.235 -43.355 122.565 ;
        RECT -43.685 120.875 -43.355 121.205 ;
        RECT -43.685 119.515 -43.355 119.845 ;
        RECT -43.685 118.155 -43.355 118.485 ;
        RECT -43.685 116.795 -43.355 117.125 ;
        RECT -43.685 115.435 -43.355 115.765 ;
        RECT -43.685 114.075 -43.355 114.405 ;
        RECT -43.685 112.715 -43.355 113.045 ;
        RECT -43.685 111.355 -43.355 111.685 ;
        RECT -43.685 109.995 -43.355 110.325 ;
        RECT -43.685 108.635 -43.355 108.965 ;
        RECT -43.685 107.275 -43.355 107.605 ;
        RECT -43.685 105.915 -43.355 106.245 ;
        RECT -43.685 104.555 -43.355 104.885 ;
        RECT -43.685 103.195 -43.355 103.525 ;
        RECT -43.685 101.835 -43.355 102.165 ;
        RECT -43.685 100.475 -43.355 100.805 ;
        RECT -43.685 99.115 -43.355 99.445 ;
        RECT -43.685 97.755 -43.355 98.085 ;
        RECT -43.685 96.395 -43.355 96.725 ;
        RECT -43.685 95.035 -43.355 95.365 ;
        RECT -43.685 93.675 -43.355 94.005 ;
        RECT -43.685 92.315 -43.355 92.645 ;
        RECT -43.685 90.955 -43.355 91.285 ;
        RECT -43.685 89.595 -43.355 89.925 ;
        RECT -43.685 88.235 -43.355 88.565 ;
        RECT -43.685 86.875 -43.355 87.205 ;
        RECT -43.685 85.515 -43.355 85.845 ;
        RECT -43.685 84.155 -43.355 84.485 ;
        RECT -43.685 82.795 -43.355 83.125 ;
        RECT -43.685 81.435 -43.355 81.765 ;
        RECT -43.685 80.075 -43.355 80.405 ;
        RECT -43.685 78.715 -43.355 79.045 ;
        RECT -43.685 77.355 -43.355 77.685 ;
        RECT -43.685 75.995 -43.355 76.325 ;
        RECT -43.685 74.635 -43.355 74.965 ;
        RECT -43.685 73.275 -43.355 73.605 ;
        RECT -43.685 48.795 -43.355 49.125 ;
        RECT -43.685 47.435 -43.355 47.765 ;
        RECT -43.685 46.075 -43.355 46.405 ;
        RECT -43.685 44.715 -43.355 45.045 ;
        RECT -43.685 43.355 -43.355 43.685 ;
        RECT -43.685 41.995 -43.355 42.325 ;
        RECT -43.685 40.635 -43.355 40.965 ;
        RECT -43.685 39.275 -43.355 39.605 ;
        RECT -43.685 37.915 -43.355 38.245 ;
        RECT -43.685 36.555 -43.355 36.885 ;
        RECT -43.685 35.195 -43.355 35.525 ;
        RECT -43.685 33.835 -43.355 34.165 ;
        RECT -43.685 32.475 -43.355 32.805 ;
        RECT -43.685 31.115 -43.355 31.445 ;
        RECT -43.685 29.755 -43.355 30.085 ;
        RECT -43.685 28.395 -43.355 28.725 ;
        RECT -43.685 27.035 -43.355 27.365 ;
        RECT -43.685 25.675 -43.355 26.005 ;
        RECT -43.685 24.315 -43.355 24.645 ;
        RECT -43.685 22.955 -43.355 23.285 ;
        RECT -43.685 21.595 -43.355 21.925 ;
        RECT -43.685 20.235 -43.355 20.565 ;
        RECT -43.685 18.875 -43.355 19.205 ;
        RECT -43.685 17.515 -43.355 17.845 ;
        RECT -43.685 16.155 -43.355 16.485 ;
        RECT -43.685 14.795 -43.355 15.125 ;
        RECT -43.685 13.435 -43.355 13.765 ;
        RECT -43.685 12.075 -43.355 12.405 ;
        RECT -43.685 10.715 -43.355 11.045 ;
        RECT -43.685 9.355 -43.355 9.685 ;
        RECT -43.685 7.995 -43.355 8.325 ;
        RECT -43.685 6.635 -43.355 6.965 ;
        RECT -43.685 5.275 -43.355 5.605 ;
        RECT -43.685 3.915 -43.355 4.245 ;
        RECT -43.685 2.555 -43.355 2.885 ;
        RECT -43.685 1.195 -43.355 1.525 ;
        RECT -43.685 -0.165 -43.355 0.165 ;
        RECT -43.685 -1.525 -43.355 -1.195 ;
        RECT -43.685 -2.885 -43.355 -2.555 ;
        RECT -43.685 -4.245 -43.355 -3.915 ;
        RECT -43.685 -5.605 -43.355 -5.275 ;
        RECT -43.685 -8.325 -43.355 -7.995 ;
        RECT -43.685 -12.405 -43.355 -12.075 ;
        RECT -43.685 -13.765 -43.355 -13.435 ;
        RECT -43.685 -15.125 -43.355 -14.795 ;
        RECT -43.685 -16.485 -43.355 -16.155 ;
        RECT -43.685 -17.845 -43.355 -17.515 ;
        RECT -43.685 -19.205 -43.355 -18.875 ;
        RECT -43.685 -20.565 -43.355 -20.235 ;
        RECT -43.685 -21.925 -43.355 -21.595 ;
        RECT -43.685 -27.365 -43.355 -27.035 ;
        RECT -43.685 -28.725 -43.355 -28.395 ;
        RECT -43.685 -30.085 -43.355 -29.755 ;
        RECT -43.685 -31.445 -43.355 -31.115 ;
        RECT -43.685 -32.805 -43.355 -32.475 ;
        RECT -43.685 -34.165 -43.355 -33.835 ;
        RECT -43.685 -35.525 -43.355 -35.195 ;
        RECT -43.685 -36.885 -43.355 -36.555 ;
        RECT -43.685 -38.245 -43.355 -37.915 ;
        RECT -43.685 -39.605 -43.355 -39.275 ;
        RECT -43.685 -40.965 -43.355 -40.635 ;
        RECT -43.685 -42.325 -43.355 -41.995 ;
        RECT -43.685 -43.685 -43.355 -43.355 ;
        RECT -43.685 -45.045 -43.355 -44.715 ;
        RECT -43.685 -46.405 -43.355 -46.075 ;
        RECT -43.685 -47.765 -43.355 -47.435 ;
        RECT -43.685 -49.125 -43.355 -48.795 ;
        RECT -43.685 -50.485 -43.355 -50.155 ;
        RECT -43.685 -51.845 -43.355 -51.515 ;
        RECT -43.685 -53.205 -43.355 -52.875 ;
        RECT -43.685 -54.565 -43.355 -54.235 ;
        RECT -43.685 -55.925 -43.355 -55.595 ;
        RECT -43.685 -57.285 -43.355 -56.955 ;
        RECT -43.685 -58.645 -43.355 -58.315 ;
        RECT -43.685 -60.005 -43.355 -59.675 ;
        RECT -43.685 -61.365 -43.355 -61.035 ;
        RECT -43.685 -62.725 -43.355 -62.395 ;
        RECT -43.685 -64.085 -43.355 -63.755 ;
        RECT -43.685 -65.445 -43.355 -65.115 ;
        RECT -43.685 -66.805 -43.355 -66.475 ;
        RECT -43.685 -68.165 -43.355 -67.835 ;
        RECT -43.685 -69.525 -43.355 -69.195 ;
        RECT -43.685 -72.245 -43.355 -71.915 ;
        RECT -43.685 -73.605 -43.355 -73.275 ;
        RECT -43.685 -74.965 -43.355 -74.635 ;
        RECT -43.685 -76.325 -43.355 -75.995 ;
        RECT -43.685 -78.29 -43.355 -77.96 ;
        RECT -43.685 -79.045 -43.355 -78.715 ;
        RECT -43.685 -81.765 -43.355 -81.435 ;
        RECT -43.685 -83.125 -43.355 -82.795 ;
        RECT -43.685 -84.485 -43.355 -84.155 ;
        RECT -43.685 -86.43 -43.355 -86.1 ;
        RECT -43.685 -87.205 -43.355 -86.875 ;
        RECT -43.685 -88.565 -43.355 -88.235 ;
        RECT -43.685 -89.925 -43.355 -89.595 ;
        RECT -43.68 -91.28 -43.36 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 -153.845 -43.355 -153.515 ;
        RECT -43.685 -155.285 -43.355 -154.955 ;
        RECT -43.685 -156.565 -43.355 -156.235 ;
        RECT -43.685 -157.925 -43.355 -157.595 ;
        RECT -43.685 -160.17 -43.355 -159.04 ;
        RECT -43.68 -160.285 -43.36 -153.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 127.225 -41.995 128.355 ;
        RECT -42.325 124.955 -41.995 125.285 ;
        RECT -42.325 123.595 -41.995 123.925 ;
        RECT -42.325 122.235 -41.995 122.565 ;
        RECT -42.325 120.875 -41.995 121.205 ;
        RECT -42.325 119.515 -41.995 119.845 ;
        RECT -42.325 118.155 -41.995 118.485 ;
        RECT -42.325 116.795 -41.995 117.125 ;
        RECT -42.325 115.435 -41.995 115.765 ;
        RECT -42.325 114.075 -41.995 114.405 ;
        RECT -42.325 112.715 -41.995 113.045 ;
        RECT -42.325 111.355 -41.995 111.685 ;
        RECT -42.325 109.995 -41.995 110.325 ;
        RECT -42.325 108.635 -41.995 108.965 ;
        RECT -42.325 107.275 -41.995 107.605 ;
        RECT -42.325 105.915 -41.995 106.245 ;
        RECT -42.325 104.555 -41.995 104.885 ;
        RECT -42.325 103.195 -41.995 103.525 ;
        RECT -42.325 101.835 -41.995 102.165 ;
        RECT -42.325 100.475 -41.995 100.805 ;
        RECT -42.325 99.115 -41.995 99.445 ;
        RECT -42.325 97.755 -41.995 98.085 ;
        RECT -42.325 96.395 -41.995 96.725 ;
        RECT -42.325 95.035 -41.995 95.365 ;
        RECT -42.325 93.675 -41.995 94.005 ;
        RECT -42.325 92.315 -41.995 92.645 ;
        RECT -42.325 90.955 -41.995 91.285 ;
        RECT -42.325 89.595 -41.995 89.925 ;
        RECT -42.325 88.235 -41.995 88.565 ;
        RECT -42.325 86.875 -41.995 87.205 ;
        RECT -42.325 85.515 -41.995 85.845 ;
        RECT -42.325 84.155 -41.995 84.485 ;
        RECT -42.325 82.795 -41.995 83.125 ;
        RECT -42.325 81.435 -41.995 81.765 ;
        RECT -42.325 80.075 -41.995 80.405 ;
        RECT -42.325 78.715 -41.995 79.045 ;
        RECT -42.325 77.355 -41.995 77.685 ;
        RECT -42.325 75.995 -41.995 76.325 ;
        RECT -42.325 74.635 -41.995 74.965 ;
        RECT -42.325 73.275 -41.995 73.605 ;
        RECT -42.325 71.915 -41.995 72.245 ;
        RECT -42.325 70.555 -41.995 70.885 ;
        RECT -42.325 69.195 -41.995 69.525 ;
        RECT -42.325 67.835 -41.995 68.165 ;
        RECT -42.325 66.475 -41.995 66.805 ;
        RECT -42.325 65.115 -41.995 65.445 ;
        RECT -42.325 63.755 -41.995 64.085 ;
        RECT -42.325 62.395 -41.995 62.725 ;
        RECT -42.325 61.035 -41.995 61.365 ;
        RECT -42.325 59.675 -41.995 60.005 ;
        RECT -42.325 58.315 -41.995 58.645 ;
        RECT -42.325 56.955 -41.995 57.285 ;
        RECT -42.325 55.595 -41.995 55.925 ;
        RECT -42.325 54.235 -41.995 54.565 ;
        RECT -42.325 52.875 -41.995 53.205 ;
        RECT -42.325 51.515 -41.995 51.845 ;
        RECT -42.325 50.155 -41.995 50.485 ;
        RECT -42.325 48.795 -41.995 49.125 ;
        RECT -42.325 47.435 -41.995 47.765 ;
        RECT -42.325 46.075 -41.995 46.405 ;
        RECT -42.325 44.715 -41.995 45.045 ;
        RECT -42.325 43.355 -41.995 43.685 ;
        RECT -42.325 41.995 -41.995 42.325 ;
        RECT -42.325 40.635 -41.995 40.965 ;
        RECT -42.325 39.275 -41.995 39.605 ;
        RECT -42.325 37.915 -41.995 38.245 ;
        RECT -42.325 36.555 -41.995 36.885 ;
        RECT -42.325 35.195 -41.995 35.525 ;
        RECT -42.325 33.835 -41.995 34.165 ;
        RECT -42.325 32.475 -41.995 32.805 ;
        RECT -42.325 31.115 -41.995 31.445 ;
        RECT -42.325 29.755 -41.995 30.085 ;
        RECT -42.325 28.395 -41.995 28.725 ;
        RECT -42.325 27.035 -41.995 27.365 ;
        RECT -42.325 25.675 -41.995 26.005 ;
        RECT -42.325 24.315 -41.995 24.645 ;
        RECT -42.325 22.955 -41.995 23.285 ;
        RECT -42.325 21.595 -41.995 21.925 ;
        RECT -42.325 20.235 -41.995 20.565 ;
        RECT -42.325 18.875 -41.995 19.205 ;
        RECT -42.325 17.515 -41.995 17.845 ;
        RECT -42.325 16.155 -41.995 16.485 ;
        RECT -42.325 14.795 -41.995 15.125 ;
        RECT -42.325 13.435 -41.995 13.765 ;
        RECT -42.325 12.075 -41.995 12.405 ;
        RECT -42.325 10.715 -41.995 11.045 ;
        RECT -42.325 9.355 -41.995 9.685 ;
        RECT -42.325 7.995 -41.995 8.325 ;
        RECT -42.325 6.635 -41.995 6.965 ;
        RECT -42.325 5.275 -41.995 5.605 ;
        RECT -42.325 3.915 -41.995 4.245 ;
        RECT -42.325 2.555 -41.995 2.885 ;
        RECT -42.325 1.195 -41.995 1.525 ;
        RECT -42.325 -0.165 -41.995 0.165 ;
        RECT -42.325 -1.525 -41.995 -1.195 ;
        RECT -42.325 -2.885 -41.995 -2.555 ;
        RECT -42.325 -4.245 -41.995 -3.915 ;
        RECT -42.325 -5.605 -41.995 -5.275 ;
        RECT -42.325 -8.325 -41.995 -7.995 ;
        RECT -42.325 -12.405 -41.995 -12.075 ;
        RECT -42.325 -13.765 -41.995 -13.435 ;
        RECT -42.325 -15.125 -41.995 -14.795 ;
        RECT -42.325 -16.485 -41.995 -16.155 ;
        RECT -42.325 -17.845 -41.995 -17.515 ;
        RECT -42.325 -19.205 -41.995 -18.875 ;
        RECT -42.325 -20.565 -41.995 -20.235 ;
        RECT -42.325 -21.925 -41.995 -21.595 ;
        RECT -42.325 -27.365 -41.995 -27.035 ;
        RECT -42.325 -28.725 -41.995 -28.395 ;
        RECT -42.325 -30.085 -41.995 -29.755 ;
        RECT -42.325 -31.445 -41.995 -31.115 ;
        RECT -42.325 -32.805 -41.995 -32.475 ;
        RECT -42.325 -34.165 -41.995 -33.835 ;
        RECT -42.325 -35.525 -41.995 -35.195 ;
        RECT -42.325 -36.885 -41.995 -36.555 ;
        RECT -42.325 -38.245 -41.995 -37.915 ;
        RECT -42.325 -39.605 -41.995 -39.275 ;
        RECT -42.325 -40.965 -41.995 -40.635 ;
        RECT -42.325 -42.325 -41.995 -41.995 ;
        RECT -42.325 -43.685 -41.995 -43.355 ;
        RECT -42.325 -45.045 -41.995 -44.715 ;
        RECT -42.325 -46.405 -41.995 -46.075 ;
        RECT -42.325 -47.765 -41.995 -47.435 ;
        RECT -42.325 -49.125 -41.995 -48.795 ;
        RECT -42.325 -50.485 -41.995 -50.155 ;
        RECT -42.325 -51.845 -41.995 -51.515 ;
        RECT -42.325 -53.205 -41.995 -52.875 ;
        RECT -42.325 -54.565 -41.995 -54.235 ;
        RECT -42.325 -55.925 -41.995 -55.595 ;
        RECT -42.325 -57.285 -41.995 -56.955 ;
        RECT -42.325 -58.645 -41.995 -58.315 ;
        RECT -42.325 -60.005 -41.995 -59.675 ;
        RECT -42.325 -61.365 -41.995 -61.035 ;
        RECT -42.325 -62.725 -41.995 -62.395 ;
        RECT -42.325 -64.085 -41.995 -63.755 ;
        RECT -42.325 -65.445 -41.995 -65.115 ;
        RECT -42.325 -66.805 -41.995 -66.475 ;
        RECT -42.325 -68.165 -41.995 -67.835 ;
        RECT -42.325 -69.525 -41.995 -69.195 ;
        RECT -42.325 -72.245 -41.995 -71.915 ;
        RECT -42.325 -73.605 -41.995 -73.275 ;
        RECT -42.325 -74.965 -41.995 -74.635 ;
        RECT -42.325 -76.325 -41.995 -75.995 ;
        RECT -42.325 -78.29 -41.995 -77.96 ;
        RECT -42.325 -79.045 -41.995 -78.715 ;
        RECT -42.325 -81.765 -41.995 -81.435 ;
        RECT -42.325 -83.125 -41.995 -82.795 ;
        RECT -42.325 -84.485 -41.995 -84.155 ;
        RECT -42.325 -86.43 -41.995 -86.1 ;
        RECT -42.325 -87.205 -41.995 -86.875 ;
        RECT -42.325 -88.565 -41.995 -88.235 ;
        RECT -42.325 -89.925 -41.995 -89.595 ;
        RECT -42.325 -92.645 -41.995 -92.315 ;
        RECT -42.325 -94.005 -41.995 -93.675 ;
        RECT -42.325 -95.365 -41.995 -95.035 ;
        RECT -42.325 -96.725 -41.995 -96.395 ;
        RECT -42.325 -98.085 -41.995 -97.755 ;
        RECT -42.325 -102.165 -41.995 -101.835 ;
        RECT -42.325 -103.525 -41.995 -103.195 ;
        RECT -42.325 -104.885 -41.995 -104.555 ;
        RECT -42.325 -106.245 -41.995 -105.915 ;
        RECT -42.325 -107.605 -41.995 -107.275 ;
        RECT -42.325 -108.965 -41.995 -108.635 ;
        RECT -42.325 -110.325 -41.995 -109.995 ;
        RECT -42.325 -111.685 -41.995 -111.355 ;
        RECT -42.325 -113.045 -41.995 -112.715 ;
        RECT -42.325 -114.405 -41.995 -114.075 ;
        RECT -42.325 -115.765 -41.995 -115.435 ;
        RECT -42.325 -117.125 -41.995 -116.795 ;
        RECT -42.325 -118.485 -41.995 -118.155 ;
        RECT -42.325 -119.845 -41.995 -119.515 ;
        RECT -42.325 -121.205 -41.995 -120.875 ;
        RECT -42.325 -122.565 -41.995 -122.235 ;
        RECT -42.325 -123.925 -41.995 -123.595 ;
        RECT -42.325 -125.285 -41.995 -124.955 ;
        RECT -42.325 -126.645 -41.995 -126.315 ;
        RECT -42.325 -128.005 -41.995 -127.675 ;
        RECT -42.325 -129.365 -41.995 -129.035 ;
        RECT -42.325 -130.725 -41.995 -130.395 ;
        RECT -42.325 -132.085 -41.995 -131.755 ;
        RECT -42.325 -133.445 -41.995 -133.115 ;
        RECT -42.325 -134.805 -41.995 -134.475 ;
        RECT -42.325 -136.165 -41.995 -135.835 ;
        RECT -42.325 -137.525 -41.995 -137.195 ;
        RECT -42.325 -138.885 -41.995 -138.555 ;
        RECT -42.325 -140.245 -41.995 -139.915 ;
        RECT -42.325 -141.605 -41.995 -141.275 ;
        RECT -42.325 -142.965 -41.995 -142.635 ;
        RECT -42.325 -144.325 -41.995 -143.995 ;
        RECT -42.325 -145.685 -41.995 -145.355 ;
        RECT -42.325 -147.045 -41.995 -146.715 ;
        RECT -42.325 -149.765 -41.995 -149.435 ;
        RECT -42.325 -153.845 -41.995 -153.515 ;
        RECT -42.325 -155.285 -41.995 -154.955 ;
        RECT -42.325 -156.565 -41.995 -156.235 ;
        RECT -42.325 -157.925 -41.995 -157.595 ;
        RECT -42.325 -160.17 -41.995 -159.04 ;
        RECT -42.32 -160.285 -42 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.965 127.225 -40.635 128.355 ;
        RECT -40.965 124.955 -40.635 125.285 ;
        RECT -40.965 123.595 -40.635 123.925 ;
        RECT -40.965 122.235 -40.635 122.565 ;
        RECT -40.965 120.875 -40.635 121.205 ;
        RECT -40.965 119.515 -40.635 119.845 ;
        RECT -40.965 118.155 -40.635 118.485 ;
        RECT -40.965 116.795 -40.635 117.125 ;
        RECT -40.965 115.435 -40.635 115.765 ;
        RECT -40.965 114.075 -40.635 114.405 ;
        RECT -40.965 112.715 -40.635 113.045 ;
        RECT -40.965 111.355 -40.635 111.685 ;
        RECT -40.965 109.995 -40.635 110.325 ;
        RECT -40.965 108.635 -40.635 108.965 ;
        RECT -40.965 107.275 -40.635 107.605 ;
        RECT -40.965 105.915 -40.635 106.245 ;
        RECT -40.965 104.555 -40.635 104.885 ;
        RECT -40.965 103.195 -40.635 103.525 ;
        RECT -40.965 101.835 -40.635 102.165 ;
        RECT -40.965 100.475 -40.635 100.805 ;
        RECT -40.965 99.115 -40.635 99.445 ;
        RECT -40.965 97.755 -40.635 98.085 ;
        RECT -40.965 96.395 -40.635 96.725 ;
        RECT -40.965 95.035 -40.635 95.365 ;
        RECT -40.965 93.675 -40.635 94.005 ;
        RECT -40.965 92.315 -40.635 92.645 ;
        RECT -40.965 90.955 -40.635 91.285 ;
        RECT -40.965 89.595 -40.635 89.925 ;
        RECT -40.965 88.235 -40.635 88.565 ;
        RECT -40.965 86.875 -40.635 87.205 ;
        RECT -40.965 85.515 -40.635 85.845 ;
        RECT -40.965 84.155 -40.635 84.485 ;
        RECT -40.965 82.795 -40.635 83.125 ;
        RECT -40.965 81.435 -40.635 81.765 ;
        RECT -40.965 80.075 -40.635 80.405 ;
        RECT -40.965 78.715 -40.635 79.045 ;
        RECT -40.965 77.355 -40.635 77.685 ;
        RECT -40.965 75.995 -40.635 76.325 ;
        RECT -40.965 74.635 -40.635 74.965 ;
        RECT -40.965 73.275 -40.635 73.605 ;
        RECT -40.965 71.915 -40.635 72.245 ;
        RECT -40.965 70.555 -40.635 70.885 ;
        RECT -40.965 69.195 -40.635 69.525 ;
        RECT -40.965 67.835 -40.635 68.165 ;
        RECT -40.965 66.475 -40.635 66.805 ;
        RECT -40.965 65.115 -40.635 65.445 ;
        RECT -40.965 63.755 -40.635 64.085 ;
        RECT -40.965 62.395 -40.635 62.725 ;
        RECT -40.965 61.035 -40.635 61.365 ;
        RECT -40.965 59.675 -40.635 60.005 ;
        RECT -40.965 58.315 -40.635 58.645 ;
        RECT -40.965 56.955 -40.635 57.285 ;
        RECT -40.965 55.595 -40.635 55.925 ;
        RECT -40.965 54.235 -40.635 54.565 ;
        RECT -40.965 52.875 -40.635 53.205 ;
        RECT -40.965 51.515 -40.635 51.845 ;
        RECT -40.965 50.155 -40.635 50.485 ;
        RECT -40.965 48.795 -40.635 49.125 ;
        RECT -40.965 47.435 -40.635 47.765 ;
        RECT -40.965 46.075 -40.635 46.405 ;
        RECT -40.965 44.715 -40.635 45.045 ;
        RECT -40.965 43.355 -40.635 43.685 ;
        RECT -40.965 41.995 -40.635 42.325 ;
        RECT -40.965 40.635 -40.635 40.965 ;
        RECT -40.965 39.275 -40.635 39.605 ;
        RECT -40.965 37.915 -40.635 38.245 ;
        RECT -40.965 36.555 -40.635 36.885 ;
        RECT -40.965 35.195 -40.635 35.525 ;
        RECT -40.965 33.835 -40.635 34.165 ;
        RECT -40.965 32.475 -40.635 32.805 ;
        RECT -40.965 31.115 -40.635 31.445 ;
        RECT -40.965 29.755 -40.635 30.085 ;
        RECT -40.965 28.395 -40.635 28.725 ;
        RECT -40.965 27.035 -40.635 27.365 ;
        RECT -40.965 25.675 -40.635 26.005 ;
        RECT -40.965 24.315 -40.635 24.645 ;
        RECT -40.965 22.955 -40.635 23.285 ;
        RECT -40.965 21.595 -40.635 21.925 ;
        RECT -40.965 20.235 -40.635 20.565 ;
        RECT -40.965 18.875 -40.635 19.205 ;
        RECT -40.965 17.515 -40.635 17.845 ;
        RECT -40.965 16.155 -40.635 16.485 ;
        RECT -40.965 14.795 -40.635 15.125 ;
        RECT -40.965 13.435 -40.635 13.765 ;
        RECT -40.965 12.075 -40.635 12.405 ;
        RECT -40.965 10.715 -40.635 11.045 ;
        RECT -40.965 9.355 -40.635 9.685 ;
        RECT -40.965 7.995 -40.635 8.325 ;
        RECT -40.965 6.635 -40.635 6.965 ;
        RECT -40.965 5.275 -40.635 5.605 ;
        RECT -40.965 3.915 -40.635 4.245 ;
        RECT -40.965 2.555 -40.635 2.885 ;
        RECT -40.965 1.195 -40.635 1.525 ;
        RECT -40.965 -0.165 -40.635 0.165 ;
        RECT -40.965 -1.525 -40.635 -1.195 ;
        RECT -40.965 -2.885 -40.635 -2.555 ;
        RECT -40.965 -4.245 -40.635 -3.915 ;
        RECT -40.965 -8.325 -40.635 -7.995 ;
        RECT -40.965 -12.405 -40.635 -12.075 ;
        RECT -40.965 -13.765 -40.635 -13.435 ;
        RECT -40.965 -15.125 -40.635 -14.795 ;
        RECT -40.965 -16.485 -40.635 -16.155 ;
        RECT -40.965 -17.845 -40.635 -17.515 ;
        RECT -40.965 -19.205 -40.635 -18.875 ;
        RECT -40.965 -20.565 -40.635 -20.235 ;
        RECT -40.965 -21.925 -40.635 -21.595 ;
        RECT -40.965 -28.725 -40.635 -28.395 ;
        RECT -40.965 -30.085 -40.635 -29.755 ;
        RECT -40.965 -31.445 -40.635 -31.115 ;
        RECT -40.965 -32.805 -40.635 -32.475 ;
        RECT -40.965 -34.165 -40.635 -33.835 ;
        RECT -40.965 -35.525 -40.635 -35.195 ;
        RECT -40.965 -36.885 -40.635 -36.555 ;
        RECT -40.965 -38.245 -40.635 -37.915 ;
        RECT -40.965 -39.605 -40.635 -39.275 ;
        RECT -40.965 -40.965 -40.635 -40.635 ;
        RECT -40.965 -42.325 -40.635 -41.995 ;
        RECT -40.965 -43.685 -40.635 -43.355 ;
        RECT -40.965 -45.045 -40.635 -44.715 ;
        RECT -40.965 -46.405 -40.635 -46.075 ;
        RECT -40.965 -47.765 -40.635 -47.435 ;
        RECT -40.965 -49.125 -40.635 -48.795 ;
        RECT -40.965 -50.485 -40.635 -50.155 ;
        RECT -40.965 -51.845 -40.635 -51.515 ;
        RECT -40.965 -53.205 -40.635 -52.875 ;
        RECT -40.965 -54.565 -40.635 -54.235 ;
        RECT -40.965 -55.925 -40.635 -55.595 ;
        RECT -40.965 -57.285 -40.635 -56.955 ;
        RECT -40.965 -58.645 -40.635 -58.315 ;
        RECT -40.965 -60.005 -40.635 -59.675 ;
        RECT -40.965 -61.365 -40.635 -61.035 ;
        RECT -40.965 -62.725 -40.635 -62.395 ;
        RECT -40.965 -64.085 -40.635 -63.755 ;
        RECT -40.965 -65.445 -40.635 -65.115 ;
        RECT -40.965 -66.805 -40.635 -66.475 ;
        RECT -40.965 -68.165 -40.635 -67.835 ;
        RECT -40.965 -69.525 -40.635 -69.195 ;
        RECT -40.965 -72.245 -40.635 -71.915 ;
        RECT -40.965 -73.605 -40.635 -73.275 ;
        RECT -40.965 -74.965 -40.635 -74.635 ;
        RECT -40.965 -76.325 -40.635 -75.995 ;
        RECT -40.965 -78.29 -40.635 -77.96 ;
        RECT -40.965 -79.045 -40.635 -78.715 ;
        RECT -40.965 -81.765 -40.635 -81.435 ;
        RECT -40.965 -83.125 -40.635 -82.795 ;
        RECT -40.965 -84.485 -40.635 -84.155 ;
        RECT -40.965 -86.43 -40.635 -86.1 ;
        RECT -40.965 -87.205 -40.635 -86.875 ;
        RECT -40.965 -88.565 -40.635 -88.235 ;
        RECT -40.965 -89.925 -40.635 -89.595 ;
        RECT -40.965 -92.645 -40.635 -92.315 ;
        RECT -40.965 -94.005 -40.635 -93.675 ;
        RECT -40.965 -95.365 -40.635 -95.035 ;
        RECT -40.965 -96.725 -40.635 -96.395 ;
        RECT -40.965 -98.085 -40.635 -97.755 ;
        RECT -40.965 -102.165 -40.635 -101.835 ;
        RECT -40.965 -103.525 -40.635 -103.195 ;
        RECT -40.965 -104.885 -40.635 -104.555 ;
        RECT -40.965 -106.245 -40.635 -105.915 ;
        RECT -40.965 -107.605 -40.635 -107.275 ;
        RECT -40.965 -108.965 -40.635 -108.635 ;
        RECT -40.965 -110.325 -40.635 -109.995 ;
        RECT -40.965 -111.685 -40.635 -111.355 ;
        RECT -40.965 -113.045 -40.635 -112.715 ;
        RECT -40.965 -114.405 -40.635 -114.075 ;
        RECT -40.965 -115.765 -40.635 -115.435 ;
        RECT -40.965 -117.125 -40.635 -116.795 ;
        RECT -40.965 -118.485 -40.635 -118.155 ;
        RECT -40.965 -119.845 -40.635 -119.515 ;
        RECT -40.965 -121.205 -40.635 -120.875 ;
        RECT -40.965 -122.565 -40.635 -122.235 ;
        RECT -40.965 -123.925 -40.635 -123.595 ;
        RECT -40.965 -125.285 -40.635 -124.955 ;
        RECT -40.965 -126.645 -40.635 -126.315 ;
        RECT -40.965 -128.005 -40.635 -127.675 ;
        RECT -40.965 -130.725 -40.635 -130.395 ;
        RECT -40.965 -132.085 -40.635 -131.755 ;
        RECT -40.965 -133.445 -40.635 -133.115 ;
        RECT -40.965 -134.805 -40.635 -134.475 ;
        RECT -40.965 -137.525 -40.635 -137.195 ;
        RECT -40.965 -138.885 -40.635 -138.555 ;
        RECT -40.965 -140.245 -40.635 -139.915 ;
        RECT -40.965 -141.605 -40.635 -141.275 ;
        RECT -40.965 -142.965 -40.635 -142.635 ;
        RECT -40.965 -144.325 -40.635 -143.995 ;
        RECT -40.965 -145.685 -40.635 -145.355 ;
        RECT -40.965 -147.045 -40.635 -146.715 ;
        RECT -40.965 -149.765 -40.635 -149.435 ;
        RECT -40.965 -153.845 -40.635 -153.515 ;
        RECT -40.965 -156.565 -40.635 -156.235 ;
        RECT -40.965 -157.925 -40.635 -157.595 ;
        RECT -40.965 -160.17 -40.635 -159.04 ;
        RECT -40.96 -160.285 -40.64 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.605 127.225 -39.275 128.355 ;
        RECT -39.605 124.955 -39.275 125.285 ;
        RECT -39.605 123.595 -39.275 123.925 ;
        RECT -39.605 122.235 -39.275 122.565 ;
        RECT -39.605 120.875 -39.275 121.205 ;
        RECT -39.605 119.515 -39.275 119.845 ;
        RECT -39.605 118.155 -39.275 118.485 ;
        RECT -39.605 116.795 -39.275 117.125 ;
        RECT -39.605 115.435 -39.275 115.765 ;
        RECT -39.605 114.075 -39.275 114.405 ;
        RECT -39.605 112.715 -39.275 113.045 ;
        RECT -39.605 111.355 -39.275 111.685 ;
        RECT -39.605 109.995 -39.275 110.325 ;
        RECT -39.605 108.635 -39.275 108.965 ;
        RECT -39.605 107.275 -39.275 107.605 ;
        RECT -39.605 105.915 -39.275 106.245 ;
        RECT -39.605 104.555 -39.275 104.885 ;
        RECT -39.605 103.195 -39.275 103.525 ;
        RECT -39.605 101.835 -39.275 102.165 ;
        RECT -39.605 100.475 -39.275 100.805 ;
        RECT -39.605 99.115 -39.275 99.445 ;
        RECT -39.605 97.755 -39.275 98.085 ;
        RECT -39.605 96.395 -39.275 96.725 ;
        RECT -39.605 95.035 -39.275 95.365 ;
        RECT -39.605 93.675 -39.275 94.005 ;
        RECT -39.605 92.315 -39.275 92.645 ;
        RECT -39.605 90.955 -39.275 91.285 ;
        RECT -39.605 89.595 -39.275 89.925 ;
        RECT -39.605 88.235 -39.275 88.565 ;
        RECT -39.605 86.875 -39.275 87.205 ;
        RECT -39.605 85.515 -39.275 85.845 ;
        RECT -39.605 84.155 -39.275 84.485 ;
        RECT -39.605 82.795 -39.275 83.125 ;
        RECT -39.605 81.435 -39.275 81.765 ;
        RECT -39.605 80.075 -39.275 80.405 ;
        RECT -39.605 78.715 -39.275 79.045 ;
        RECT -39.605 77.355 -39.275 77.685 ;
        RECT -39.605 75.995 -39.275 76.325 ;
        RECT -39.605 74.635 -39.275 74.965 ;
        RECT -39.605 73.275 -39.275 73.605 ;
        RECT -39.605 71.915 -39.275 72.245 ;
        RECT -39.605 70.555 -39.275 70.885 ;
        RECT -39.605 69.195 -39.275 69.525 ;
        RECT -39.605 67.835 -39.275 68.165 ;
        RECT -39.605 66.475 -39.275 66.805 ;
        RECT -39.605 65.115 -39.275 65.445 ;
        RECT -39.605 63.755 -39.275 64.085 ;
        RECT -39.605 62.395 -39.275 62.725 ;
        RECT -39.605 61.035 -39.275 61.365 ;
        RECT -39.605 59.675 -39.275 60.005 ;
        RECT -39.605 58.315 -39.275 58.645 ;
        RECT -39.605 56.955 -39.275 57.285 ;
        RECT -39.605 55.595 -39.275 55.925 ;
        RECT -39.605 54.235 -39.275 54.565 ;
        RECT -39.605 52.875 -39.275 53.205 ;
        RECT -39.605 51.515 -39.275 51.845 ;
        RECT -39.605 50.155 -39.275 50.485 ;
        RECT -39.605 48.795 -39.275 49.125 ;
        RECT -39.605 47.435 -39.275 47.765 ;
        RECT -39.605 46.075 -39.275 46.405 ;
        RECT -39.605 44.715 -39.275 45.045 ;
        RECT -39.605 43.355 -39.275 43.685 ;
        RECT -39.605 41.995 -39.275 42.325 ;
        RECT -39.605 40.635 -39.275 40.965 ;
        RECT -39.605 39.275 -39.275 39.605 ;
        RECT -39.605 37.915 -39.275 38.245 ;
        RECT -39.605 36.555 -39.275 36.885 ;
        RECT -39.605 35.195 -39.275 35.525 ;
        RECT -39.605 33.835 -39.275 34.165 ;
        RECT -39.605 32.475 -39.275 32.805 ;
        RECT -39.605 31.115 -39.275 31.445 ;
        RECT -39.605 29.755 -39.275 30.085 ;
        RECT -39.605 28.395 -39.275 28.725 ;
        RECT -39.605 27.035 -39.275 27.365 ;
        RECT -39.605 25.675 -39.275 26.005 ;
        RECT -39.605 24.315 -39.275 24.645 ;
        RECT -39.605 22.955 -39.275 23.285 ;
        RECT -39.605 21.595 -39.275 21.925 ;
        RECT -39.605 20.235 -39.275 20.565 ;
        RECT -39.605 18.875 -39.275 19.205 ;
        RECT -39.605 17.515 -39.275 17.845 ;
        RECT -39.605 16.155 -39.275 16.485 ;
        RECT -39.605 14.795 -39.275 15.125 ;
        RECT -39.605 13.435 -39.275 13.765 ;
        RECT -39.605 12.075 -39.275 12.405 ;
        RECT -39.605 10.715 -39.275 11.045 ;
        RECT -39.605 9.355 -39.275 9.685 ;
        RECT -39.605 7.995 -39.275 8.325 ;
        RECT -39.605 6.635 -39.275 6.965 ;
        RECT -39.605 5.275 -39.275 5.605 ;
        RECT -39.605 3.915 -39.275 4.245 ;
        RECT -39.605 2.555 -39.275 2.885 ;
        RECT -39.605 1.195 -39.275 1.525 ;
        RECT -39.605 -0.165 -39.275 0.165 ;
        RECT -39.605 -1.525 -39.275 -1.195 ;
        RECT -39.605 -2.885 -39.275 -2.555 ;
        RECT -39.605 -8.325 -39.275 -7.995 ;
        RECT -39.605 -12.405 -39.275 -12.075 ;
        RECT -39.605 -13.765 -39.275 -13.435 ;
        RECT -39.605 -15.125 -39.275 -14.795 ;
        RECT -39.605 -16.485 -39.275 -16.155 ;
        RECT -39.605 -17.845 -39.275 -17.515 ;
        RECT -39.605 -19.205 -39.275 -18.875 ;
        RECT -39.605 -20.565 -39.275 -20.235 ;
        RECT -39.605 -21.925 -39.275 -21.595 ;
        RECT -39.605 -28.725 -39.275 -28.395 ;
        RECT -39.605 -30.085 -39.275 -29.755 ;
        RECT -39.605 -31.445 -39.275 -31.115 ;
        RECT -39.605 -32.805 -39.275 -32.475 ;
        RECT -39.605 -34.165 -39.275 -33.835 ;
        RECT -39.605 -35.525 -39.275 -35.195 ;
        RECT -39.605 -36.885 -39.275 -36.555 ;
        RECT -39.605 -38.245 -39.275 -37.915 ;
        RECT -39.605 -39.605 -39.275 -39.275 ;
        RECT -39.605 -40.965 -39.275 -40.635 ;
        RECT -39.605 -42.325 -39.275 -41.995 ;
        RECT -39.605 -43.685 -39.275 -43.355 ;
        RECT -39.605 -45.045 -39.275 -44.715 ;
        RECT -39.605 -47.765 -39.275 -47.435 ;
        RECT -39.605 -49.125 -39.275 -48.795 ;
        RECT -39.605 -50.485 -39.275 -50.155 ;
        RECT -39.605 -51.845 -39.275 -51.515 ;
        RECT -39.605 -53.205 -39.275 -52.875 ;
        RECT -39.605 -54.565 -39.275 -54.235 ;
        RECT -39.605 -55.925 -39.275 -55.595 ;
        RECT -39.605 -57.285 -39.275 -56.955 ;
        RECT -39.605 -58.645 -39.275 -58.315 ;
        RECT -39.605 -60.005 -39.275 -59.675 ;
        RECT -39.605 -61.365 -39.275 -61.035 ;
        RECT -39.605 -62.725 -39.275 -62.395 ;
        RECT -39.605 -64.085 -39.275 -63.755 ;
        RECT -39.605 -65.445 -39.275 -65.115 ;
        RECT -39.605 -66.805 -39.275 -66.475 ;
        RECT -39.605 -68.165 -39.275 -67.835 ;
        RECT -39.605 -69.525 -39.275 -69.195 ;
        RECT -39.605 -72.245 -39.275 -71.915 ;
        RECT -39.605 -73.605 -39.275 -73.275 ;
        RECT -39.605 -74.965 -39.275 -74.635 ;
        RECT -39.605 -76.325 -39.275 -75.995 ;
        RECT -39.605 -78.29 -39.275 -77.96 ;
        RECT -39.605 -79.045 -39.275 -78.715 ;
        RECT -39.605 -81.765 -39.275 -81.435 ;
        RECT -39.605 -83.125 -39.275 -82.795 ;
        RECT -39.605 -84.485 -39.275 -84.155 ;
        RECT -39.605 -86.43 -39.275 -86.1 ;
        RECT -39.605 -87.205 -39.275 -86.875 ;
        RECT -39.605 -88.565 -39.275 -88.235 ;
        RECT -39.605 -89.925 -39.275 -89.595 ;
        RECT -39.605 -92.645 -39.275 -92.315 ;
        RECT -39.605 -94.005 -39.275 -93.675 ;
        RECT -39.605 -95.365 -39.275 -95.035 ;
        RECT -39.605 -96.725 -39.275 -96.395 ;
        RECT -39.605 -98.085 -39.275 -97.755 ;
        RECT -39.605 -102.165 -39.275 -101.835 ;
        RECT -39.605 -103.525 -39.275 -103.195 ;
        RECT -39.605 -104.885 -39.275 -104.555 ;
        RECT -39.605 -106.245 -39.275 -105.915 ;
        RECT -39.605 -107.605 -39.275 -107.275 ;
        RECT -39.605 -108.965 -39.275 -108.635 ;
        RECT -39.605 -110.325 -39.275 -109.995 ;
        RECT -39.605 -113.045 -39.275 -112.715 ;
        RECT -39.605 -114.405 -39.275 -114.075 ;
        RECT -39.605 -115.765 -39.275 -115.435 ;
        RECT -39.605 -117.125 -39.275 -116.795 ;
        RECT -39.605 -118.485 -39.275 -118.155 ;
        RECT -39.605 -119.845 -39.275 -119.515 ;
        RECT -39.605 -121.205 -39.275 -120.875 ;
        RECT -39.605 -122.565 -39.275 -122.235 ;
        RECT -39.605 -123.925 -39.275 -123.595 ;
        RECT -39.605 -125.285 -39.275 -124.955 ;
        RECT -39.605 -126.645 -39.275 -126.315 ;
        RECT -39.605 -128.005 -39.275 -127.675 ;
        RECT -39.605 -130.725 -39.275 -130.395 ;
        RECT -39.605 -132.085 -39.275 -131.755 ;
        RECT -39.605 -134.805 -39.275 -134.475 ;
        RECT -39.605 -137.525 -39.275 -137.195 ;
        RECT -39.605 -138.885 -39.275 -138.555 ;
        RECT -39.605 -140.245 -39.275 -139.915 ;
        RECT -39.605 -141.605 -39.275 -141.275 ;
        RECT -39.605 -142.965 -39.275 -142.635 ;
        RECT -39.605 -144.325 -39.275 -143.995 ;
        RECT -39.605 -145.685 -39.275 -145.355 ;
        RECT -39.605 -147.045 -39.275 -146.715 ;
        RECT -39.605 -149.765 -39.275 -149.435 ;
        RECT -39.6 -151.8 -39.28 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.245 120.875 -37.915 121.205 ;
        RECT -38.245 119.515 -37.915 119.845 ;
        RECT -38.245 118.155 -37.915 118.485 ;
        RECT -38.245 116.795 -37.915 117.125 ;
        RECT -38.245 115.435 -37.915 115.765 ;
        RECT -38.245 114.075 -37.915 114.405 ;
        RECT -38.245 112.715 -37.915 113.045 ;
        RECT -38.245 111.355 -37.915 111.685 ;
        RECT -38.245 109.995 -37.915 110.325 ;
        RECT -38.245 108.635 -37.915 108.965 ;
        RECT -38.245 107.275 -37.915 107.605 ;
        RECT -38.245 105.915 -37.915 106.245 ;
        RECT -38.245 104.555 -37.915 104.885 ;
        RECT -38.245 103.195 -37.915 103.525 ;
        RECT -38.245 101.835 -37.915 102.165 ;
        RECT -38.245 100.475 -37.915 100.805 ;
        RECT -38.245 99.115 -37.915 99.445 ;
        RECT -38.245 97.755 -37.915 98.085 ;
        RECT -38.245 96.395 -37.915 96.725 ;
        RECT -38.245 95.035 -37.915 95.365 ;
        RECT -38.245 93.675 -37.915 94.005 ;
        RECT -38.245 92.315 -37.915 92.645 ;
        RECT -38.245 90.955 -37.915 91.285 ;
        RECT -38.245 89.595 -37.915 89.925 ;
        RECT -38.245 88.235 -37.915 88.565 ;
        RECT -38.245 86.875 -37.915 87.205 ;
        RECT -38.245 85.515 -37.915 85.845 ;
        RECT -38.245 84.155 -37.915 84.485 ;
        RECT -38.245 82.795 -37.915 83.125 ;
        RECT -38.245 81.435 -37.915 81.765 ;
        RECT -38.245 80.075 -37.915 80.405 ;
        RECT -38.245 78.715 -37.915 79.045 ;
        RECT -38.245 77.355 -37.915 77.685 ;
        RECT -38.245 75.995 -37.915 76.325 ;
        RECT -38.245 74.635 -37.915 74.965 ;
        RECT -38.245 73.275 -37.915 73.605 ;
        RECT -38.245 71.915 -37.915 72.245 ;
        RECT -38.245 70.555 -37.915 70.885 ;
        RECT -38.245 69.195 -37.915 69.525 ;
        RECT -38.245 67.835 -37.915 68.165 ;
        RECT -38.245 66.475 -37.915 66.805 ;
        RECT -38.245 65.115 -37.915 65.445 ;
        RECT -38.245 63.755 -37.915 64.085 ;
        RECT -38.245 62.395 -37.915 62.725 ;
        RECT -38.245 61.035 -37.915 61.365 ;
        RECT -38.245 59.675 -37.915 60.005 ;
        RECT -38.245 58.315 -37.915 58.645 ;
        RECT -38.245 56.955 -37.915 57.285 ;
        RECT -38.245 55.595 -37.915 55.925 ;
        RECT -38.245 54.235 -37.915 54.565 ;
        RECT -38.245 52.875 -37.915 53.205 ;
        RECT -38.245 51.515 -37.915 51.845 ;
        RECT -38.245 50.155 -37.915 50.485 ;
        RECT -38.245 48.795 -37.915 49.125 ;
        RECT -38.245 47.435 -37.915 47.765 ;
        RECT -38.245 46.075 -37.915 46.405 ;
        RECT -38.245 44.715 -37.915 45.045 ;
        RECT -38.245 43.355 -37.915 43.685 ;
        RECT -38.245 41.995 -37.915 42.325 ;
        RECT -38.245 40.635 -37.915 40.965 ;
        RECT -38.245 39.275 -37.915 39.605 ;
        RECT -38.245 37.915 -37.915 38.245 ;
        RECT -38.245 36.555 -37.915 36.885 ;
        RECT -38.245 35.195 -37.915 35.525 ;
        RECT -38.245 33.835 -37.915 34.165 ;
        RECT -38.245 32.475 -37.915 32.805 ;
        RECT -38.245 31.115 -37.915 31.445 ;
        RECT -38.245 29.755 -37.915 30.085 ;
        RECT -38.245 28.395 -37.915 28.725 ;
        RECT -38.245 27.035 -37.915 27.365 ;
        RECT -38.245 25.675 -37.915 26.005 ;
        RECT -38.245 24.315 -37.915 24.645 ;
        RECT -38.245 22.955 -37.915 23.285 ;
        RECT -38.245 21.595 -37.915 21.925 ;
        RECT -38.245 20.235 -37.915 20.565 ;
        RECT -38.245 18.875 -37.915 19.205 ;
        RECT -38.245 17.515 -37.915 17.845 ;
        RECT -38.245 16.155 -37.915 16.485 ;
        RECT -38.245 14.795 -37.915 15.125 ;
        RECT -38.245 13.435 -37.915 13.765 ;
        RECT -38.245 12.075 -37.915 12.405 ;
        RECT -38.245 10.715 -37.915 11.045 ;
        RECT -38.245 9.355 -37.915 9.685 ;
        RECT -38.245 7.995 -37.915 8.325 ;
        RECT -38.245 6.635 -37.915 6.965 ;
        RECT -38.245 5.275 -37.915 5.605 ;
        RECT -38.245 3.915 -37.915 4.245 ;
        RECT -38.245 2.555 -37.915 2.885 ;
        RECT -38.245 1.195 -37.915 1.525 ;
        RECT -38.245 -0.165 -37.915 0.165 ;
        RECT -38.245 -1.525 -37.915 -1.195 ;
        RECT -38.245 -8.325 -37.915 -7.995 ;
        RECT -38.245 -12.405 -37.915 -12.075 ;
        RECT -38.245 -13.765 -37.915 -13.435 ;
        RECT -38.245 -15.125 -37.915 -14.795 ;
        RECT -38.245 -16.485 -37.915 -16.155 ;
        RECT -38.245 -17.845 -37.915 -17.515 ;
        RECT -38.245 -19.205 -37.915 -18.875 ;
        RECT -38.245 -20.565 -37.915 -20.235 ;
        RECT -38.245 -21.925 -37.915 -21.595 ;
        RECT -38.245 -28.725 -37.915 -28.395 ;
        RECT -38.245 -30.085 -37.915 -29.755 ;
        RECT -38.245 -31.445 -37.915 -31.115 ;
        RECT -38.245 -32.805 -37.915 -32.475 ;
        RECT -38.245 -34.165 -37.915 -33.835 ;
        RECT -38.245 -35.525 -37.915 -35.195 ;
        RECT -38.245 -36.885 -37.915 -36.555 ;
        RECT -38.245 -38.245 -37.915 -37.915 ;
        RECT -38.245 -39.605 -37.915 -39.275 ;
        RECT -38.245 -40.965 -37.915 -40.635 ;
        RECT -38.245 -42.325 -37.915 -41.995 ;
        RECT -38.245 -43.685 -37.915 -43.355 ;
        RECT -38.245 -45.045 -37.915 -44.715 ;
        RECT -38.245 -47.765 -37.915 -47.435 ;
        RECT -38.245 -49.125 -37.915 -48.795 ;
        RECT -38.245 -50.485 -37.915 -50.155 ;
        RECT -38.245 -51.845 -37.915 -51.515 ;
        RECT -38.245 -53.205 -37.915 -52.875 ;
        RECT -38.245 -54.565 -37.915 -54.235 ;
        RECT -38.245 -55.925 -37.915 -55.595 ;
        RECT -38.245 -57.285 -37.915 -56.955 ;
        RECT -38.245 -58.645 -37.915 -58.315 ;
        RECT -38.245 -60.005 -37.915 -59.675 ;
        RECT -38.245 -61.365 -37.915 -61.035 ;
        RECT -38.245 -62.725 -37.915 -62.395 ;
        RECT -38.245 -64.085 -37.915 -63.755 ;
        RECT -38.245 -65.445 -37.915 -65.115 ;
        RECT -38.245 -66.805 -37.915 -66.475 ;
        RECT -38.245 -68.165 -37.915 -67.835 ;
        RECT -38.245 -69.525 -37.915 -69.195 ;
        RECT -38.245 -72.245 -37.915 -71.915 ;
        RECT -38.245 -73.605 -37.915 -73.275 ;
        RECT -38.245 -74.965 -37.915 -74.635 ;
        RECT -38.245 -76.325 -37.915 -75.995 ;
        RECT -38.245 -78.29 -37.915 -77.96 ;
        RECT -38.245 -79.045 -37.915 -78.715 ;
        RECT -38.245 -81.765 -37.915 -81.435 ;
        RECT -38.245 -83.125 -37.915 -82.795 ;
        RECT -38.245 -84.485 -37.915 -84.155 ;
        RECT -38.245 -86.43 -37.915 -86.1 ;
        RECT -38.245 -87.205 -37.915 -86.875 ;
        RECT -38.245 -88.565 -37.915 -88.235 ;
        RECT -38.245 -89.925 -37.915 -89.595 ;
        RECT -38.245 -92.645 -37.915 -92.315 ;
        RECT -38.245 -94.005 -37.915 -93.675 ;
        RECT -38.245 -95.365 -37.915 -95.035 ;
        RECT -38.245 -96.725 -37.915 -96.395 ;
        RECT -38.245 -98.085 -37.915 -97.755 ;
        RECT -38.245 -102.165 -37.915 -101.835 ;
        RECT -38.245 -103.525 -37.915 -103.195 ;
        RECT -38.245 -104.885 -37.915 -104.555 ;
        RECT -38.245 -106.245 -37.915 -105.915 ;
        RECT -38.245 -107.605 -37.915 -107.275 ;
        RECT -38.245 -108.965 -37.915 -108.635 ;
        RECT -38.245 -113.045 -37.915 -112.715 ;
        RECT -38.245 -114.405 -37.915 -114.075 ;
        RECT -38.245 -115.765 -37.915 -115.435 ;
        RECT -38.245 -117.125 -37.915 -116.795 ;
        RECT -38.245 -118.485 -37.915 -118.155 ;
        RECT -38.245 -119.845 -37.915 -119.515 ;
        RECT -38.245 -121.205 -37.915 -120.875 ;
        RECT -38.245 -122.565 -37.915 -122.235 ;
        RECT -38.245 -123.925 -37.915 -123.595 ;
        RECT -38.245 -125.285 -37.915 -124.955 ;
        RECT -38.245 -126.645 -37.915 -126.315 ;
        RECT -38.245 -128.005 -37.915 -127.675 ;
        RECT -38.245 -130.725 -37.915 -130.395 ;
        RECT -38.245 -132.085 -37.915 -131.755 ;
        RECT -38.245 -134.805 -37.915 -134.475 ;
        RECT -38.245 -136.165 -37.915 -135.835 ;
        RECT -38.245 -137.525 -37.915 -137.195 ;
        RECT -38.245 -138.885 -37.915 -138.555 ;
        RECT -38.245 -140.245 -37.915 -139.915 ;
        RECT -38.245 -141.605 -37.915 -141.275 ;
        RECT -38.245 -142.965 -37.915 -142.635 ;
        RECT -38.245 -144.325 -37.915 -143.995 ;
        RECT -38.245 -145.685 -37.915 -145.355 ;
        RECT -38.245 -147.045 -37.915 -146.715 ;
        RECT -38.245 -149.765 -37.915 -149.435 ;
        RECT -38.245 -152.485 -37.915 -152.155 ;
        RECT -38.245 -153.845 -37.915 -153.515 ;
        RECT -38.245 -155.285 -37.915 -154.955 ;
        RECT -38.245 -156.565 -37.915 -156.235 ;
        RECT -38.245 -157.925 -37.915 -157.595 ;
        RECT -38.245 -160.17 -37.915 -159.04 ;
        RECT -38.24 -160.285 -37.92 128.47 ;
        RECT -38.245 127.225 -37.915 128.355 ;
        RECT -38.245 124.955 -37.915 125.285 ;
        RECT -38.245 123.595 -37.915 123.925 ;
        RECT -38.245 122.235 -37.915 122.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 127.225 -51.515 128.355 ;
        RECT -51.845 124.955 -51.515 125.285 ;
        RECT -51.845 123.595 -51.515 123.925 ;
        RECT -51.845 122.235 -51.515 122.565 ;
        RECT -51.845 120.875 -51.515 121.205 ;
        RECT -51.845 119.515 -51.515 119.845 ;
        RECT -51.845 118.155 -51.515 118.485 ;
        RECT -51.845 116.795 -51.515 117.125 ;
        RECT -51.845 115.435 -51.515 115.765 ;
        RECT -51.845 114.075 -51.515 114.405 ;
        RECT -51.845 112.715 -51.515 113.045 ;
        RECT -51.845 111.355 -51.515 111.685 ;
        RECT -51.845 109.995 -51.515 110.325 ;
        RECT -51.845 108.635 -51.515 108.965 ;
        RECT -51.845 107.275 -51.515 107.605 ;
        RECT -51.845 105.915 -51.515 106.245 ;
        RECT -51.845 104.555 -51.515 104.885 ;
        RECT -51.845 103.195 -51.515 103.525 ;
        RECT -51.845 101.835 -51.515 102.165 ;
        RECT -51.845 100.475 -51.515 100.805 ;
        RECT -51.845 99.115 -51.515 99.445 ;
        RECT -51.845 97.755 -51.515 98.085 ;
        RECT -51.845 96.395 -51.515 96.725 ;
        RECT -51.845 95.035 -51.515 95.365 ;
        RECT -51.845 93.675 -51.515 94.005 ;
        RECT -51.845 92.315 -51.515 92.645 ;
        RECT -51.845 90.955 -51.515 91.285 ;
        RECT -51.845 89.595 -51.515 89.925 ;
        RECT -51.845 88.235 -51.515 88.565 ;
        RECT -51.845 86.875 -51.515 87.205 ;
        RECT -51.845 85.515 -51.515 85.845 ;
        RECT -51.845 84.155 -51.515 84.485 ;
        RECT -51.845 82.795 -51.515 83.125 ;
        RECT -51.845 81.435 -51.515 81.765 ;
        RECT -51.845 80.075 -51.515 80.405 ;
        RECT -51.845 78.715 -51.515 79.045 ;
        RECT -51.845 77.355 -51.515 77.685 ;
        RECT -51.845 75.995 -51.515 76.325 ;
        RECT -51.845 74.635 -51.515 74.965 ;
        RECT -51.845 73.275 -51.515 73.605 ;
        RECT -51.84 73.275 -51.52 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 48.795 -51.515 49.125 ;
        RECT -51.845 47.435 -51.515 47.765 ;
        RECT -51.845 46.075 -51.515 46.405 ;
        RECT -51.845 44.715 -51.515 45.045 ;
        RECT -51.845 43.355 -51.515 43.685 ;
        RECT -51.845 40.635 -51.515 40.965 ;
        RECT -51.845 39.275 -51.515 39.605 ;
        RECT -51.845 35.195 -51.515 35.525 ;
        RECT -51.845 33.835 -51.515 34.165 ;
        RECT -51.845 32.475 -51.515 32.805 ;
        RECT -51.845 31.115 -51.515 31.445 ;
        RECT -51.845 29.755 -51.515 30.085 ;
        RECT -51.845 28.395 -51.515 28.725 ;
        RECT -51.845 27.035 -51.515 27.365 ;
        RECT -51.845 25.675 -51.515 26.005 ;
        RECT -51.845 24.315 -51.515 24.645 ;
        RECT -51.845 22.955 -51.515 23.285 ;
        RECT -51.845 21.595 -51.515 21.925 ;
        RECT -51.845 20.235 -51.515 20.565 ;
        RECT -51.845 18.875 -51.515 19.205 ;
        RECT -51.845 17.515 -51.515 17.845 ;
        RECT -51.845 16.155 -51.515 16.485 ;
        RECT -51.845 14.795 -51.515 15.125 ;
        RECT -51.845 13.435 -51.515 13.765 ;
        RECT -51.845 12.075 -51.515 12.405 ;
        RECT -51.845 10.715 -51.515 11.045 ;
        RECT -51.845 9.355 -51.515 9.685 ;
        RECT -51.845 7.995 -51.515 8.325 ;
        RECT -51.845 6.635 -51.515 6.965 ;
        RECT -51.845 5.275 -51.515 5.605 ;
        RECT -51.845 3.915 -51.515 4.245 ;
        RECT -51.845 2.555 -51.515 2.885 ;
        RECT -51.845 1.195 -51.515 1.525 ;
        RECT -51.845 -0.165 -51.515 0.165 ;
        RECT -51.845 -1.525 -51.515 -1.195 ;
        RECT -51.845 -2.885 -51.515 -2.555 ;
        RECT -51.845 -4.245 -51.515 -3.915 ;
        RECT -51.845 -5.605 -51.515 -5.275 ;
        RECT -51.845 -6.965 -51.515 -6.635 ;
        RECT -51.845 -8.325 -51.515 -7.995 ;
        RECT -51.845 -9.685 -51.515 -9.355 ;
        RECT -51.845 -12.405 -51.515 -12.075 ;
        RECT -51.845 -13.765 -51.515 -13.435 ;
        RECT -51.845 -15.125 -51.515 -14.795 ;
        RECT -51.845 -16.485 -51.515 -16.155 ;
        RECT -51.845 -17.845 -51.515 -17.515 ;
        RECT -51.845 -19.205 -51.515 -18.875 ;
        RECT -51.845 -20.565 -51.515 -20.235 ;
        RECT -51.845 -21.925 -51.515 -21.595 ;
        RECT -51.845 -24.645 -51.515 -24.315 ;
        RECT -51.845 -26.005 -51.515 -25.675 ;
        RECT -51.845 -27.365 -51.515 -27.035 ;
        RECT -51.845 -28.725 -51.515 -28.395 ;
        RECT -51.845 -30.085 -51.515 -29.755 ;
        RECT -51.845 -31.445 -51.515 -31.115 ;
        RECT -51.845 -32.805 -51.515 -32.475 ;
        RECT -51.845 -34.165 -51.515 -33.835 ;
        RECT -51.845 -35.525 -51.515 -35.195 ;
        RECT -51.845 -36.885 -51.515 -36.555 ;
        RECT -51.845 -38.245 -51.515 -37.915 ;
        RECT -51.845 -39.605 -51.515 -39.275 ;
        RECT -51.845 -40.965 -51.515 -40.635 ;
        RECT -51.845 -42.325 -51.515 -41.995 ;
        RECT -51.845 -43.685 -51.515 -43.355 ;
        RECT -51.845 -45.045 -51.515 -44.715 ;
        RECT -51.845 -46.405 -51.515 -46.075 ;
        RECT -51.845 -47.765 -51.515 -47.435 ;
        RECT -51.845 -49.125 -51.515 -48.795 ;
        RECT -51.845 -50.485 -51.515 -50.155 ;
        RECT -51.845 -51.845 -51.515 -51.515 ;
        RECT -51.845 -53.205 -51.515 -52.875 ;
        RECT -51.845 -54.565 -51.515 -54.235 ;
        RECT -51.845 -55.925 -51.515 -55.595 ;
        RECT -51.845 -57.285 -51.515 -56.955 ;
        RECT -51.845 -58.645 -51.515 -58.315 ;
        RECT -51.845 -60.005 -51.515 -59.675 ;
        RECT -51.845 -61.365 -51.515 -61.035 ;
        RECT -51.845 -62.725 -51.515 -62.395 ;
        RECT -51.845 -64.085 -51.515 -63.755 ;
        RECT -51.845 -65.445 -51.515 -65.115 ;
        RECT -51.845 -66.805 -51.515 -66.475 ;
        RECT -51.845 -68.165 -51.515 -67.835 ;
        RECT -51.845 -69.525 -51.515 -69.195 ;
        RECT -51.845 -72.245 -51.515 -71.915 ;
        RECT -51.845 -73.605 -51.515 -73.275 ;
        RECT -51.845 -74.965 -51.515 -74.635 ;
        RECT -51.845 -76.325 -51.515 -75.995 ;
        RECT -51.845 -78.29 -51.515 -77.96 ;
        RECT -51.845 -79.045 -51.515 -78.715 ;
        RECT -51.845 -81.765 -51.515 -81.435 ;
        RECT -51.845 -83.125 -51.515 -82.795 ;
        RECT -51.845 -84.485 -51.515 -84.155 ;
        RECT -51.845 -86.43 -51.515 -86.1 ;
        RECT -51.845 -87.205 -51.515 -86.875 ;
        RECT -51.845 -88.565 -51.515 -88.235 ;
        RECT -51.845 -89.925 -51.515 -89.595 ;
        RECT -51.845 -92.645 -51.515 -92.315 ;
        RECT -51.845 -94.005 -51.515 -93.675 ;
        RECT -51.845 -95.365 -51.515 -95.035 ;
        RECT -51.845 -96.725 -51.515 -96.395 ;
        RECT -51.845 -98.085 -51.515 -97.755 ;
        RECT -51.845 -102.165 -51.515 -101.835 ;
        RECT -51.845 -103.525 -51.515 -103.195 ;
        RECT -51.845 -104.885 -51.515 -104.555 ;
        RECT -51.845 -106.245 -51.515 -105.915 ;
        RECT -51.845 -107.605 -51.515 -107.275 ;
        RECT -51.845 -108.965 -51.515 -108.635 ;
        RECT -51.845 -110.325 -51.515 -109.995 ;
        RECT -51.845 -111.685 -51.515 -111.355 ;
        RECT -51.845 -113.045 -51.515 -112.715 ;
        RECT -51.845 -114.405 -51.515 -114.075 ;
        RECT -51.845 -115.765 -51.515 -115.435 ;
        RECT -51.845 -117.125 -51.515 -116.795 ;
        RECT -51.845 -118.485 -51.515 -118.155 ;
        RECT -51.845 -119.845 -51.515 -119.515 ;
        RECT -51.845 -121.205 -51.515 -120.875 ;
        RECT -51.845 -122.565 -51.515 -122.235 ;
        RECT -51.845 -123.925 -51.515 -123.595 ;
        RECT -51.845 -125.285 -51.515 -124.955 ;
        RECT -51.845 -126.645 -51.515 -126.315 ;
        RECT -51.845 -128.005 -51.515 -127.675 ;
        RECT -51.845 -129.365 -51.515 -129.035 ;
        RECT -51.845 -130.725 -51.515 -130.395 ;
        RECT -51.845 -132.085 -51.515 -131.755 ;
        RECT -51.845 -133.445 -51.515 -133.115 ;
        RECT -51.845 -134.805 -51.515 -134.475 ;
        RECT -51.845 -136.165 -51.515 -135.835 ;
        RECT -51.845 -137.525 -51.515 -137.195 ;
        RECT -51.845 -138.885 -51.515 -138.555 ;
        RECT -51.845 -140.245 -51.515 -139.915 ;
        RECT -51.845 -141.605 -51.515 -141.275 ;
        RECT -51.845 -142.965 -51.515 -142.635 ;
        RECT -51.845 -144.325 -51.515 -143.995 ;
        RECT -51.845 -145.685 -51.515 -145.355 ;
        RECT -51.845 -147.045 -51.515 -146.715 ;
        RECT -51.845 -149.765 -51.515 -149.435 ;
        RECT -51.845 -153.845 -51.515 -153.515 ;
        RECT -51.845 -155.285 -51.515 -154.955 ;
        RECT -51.845 -156.565 -51.515 -156.235 ;
        RECT -51.845 -157.925 -51.515 -157.595 ;
        RECT -51.845 -160.17 -51.515 -159.04 ;
        RECT -51.84 -160.285 -51.52 49.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 127.225 -50.155 128.355 ;
        RECT -50.485 124.955 -50.155 125.285 ;
        RECT -50.485 123.595 -50.155 123.925 ;
        RECT -50.485 122.235 -50.155 122.565 ;
        RECT -50.485 120.875 -50.155 121.205 ;
        RECT -50.485 119.515 -50.155 119.845 ;
        RECT -50.485 118.155 -50.155 118.485 ;
        RECT -50.485 116.795 -50.155 117.125 ;
        RECT -50.485 115.435 -50.155 115.765 ;
        RECT -50.485 114.075 -50.155 114.405 ;
        RECT -50.485 112.715 -50.155 113.045 ;
        RECT -50.485 111.355 -50.155 111.685 ;
        RECT -50.485 109.995 -50.155 110.325 ;
        RECT -50.485 108.635 -50.155 108.965 ;
        RECT -50.485 107.275 -50.155 107.605 ;
        RECT -50.485 105.915 -50.155 106.245 ;
        RECT -50.485 104.555 -50.155 104.885 ;
        RECT -50.485 103.195 -50.155 103.525 ;
        RECT -50.485 101.835 -50.155 102.165 ;
        RECT -50.485 100.475 -50.155 100.805 ;
        RECT -50.485 99.115 -50.155 99.445 ;
        RECT -50.485 97.755 -50.155 98.085 ;
        RECT -50.485 96.395 -50.155 96.725 ;
        RECT -50.485 95.035 -50.155 95.365 ;
        RECT -50.485 93.675 -50.155 94.005 ;
        RECT -50.485 92.315 -50.155 92.645 ;
        RECT -50.485 90.955 -50.155 91.285 ;
        RECT -50.485 89.595 -50.155 89.925 ;
        RECT -50.485 88.235 -50.155 88.565 ;
        RECT -50.485 86.875 -50.155 87.205 ;
        RECT -50.485 85.515 -50.155 85.845 ;
        RECT -50.485 84.155 -50.155 84.485 ;
        RECT -50.485 82.795 -50.155 83.125 ;
        RECT -50.485 81.435 -50.155 81.765 ;
        RECT -50.485 80.075 -50.155 80.405 ;
        RECT -50.485 78.715 -50.155 79.045 ;
        RECT -50.485 77.355 -50.155 77.685 ;
        RECT -50.485 75.995 -50.155 76.325 ;
        RECT -50.485 74.635 -50.155 74.965 ;
        RECT -50.485 73.275 -50.155 73.605 ;
        RECT -50.48 73.275 -50.16 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 48.795 -50.155 49.125 ;
        RECT -50.485 47.435 -50.155 47.765 ;
        RECT -50.485 46.075 -50.155 46.405 ;
        RECT -50.485 44.715 -50.155 45.045 ;
        RECT -50.485 43.355 -50.155 43.685 ;
        RECT -50.485 40.635 -50.155 40.965 ;
        RECT -50.485 39.275 -50.155 39.605 ;
        RECT -50.485 35.195 -50.155 35.525 ;
        RECT -50.485 33.835 -50.155 34.165 ;
        RECT -50.485 32.475 -50.155 32.805 ;
        RECT -50.485 31.115 -50.155 31.445 ;
        RECT -50.485 29.755 -50.155 30.085 ;
        RECT -50.485 28.395 -50.155 28.725 ;
        RECT -50.485 27.035 -50.155 27.365 ;
        RECT -50.485 25.675 -50.155 26.005 ;
        RECT -50.485 24.315 -50.155 24.645 ;
        RECT -50.485 22.955 -50.155 23.285 ;
        RECT -50.485 21.595 -50.155 21.925 ;
        RECT -50.485 20.235 -50.155 20.565 ;
        RECT -50.485 18.875 -50.155 19.205 ;
        RECT -50.485 17.515 -50.155 17.845 ;
        RECT -50.485 16.155 -50.155 16.485 ;
        RECT -50.485 14.795 -50.155 15.125 ;
        RECT -50.485 13.435 -50.155 13.765 ;
        RECT -50.485 12.075 -50.155 12.405 ;
        RECT -50.485 10.715 -50.155 11.045 ;
        RECT -50.485 9.355 -50.155 9.685 ;
        RECT -50.485 7.995 -50.155 8.325 ;
        RECT -50.485 6.635 -50.155 6.965 ;
        RECT -50.485 5.275 -50.155 5.605 ;
        RECT -50.485 3.915 -50.155 4.245 ;
        RECT -50.485 2.555 -50.155 2.885 ;
        RECT -50.485 1.195 -50.155 1.525 ;
        RECT -50.485 -0.165 -50.155 0.165 ;
        RECT -50.485 -1.525 -50.155 -1.195 ;
        RECT -50.485 -2.885 -50.155 -2.555 ;
        RECT -50.485 -4.245 -50.155 -3.915 ;
        RECT -50.485 -5.605 -50.155 -5.275 ;
        RECT -50.485 -6.965 -50.155 -6.635 ;
        RECT -50.485 -8.325 -50.155 -7.995 ;
        RECT -50.485 -9.685 -50.155 -9.355 ;
        RECT -50.485 -12.405 -50.155 -12.075 ;
        RECT -50.485 -13.765 -50.155 -13.435 ;
        RECT -50.485 -15.125 -50.155 -14.795 ;
        RECT -50.485 -16.485 -50.155 -16.155 ;
        RECT -50.485 -17.845 -50.155 -17.515 ;
        RECT -50.485 -19.205 -50.155 -18.875 ;
        RECT -50.485 -20.565 -50.155 -20.235 ;
        RECT -50.485 -21.925 -50.155 -21.595 ;
        RECT -50.485 -24.645 -50.155 -24.315 ;
        RECT -50.485 -26.005 -50.155 -25.675 ;
        RECT -50.485 -27.365 -50.155 -27.035 ;
        RECT -50.485 -28.725 -50.155 -28.395 ;
        RECT -50.485 -30.085 -50.155 -29.755 ;
        RECT -50.485 -31.445 -50.155 -31.115 ;
        RECT -50.485 -32.805 -50.155 -32.475 ;
        RECT -50.485 -34.165 -50.155 -33.835 ;
        RECT -50.485 -35.525 -50.155 -35.195 ;
        RECT -50.485 -36.885 -50.155 -36.555 ;
        RECT -50.485 -38.245 -50.155 -37.915 ;
        RECT -50.485 -39.605 -50.155 -39.275 ;
        RECT -50.485 -40.965 -50.155 -40.635 ;
        RECT -50.485 -42.325 -50.155 -41.995 ;
        RECT -50.485 -43.685 -50.155 -43.355 ;
        RECT -50.485 -45.045 -50.155 -44.715 ;
        RECT -50.485 -46.405 -50.155 -46.075 ;
        RECT -50.485 -47.765 -50.155 -47.435 ;
        RECT -50.485 -49.125 -50.155 -48.795 ;
        RECT -50.485 -50.485 -50.155 -50.155 ;
        RECT -50.485 -51.845 -50.155 -51.515 ;
        RECT -50.485 -53.205 -50.155 -52.875 ;
        RECT -50.485 -54.565 -50.155 -54.235 ;
        RECT -50.485 -55.925 -50.155 -55.595 ;
        RECT -50.485 -57.285 -50.155 -56.955 ;
        RECT -50.485 -58.645 -50.155 -58.315 ;
        RECT -50.485 -60.005 -50.155 -59.675 ;
        RECT -50.485 -61.365 -50.155 -61.035 ;
        RECT -50.485 -62.725 -50.155 -62.395 ;
        RECT -50.485 -64.085 -50.155 -63.755 ;
        RECT -50.485 -65.445 -50.155 -65.115 ;
        RECT -50.485 -66.805 -50.155 -66.475 ;
        RECT -50.485 -68.165 -50.155 -67.835 ;
        RECT -50.485 -69.525 -50.155 -69.195 ;
        RECT -50.485 -72.245 -50.155 -71.915 ;
        RECT -50.485 -73.605 -50.155 -73.275 ;
        RECT -50.485 -74.965 -50.155 -74.635 ;
        RECT -50.485 -76.325 -50.155 -75.995 ;
        RECT -50.485 -78.29 -50.155 -77.96 ;
        RECT -50.485 -79.045 -50.155 -78.715 ;
        RECT -50.485 -81.765 -50.155 -81.435 ;
        RECT -50.485 -83.125 -50.155 -82.795 ;
        RECT -50.485 -84.485 -50.155 -84.155 ;
        RECT -50.485 -86.43 -50.155 -86.1 ;
        RECT -50.485 -87.205 -50.155 -86.875 ;
        RECT -50.485 -88.565 -50.155 -88.235 ;
        RECT -50.485 -89.925 -50.155 -89.595 ;
        RECT -50.485 -92.645 -50.155 -92.315 ;
        RECT -50.485 -94.005 -50.155 -93.675 ;
        RECT -50.485 -95.365 -50.155 -95.035 ;
        RECT -50.485 -96.725 -50.155 -96.395 ;
        RECT -50.485 -98.085 -50.155 -97.755 ;
        RECT -50.485 -102.165 -50.155 -101.835 ;
        RECT -50.485 -103.525 -50.155 -103.195 ;
        RECT -50.485 -104.885 -50.155 -104.555 ;
        RECT -50.485 -106.245 -50.155 -105.915 ;
        RECT -50.485 -107.605 -50.155 -107.275 ;
        RECT -50.485 -108.965 -50.155 -108.635 ;
        RECT -50.485 -110.325 -50.155 -109.995 ;
        RECT -50.485 -111.685 -50.155 -111.355 ;
        RECT -50.485 -113.045 -50.155 -112.715 ;
        RECT -50.485 -114.405 -50.155 -114.075 ;
        RECT -50.485 -115.765 -50.155 -115.435 ;
        RECT -50.485 -117.125 -50.155 -116.795 ;
        RECT -50.485 -118.485 -50.155 -118.155 ;
        RECT -50.485 -119.845 -50.155 -119.515 ;
        RECT -50.485 -121.205 -50.155 -120.875 ;
        RECT -50.485 -122.565 -50.155 -122.235 ;
        RECT -50.485 -123.925 -50.155 -123.595 ;
        RECT -50.485 -125.285 -50.155 -124.955 ;
        RECT -50.485 -126.645 -50.155 -126.315 ;
        RECT -50.485 -128.005 -50.155 -127.675 ;
        RECT -50.485 -129.365 -50.155 -129.035 ;
        RECT -50.485 -130.725 -50.155 -130.395 ;
        RECT -50.485 -132.085 -50.155 -131.755 ;
        RECT -50.485 -133.445 -50.155 -133.115 ;
        RECT -50.485 -134.805 -50.155 -134.475 ;
        RECT -50.485 -136.165 -50.155 -135.835 ;
        RECT -50.485 -137.525 -50.155 -137.195 ;
        RECT -50.485 -138.885 -50.155 -138.555 ;
        RECT -50.485 -140.245 -50.155 -139.915 ;
        RECT -50.485 -141.605 -50.155 -141.275 ;
        RECT -50.485 -142.965 -50.155 -142.635 ;
        RECT -50.485 -144.325 -50.155 -143.995 ;
        RECT -50.485 -145.685 -50.155 -145.355 ;
        RECT -50.485 -147.045 -50.155 -146.715 ;
        RECT -50.485 -149.765 -50.155 -149.435 ;
        RECT -50.485 -152.485 -50.155 -152.155 ;
        RECT -50.485 -153.845 -50.155 -153.515 ;
        RECT -50.485 -155.285 -50.155 -154.955 ;
        RECT -50.485 -156.565 -50.155 -156.235 ;
        RECT -50.485 -157.925 -50.155 -157.595 ;
        RECT -50.485 -160.17 -50.155 -159.04 ;
        RECT -50.48 -160.285 -50.16 49.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 127.225 -48.795 128.355 ;
        RECT -49.125 124.955 -48.795 125.285 ;
        RECT -49.125 123.595 -48.795 123.925 ;
        RECT -49.125 122.235 -48.795 122.565 ;
        RECT -49.125 120.875 -48.795 121.205 ;
        RECT -49.125 119.515 -48.795 119.845 ;
        RECT -49.125 118.155 -48.795 118.485 ;
        RECT -49.125 116.795 -48.795 117.125 ;
        RECT -49.125 115.435 -48.795 115.765 ;
        RECT -49.125 114.075 -48.795 114.405 ;
        RECT -49.125 112.715 -48.795 113.045 ;
        RECT -49.125 111.355 -48.795 111.685 ;
        RECT -49.125 109.995 -48.795 110.325 ;
        RECT -49.125 108.635 -48.795 108.965 ;
        RECT -49.125 107.275 -48.795 107.605 ;
        RECT -49.125 105.915 -48.795 106.245 ;
        RECT -49.125 104.555 -48.795 104.885 ;
        RECT -49.125 103.195 -48.795 103.525 ;
        RECT -49.125 101.835 -48.795 102.165 ;
        RECT -49.125 100.475 -48.795 100.805 ;
        RECT -49.125 99.115 -48.795 99.445 ;
        RECT -49.125 97.755 -48.795 98.085 ;
        RECT -49.125 96.395 -48.795 96.725 ;
        RECT -49.125 95.035 -48.795 95.365 ;
        RECT -49.125 93.675 -48.795 94.005 ;
        RECT -49.125 92.315 -48.795 92.645 ;
        RECT -49.125 90.955 -48.795 91.285 ;
        RECT -49.125 89.595 -48.795 89.925 ;
        RECT -49.125 88.235 -48.795 88.565 ;
        RECT -49.125 86.875 -48.795 87.205 ;
        RECT -49.125 85.515 -48.795 85.845 ;
        RECT -49.125 84.155 -48.795 84.485 ;
        RECT -49.125 82.795 -48.795 83.125 ;
        RECT -49.125 81.435 -48.795 81.765 ;
        RECT -49.125 80.075 -48.795 80.405 ;
        RECT -49.125 78.715 -48.795 79.045 ;
        RECT -49.125 77.355 -48.795 77.685 ;
        RECT -49.125 75.995 -48.795 76.325 ;
        RECT -49.125 74.635 -48.795 74.965 ;
        RECT -49.125 73.275 -48.795 73.605 ;
        RECT -49.12 73.275 -48.8 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 48.795 -48.795 49.125 ;
        RECT -49.125 47.435 -48.795 47.765 ;
        RECT -49.125 46.075 -48.795 46.405 ;
        RECT -49.125 44.715 -48.795 45.045 ;
        RECT -49.125 43.355 -48.795 43.685 ;
        RECT -49.125 40.635 -48.795 40.965 ;
        RECT -49.125 39.275 -48.795 39.605 ;
        RECT -49.125 35.195 -48.795 35.525 ;
        RECT -49.125 33.835 -48.795 34.165 ;
        RECT -49.125 32.475 -48.795 32.805 ;
        RECT -49.125 31.115 -48.795 31.445 ;
        RECT -49.125 29.755 -48.795 30.085 ;
        RECT -49.125 28.395 -48.795 28.725 ;
        RECT -49.125 27.035 -48.795 27.365 ;
        RECT -49.125 25.675 -48.795 26.005 ;
        RECT -49.125 24.315 -48.795 24.645 ;
        RECT -49.125 22.955 -48.795 23.285 ;
        RECT -49.125 21.595 -48.795 21.925 ;
        RECT -49.125 20.235 -48.795 20.565 ;
        RECT -49.125 18.875 -48.795 19.205 ;
        RECT -49.125 17.515 -48.795 17.845 ;
        RECT -49.125 16.155 -48.795 16.485 ;
        RECT -49.125 14.795 -48.795 15.125 ;
        RECT -49.125 13.435 -48.795 13.765 ;
        RECT -49.125 12.075 -48.795 12.405 ;
        RECT -49.125 10.715 -48.795 11.045 ;
        RECT -49.125 9.355 -48.795 9.685 ;
        RECT -49.125 7.995 -48.795 8.325 ;
        RECT -49.125 6.635 -48.795 6.965 ;
        RECT -49.125 5.275 -48.795 5.605 ;
        RECT -49.125 3.915 -48.795 4.245 ;
        RECT -49.125 2.555 -48.795 2.885 ;
        RECT -49.125 1.195 -48.795 1.525 ;
        RECT -49.125 -0.165 -48.795 0.165 ;
        RECT -49.125 -1.525 -48.795 -1.195 ;
        RECT -49.125 -2.885 -48.795 -2.555 ;
        RECT -49.125 -4.245 -48.795 -3.915 ;
        RECT -49.125 -5.605 -48.795 -5.275 ;
        RECT -49.125 -6.965 -48.795 -6.635 ;
        RECT -49.125 -8.325 -48.795 -7.995 ;
        RECT -49.125 -9.685 -48.795 -9.355 ;
        RECT -49.125 -12.405 -48.795 -12.075 ;
        RECT -49.125 -13.765 -48.795 -13.435 ;
        RECT -49.125 -15.125 -48.795 -14.795 ;
        RECT -49.125 -16.485 -48.795 -16.155 ;
        RECT -49.125 -17.845 -48.795 -17.515 ;
        RECT -49.125 -19.205 -48.795 -18.875 ;
        RECT -49.125 -20.565 -48.795 -20.235 ;
        RECT -49.125 -21.925 -48.795 -21.595 ;
        RECT -49.125 -26.005 -48.795 -25.675 ;
        RECT -49.125 -27.365 -48.795 -27.035 ;
        RECT -49.125 -28.725 -48.795 -28.395 ;
        RECT -49.125 -30.085 -48.795 -29.755 ;
        RECT -49.125 -31.445 -48.795 -31.115 ;
        RECT -49.125 -32.805 -48.795 -32.475 ;
        RECT -49.125 -34.165 -48.795 -33.835 ;
        RECT -49.125 -35.525 -48.795 -35.195 ;
        RECT -49.125 -36.885 -48.795 -36.555 ;
        RECT -49.125 -38.245 -48.795 -37.915 ;
        RECT -49.125 -39.605 -48.795 -39.275 ;
        RECT -49.125 -40.965 -48.795 -40.635 ;
        RECT -49.125 -42.325 -48.795 -41.995 ;
        RECT -49.125 -43.685 -48.795 -43.355 ;
        RECT -49.125 -45.045 -48.795 -44.715 ;
        RECT -49.125 -46.405 -48.795 -46.075 ;
        RECT -49.125 -47.765 -48.795 -47.435 ;
        RECT -49.125 -49.125 -48.795 -48.795 ;
        RECT -49.125 -50.485 -48.795 -50.155 ;
        RECT -49.125 -51.845 -48.795 -51.515 ;
        RECT -49.125 -53.205 -48.795 -52.875 ;
        RECT -49.125 -54.565 -48.795 -54.235 ;
        RECT -49.125 -55.925 -48.795 -55.595 ;
        RECT -49.125 -57.285 -48.795 -56.955 ;
        RECT -49.125 -58.645 -48.795 -58.315 ;
        RECT -49.125 -60.005 -48.795 -59.675 ;
        RECT -49.125 -61.365 -48.795 -61.035 ;
        RECT -49.125 -62.725 -48.795 -62.395 ;
        RECT -49.125 -64.085 -48.795 -63.755 ;
        RECT -49.125 -65.445 -48.795 -65.115 ;
        RECT -49.125 -66.805 -48.795 -66.475 ;
        RECT -49.125 -68.165 -48.795 -67.835 ;
        RECT -49.125 -69.525 -48.795 -69.195 ;
        RECT -49.125 -72.245 -48.795 -71.915 ;
        RECT -49.125 -73.605 -48.795 -73.275 ;
        RECT -49.125 -74.965 -48.795 -74.635 ;
        RECT -49.125 -76.325 -48.795 -75.995 ;
        RECT -49.125 -78.29 -48.795 -77.96 ;
        RECT -49.125 -79.045 -48.795 -78.715 ;
        RECT -49.125 -81.765 -48.795 -81.435 ;
        RECT -49.125 -83.125 -48.795 -82.795 ;
        RECT -49.125 -84.485 -48.795 -84.155 ;
        RECT -49.125 -86.43 -48.795 -86.1 ;
        RECT -49.125 -87.205 -48.795 -86.875 ;
        RECT -49.125 -88.565 -48.795 -88.235 ;
        RECT -49.125 -89.925 -48.795 -89.595 ;
        RECT -49.12 -91.28 -48.8 49.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 -153.845 -48.795 -153.515 ;
        RECT -49.125 -155.285 -48.795 -154.955 ;
        RECT -49.125 -156.565 -48.795 -156.235 ;
        RECT -49.125 -157.925 -48.795 -157.595 ;
        RECT -49.125 -160.17 -48.795 -159.04 ;
        RECT -49.12 -160.285 -48.8 -153.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 127.225 -47.435 128.355 ;
        RECT -47.765 124.955 -47.435 125.285 ;
        RECT -47.765 123.595 -47.435 123.925 ;
        RECT -47.765 122.235 -47.435 122.565 ;
        RECT -47.765 120.875 -47.435 121.205 ;
        RECT -47.765 119.515 -47.435 119.845 ;
        RECT -47.765 118.155 -47.435 118.485 ;
        RECT -47.765 116.795 -47.435 117.125 ;
        RECT -47.765 115.435 -47.435 115.765 ;
        RECT -47.765 114.075 -47.435 114.405 ;
        RECT -47.765 112.715 -47.435 113.045 ;
        RECT -47.765 111.355 -47.435 111.685 ;
        RECT -47.765 109.995 -47.435 110.325 ;
        RECT -47.765 108.635 -47.435 108.965 ;
        RECT -47.765 107.275 -47.435 107.605 ;
        RECT -47.765 105.915 -47.435 106.245 ;
        RECT -47.765 104.555 -47.435 104.885 ;
        RECT -47.765 103.195 -47.435 103.525 ;
        RECT -47.765 101.835 -47.435 102.165 ;
        RECT -47.765 100.475 -47.435 100.805 ;
        RECT -47.765 99.115 -47.435 99.445 ;
        RECT -47.765 97.755 -47.435 98.085 ;
        RECT -47.765 96.395 -47.435 96.725 ;
        RECT -47.765 95.035 -47.435 95.365 ;
        RECT -47.765 93.675 -47.435 94.005 ;
        RECT -47.765 92.315 -47.435 92.645 ;
        RECT -47.765 90.955 -47.435 91.285 ;
        RECT -47.765 89.595 -47.435 89.925 ;
        RECT -47.765 88.235 -47.435 88.565 ;
        RECT -47.765 86.875 -47.435 87.205 ;
        RECT -47.765 85.515 -47.435 85.845 ;
        RECT -47.765 84.155 -47.435 84.485 ;
        RECT -47.765 82.795 -47.435 83.125 ;
        RECT -47.765 81.435 -47.435 81.765 ;
        RECT -47.765 80.075 -47.435 80.405 ;
        RECT -47.765 78.715 -47.435 79.045 ;
        RECT -47.765 77.355 -47.435 77.685 ;
        RECT -47.765 75.995 -47.435 76.325 ;
        RECT -47.765 74.635 -47.435 74.965 ;
        RECT -47.765 73.275 -47.435 73.605 ;
        RECT -47.765 72.445 -47.435 72.775 ;
        RECT -47.765 70.395 -47.435 70.725 ;
        RECT -47.765 68.035 -47.435 68.365 ;
        RECT -47.765 66.885 -47.435 67.215 ;
        RECT -47.765 64.875 -47.435 65.205 ;
        RECT -47.765 63.725 -47.435 64.055 ;
        RECT -47.765 61.715 -47.435 62.045 ;
        RECT -47.765 60.395 -47.435 60.725 ;
        RECT -47.765 58.555 -47.435 58.885 ;
        RECT -47.765 57.405 -47.435 57.735 ;
        RECT -47.765 55.395 -47.435 55.725 ;
        RECT -47.765 54.245 -47.435 54.575 ;
        RECT -47.765 51.885 -47.435 52.215 ;
        RECT -47.765 49.83 -47.435 50.16 ;
        RECT -47.765 48.795 -47.435 49.125 ;
        RECT -47.765 47.435 -47.435 47.765 ;
        RECT -47.765 46.075 -47.435 46.405 ;
        RECT -47.765 44.715 -47.435 45.045 ;
        RECT -47.765 43.355 -47.435 43.685 ;
        RECT -47.765 41.995 -47.435 42.325 ;
        RECT -47.765 40.635 -47.435 40.965 ;
        RECT -47.765 39.275 -47.435 39.605 ;
        RECT -47.765 37.915 -47.435 38.245 ;
        RECT -47.765 36.555 -47.435 36.885 ;
        RECT -47.765 35.195 -47.435 35.525 ;
        RECT -47.765 33.835 -47.435 34.165 ;
        RECT -47.765 32.475 -47.435 32.805 ;
        RECT -47.765 31.115 -47.435 31.445 ;
        RECT -47.765 29.755 -47.435 30.085 ;
        RECT -47.765 28.395 -47.435 28.725 ;
        RECT -47.765 27.035 -47.435 27.365 ;
        RECT -47.765 25.675 -47.435 26.005 ;
        RECT -47.765 24.315 -47.435 24.645 ;
        RECT -47.765 22.955 -47.435 23.285 ;
        RECT -47.765 21.595 -47.435 21.925 ;
        RECT -47.765 20.235 -47.435 20.565 ;
        RECT -47.765 18.875 -47.435 19.205 ;
        RECT -47.765 17.515 -47.435 17.845 ;
        RECT -47.765 16.155 -47.435 16.485 ;
        RECT -47.765 14.795 -47.435 15.125 ;
        RECT -47.765 13.435 -47.435 13.765 ;
        RECT -47.765 12.075 -47.435 12.405 ;
        RECT -47.765 10.715 -47.435 11.045 ;
        RECT -47.765 9.355 -47.435 9.685 ;
        RECT -47.765 7.995 -47.435 8.325 ;
        RECT -47.765 6.635 -47.435 6.965 ;
        RECT -47.765 5.275 -47.435 5.605 ;
        RECT -47.765 3.915 -47.435 4.245 ;
        RECT -47.765 2.555 -47.435 2.885 ;
        RECT -47.765 1.195 -47.435 1.525 ;
        RECT -47.765 -0.165 -47.435 0.165 ;
        RECT -47.765 -1.525 -47.435 -1.195 ;
        RECT -47.765 -2.885 -47.435 -2.555 ;
        RECT -47.765 -4.245 -47.435 -3.915 ;
        RECT -47.765 -5.605 -47.435 -5.275 ;
        RECT -47.765 -6.965 -47.435 -6.635 ;
        RECT -47.765 -8.325 -47.435 -7.995 ;
        RECT -47.765 -9.685 -47.435 -9.355 ;
        RECT -47.765 -12.405 -47.435 -12.075 ;
        RECT -47.765 -13.765 -47.435 -13.435 ;
        RECT -47.765 -15.125 -47.435 -14.795 ;
        RECT -47.765 -16.485 -47.435 -16.155 ;
        RECT -47.765 -17.845 -47.435 -17.515 ;
        RECT -47.765 -19.205 -47.435 -18.875 ;
        RECT -47.765 -20.565 -47.435 -20.235 ;
        RECT -47.765 -21.925 -47.435 -21.595 ;
        RECT -47.765 -26.005 -47.435 -25.675 ;
        RECT -47.765 -27.365 -47.435 -27.035 ;
        RECT -47.765 -28.725 -47.435 -28.395 ;
        RECT -47.765 -30.085 -47.435 -29.755 ;
        RECT -47.765 -31.445 -47.435 -31.115 ;
        RECT -47.765 -32.805 -47.435 -32.475 ;
        RECT -47.765 -34.165 -47.435 -33.835 ;
        RECT -47.765 -35.525 -47.435 -35.195 ;
        RECT -47.765 -36.885 -47.435 -36.555 ;
        RECT -47.765 -38.245 -47.435 -37.915 ;
        RECT -47.765 -39.605 -47.435 -39.275 ;
        RECT -47.765 -40.965 -47.435 -40.635 ;
        RECT -47.765 -42.325 -47.435 -41.995 ;
        RECT -47.765 -43.685 -47.435 -43.355 ;
        RECT -47.765 -45.045 -47.435 -44.715 ;
        RECT -47.765 -46.405 -47.435 -46.075 ;
        RECT -47.765 -47.765 -47.435 -47.435 ;
        RECT -47.765 -49.125 -47.435 -48.795 ;
        RECT -47.765 -50.485 -47.435 -50.155 ;
        RECT -47.765 -51.845 -47.435 -51.515 ;
        RECT -47.765 -53.205 -47.435 -52.875 ;
        RECT -47.765 -54.565 -47.435 -54.235 ;
        RECT -47.765 -55.925 -47.435 -55.595 ;
        RECT -47.765 -57.285 -47.435 -56.955 ;
        RECT -47.765 -58.645 -47.435 -58.315 ;
        RECT -47.765 -60.005 -47.435 -59.675 ;
        RECT -47.765 -61.365 -47.435 -61.035 ;
        RECT -47.765 -62.725 -47.435 -62.395 ;
        RECT -47.765 -64.085 -47.435 -63.755 ;
        RECT -47.765 -65.445 -47.435 -65.115 ;
        RECT -47.765 -66.805 -47.435 -66.475 ;
        RECT -47.765 -68.165 -47.435 -67.835 ;
        RECT -47.765 -69.525 -47.435 -69.195 ;
        RECT -47.765 -72.245 -47.435 -71.915 ;
        RECT -47.765 -73.605 -47.435 -73.275 ;
        RECT -47.765 -74.965 -47.435 -74.635 ;
        RECT -47.765 -76.325 -47.435 -75.995 ;
        RECT -47.765 -78.29 -47.435 -77.96 ;
        RECT -47.765 -79.045 -47.435 -78.715 ;
        RECT -47.765 -81.765 -47.435 -81.435 ;
        RECT -47.765 -83.125 -47.435 -82.795 ;
        RECT -47.765 -84.485 -47.435 -84.155 ;
        RECT -47.765 -86.43 -47.435 -86.1 ;
        RECT -47.765 -87.205 -47.435 -86.875 ;
        RECT -47.765 -88.565 -47.435 -88.235 ;
        RECT -47.765 -89.925 -47.435 -89.595 ;
        RECT -47.76 -91.28 -47.44 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 -153.845 -47.435 -153.515 ;
        RECT -47.765 -155.285 -47.435 -154.955 ;
        RECT -47.765 -156.565 -47.435 -156.235 ;
        RECT -47.765 -157.925 -47.435 -157.595 ;
        RECT -47.765 -160.17 -47.435 -159.04 ;
        RECT -47.76 -160.285 -47.44 -152.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 127.225 -46.075 128.355 ;
        RECT -46.405 124.955 -46.075 125.285 ;
        RECT -46.405 123.595 -46.075 123.925 ;
        RECT -46.405 122.235 -46.075 122.565 ;
        RECT -46.405 120.875 -46.075 121.205 ;
        RECT -46.405 119.515 -46.075 119.845 ;
        RECT -46.405 118.155 -46.075 118.485 ;
        RECT -46.405 116.795 -46.075 117.125 ;
        RECT -46.405 115.435 -46.075 115.765 ;
        RECT -46.405 114.075 -46.075 114.405 ;
        RECT -46.405 112.715 -46.075 113.045 ;
        RECT -46.405 111.355 -46.075 111.685 ;
        RECT -46.405 109.995 -46.075 110.325 ;
        RECT -46.405 108.635 -46.075 108.965 ;
        RECT -46.405 107.275 -46.075 107.605 ;
        RECT -46.405 105.915 -46.075 106.245 ;
        RECT -46.405 104.555 -46.075 104.885 ;
        RECT -46.405 103.195 -46.075 103.525 ;
        RECT -46.405 101.835 -46.075 102.165 ;
        RECT -46.405 100.475 -46.075 100.805 ;
        RECT -46.405 99.115 -46.075 99.445 ;
        RECT -46.405 97.755 -46.075 98.085 ;
        RECT -46.405 96.395 -46.075 96.725 ;
        RECT -46.405 95.035 -46.075 95.365 ;
        RECT -46.405 93.675 -46.075 94.005 ;
        RECT -46.405 92.315 -46.075 92.645 ;
        RECT -46.405 90.955 -46.075 91.285 ;
        RECT -46.405 89.595 -46.075 89.925 ;
        RECT -46.405 88.235 -46.075 88.565 ;
        RECT -46.405 86.875 -46.075 87.205 ;
        RECT -46.405 85.515 -46.075 85.845 ;
        RECT -46.405 84.155 -46.075 84.485 ;
        RECT -46.405 82.795 -46.075 83.125 ;
        RECT -46.405 81.435 -46.075 81.765 ;
        RECT -46.405 80.075 -46.075 80.405 ;
        RECT -46.405 78.715 -46.075 79.045 ;
        RECT -46.405 77.355 -46.075 77.685 ;
        RECT -46.405 75.995 -46.075 76.325 ;
        RECT -46.405 74.635 -46.075 74.965 ;
        RECT -46.405 73.275 -46.075 73.605 ;
        RECT -46.405 72.445 -46.075 72.775 ;
        RECT -46.405 70.395 -46.075 70.725 ;
        RECT -46.405 68.035 -46.075 68.365 ;
        RECT -46.405 66.885 -46.075 67.215 ;
        RECT -46.405 64.875 -46.075 65.205 ;
        RECT -46.405 63.725 -46.075 64.055 ;
        RECT -46.405 61.715 -46.075 62.045 ;
        RECT -46.405 60.395 -46.075 60.725 ;
        RECT -46.405 58.555 -46.075 58.885 ;
        RECT -46.405 57.405 -46.075 57.735 ;
        RECT -46.405 55.395 -46.075 55.725 ;
        RECT -46.405 54.245 -46.075 54.575 ;
        RECT -46.405 51.885 -46.075 52.215 ;
        RECT -46.405 49.83 -46.075 50.16 ;
        RECT -46.405 48.795 -46.075 49.125 ;
        RECT -46.405 47.435 -46.075 47.765 ;
        RECT -46.405 46.075 -46.075 46.405 ;
        RECT -46.405 44.715 -46.075 45.045 ;
        RECT -46.405 43.355 -46.075 43.685 ;
        RECT -46.405 41.995 -46.075 42.325 ;
        RECT -46.405 40.635 -46.075 40.965 ;
        RECT -46.405 39.275 -46.075 39.605 ;
        RECT -46.405 37.915 -46.075 38.245 ;
        RECT -46.405 36.555 -46.075 36.885 ;
        RECT -46.405 35.195 -46.075 35.525 ;
        RECT -46.405 33.835 -46.075 34.165 ;
        RECT -46.405 32.475 -46.075 32.805 ;
        RECT -46.405 31.115 -46.075 31.445 ;
        RECT -46.405 29.755 -46.075 30.085 ;
        RECT -46.405 28.395 -46.075 28.725 ;
        RECT -46.405 27.035 -46.075 27.365 ;
        RECT -46.405 25.675 -46.075 26.005 ;
        RECT -46.405 24.315 -46.075 24.645 ;
        RECT -46.405 22.955 -46.075 23.285 ;
        RECT -46.405 21.595 -46.075 21.925 ;
        RECT -46.405 20.235 -46.075 20.565 ;
        RECT -46.405 18.875 -46.075 19.205 ;
        RECT -46.405 17.515 -46.075 17.845 ;
        RECT -46.405 16.155 -46.075 16.485 ;
        RECT -46.405 14.795 -46.075 15.125 ;
        RECT -46.405 13.435 -46.075 13.765 ;
        RECT -46.405 12.075 -46.075 12.405 ;
        RECT -46.405 10.715 -46.075 11.045 ;
        RECT -46.405 9.355 -46.075 9.685 ;
        RECT -46.405 7.995 -46.075 8.325 ;
        RECT -46.405 6.635 -46.075 6.965 ;
        RECT -46.405 5.275 -46.075 5.605 ;
        RECT -46.405 3.915 -46.075 4.245 ;
        RECT -46.405 2.555 -46.075 2.885 ;
        RECT -46.405 1.195 -46.075 1.525 ;
        RECT -46.405 -0.165 -46.075 0.165 ;
        RECT -46.405 -1.525 -46.075 -1.195 ;
        RECT -46.405 -2.885 -46.075 -2.555 ;
        RECT -46.405 -4.245 -46.075 -3.915 ;
        RECT -46.405 -5.605 -46.075 -5.275 ;
        RECT -46.405 -6.965 -46.075 -6.635 ;
        RECT -46.405 -8.325 -46.075 -7.995 ;
        RECT -46.405 -9.685 -46.075 -9.355 ;
        RECT -46.405 -12.405 -46.075 -12.075 ;
        RECT -46.405 -13.765 -46.075 -13.435 ;
        RECT -46.405 -15.125 -46.075 -14.795 ;
        RECT -46.405 -16.485 -46.075 -16.155 ;
        RECT -46.405 -17.845 -46.075 -17.515 ;
        RECT -46.405 -19.205 -46.075 -18.875 ;
        RECT -46.405 -20.565 -46.075 -20.235 ;
        RECT -46.405 -21.925 -46.075 -21.595 ;
        RECT -46.405 -26.005 -46.075 -25.675 ;
        RECT -46.405 -27.365 -46.075 -27.035 ;
        RECT -46.405 -28.725 -46.075 -28.395 ;
        RECT -46.405 -30.085 -46.075 -29.755 ;
        RECT -46.405 -31.445 -46.075 -31.115 ;
        RECT -46.405 -32.805 -46.075 -32.475 ;
        RECT -46.405 -34.165 -46.075 -33.835 ;
        RECT -46.405 -35.525 -46.075 -35.195 ;
        RECT -46.405 -36.885 -46.075 -36.555 ;
        RECT -46.405 -38.245 -46.075 -37.915 ;
        RECT -46.405 -39.605 -46.075 -39.275 ;
        RECT -46.405 -40.965 -46.075 -40.635 ;
        RECT -46.405 -42.325 -46.075 -41.995 ;
        RECT -46.405 -43.685 -46.075 -43.355 ;
        RECT -46.405 -45.045 -46.075 -44.715 ;
        RECT -46.405 -46.405 -46.075 -46.075 ;
        RECT -46.405 -47.765 -46.075 -47.435 ;
        RECT -46.405 -49.125 -46.075 -48.795 ;
        RECT -46.405 -50.485 -46.075 -50.155 ;
        RECT -46.405 -51.845 -46.075 -51.515 ;
        RECT -46.405 -53.205 -46.075 -52.875 ;
        RECT -46.405 -54.565 -46.075 -54.235 ;
        RECT -46.405 -55.925 -46.075 -55.595 ;
        RECT -46.405 -57.285 -46.075 -56.955 ;
        RECT -46.405 -58.645 -46.075 -58.315 ;
        RECT -46.405 -60.005 -46.075 -59.675 ;
        RECT -46.405 -61.365 -46.075 -61.035 ;
        RECT -46.405 -62.725 -46.075 -62.395 ;
        RECT -46.405 -64.085 -46.075 -63.755 ;
        RECT -46.405 -65.445 -46.075 -65.115 ;
        RECT -46.405 -66.805 -46.075 -66.475 ;
        RECT -46.405 -68.165 -46.075 -67.835 ;
        RECT -46.405 -69.525 -46.075 -69.195 ;
        RECT -46.405 -72.245 -46.075 -71.915 ;
        RECT -46.405 -73.605 -46.075 -73.275 ;
        RECT -46.405 -74.965 -46.075 -74.635 ;
        RECT -46.405 -76.325 -46.075 -75.995 ;
        RECT -46.405 -78.29 -46.075 -77.96 ;
        RECT -46.405 -79.045 -46.075 -78.715 ;
        RECT -46.405 -81.765 -46.075 -81.435 ;
        RECT -46.405 -83.125 -46.075 -82.795 ;
        RECT -46.405 -84.485 -46.075 -84.155 ;
        RECT -46.405 -86.43 -46.075 -86.1 ;
        RECT -46.405 -87.205 -46.075 -86.875 ;
        RECT -46.405 -88.565 -46.075 -88.235 ;
        RECT -46.405 -89.925 -46.075 -89.595 ;
        RECT -46.405 -92.645 -46.075 -92.315 ;
        RECT -46.405 -94.005 -46.075 -93.675 ;
        RECT -46.405 -95.365 -46.075 -95.035 ;
        RECT -46.405 -96.725 -46.075 -96.395 ;
        RECT -46.405 -98.085 -46.075 -97.755 ;
        RECT -46.405 -102.165 -46.075 -101.835 ;
        RECT -46.405 -103.525 -46.075 -103.195 ;
        RECT -46.405 -104.885 -46.075 -104.555 ;
        RECT -46.405 -106.245 -46.075 -105.915 ;
        RECT -46.405 -107.605 -46.075 -107.275 ;
        RECT -46.405 -108.965 -46.075 -108.635 ;
        RECT -46.405 -110.325 -46.075 -109.995 ;
        RECT -46.405 -111.685 -46.075 -111.355 ;
        RECT -46.405 -113.045 -46.075 -112.715 ;
        RECT -46.405 -114.405 -46.075 -114.075 ;
        RECT -46.405 -115.765 -46.075 -115.435 ;
        RECT -46.405 -117.125 -46.075 -116.795 ;
        RECT -46.405 -118.485 -46.075 -118.155 ;
        RECT -46.405 -119.845 -46.075 -119.515 ;
        RECT -46.405 -121.205 -46.075 -120.875 ;
        RECT -46.405 -122.565 -46.075 -122.235 ;
        RECT -46.405 -123.925 -46.075 -123.595 ;
        RECT -46.405 -125.285 -46.075 -124.955 ;
        RECT -46.405 -126.645 -46.075 -126.315 ;
        RECT -46.405 -128.005 -46.075 -127.675 ;
        RECT -46.405 -129.365 -46.075 -129.035 ;
        RECT -46.405 -130.725 -46.075 -130.395 ;
        RECT -46.405 -132.085 -46.075 -131.755 ;
        RECT -46.405 -133.445 -46.075 -133.115 ;
        RECT -46.405 -134.805 -46.075 -134.475 ;
        RECT -46.405 -136.165 -46.075 -135.835 ;
        RECT -46.405 -137.525 -46.075 -137.195 ;
        RECT -46.405 -138.885 -46.075 -138.555 ;
        RECT -46.405 -140.245 -46.075 -139.915 ;
        RECT -46.405 -141.605 -46.075 -141.275 ;
        RECT -46.405 -142.965 -46.075 -142.635 ;
        RECT -46.405 -144.325 -46.075 -143.995 ;
        RECT -46.405 -145.685 -46.075 -145.355 ;
        RECT -46.405 -147.045 -46.075 -146.715 ;
        RECT -46.405 -149.765 -46.075 -149.435 ;
        RECT -46.4 -151.8 -46.08 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 -8.325 -44.715 -7.995 ;
        RECT -45.045 -12.405 -44.715 -12.075 ;
        RECT -45.045 -13.765 -44.715 -13.435 ;
        RECT -45.045 -15.125 -44.715 -14.795 ;
        RECT -45.045 -16.485 -44.715 -16.155 ;
        RECT -45.045 -17.845 -44.715 -17.515 ;
        RECT -45.045 -19.205 -44.715 -18.875 ;
        RECT -45.045 -20.565 -44.715 -20.235 ;
        RECT -45.045 -21.925 -44.715 -21.595 ;
        RECT -45.045 -26.005 -44.715 -25.675 ;
        RECT -45.045 -27.365 -44.715 -27.035 ;
        RECT -45.045 -28.725 -44.715 -28.395 ;
        RECT -45.045 -30.085 -44.715 -29.755 ;
        RECT -45.045 -31.445 -44.715 -31.115 ;
        RECT -45.045 -32.805 -44.715 -32.475 ;
        RECT -45.045 -34.165 -44.715 -33.835 ;
        RECT -45.045 -35.525 -44.715 -35.195 ;
        RECT -45.045 -36.885 -44.715 -36.555 ;
        RECT -45.045 -38.245 -44.715 -37.915 ;
        RECT -45.045 -39.605 -44.715 -39.275 ;
        RECT -45.045 -40.965 -44.715 -40.635 ;
        RECT -45.045 -42.325 -44.715 -41.995 ;
        RECT -45.045 -43.685 -44.715 -43.355 ;
        RECT -45.045 -45.045 -44.715 -44.715 ;
        RECT -45.045 -46.405 -44.715 -46.075 ;
        RECT -45.045 -47.765 -44.715 -47.435 ;
        RECT -45.045 -49.125 -44.715 -48.795 ;
        RECT -45.045 -50.485 -44.715 -50.155 ;
        RECT -45.045 -51.845 -44.715 -51.515 ;
        RECT -45.045 -53.205 -44.715 -52.875 ;
        RECT -45.045 -54.565 -44.715 -54.235 ;
        RECT -45.045 -55.925 -44.715 -55.595 ;
        RECT -45.045 -57.285 -44.715 -56.955 ;
        RECT -45.045 -58.645 -44.715 -58.315 ;
        RECT -45.045 -60.005 -44.715 -59.675 ;
        RECT -45.045 -61.365 -44.715 -61.035 ;
        RECT -45.045 -62.725 -44.715 -62.395 ;
        RECT -45.045 -64.085 -44.715 -63.755 ;
        RECT -45.045 -65.445 -44.715 -65.115 ;
        RECT -45.045 -66.805 -44.715 -66.475 ;
        RECT -45.045 -68.165 -44.715 -67.835 ;
        RECT -45.045 -69.525 -44.715 -69.195 ;
        RECT -45.045 -72.245 -44.715 -71.915 ;
        RECT -45.045 -73.605 -44.715 -73.275 ;
        RECT -45.045 -74.965 -44.715 -74.635 ;
        RECT -45.045 -76.325 -44.715 -75.995 ;
        RECT -45.045 -78.29 -44.715 -77.96 ;
        RECT -45.045 -79.045 -44.715 -78.715 ;
        RECT -45.045 -81.765 -44.715 -81.435 ;
        RECT -45.045 -83.125 -44.715 -82.795 ;
        RECT -45.045 -84.485 -44.715 -84.155 ;
        RECT -45.045 -86.43 -44.715 -86.1 ;
        RECT -45.045 -87.205 -44.715 -86.875 ;
        RECT -45.045 -88.565 -44.715 -88.235 ;
        RECT -45.045 -89.925 -44.715 -89.595 ;
        RECT -45.045 -92.645 -44.715 -92.315 ;
        RECT -45.045 -94.005 -44.715 -93.675 ;
        RECT -45.045 -95.365 -44.715 -95.035 ;
        RECT -45.045 -96.725 -44.715 -96.395 ;
        RECT -45.045 -98.085 -44.715 -97.755 ;
        RECT -45.045 -102.165 -44.715 -101.835 ;
        RECT -45.045 -103.525 -44.715 -103.195 ;
        RECT -45.045 -104.885 -44.715 -104.555 ;
        RECT -45.045 -106.245 -44.715 -105.915 ;
        RECT -45.045 -107.605 -44.715 -107.275 ;
        RECT -45.045 -108.965 -44.715 -108.635 ;
        RECT -45.045 -110.325 -44.715 -109.995 ;
        RECT -45.045 -111.685 -44.715 -111.355 ;
        RECT -45.045 -113.045 -44.715 -112.715 ;
        RECT -45.045 -114.405 -44.715 -114.075 ;
        RECT -45.045 -115.765 -44.715 -115.435 ;
        RECT -45.045 -117.125 -44.715 -116.795 ;
        RECT -45.045 -118.485 -44.715 -118.155 ;
        RECT -45.045 -119.845 -44.715 -119.515 ;
        RECT -45.045 -121.205 -44.715 -120.875 ;
        RECT -45.045 -122.565 -44.715 -122.235 ;
        RECT -45.045 -123.925 -44.715 -123.595 ;
        RECT -45.045 -125.285 -44.715 -124.955 ;
        RECT -45.045 -126.645 -44.715 -126.315 ;
        RECT -45.045 -128.005 -44.715 -127.675 ;
        RECT -45.045 -129.365 -44.715 -129.035 ;
        RECT -45.045 -130.725 -44.715 -130.395 ;
        RECT -45.045 -132.085 -44.715 -131.755 ;
        RECT -45.045 -133.445 -44.715 -133.115 ;
        RECT -45.045 -134.805 -44.715 -134.475 ;
        RECT -45.045 -136.165 -44.715 -135.835 ;
        RECT -45.045 -137.525 -44.715 -137.195 ;
        RECT -45.045 -138.885 -44.715 -138.555 ;
        RECT -45.045 -140.245 -44.715 -139.915 ;
        RECT -45.045 -141.605 -44.715 -141.275 ;
        RECT -45.045 -142.965 -44.715 -142.635 ;
        RECT -45.045 -144.325 -44.715 -143.995 ;
        RECT -45.045 -145.685 -44.715 -145.355 ;
        RECT -45.045 -147.045 -44.715 -146.715 ;
        RECT -45.045 -149.765 -44.715 -149.435 ;
        RECT -45.045 -152.485 -44.715 -152.155 ;
        RECT -45.045 -153.845 -44.715 -153.515 ;
        RECT -45.045 -155.285 -44.715 -154.955 ;
        RECT -45.045 -156.565 -44.715 -156.235 ;
        RECT -45.045 -157.925 -44.715 -157.595 ;
        RECT -45.045 -160.17 -44.715 -159.04 ;
        RECT -45.04 -160.285 -44.72 128.47 ;
        RECT -45.045 127.225 -44.715 128.355 ;
        RECT -45.045 124.955 -44.715 125.285 ;
        RECT -45.045 123.595 -44.715 123.925 ;
        RECT -45.045 122.235 -44.715 122.565 ;
        RECT -45.045 120.875 -44.715 121.205 ;
        RECT -45.045 119.515 -44.715 119.845 ;
        RECT -45.045 118.155 -44.715 118.485 ;
        RECT -45.045 116.795 -44.715 117.125 ;
        RECT -45.045 115.435 -44.715 115.765 ;
        RECT -45.045 114.075 -44.715 114.405 ;
        RECT -45.045 112.715 -44.715 113.045 ;
        RECT -45.045 111.355 -44.715 111.685 ;
        RECT -45.045 109.995 -44.715 110.325 ;
        RECT -45.045 108.635 -44.715 108.965 ;
        RECT -45.045 107.275 -44.715 107.605 ;
        RECT -45.045 105.915 -44.715 106.245 ;
        RECT -45.045 104.555 -44.715 104.885 ;
        RECT -45.045 103.195 -44.715 103.525 ;
        RECT -45.045 101.835 -44.715 102.165 ;
        RECT -45.045 100.475 -44.715 100.805 ;
        RECT -45.045 99.115 -44.715 99.445 ;
        RECT -45.045 97.755 -44.715 98.085 ;
        RECT -45.045 96.395 -44.715 96.725 ;
        RECT -45.045 95.035 -44.715 95.365 ;
        RECT -45.045 93.675 -44.715 94.005 ;
        RECT -45.045 92.315 -44.715 92.645 ;
        RECT -45.045 90.955 -44.715 91.285 ;
        RECT -45.045 89.595 -44.715 89.925 ;
        RECT -45.045 88.235 -44.715 88.565 ;
        RECT -45.045 86.875 -44.715 87.205 ;
        RECT -45.045 85.515 -44.715 85.845 ;
        RECT -45.045 84.155 -44.715 84.485 ;
        RECT -45.045 82.795 -44.715 83.125 ;
        RECT -45.045 81.435 -44.715 81.765 ;
        RECT -45.045 80.075 -44.715 80.405 ;
        RECT -45.045 78.715 -44.715 79.045 ;
        RECT -45.045 77.355 -44.715 77.685 ;
        RECT -45.045 75.995 -44.715 76.325 ;
        RECT -45.045 74.635 -44.715 74.965 ;
        RECT -45.045 73.275 -44.715 73.605 ;
        RECT -45.045 72.445 -44.715 72.775 ;
        RECT -45.045 70.395 -44.715 70.725 ;
        RECT -45.045 68.035 -44.715 68.365 ;
        RECT -45.045 66.885 -44.715 67.215 ;
        RECT -45.045 64.875 -44.715 65.205 ;
        RECT -45.045 63.725 -44.715 64.055 ;
        RECT -45.045 61.715 -44.715 62.045 ;
        RECT -45.045 60.395 -44.715 60.725 ;
        RECT -45.045 58.555 -44.715 58.885 ;
        RECT -45.045 57.405 -44.715 57.735 ;
        RECT -45.045 55.395 -44.715 55.725 ;
        RECT -45.045 54.245 -44.715 54.575 ;
        RECT -45.045 51.885 -44.715 52.215 ;
        RECT -45.045 49.83 -44.715 50.16 ;
        RECT -45.045 48.795 -44.715 49.125 ;
        RECT -45.045 47.435 -44.715 47.765 ;
        RECT -45.045 46.075 -44.715 46.405 ;
        RECT -45.045 44.715 -44.715 45.045 ;
        RECT -45.045 43.355 -44.715 43.685 ;
        RECT -45.045 41.995 -44.715 42.325 ;
        RECT -45.045 40.635 -44.715 40.965 ;
        RECT -45.045 39.275 -44.715 39.605 ;
        RECT -45.045 37.915 -44.715 38.245 ;
        RECT -45.045 36.555 -44.715 36.885 ;
        RECT -45.045 35.195 -44.715 35.525 ;
        RECT -45.045 33.835 -44.715 34.165 ;
        RECT -45.045 32.475 -44.715 32.805 ;
        RECT -45.045 31.115 -44.715 31.445 ;
        RECT -45.045 29.755 -44.715 30.085 ;
        RECT -45.045 28.395 -44.715 28.725 ;
        RECT -45.045 27.035 -44.715 27.365 ;
        RECT -45.045 25.675 -44.715 26.005 ;
        RECT -45.045 24.315 -44.715 24.645 ;
        RECT -45.045 22.955 -44.715 23.285 ;
        RECT -45.045 21.595 -44.715 21.925 ;
        RECT -45.045 20.235 -44.715 20.565 ;
        RECT -45.045 18.875 -44.715 19.205 ;
        RECT -45.045 17.515 -44.715 17.845 ;
        RECT -45.045 16.155 -44.715 16.485 ;
        RECT -45.045 14.795 -44.715 15.125 ;
        RECT -45.045 13.435 -44.715 13.765 ;
        RECT -45.045 12.075 -44.715 12.405 ;
        RECT -45.045 10.715 -44.715 11.045 ;
        RECT -45.045 9.355 -44.715 9.685 ;
        RECT -45.045 7.995 -44.715 8.325 ;
        RECT -45.045 6.635 -44.715 6.965 ;
        RECT -45.045 5.275 -44.715 5.605 ;
        RECT -45.045 3.915 -44.715 4.245 ;
        RECT -45.045 2.555 -44.715 2.885 ;
        RECT -45.045 1.195 -44.715 1.525 ;
        RECT -45.045 -0.165 -44.715 0.165 ;
        RECT -45.045 -1.525 -44.715 -1.195 ;
        RECT -45.045 -2.885 -44.715 -2.555 ;
        RECT -45.045 -4.245 -44.715 -3.915 ;
        RECT -45.045 -5.605 -44.715 -5.275 ;
        RECT -45.045 -6.965 -44.715 -6.635 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 -153.845 -59.675 -153.515 ;
        RECT -60.005 -155.285 -59.675 -154.955 ;
        RECT -60.005 -156.565 -59.675 -156.235 ;
        RECT -60.005 -157.925 -59.675 -157.595 ;
        RECT -60.005 -160.17 -59.675 -159.04 ;
        RECT -60 -160.285 -59.68 -152.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.645 127.225 -58.315 128.355 ;
        RECT -58.645 124.955 -58.315 125.285 ;
        RECT -58.645 123.595 -58.315 123.925 ;
        RECT -58.645 122.235 -58.315 122.565 ;
        RECT -58.645 120.875 -58.315 121.205 ;
        RECT -58.645 119.515 -58.315 119.845 ;
        RECT -58.645 118.155 -58.315 118.485 ;
        RECT -58.645 116.795 -58.315 117.125 ;
        RECT -58.645 115.435 -58.315 115.765 ;
        RECT -58.645 114.075 -58.315 114.405 ;
        RECT -58.645 112.715 -58.315 113.045 ;
        RECT -58.645 111.355 -58.315 111.685 ;
        RECT -58.645 109.995 -58.315 110.325 ;
        RECT -58.645 108.635 -58.315 108.965 ;
        RECT -58.645 107.275 -58.315 107.605 ;
        RECT -58.645 105.915 -58.315 106.245 ;
        RECT -58.645 104.555 -58.315 104.885 ;
        RECT -58.645 103.195 -58.315 103.525 ;
        RECT -58.645 101.835 -58.315 102.165 ;
        RECT -58.645 100.475 -58.315 100.805 ;
        RECT -58.645 99.115 -58.315 99.445 ;
        RECT -58.645 97.755 -58.315 98.085 ;
        RECT -58.645 96.395 -58.315 96.725 ;
        RECT -58.645 95.035 -58.315 95.365 ;
        RECT -58.645 93.675 -58.315 94.005 ;
        RECT -58.645 92.315 -58.315 92.645 ;
        RECT -58.645 90.955 -58.315 91.285 ;
        RECT -58.645 89.595 -58.315 89.925 ;
        RECT -58.645 88.235 -58.315 88.565 ;
        RECT -58.645 86.875 -58.315 87.205 ;
        RECT -58.645 85.515 -58.315 85.845 ;
        RECT -58.645 84.155 -58.315 84.485 ;
        RECT -58.645 82.795 -58.315 83.125 ;
        RECT -58.645 81.435 -58.315 81.765 ;
        RECT -58.645 80.075 -58.315 80.405 ;
        RECT -58.645 78.715 -58.315 79.045 ;
        RECT -58.645 77.355 -58.315 77.685 ;
        RECT -58.645 75.995 -58.315 76.325 ;
        RECT -58.645 74.635 -58.315 74.965 ;
        RECT -58.645 73.275 -58.315 73.605 ;
        RECT -58.645 72.445 -58.315 72.775 ;
        RECT -58.645 70.395 -58.315 70.725 ;
        RECT -58.645 68.035 -58.315 68.365 ;
        RECT -58.645 66.885 -58.315 67.215 ;
        RECT -58.645 64.875 -58.315 65.205 ;
        RECT -58.645 63.725 -58.315 64.055 ;
        RECT -58.645 61.715 -58.315 62.045 ;
        RECT -58.645 60.395 -58.315 60.725 ;
        RECT -58.645 58.555 -58.315 58.885 ;
        RECT -58.645 57.405 -58.315 57.735 ;
        RECT -58.645 55.395 -58.315 55.725 ;
        RECT -58.645 54.245 -58.315 54.575 ;
        RECT -58.645 51.885 -58.315 52.215 ;
        RECT -58.645 49.83 -58.315 50.16 ;
        RECT -58.645 48.795 -58.315 49.125 ;
        RECT -58.645 47.435 -58.315 47.765 ;
        RECT -58.645 46.075 -58.315 46.405 ;
        RECT -58.645 44.715 -58.315 45.045 ;
        RECT -58.645 43.355 -58.315 43.685 ;
        RECT -58.645 41.995 -58.315 42.325 ;
        RECT -58.645 40.635 -58.315 40.965 ;
        RECT -58.645 39.275 -58.315 39.605 ;
        RECT -58.645 37.915 -58.315 38.245 ;
        RECT -58.645 36.555 -58.315 36.885 ;
        RECT -58.645 35.195 -58.315 35.525 ;
        RECT -58.645 33.835 -58.315 34.165 ;
        RECT -58.645 32.475 -58.315 32.805 ;
        RECT -58.645 31.115 -58.315 31.445 ;
        RECT -58.645 29.755 -58.315 30.085 ;
        RECT -58.645 28.395 -58.315 28.725 ;
        RECT -58.645 27.035 -58.315 27.365 ;
        RECT -58.645 25.675 -58.315 26.005 ;
        RECT -58.645 24.315 -58.315 24.645 ;
        RECT -58.645 22.955 -58.315 23.285 ;
        RECT -58.645 21.595 -58.315 21.925 ;
        RECT -58.645 20.235 -58.315 20.565 ;
        RECT -58.645 18.875 -58.315 19.205 ;
        RECT -58.645 17.515 -58.315 17.845 ;
        RECT -58.645 16.155 -58.315 16.485 ;
        RECT -58.645 14.795 -58.315 15.125 ;
        RECT -58.645 13.435 -58.315 13.765 ;
        RECT -58.645 12.075 -58.315 12.405 ;
        RECT -58.645 10.715 -58.315 11.045 ;
        RECT -58.645 9.355 -58.315 9.685 ;
        RECT -58.645 7.995 -58.315 8.325 ;
        RECT -58.645 6.635 -58.315 6.965 ;
        RECT -58.645 5.275 -58.315 5.605 ;
        RECT -58.645 3.915 -58.315 4.245 ;
        RECT -58.645 2.555 -58.315 2.885 ;
        RECT -58.645 1.195 -58.315 1.525 ;
        RECT -58.645 -0.165 -58.315 0.165 ;
        RECT -58.645 -1.525 -58.315 -1.195 ;
        RECT -58.645 -2.885 -58.315 -2.555 ;
        RECT -58.645 -4.245 -58.315 -3.915 ;
        RECT -58.645 -5.605 -58.315 -5.275 ;
        RECT -58.645 -6.965 -58.315 -6.635 ;
        RECT -58.645 -8.325 -58.315 -7.995 ;
        RECT -58.645 -9.685 -58.315 -9.355 ;
        RECT -58.645 -11.045 -58.315 -10.715 ;
        RECT -58.645 -12.405 -58.315 -12.075 ;
        RECT -58.645 -13.765 -58.315 -13.435 ;
        RECT -58.645 -15.125 -58.315 -14.795 ;
        RECT -58.645 -16.485 -58.315 -16.155 ;
        RECT -58.645 -17.845 -58.315 -17.515 ;
        RECT -58.645 -19.205 -58.315 -18.875 ;
        RECT -58.645 -20.565 -58.315 -20.235 ;
        RECT -58.645 -21.925 -58.315 -21.595 ;
        RECT -58.645 -23.285 -58.315 -22.955 ;
        RECT -58.645 -24.645 -58.315 -24.315 ;
        RECT -58.645 -26.005 -58.315 -25.675 ;
        RECT -58.645 -27.365 -58.315 -27.035 ;
        RECT -58.645 -28.725 -58.315 -28.395 ;
        RECT -58.645 -30.085 -58.315 -29.755 ;
        RECT -58.645 -31.445 -58.315 -31.115 ;
        RECT -58.645 -32.805 -58.315 -32.475 ;
        RECT -58.645 -34.165 -58.315 -33.835 ;
        RECT -58.645 -35.525 -58.315 -35.195 ;
        RECT -58.645 -36.885 -58.315 -36.555 ;
        RECT -58.645 -38.245 -58.315 -37.915 ;
        RECT -58.645 -39.605 -58.315 -39.275 ;
        RECT -58.645 -40.965 -58.315 -40.635 ;
        RECT -58.645 -42.325 -58.315 -41.995 ;
        RECT -58.645 -43.685 -58.315 -43.355 ;
        RECT -58.645 -45.045 -58.315 -44.715 ;
        RECT -58.645 -46.405 -58.315 -46.075 ;
        RECT -58.645 -47.765 -58.315 -47.435 ;
        RECT -58.645 -49.125 -58.315 -48.795 ;
        RECT -58.645 -50.485 -58.315 -50.155 ;
        RECT -58.645 -51.845 -58.315 -51.515 ;
        RECT -58.645 -53.205 -58.315 -52.875 ;
        RECT -58.645 -54.565 -58.315 -54.235 ;
        RECT -58.645 -55.925 -58.315 -55.595 ;
        RECT -58.645 -57.285 -58.315 -56.955 ;
        RECT -58.645 -58.645 -58.315 -58.315 ;
        RECT -58.645 -60.005 -58.315 -59.675 ;
        RECT -58.645 -61.365 -58.315 -61.035 ;
        RECT -58.645 -62.725 -58.315 -62.395 ;
        RECT -58.645 -64.085 -58.315 -63.755 ;
        RECT -58.645 -65.445 -58.315 -65.115 ;
        RECT -58.645 -66.805 -58.315 -66.475 ;
        RECT -58.645 -68.165 -58.315 -67.835 ;
        RECT -58.645 -69.525 -58.315 -69.195 ;
        RECT -58.645 -70.885 -58.315 -70.555 ;
        RECT -58.645 -72.245 -58.315 -71.915 ;
        RECT -58.645 -73.605 -58.315 -73.275 ;
        RECT -58.645 -74.965 -58.315 -74.635 ;
        RECT -58.645 -76.325 -58.315 -75.995 ;
        RECT -58.645 -77.685 -58.315 -77.355 ;
        RECT -58.645 -79.045 -58.315 -78.715 ;
        RECT -58.645 -80.405 -58.315 -80.075 ;
        RECT -58.645 -81.765 -58.315 -81.435 ;
        RECT -58.645 -83.125 -58.315 -82.795 ;
        RECT -58.645 -84.485 -58.315 -84.155 ;
        RECT -58.645 -85.845 -58.315 -85.515 ;
        RECT -58.645 -87.205 -58.315 -86.875 ;
        RECT -58.645 -88.565 -58.315 -88.235 ;
        RECT -58.645 -89.925 -58.315 -89.595 ;
        RECT -58.645 -91.285 -58.315 -90.955 ;
        RECT -58.645 -94.005 -58.315 -93.675 ;
        RECT -58.645 -95.365 -58.315 -95.035 ;
        RECT -58.645 -96.725 -58.315 -96.395 ;
        RECT -58.645 -98.085 -58.315 -97.755 ;
        RECT -58.645 -99.445 -58.315 -99.115 ;
        RECT -58.645 -100.805 -58.315 -100.475 ;
        RECT -58.645 -102.165 -58.315 -101.835 ;
        RECT -58.645 -103.525 -58.315 -103.195 ;
        RECT -58.645 -104.885 -58.315 -104.555 ;
        RECT -58.645 -106.245 -58.315 -105.915 ;
        RECT -58.645 -107.605 -58.315 -107.275 ;
        RECT -58.645 -108.965 -58.315 -108.635 ;
        RECT -58.645 -110.325 -58.315 -109.995 ;
        RECT -58.645 -111.685 -58.315 -111.355 ;
        RECT -58.645 -113.045 -58.315 -112.715 ;
        RECT -58.645 -114.405 -58.315 -114.075 ;
        RECT -58.645 -115.765 -58.315 -115.435 ;
        RECT -58.645 -117.125 -58.315 -116.795 ;
        RECT -58.645 -118.485 -58.315 -118.155 ;
        RECT -58.645 -119.845 -58.315 -119.515 ;
        RECT -58.645 -121.205 -58.315 -120.875 ;
        RECT -58.645 -122.565 -58.315 -122.235 ;
        RECT -58.645 -123.925 -58.315 -123.595 ;
        RECT -58.645 -125.285 -58.315 -124.955 ;
        RECT -58.645 -126.645 -58.315 -126.315 ;
        RECT -58.645 -128.005 -58.315 -127.675 ;
        RECT -58.645 -129.365 -58.315 -129.035 ;
        RECT -58.645 -130.725 -58.315 -130.395 ;
        RECT -58.645 -132.085 -58.315 -131.755 ;
        RECT -58.645 -133.445 -58.315 -133.115 ;
        RECT -58.645 -134.805 -58.315 -134.475 ;
        RECT -58.645 -136.165 -58.315 -135.835 ;
        RECT -58.645 -137.525 -58.315 -137.195 ;
        RECT -58.645 -138.885 -58.315 -138.555 ;
        RECT -58.645 -140.245 -58.315 -139.915 ;
        RECT -58.645 -141.605 -58.315 -141.275 ;
        RECT -58.645 -142.965 -58.315 -142.635 ;
        RECT -58.645 -144.325 -58.315 -143.995 ;
        RECT -58.645 -145.685 -58.315 -145.355 ;
        RECT -58.645 -147.045 -58.315 -146.715 ;
        RECT -58.645 -149.765 -58.315 -149.435 ;
        RECT -58.64 -151.8 -58.32 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.285 127.225 -56.955 128.355 ;
        RECT -57.285 124.955 -56.955 125.285 ;
        RECT -57.285 123.595 -56.955 123.925 ;
        RECT -57.285 122.235 -56.955 122.565 ;
        RECT -57.285 120.875 -56.955 121.205 ;
        RECT -57.285 119.515 -56.955 119.845 ;
        RECT -57.285 118.155 -56.955 118.485 ;
        RECT -57.285 116.795 -56.955 117.125 ;
        RECT -57.285 115.435 -56.955 115.765 ;
        RECT -57.285 114.075 -56.955 114.405 ;
        RECT -57.285 112.715 -56.955 113.045 ;
        RECT -57.285 111.355 -56.955 111.685 ;
        RECT -57.285 109.995 -56.955 110.325 ;
        RECT -57.285 108.635 -56.955 108.965 ;
        RECT -57.285 107.275 -56.955 107.605 ;
        RECT -57.285 105.915 -56.955 106.245 ;
        RECT -57.285 104.555 -56.955 104.885 ;
        RECT -57.285 103.195 -56.955 103.525 ;
        RECT -57.285 101.835 -56.955 102.165 ;
        RECT -57.285 100.475 -56.955 100.805 ;
        RECT -57.285 99.115 -56.955 99.445 ;
        RECT -57.285 97.755 -56.955 98.085 ;
        RECT -57.285 96.395 -56.955 96.725 ;
        RECT -57.285 95.035 -56.955 95.365 ;
        RECT -57.285 93.675 -56.955 94.005 ;
        RECT -57.285 92.315 -56.955 92.645 ;
        RECT -57.285 90.955 -56.955 91.285 ;
        RECT -57.285 89.595 -56.955 89.925 ;
        RECT -57.285 88.235 -56.955 88.565 ;
        RECT -57.285 86.875 -56.955 87.205 ;
        RECT -57.285 85.515 -56.955 85.845 ;
        RECT -57.285 84.155 -56.955 84.485 ;
        RECT -57.285 82.795 -56.955 83.125 ;
        RECT -57.285 81.435 -56.955 81.765 ;
        RECT -57.285 80.075 -56.955 80.405 ;
        RECT -57.285 78.715 -56.955 79.045 ;
        RECT -57.285 77.355 -56.955 77.685 ;
        RECT -57.285 75.995 -56.955 76.325 ;
        RECT -57.285 74.635 -56.955 74.965 ;
        RECT -57.285 73.275 -56.955 73.605 ;
        RECT -57.285 72.445 -56.955 72.775 ;
        RECT -57.285 70.395 -56.955 70.725 ;
        RECT -57.285 68.035 -56.955 68.365 ;
        RECT -57.285 66.885 -56.955 67.215 ;
        RECT -57.285 64.875 -56.955 65.205 ;
        RECT -57.285 63.725 -56.955 64.055 ;
        RECT -57.285 61.715 -56.955 62.045 ;
        RECT -57.285 60.395 -56.955 60.725 ;
        RECT -57.285 58.555 -56.955 58.885 ;
        RECT -57.285 57.405 -56.955 57.735 ;
        RECT -57.285 55.395 -56.955 55.725 ;
        RECT -57.285 54.245 -56.955 54.575 ;
        RECT -57.285 51.885 -56.955 52.215 ;
        RECT -57.285 49.83 -56.955 50.16 ;
        RECT -57.285 48.795 -56.955 49.125 ;
        RECT -57.285 47.435 -56.955 47.765 ;
        RECT -57.285 46.075 -56.955 46.405 ;
        RECT -57.285 44.715 -56.955 45.045 ;
        RECT -57.285 43.355 -56.955 43.685 ;
        RECT -57.285 41.995 -56.955 42.325 ;
        RECT -57.285 40.635 -56.955 40.965 ;
        RECT -57.285 39.275 -56.955 39.605 ;
        RECT -57.285 37.915 -56.955 38.245 ;
        RECT -57.285 36.555 -56.955 36.885 ;
        RECT -57.285 35.195 -56.955 35.525 ;
        RECT -57.285 33.835 -56.955 34.165 ;
        RECT -57.285 32.475 -56.955 32.805 ;
        RECT -57.285 31.115 -56.955 31.445 ;
        RECT -57.285 29.755 -56.955 30.085 ;
        RECT -57.285 28.395 -56.955 28.725 ;
        RECT -57.285 27.035 -56.955 27.365 ;
        RECT -57.285 25.675 -56.955 26.005 ;
        RECT -57.285 24.315 -56.955 24.645 ;
        RECT -57.285 22.955 -56.955 23.285 ;
        RECT -57.285 21.595 -56.955 21.925 ;
        RECT -57.285 20.235 -56.955 20.565 ;
        RECT -57.285 18.875 -56.955 19.205 ;
        RECT -57.285 17.515 -56.955 17.845 ;
        RECT -57.285 16.155 -56.955 16.485 ;
        RECT -57.285 14.795 -56.955 15.125 ;
        RECT -57.285 13.435 -56.955 13.765 ;
        RECT -57.285 12.075 -56.955 12.405 ;
        RECT -57.285 10.715 -56.955 11.045 ;
        RECT -57.285 9.355 -56.955 9.685 ;
        RECT -57.285 7.995 -56.955 8.325 ;
        RECT -57.285 6.635 -56.955 6.965 ;
        RECT -57.285 5.275 -56.955 5.605 ;
        RECT -57.285 3.915 -56.955 4.245 ;
        RECT -57.285 2.555 -56.955 2.885 ;
        RECT -57.285 1.195 -56.955 1.525 ;
        RECT -57.285 -0.165 -56.955 0.165 ;
        RECT -57.285 -1.525 -56.955 -1.195 ;
        RECT -57.285 -2.885 -56.955 -2.555 ;
        RECT -57.285 -4.245 -56.955 -3.915 ;
        RECT -57.285 -5.605 -56.955 -5.275 ;
        RECT -57.285 -6.965 -56.955 -6.635 ;
        RECT -57.285 -8.325 -56.955 -7.995 ;
        RECT -57.285 -9.685 -56.955 -9.355 ;
        RECT -57.285 -11.045 -56.955 -10.715 ;
        RECT -57.285 -12.405 -56.955 -12.075 ;
        RECT -57.285 -13.765 -56.955 -13.435 ;
        RECT -57.285 -15.125 -56.955 -14.795 ;
        RECT -57.285 -16.485 -56.955 -16.155 ;
        RECT -57.285 -17.845 -56.955 -17.515 ;
        RECT -57.285 -19.205 -56.955 -18.875 ;
        RECT -57.285 -20.565 -56.955 -20.235 ;
        RECT -57.285 -21.925 -56.955 -21.595 ;
        RECT -57.285 -23.285 -56.955 -22.955 ;
        RECT -57.285 -24.645 -56.955 -24.315 ;
        RECT -57.285 -26.005 -56.955 -25.675 ;
        RECT -57.285 -27.365 -56.955 -27.035 ;
        RECT -57.285 -28.725 -56.955 -28.395 ;
        RECT -57.285 -30.085 -56.955 -29.755 ;
        RECT -57.285 -31.445 -56.955 -31.115 ;
        RECT -57.285 -32.805 -56.955 -32.475 ;
        RECT -57.285 -34.165 -56.955 -33.835 ;
        RECT -57.285 -35.525 -56.955 -35.195 ;
        RECT -57.285 -36.885 -56.955 -36.555 ;
        RECT -57.285 -38.245 -56.955 -37.915 ;
        RECT -57.285 -39.605 -56.955 -39.275 ;
        RECT -57.285 -40.965 -56.955 -40.635 ;
        RECT -57.285 -42.325 -56.955 -41.995 ;
        RECT -57.285 -43.685 -56.955 -43.355 ;
        RECT -57.285 -45.045 -56.955 -44.715 ;
        RECT -57.285 -46.405 -56.955 -46.075 ;
        RECT -57.285 -47.765 -56.955 -47.435 ;
        RECT -57.285 -49.125 -56.955 -48.795 ;
        RECT -57.285 -50.485 -56.955 -50.155 ;
        RECT -57.285 -51.845 -56.955 -51.515 ;
        RECT -57.285 -53.205 -56.955 -52.875 ;
        RECT -57.285 -54.565 -56.955 -54.235 ;
        RECT -57.285 -55.925 -56.955 -55.595 ;
        RECT -57.285 -57.285 -56.955 -56.955 ;
        RECT -57.285 -58.645 -56.955 -58.315 ;
        RECT -57.285 -60.005 -56.955 -59.675 ;
        RECT -57.285 -61.365 -56.955 -61.035 ;
        RECT -57.285 -62.725 -56.955 -62.395 ;
        RECT -57.285 -64.085 -56.955 -63.755 ;
        RECT -57.285 -65.445 -56.955 -65.115 ;
        RECT -57.285 -66.805 -56.955 -66.475 ;
        RECT -57.285 -68.165 -56.955 -67.835 ;
        RECT -57.285 -69.525 -56.955 -69.195 ;
        RECT -57.285 -70.885 -56.955 -70.555 ;
        RECT -57.285 -72.245 -56.955 -71.915 ;
        RECT -57.285 -73.605 -56.955 -73.275 ;
        RECT -57.285 -74.965 -56.955 -74.635 ;
        RECT -57.285 -76.325 -56.955 -75.995 ;
        RECT -57.285 -77.685 -56.955 -77.355 ;
        RECT -57.285 -79.045 -56.955 -78.715 ;
        RECT -57.285 -80.405 -56.955 -80.075 ;
        RECT -57.285 -81.765 -56.955 -81.435 ;
        RECT -57.285 -83.125 -56.955 -82.795 ;
        RECT -57.285 -84.485 -56.955 -84.155 ;
        RECT -57.285 -85.845 -56.955 -85.515 ;
        RECT -57.285 -87.205 -56.955 -86.875 ;
        RECT -57.285 -88.565 -56.955 -88.235 ;
        RECT -57.285 -89.925 -56.955 -89.595 ;
        RECT -57.285 -91.285 -56.955 -90.955 ;
        RECT -57.285 -94.005 -56.955 -93.675 ;
        RECT -57.285 -95.365 -56.955 -95.035 ;
        RECT -57.285 -96.725 -56.955 -96.395 ;
        RECT -57.285 -98.085 -56.955 -97.755 ;
        RECT -57.285 -99.445 -56.955 -99.115 ;
        RECT -57.285 -100.805 -56.955 -100.475 ;
        RECT -57.285 -102.165 -56.955 -101.835 ;
        RECT -57.285 -103.525 -56.955 -103.195 ;
        RECT -57.285 -104.885 -56.955 -104.555 ;
        RECT -57.285 -106.245 -56.955 -105.915 ;
        RECT -57.285 -107.605 -56.955 -107.275 ;
        RECT -57.285 -108.965 -56.955 -108.635 ;
        RECT -57.285 -110.325 -56.955 -109.995 ;
        RECT -57.285 -111.685 -56.955 -111.355 ;
        RECT -57.285 -113.045 -56.955 -112.715 ;
        RECT -57.285 -114.405 -56.955 -114.075 ;
        RECT -57.285 -115.765 -56.955 -115.435 ;
        RECT -57.285 -117.125 -56.955 -116.795 ;
        RECT -57.285 -118.485 -56.955 -118.155 ;
        RECT -57.285 -119.845 -56.955 -119.515 ;
        RECT -57.285 -121.205 -56.955 -120.875 ;
        RECT -57.285 -122.565 -56.955 -122.235 ;
        RECT -57.285 -123.925 -56.955 -123.595 ;
        RECT -57.285 -125.285 -56.955 -124.955 ;
        RECT -57.285 -126.645 -56.955 -126.315 ;
        RECT -57.285 -128.005 -56.955 -127.675 ;
        RECT -57.285 -129.365 -56.955 -129.035 ;
        RECT -57.285 -130.725 -56.955 -130.395 ;
        RECT -57.285 -132.085 -56.955 -131.755 ;
        RECT -57.285 -133.445 -56.955 -133.115 ;
        RECT -57.285 -134.805 -56.955 -134.475 ;
        RECT -57.285 -136.165 -56.955 -135.835 ;
        RECT -57.285 -137.525 -56.955 -137.195 ;
        RECT -57.285 -138.885 -56.955 -138.555 ;
        RECT -57.285 -140.245 -56.955 -139.915 ;
        RECT -57.285 -141.605 -56.955 -141.275 ;
        RECT -57.285 -142.965 -56.955 -142.635 ;
        RECT -57.285 -144.325 -56.955 -143.995 ;
        RECT -57.285 -145.685 -56.955 -145.355 ;
        RECT -57.285 -147.045 -56.955 -146.715 ;
        RECT -57.285 -149.765 -56.955 -149.435 ;
        RECT -57.285 -152.485 -56.955 -152.155 ;
        RECT -57.285 -153.845 -56.955 -153.515 ;
        RECT -57.285 -155.285 -56.955 -154.955 ;
        RECT -57.285 -156.565 -56.955 -156.235 ;
        RECT -57.285 -157.925 -56.955 -157.595 ;
        RECT -57.285 -160.17 -56.955 -159.04 ;
        RECT -57.28 -160.285 -56.96 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 127.225 -55.595 128.355 ;
        RECT -55.925 124.955 -55.595 125.285 ;
        RECT -55.925 123.595 -55.595 123.925 ;
        RECT -55.925 122.235 -55.595 122.565 ;
        RECT -55.925 120.875 -55.595 121.205 ;
        RECT -55.925 119.515 -55.595 119.845 ;
        RECT -55.925 118.155 -55.595 118.485 ;
        RECT -55.925 116.795 -55.595 117.125 ;
        RECT -55.925 115.435 -55.595 115.765 ;
        RECT -55.925 114.075 -55.595 114.405 ;
        RECT -55.925 112.715 -55.595 113.045 ;
        RECT -55.925 111.355 -55.595 111.685 ;
        RECT -55.925 109.995 -55.595 110.325 ;
        RECT -55.925 108.635 -55.595 108.965 ;
        RECT -55.925 107.275 -55.595 107.605 ;
        RECT -55.925 105.915 -55.595 106.245 ;
        RECT -55.925 104.555 -55.595 104.885 ;
        RECT -55.925 103.195 -55.595 103.525 ;
        RECT -55.925 101.835 -55.595 102.165 ;
        RECT -55.925 100.475 -55.595 100.805 ;
        RECT -55.925 99.115 -55.595 99.445 ;
        RECT -55.925 97.755 -55.595 98.085 ;
        RECT -55.925 96.395 -55.595 96.725 ;
        RECT -55.925 95.035 -55.595 95.365 ;
        RECT -55.925 93.675 -55.595 94.005 ;
        RECT -55.925 92.315 -55.595 92.645 ;
        RECT -55.925 90.955 -55.595 91.285 ;
        RECT -55.925 89.595 -55.595 89.925 ;
        RECT -55.925 88.235 -55.595 88.565 ;
        RECT -55.925 86.875 -55.595 87.205 ;
        RECT -55.925 85.515 -55.595 85.845 ;
        RECT -55.925 84.155 -55.595 84.485 ;
        RECT -55.925 82.795 -55.595 83.125 ;
        RECT -55.925 81.435 -55.595 81.765 ;
        RECT -55.925 80.075 -55.595 80.405 ;
        RECT -55.925 78.715 -55.595 79.045 ;
        RECT -55.925 77.355 -55.595 77.685 ;
        RECT -55.925 75.995 -55.595 76.325 ;
        RECT -55.925 74.635 -55.595 74.965 ;
        RECT -55.925 73.275 -55.595 73.605 ;
        RECT -55.925 72.445 -55.595 72.775 ;
        RECT -55.925 70.395 -55.595 70.725 ;
        RECT -55.925 68.035 -55.595 68.365 ;
        RECT -55.925 66.885 -55.595 67.215 ;
        RECT -55.925 64.875 -55.595 65.205 ;
        RECT -55.925 63.725 -55.595 64.055 ;
        RECT -55.925 61.715 -55.595 62.045 ;
        RECT -55.925 60.395 -55.595 60.725 ;
        RECT -55.925 58.555 -55.595 58.885 ;
        RECT -55.925 57.405 -55.595 57.735 ;
        RECT -55.925 55.395 -55.595 55.725 ;
        RECT -55.925 54.245 -55.595 54.575 ;
        RECT -55.925 51.885 -55.595 52.215 ;
        RECT -55.925 49.83 -55.595 50.16 ;
        RECT -55.925 48.795 -55.595 49.125 ;
        RECT -55.925 47.435 -55.595 47.765 ;
        RECT -55.925 46.075 -55.595 46.405 ;
        RECT -55.925 44.715 -55.595 45.045 ;
        RECT -55.925 43.355 -55.595 43.685 ;
        RECT -55.925 41.995 -55.595 42.325 ;
        RECT -55.925 40.635 -55.595 40.965 ;
        RECT -55.925 39.275 -55.595 39.605 ;
        RECT -55.92 37.92 -55.6 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 -102.165 -55.595 -101.835 ;
        RECT -55.925 -103.525 -55.595 -103.195 ;
        RECT -55.925 -104.885 -55.595 -104.555 ;
        RECT -55.925 -106.245 -55.595 -105.915 ;
        RECT -55.925 -107.605 -55.595 -107.275 ;
        RECT -55.925 -108.965 -55.595 -108.635 ;
        RECT -55.925 -110.325 -55.595 -109.995 ;
        RECT -55.925 -111.685 -55.595 -111.355 ;
        RECT -55.925 -113.045 -55.595 -112.715 ;
        RECT -55.925 -114.405 -55.595 -114.075 ;
        RECT -55.925 -115.765 -55.595 -115.435 ;
        RECT -55.925 -117.125 -55.595 -116.795 ;
        RECT -55.925 -118.485 -55.595 -118.155 ;
        RECT -55.925 -119.845 -55.595 -119.515 ;
        RECT -55.925 -121.205 -55.595 -120.875 ;
        RECT -55.925 -122.565 -55.595 -122.235 ;
        RECT -55.925 -123.925 -55.595 -123.595 ;
        RECT -55.925 -125.285 -55.595 -124.955 ;
        RECT -55.925 -126.645 -55.595 -126.315 ;
        RECT -55.925 -128.005 -55.595 -127.675 ;
        RECT -55.925 -129.365 -55.595 -129.035 ;
        RECT -55.925 -130.725 -55.595 -130.395 ;
        RECT -55.925 -132.085 -55.595 -131.755 ;
        RECT -55.925 -133.445 -55.595 -133.115 ;
        RECT -55.925 -134.805 -55.595 -134.475 ;
        RECT -55.925 -136.165 -55.595 -135.835 ;
        RECT -55.925 -137.525 -55.595 -137.195 ;
        RECT -55.925 -138.885 -55.595 -138.555 ;
        RECT -55.925 -140.245 -55.595 -139.915 ;
        RECT -55.925 -141.605 -55.595 -141.275 ;
        RECT -55.925 -142.965 -55.595 -142.635 ;
        RECT -55.925 -144.325 -55.595 -143.995 ;
        RECT -55.925 -145.685 -55.595 -145.355 ;
        RECT -55.925 -147.045 -55.595 -146.715 ;
        RECT -55.925 -149.765 -55.595 -149.435 ;
        RECT -55.925 -152.485 -55.595 -152.155 ;
        RECT -55.925 -153.845 -55.595 -153.515 ;
        RECT -55.925 -155.285 -55.595 -154.955 ;
        RECT -55.925 -156.565 -55.595 -156.235 ;
        RECT -55.925 -157.925 -55.595 -157.595 ;
        RECT -55.925 -160.17 -55.595 -159.04 ;
        RECT -55.92 -160.285 -55.6 -101.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 127.225 -54.235 128.355 ;
        RECT -54.565 124.955 -54.235 125.285 ;
        RECT -54.565 123.595 -54.235 123.925 ;
        RECT -54.565 122.235 -54.235 122.565 ;
        RECT -54.565 120.875 -54.235 121.205 ;
        RECT -54.565 119.515 -54.235 119.845 ;
        RECT -54.565 118.155 -54.235 118.485 ;
        RECT -54.565 116.795 -54.235 117.125 ;
        RECT -54.565 115.435 -54.235 115.765 ;
        RECT -54.565 114.075 -54.235 114.405 ;
        RECT -54.565 112.715 -54.235 113.045 ;
        RECT -54.565 111.355 -54.235 111.685 ;
        RECT -54.565 109.995 -54.235 110.325 ;
        RECT -54.565 108.635 -54.235 108.965 ;
        RECT -54.565 107.275 -54.235 107.605 ;
        RECT -54.565 105.915 -54.235 106.245 ;
        RECT -54.565 104.555 -54.235 104.885 ;
        RECT -54.565 103.195 -54.235 103.525 ;
        RECT -54.565 101.835 -54.235 102.165 ;
        RECT -54.565 100.475 -54.235 100.805 ;
        RECT -54.565 99.115 -54.235 99.445 ;
        RECT -54.565 97.755 -54.235 98.085 ;
        RECT -54.565 96.395 -54.235 96.725 ;
        RECT -54.565 95.035 -54.235 95.365 ;
        RECT -54.565 93.675 -54.235 94.005 ;
        RECT -54.565 92.315 -54.235 92.645 ;
        RECT -54.565 90.955 -54.235 91.285 ;
        RECT -54.565 89.595 -54.235 89.925 ;
        RECT -54.565 88.235 -54.235 88.565 ;
        RECT -54.565 86.875 -54.235 87.205 ;
        RECT -54.565 85.515 -54.235 85.845 ;
        RECT -54.565 84.155 -54.235 84.485 ;
        RECT -54.565 82.795 -54.235 83.125 ;
        RECT -54.565 81.435 -54.235 81.765 ;
        RECT -54.565 80.075 -54.235 80.405 ;
        RECT -54.565 78.715 -54.235 79.045 ;
        RECT -54.565 77.355 -54.235 77.685 ;
        RECT -54.565 75.995 -54.235 76.325 ;
        RECT -54.565 74.635 -54.235 74.965 ;
        RECT -54.565 73.275 -54.235 73.605 ;
        RECT -54.56 73.275 -54.24 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 48.795 -54.235 49.125 ;
        RECT -54.565 47.435 -54.235 47.765 ;
        RECT -54.565 46.075 -54.235 46.405 ;
        RECT -54.565 44.715 -54.235 45.045 ;
        RECT -54.565 43.355 -54.235 43.685 ;
        RECT -54.565 40.635 -54.235 40.965 ;
        RECT -54.565 39.275 -54.235 39.605 ;
        RECT -54.565 35.195 -54.235 35.525 ;
        RECT -54.565 33.835 -54.235 34.165 ;
        RECT -54.565 32.475 -54.235 32.805 ;
        RECT -54.565 31.115 -54.235 31.445 ;
        RECT -54.565 29.755 -54.235 30.085 ;
        RECT -54.565 28.395 -54.235 28.725 ;
        RECT -54.565 27.035 -54.235 27.365 ;
        RECT -54.565 25.675 -54.235 26.005 ;
        RECT -54.565 24.315 -54.235 24.645 ;
        RECT -54.565 22.955 -54.235 23.285 ;
        RECT -54.565 21.595 -54.235 21.925 ;
        RECT -54.565 20.235 -54.235 20.565 ;
        RECT -54.565 18.875 -54.235 19.205 ;
        RECT -54.565 17.515 -54.235 17.845 ;
        RECT -54.565 16.155 -54.235 16.485 ;
        RECT -54.565 14.795 -54.235 15.125 ;
        RECT -54.565 13.435 -54.235 13.765 ;
        RECT -54.565 12.075 -54.235 12.405 ;
        RECT -54.565 10.715 -54.235 11.045 ;
        RECT -54.565 9.355 -54.235 9.685 ;
        RECT -54.565 7.995 -54.235 8.325 ;
        RECT -54.565 6.635 -54.235 6.965 ;
        RECT -54.565 5.275 -54.235 5.605 ;
        RECT -54.565 3.915 -54.235 4.245 ;
        RECT -54.565 2.555 -54.235 2.885 ;
        RECT -54.565 1.195 -54.235 1.525 ;
        RECT -54.565 -0.165 -54.235 0.165 ;
        RECT -54.565 -1.525 -54.235 -1.195 ;
        RECT -54.565 -2.885 -54.235 -2.555 ;
        RECT -54.565 -4.245 -54.235 -3.915 ;
        RECT -54.565 -5.605 -54.235 -5.275 ;
        RECT -54.565 -6.965 -54.235 -6.635 ;
        RECT -54.565 -8.325 -54.235 -7.995 ;
        RECT -54.565 -9.685 -54.235 -9.355 ;
        RECT -54.565 -12.405 -54.235 -12.075 ;
        RECT -54.565 -13.765 -54.235 -13.435 ;
        RECT -54.565 -15.125 -54.235 -14.795 ;
        RECT -54.565 -16.485 -54.235 -16.155 ;
        RECT -54.565 -17.845 -54.235 -17.515 ;
        RECT -54.565 -19.205 -54.235 -18.875 ;
        RECT -54.565 -20.565 -54.235 -20.235 ;
        RECT -54.565 -21.925 -54.235 -21.595 ;
        RECT -54.565 -23.285 -54.235 -22.955 ;
        RECT -54.565 -24.645 -54.235 -24.315 ;
        RECT -54.565 -26.005 -54.235 -25.675 ;
        RECT -54.565 -27.365 -54.235 -27.035 ;
        RECT -54.565 -28.725 -54.235 -28.395 ;
        RECT -54.565 -30.085 -54.235 -29.755 ;
        RECT -54.565 -31.445 -54.235 -31.115 ;
        RECT -54.565 -32.805 -54.235 -32.475 ;
        RECT -54.565 -34.165 -54.235 -33.835 ;
        RECT -54.565 -35.525 -54.235 -35.195 ;
        RECT -54.565 -36.885 -54.235 -36.555 ;
        RECT -54.565 -38.245 -54.235 -37.915 ;
        RECT -54.565 -39.605 -54.235 -39.275 ;
        RECT -54.565 -40.965 -54.235 -40.635 ;
        RECT -54.565 -42.325 -54.235 -41.995 ;
        RECT -54.565 -43.685 -54.235 -43.355 ;
        RECT -54.565 -45.045 -54.235 -44.715 ;
        RECT -54.565 -46.405 -54.235 -46.075 ;
        RECT -54.565 -47.765 -54.235 -47.435 ;
        RECT -54.565 -49.125 -54.235 -48.795 ;
        RECT -54.565 -50.485 -54.235 -50.155 ;
        RECT -54.565 -51.845 -54.235 -51.515 ;
        RECT -54.565 -53.205 -54.235 -52.875 ;
        RECT -54.565 -54.565 -54.235 -54.235 ;
        RECT -54.565 -55.925 -54.235 -55.595 ;
        RECT -54.565 -57.285 -54.235 -56.955 ;
        RECT -54.565 -58.645 -54.235 -58.315 ;
        RECT -54.565 -60.005 -54.235 -59.675 ;
        RECT -54.565 -61.365 -54.235 -61.035 ;
        RECT -54.565 -62.725 -54.235 -62.395 ;
        RECT -54.565 -64.085 -54.235 -63.755 ;
        RECT -54.565 -65.445 -54.235 -65.115 ;
        RECT -54.565 -66.805 -54.235 -66.475 ;
        RECT -54.565 -68.165 -54.235 -67.835 ;
        RECT -54.565 -69.525 -54.235 -69.195 ;
        RECT -54.565 -72.245 -54.235 -71.915 ;
        RECT -54.565 -73.605 -54.235 -73.275 ;
        RECT -54.565 -74.965 -54.235 -74.635 ;
        RECT -54.565 -76.325 -54.235 -75.995 ;
        RECT -54.565 -78.29 -54.235 -77.96 ;
        RECT -54.565 -79.045 -54.235 -78.715 ;
        RECT -54.565 -81.765 -54.235 -81.435 ;
        RECT -54.565 -83.125 -54.235 -82.795 ;
        RECT -54.565 -84.485 -54.235 -84.155 ;
        RECT -54.565 -86.43 -54.235 -86.1 ;
        RECT -54.565 -87.205 -54.235 -86.875 ;
        RECT -54.565 -88.565 -54.235 -88.235 ;
        RECT -54.565 -89.925 -54.235 -89.595 ;
        RECT -54.565 -94.005 -54.235 -93.675 ;
        RECT -54.565 -95.365 -54.235 -95.035 ;
        RECT -54.565 -96.725 -54.235 -96.395 ;
        RECT -54.565 -98.085 -54.235 -97.755 ;
        RECT -54.565 -102.165 -54.235 -101.835 ;
        RECT -54.565 -103.525 -54.235 -103.195 ;
        RECT -54.565 -104.885 -54.235 -104.555 ;
        RECT -54.565 -106.245 -54.235 -105.915 ;
        RECT -54.565 -107.605 -54.235 -107.275 ;
        RECT -54.565 -108.965 -54.235 -108.635 ;
        RECT -54.565 -110.325 -54.235 -109.995 ;
        RECT -54.565 -111.685 -54.235 -111.355 ;
        RECT -54.565 -113.045 -54.235 -112.715 ;
        RECT -54.565 -114.405 -54.235 -114.075 ;
        RECT -54.565 -115.765 -54.235 -115.435 ;
        RECT -54.565 -117.125 -54.235 -116.795 ;
        RECT -54.565 -118.485 -54.235 -118.155 ;
        RECT -54.565 -119.845 -54.235 -119.515 ;
        RECT -54.565 -121.205 -54.235 -120.875 ;
        RECT -54.565 -122.565 -54.235 -122.235 ;
        RECT -54.565 -123.925 -54.235 -123.595 ;
        RECT -54.565 -125.285 -54.235 -124.955 ;
        RECT -54.565 -126.645 -54.235 -126.315 ;
        RECT -54.565 -128.005 -54.235 -127.675 ;
        RECT -54.565 -129.365 -54.235 -129.035 ;
        RECT -54.565 -130.725 -54.235 -130.395 ;
        RECT -54.565 -132.085 -54.235 -131.755 ;
        RECT -54.565 -133.445 -54.235 -133.115 ;
        RECT -54.565 -134.805 -54.235 -134.475 ;
        RECT -54.565 -136.165 -54.235 -135.835 ;
        RECT -54.565 -137.525 -54.235 -137.195 ;
        RECT -54.565 -138.885 -54.235 -138.555 ;
        RECT -54.565 -140.245 -54.235 -139.915 ;
        RECT -54.565 -141.605 -54.235 -141.275 ;
        RECT -54.565 -142.965 -54.235 -142.635 ;
        RECT -54.565 -144.325 -54.235 -143.995 ;
        RECT -54.565 -145.685 -54.235 -145.355 ;
        RECT -54.565 -147.045 -54.235 -146.715 ;
        RECT -54.565 -149.765 -54.235 -149.435 ;
        RECT -54.565 -153.845 -54.235 -153.515 ;
        RECT -54.565 -155.285 -54.235 -154.955 ;
        RECT -54.565 -156.565 -54.235 -156.235 ;
        RECT -54.565 -157.925 -54.235 -157.595 ;
        RECT -54.565 -160.17 -54.235 -159.04 ;
        RECT -54.56 -160.285 -54.24 49.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 127.225 -52.875 128.355 ;
        RECT -53.205 124.955 -52.875 125.285 ;
        RECT -53.205 123.595 -52.875 123.925 ;
        RECT -53.205 122.235 -52.875 122.565 ;
        RECT -53.205 120.875 -52.875 121.205 ;
        RECT -53.205 119.515 -52.875 119.845 ;
        RECT -53.205 118.155 -52.875 118.485 ;
        RECT -53.205 116.795 -52.875 117.125 ;
        RECT -53.205 115.435 -52.875 115.765 ;
        RECT -53.205 114.075 -52.875 114.405 ;
        RECT -53.205 112.715 -52.875 113.045 ;
        RECT -53.205 111.355 -52.875 111.685 ;
        RECT -53.205 109.995 -52.875 110.325 ;
        RECT -53.205 108.635 -52.875 108.965 ;
        RECT -53.205 107.275 -52.875 107.605 ;
        RECT -53.205 105.915 -52.875 106.245 ;
        RECT -53.205 104.555 -52.875 104.885 ;
        RECT -53.205 103.195 -52.875 103.525 ;
        RECT -53.205 101.835 -52.875 102.165 ;
        RECT -53.205 100.475 -52.875 100.805 ;
        RECT -53.205 99.115 -52.875 99.445 ;
        RECT -53.205 97.755 -52.875 98.085 ;
        RECT -53.205 96.395 -52.875 96.725 ;
        RECT -53.205 95.035 -52.875 95.365 ;
        RECT -53.205 93.675 -52.875 94.005 ;
        RECT -53.205 92.315 -52.875 92.645 ;
        RECT -53.205 90.955 -52.875 91.285 ;
        RECT -53.205 89.595 -52.875 89.925 ;
        RECT -53.205 88.235 -52.875 88.565 ;
        RECT -53.205 86.875 -52.875 87.205 ;
        RECT -53.205 85.515 -52.875 85.845 ;
        RECT -53.205 84.155 -52.875 84.485 ;
        RECT -53.205 82.795 -52.875 83.125 ;
        RECT -53.205 81.435 -52.875 81.765 ;
        RECT -53.205 80.075 -52.875 80.405 ;
        RECT -53.205 78.715 -52.875 79.045 ;
        RECT -53.205 77.355 -52.875 77.685 ;
        RECT -53.205 75.995 -52.875 76.325 ;
        RECT -53.205 74.635 -52.875 74.965 ;
        RECT -53.205 73.275 -52.875 73.605 ;
        RECT -53.2 73.275 -52.88 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 -4.245 -52.875 -3.915 ;
        RECT -53.205 -5.605 -52.875 -5.275 ;
        RECT -53.205 -6.965 -52.875 -6.635 ;
        RECT -53.205 -8.325 -52.875 -7.995 ;
        RECT -53.205 -9.685 -52.875 -9.355 ;
        RECT -53.205 -12.405 -52.875 -12.075 ;
        RECT -53.205 -13.765 -52.875 -13.435 ;
        RECT -53.205 -15.125 -52.875 -14.795 ;
        RECT -53.205 -16.485 -52.875 -16.155 ;
        RECT -53.205 -17.845 -52.875 -17.515 ;
        RECT -53.205 -19.205 -52.875 -18.875 ;
        RECT -53.205 -20.565 -52.875 -20.235 ;
        RECT -53.205 -21.925 -52.875 -21.595 ;
        RECT -53.205 -24.645 -52.875 -24.315 ;
        RECT -53.205 -26.005 -52.875 -25.675 ;
        RECT -53.205 -27.365 -52.875 -27.035 ;
        RECT -53.205 -28.725 -52.875 -28.395 ;
        RECT -53.205 -30.085 -52.875 -29.755 ;
        RECT -53.205 -31.445 -52.875 -31.115 ;
        RECT -53.205 -32.805 -52.875 -32.475 ;
        RECT -53.205 -34.165 -52.875 -33.835 ;
        RECT -53.205 -35.525 -52.875 -35.195 ;
        RECT -53.205 -36.885 -52.875 -36.555 ;
        RECT -53.205 -38.245 -52.875 -37.915 ;
        RECT -53.205 -39.605 -52.875 -39.275 ;
        RECT -53.205 -40.965 -52.875 -40.635 ;
        RECT -53.205 -42.325 -52.875 -41.995 ;
        RECT -53.205 -43.685 -52.875 -43.355 ;
        RECT -53.205 -45.045 -52.875 -44.715 ;
        RECT -53.205 -46.405 -52.875 -46.075 ;
        RECT -53.205 -47.765 -52.875 -47.435 ;
        RECT -53.205 -49.125 -52.875 -48.795 ;
        RECT -53.205 -50.485 -52.875 -50.155 ;
        RECT -53.205 -51.845 -52.875 -51.515 ;
        RECT -53.205 -53.205 -52.875 -52.875 ;
        RECT -53.205 -54.565 -52.875 -54.235 ;
        RECT -53.205 -55.925 -52.875 -55.595 ;
        RECT -53.205 -57.285 -52.875 -56.955 ;
        RECT -53.205 -58.645 -52.875 -58.315 ;
        RECT -53.205 -60.005 -52.875 -59.675 ;
        RECT -53.205 -61.365 -52.875 -61.035 ;
        RECT -53.205 -62.725 -52.875 -62.395 ;
        RECT -53.205 -64.085 -52.875 -63.755 ;
        RECT -53.205 -65.445 -52.875 -65.115 ;
        RECT -53.205 -66.805 -52.875 -66.475 ;
        RECT -53.205 -68.165 -52.875 -67.835 ;
        RECT -53.205 -69.525 -52.875 -69.195 ;
        RECT -53.205 -72.245 -52.875 -71.915 ;
        RECT -53.205 -73.605 -52.875 -73.275 ;
        RECT -53.205 -74.965 -52.875 -74.635 ;
        RECT -53.205 -76.325 -52.875 -75.995 ;
        RECT -53.205 -78.29 -52.875 -77.96 ;
        RECT -53.205 -79.045 -52.875 -78.715 ;
        RECT -53.205 -81.765 -52.875 -81.435 ;
        RECT -53.205 -83.125 -52.875 -82.795 ;
        RECT -53.205 -84.485 -52.875 -84.155 ;
        RECT -53.205 -86.43 -52.875 -86.1 ;
        RECT -53.205 -87.205 -52.875 -86.875 ;
        RECT -53.205 -88.565 -52.875 -88.235 ;
        RECT -53.205 -89.925 -52.875 -89.595 ;
        RECT -53.205 -94.005 -52.875 -93.675 ;
        RECT -53.205 -95.365 -52.875 -95.035 ;
        RECT -53.205 -96.725 -52.875 -96.395 ;
        RECT -53.205 -98.085 -52.875 -97.755 ;
        RECT -53.205 -102.165 -52.875 -101.835 ;
        RECT -53.205 -103.525 -52.875 -103.195 ;
        RECT -53.205 -104.885 -52.875 -104.555 ;
        RECT -53.205 -106.245 -52.875 -105.915 ;
        RECT -53.205 -107.605 -52.875 -107.275 ;
        RECT -53.205 -108.965 -52.875 -108.635 ;
        RECT -53.205 -110.325 -52.875 -109.995 ;
        RECT -53.205 -111.685 -52.875 -111.355 ;
        RECT -53.205 -113.045 -52.875 -112.715 ;
        RECT -53.205 -114.405 -52.875 -114.075 ;
        RECT -53.205 -115.765 -52.875 -115.435 ;
        RECT -53.205 -117.125 -52.875 -116.795 ;
        RECT -53.205 -118.485 -52.875 -118.155 ;
        RECT -53.205 -119.845 -52.875 -119.515 ;
        RECT -53.205 -121.205 -52.875 -120.875 ;
        RECT -53.205 -122.565 -52.875 -122.235 ;
        RECT -53.205 -123.925 -52.875 -123.595 ;
        RECT -53.205 -125.285 -52.875 -124.955 ;
        RECT -53.205 -126.645 -52.875 -126.315 ;
        RECT -53.205 -128.005 -52.875 -127.675 ;
        RECT -53.205 -129.365 -52.875 -129.035 ;
        RECT -53.205 -130.725 -52.875 -130.395 ;
        RECT -53.205 -132.085 -52.875 -131.755 ;
        RECT -53.205 -133.445 -52.875 -133.115 ;
        RECT -53.205 -134.805 -52.875 -134.475 ;
        RECT -53.205 -136.165 -52.875 -135.835 ;
        RECT -53.205 -137.525 -52.875 -137.195 ;
        RECT -53.205 -138.885 -52.875 -138.555 ;
        RECT -53.205 -140.245 -52.875 -139.915 ;
        RECT -53.205 -141.605 -52.875 -141.275 ;
        RECT -53.205 -142.965 -52.875 -142.635 ;
        RECT -53.205 -144.325 -52.875 -143.995 ;
        RECT -53.205 -145.685 -52.875 -145.355 ;
        RECT -53.205 -147.045 -52.875 -146.715 ;
        RECT -53.205 -149.765 -52.875 -149.435 ;
        RECT -53.205 -153.845 -52.875 -153.515 ;
        RECT -53.205 -156.565 -52.875 -156.235 ;
        RECT -53.205 -157.925 -52.875 -157.595 ;
        RECT -53.205 -160.17 -52.875 -159.04 ;
        RECT -53.2 -160.285 -52.88 49.125 ;
        RECT -53.205 48.795 -52.875 49.125 ;
        RECT -53.205 47.435 -52.875 47.765 ;
        RECT -53.205 46.075 -52.875 46.405 ;
        RECT -53.205 44.715 -52.875 45.045 ;
        RECT -53.205 43.355 -52.875 43.685 ;
        RECT -53.205 40.635 -52.875 40.965 ;
        RECT -53.205 39.275 -52.875 39.605 ;
        RECT -53.205 35.195 -52.875 35.525 ;
        RECT -53.205 33.835 -52.875 34.165 ;
        RECT -53.205 32.475 -52.875 32.805 ;
        RECT -53.205 31.115 -52.875 31.445 ;
        RECT -53.205 29.755 -52.875 30.085 ;
        RECT -53.205 28.395 -52.875 28.725 ;
        RECT -53.205 27.035 -52.875 27.365 ;
        RECT -53.205 25.675 -52.875 26.005 ;
        RECT -53.205 24.315 -52.875 24.645 ;
        RECT -53.205 22.955 -52.875 23.285 ;
        RECT -53.205 21.595 -52.875 21.925 ;
        RECT -53.205 20.235 -52.875 20.565 ;
        RECT -53.205 18.875 -52.875 19.205 ;
        RECT -53.205 17.515 -52.875 17.845 ;
        RECT -53.205 16.155 -52.875 16.485 ;
        RECT -53.205 14.795 -52.875 15.125 ;
        RECT -53.205 13.435 -52.875 13.765 ;
        RECT -53.205 12.075 -52.875 12.405 ;
        RECT -53.205 10.715 -52.875 11.045 ;
        RECT -53.205 9.355 -52.875 9.685 ;
        RECT -53.205 7.995 -52.875 8.325 ;
        RECT -53.205 6.635 -52.875 6.965 ;
        RECT -53.205 5.275 -52.875 5.605 ;
        RECT -53.205 3.915 -52.875 4.245 ;
        RECT -53.205 2.555 -52.875 2.885 ;
        RECT -53.205 1.195 -52.875 1.525 ;
        RECT -53.205 -0.165 -52.875 0.165 ;
        RECT -53.205 -1.525 -52.875 -1.195 ;
        RECT -53.205 -2.885 -52.875 -2.555 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.445 127.225 -65.115 128.355 ;
        RECT -65.445 124.955 -65.115 125.285 ;
        RECT -65.445 123.595 -65.115 123.925 ;
        RECT -65.445 122.235 -65.115 122.565 ;
        RECT -65.445 120.875 -65.115 121.205 ;
        RECT -65.445 119.515 -65.115 119.845 ;
        RECT -65.445 118.155 -65.115 118.485 ;
        RECT -65.445 116.795 -65.115 117.125 ;
        RECT -65.445 115.435 -65.115 115.765 ;
        RECT -65.445 114.075 -65.115 114.405 ;
        RECT -65.445 112.715 -65.115 113.045 ;
        RECT -65.445 111.355 -65.115 111.685 ;
        RECT -65.445 109.995 -65.115 110.325 ;
        RECT -65.445 108.635 -65.115 108.965 ;
        RECT -65.445 107.275 -65.115 107.605 ;
        RECT -65.445 105.915 -65.115 106.245 ;
        RECT -65.445 104.555 -65.115 104.885 ;
        RECT -65.445 103.195 -65.115 103.525 ;
        RECT -65.445 101.835 -65.115 102.165 ;
        RECT -65.445 100.475 -65.115 100.805 ;
        RECT -65.445 99.115 -65.115 99.445 ;
        RECT -65.445 97.755 -65.115 98.085 ;
        RECT -65.445 96.395 -65.115 96.725 ;
        RECT -65.445 95.035 -65.115 95.365 ;
        RECT -65.445 93.675 -65.115 94.005 ;
        RECT -65.445 92.315 -65.115 92.645 ;
        RECT -65.445 90.955 -65.115 91.285 ;
        RECT -65.445 89.595 -65.115 89.925 ;
        RECT -65.445 88.235 -65.115 88.565 ;
        RECT -65.445 86.875 -65.115 87.205 ;
        RECT -65.445 85.515 -65.115 85.845 ;
        RECT -65.445 84.155 -65.115 84.485 ;
        RECT -65.445 82.795 -65.115 83.125 ;
        RECT -65.445 81.435 -65.115 81.765 ;
        RECT -65.445 80.075 -65.115 80.405 ;
        RECT -65.445 78.715 -65.115 79.045 ;
        RECT -65.445 77.355 -65.115 77.685 ;
        RECT -65.445 75.995 -65.115 76.325 ;
        RECT -65.445 74.635 -65.115 74.965 ;
        RECT -65.445 73.275 -65.115 73.605 ;
        RECT -65.445 71.915 -65.115 72.245 ;
        RECT -65.445 70.555 -65.115 70.885 ;
        RECT -65.445 69.195 -65.115 69.525 ;
        RECT -65.445 67.835 -65.115 68.165 ;
        RECT -65.445 66.475 -65.115 66.805 ;
        RECT -65.445 65.115 -65.115 65.445 ;
        RECT -65.445 63.755 -65.115 64.085 ;
        RECT -65.445 62.395 -65.115 62.725 ;
        RECT -65.445 61.035 -65.115 61.365 ;
        RECT -65.445 59.675 -65.115 60.005 ;
        RECT -65.445 58.315 -65.115 58.645 ;
        RECT -65.445 56.955 -65.115 57.285 ;
        RECT -65.445 55.595 -65.115 55.925 ;
        RECT -65.445 54.235 -65.115 54.565 ;
        RECT -65.445 52.875 -65.115 53.205 ;
        RECT -65.445 51.515 -65.115 51.845 ;
        RECT -65.445 50.155 -65.115 50.485 ;
        RECT -65.445 48.795 -65.115 49.125 ;
        RECT -65.445 47.435 -65.115 47.765 ;
        RECT -65.445 46.075 -65.115 46.405 ;
        RECT -65.445 44.715 -65.115 45.045 ;
        RECT -65.445 43.355 -65.115 43.685 ;
        RECT -65.445 41.995 -65.115 42.325 ;
        RECT -65.445 40.635 -65.115 40.965 ;
        RECT -65.445 39.275 -65.115 39.605 ;
        RECT -65.445 37.915 -65.115 38.245 ;
        RECT -65.445 36.555 -65.115 36.885 ;
        RECT -65.445 35.195 -65.115 35.525 ;
        RECT -65.445 33.835 -65.115 34.165 ;
        RECT -65.445 32.475 -65.115 32.805 ;
        RECT -65.445 31.115 -65.115 31.445 ;
        RECT -65.445 29.755 -65.115 30.085 ;
        RECT -65.445 28.395 -65.115 28.725 ;
        RECT -65.445 27.035 -65.115 27.365 ;
        RECT -65.445 25.675 -65.115 26.005 ;
        RECT -65.445 24.315 -65.115 24.645 ;
        RECT -65.445 22.955 -65.115 23.285 ;
        RECT -65.445 21.595 -65.115 21.925 ;
        RECT -65.445 20.235 -65.115 20.565 ;
        RECT -65.445 18.875 -65.115 19.205 ;
        RECT -65.445 17.515 -65.115 17.845 ;
        RECT -65.445 16.155 -65.115 16.485 ;
        RECT -65.445 14.795 -65.115 15.125 ;
        RECT -65.445 13.435 -65.115 13.765 ;
        RECT -65.445 12.075 -65.115 12.405 ;
        RECT -65.445 10.715 -65.115 11.045 ;
        RECT -65.445 9.355 -65.115 9.685 ;
        RECT -65.445 7.995 -65.115 8.325 ;
        RECT -65.445 6.635 -65.115 6.965 ;
        RECT -65.445 5.275 -65.115 5.605 ;
        RECT -65.445 3.915 -65.115 4.245 ;
        RECT -65.445 2.555 -65.115 2.885 ;
        RECT -65.445 1.195 -65.115 1.525 ;
        RECT -65.445 -0.165 -65.115 0.165 ;
        RECT -65.445 -1.525 -65.115 -1.195 ;
        RECT -65.445 -2.885 -65.115 -2.555 ;
        RECT -65.445 -4.245 -65.115 -3.915 ;
        RECT -65.445 -5.605 -65.115 -5.275 ;
        RECT -65.445 -6.965 -65.115 -6.635 ;
        RECT -65.445 -8.325 -65.115 -7.995 ;
        RECT -65.445 -9.685 -65.115 -9.355 ;
        RECT -65.445 -11.045 -65.115 -10.715 ;
        RECT -65.445 -12.405 -65.115 -12.075 ;
        RECT -65.445 -13.765 -65.115 -13.435 ;
        RECT -65.445 -15.125 -65.115 -14.795 ;
        RECT -65.445 -16.485 -65.115 -16.155 ;
        RECT -65.445 -17.845 -65.115 -17.515 ;
        RECT -65.445 -19.205 -65.115 -18.875 ;
        RECT -65.445 -20.565 -65.115 -20.235 ;
        RECT -65.445 -21.925 -65.115 -21.595 ;
        RECT -65.445 -23.285 -65.115 -22.955 ;
        RECT -65.445 -24.645 -65.115 -24.315 ;
        RECT -65.445 -26.005 -65.115 -25.675 ;
        RECT -65.445 -27.365 -65.115 -27.035 ;
        RECT -65.445 -28.725 -65.115 -28.395 ;
        RECT -65.445 -30.085 -65.115 -29.755 ;
        RECT -65.445 -31.445 -65.115 -31.115 ;
        RECT -65.445 -32.805 -65.115 -32.475 ;
        RECT -65.445 -34.165 -65.115 -33.835 ;
        RECT -65.445 -35.525 -65.115 -35.195 ;
        RECT -65.445 -36.885 -65.115 -36.555 ;
        RECT -65.445 -38.245 -65.115 -37.915 ;
        RECT -65.445 -39.605 -65.115 -39.275 ;
        RECT -65.445 -40.965 -65.115 -40.635 ;
        RECT -65.445 -42.325 -65.115 -41.995 ;
        RECT -65.445 -43.685 -65.115 -43.355 ;
        RECT -65.445 -45.045 -65.115 -44.715 ;
        RECT -65.445 -46.405 -65.115 -46.075 ;
        RECT -65.445 -47.765 -65.115 -47.435 ;
        RECT -65.445 -49.125 -65.115 -48.795 ;
        RECT -65.445 -50.485 -65.115 -50.155 ;
        RECT -65.445 -51.845 -65.115 -51.515 ;
        RECT -65.445 -53.205 -65.115 -52.875 ;
        RECT -65.445 -54.565 -65.115 -54.235 ;
        RECT -65.445 -55.925 -65.115 -55.595 ;
        RECT -65.445 -57.285 -65.115 -56.955 ;
        RECT -65.445 -58.645 -65.115 -58.315 ;
        RECT -65.445 -60.005 -65.115 -59.675 ;
        RECT -65.445 -61.365 -65.115 -61.035 ;
        RECT -65.445 -62.725 -65.115 -62.395 ;
        RECT -65.445 -64.085 -65.115 -63.755 ;
        RECT -65.445 -65.445 -65.115 -65.115 ;
        RECT -65.445 -66.805 -65.115 -66.475 ;
        RECT -65.445 -68.165 -65.115 -67.835 ;
        RECT -65.445 -69.525 -65.115 -69.195 ;
        RECT -65.445 -70.885 -65.115 -70.555 ;
        RECT -65.445 -72.245 -65.115 -71.915 ;
        RECT -65.445 -73.605 -65.115 -73.275 ;
        RECT -65.445 -74.965 -65.115 -74.635 ;
        RECT -65.445 -76.325 -65.115 -75.995 ;
        RECT -65.445 -77.685 -65.115 -77.355 ;
        RECT -65.445 -79.045 -65.115 -78.715 ;
        RECT -65.445 -80.405 -65.115 -80.075 ;
        RECT -65.445 -81.765 -65.115 -81.435 ;
        RECT -65.445 -83.125 -65.115 -82.795 ;
        RECT -65.445 -84.485 -65.115 -84.155 ;
        RECT -65.445 -85.845 -65.115 -85.515 ;
        RECT -65.445 -87.205 -65.115 -86.875 ;
        RECT -65.445 -88.565 -65.115 -88.235 ;
        RECT -65.445 -89.925 -65.115 -89.595 ;
        RECT -65.445 -91.285 -65.115 -90.955 ;
        RECT -65.445 -92.645 -65.115 -92.315 ;
        RECT -65.445 -94.005 -65.115 -93.675 ;
        RECT -65.445 -95.365 -65.115 -95.035 ;
        RECT -65.445 -96.725 -65.115 -96.395 ;
        RECT -65.445 -98.085 -65.115 -97.755 ;
        RECT -65.445 -99.445 -65.115 -99.115 ;
        RECT -65.445 -100.805 -65.115 -100.475 ;
        RECT -65.445 -102.165 -65.115 -101.835 ;
        RECT -65.445 -103.525 -65.115 -103.195 ;
        RECT -65.445 -104.885 -65.115 -104.555 ;
        RECT -65.445 -106.245 -65.115 -105.915 ;
        RECT -65.445 -107.605 -65.115 -107.275 ;
        RECT -65.445 -108.965 -65.115 -108.635 ;
        RECT -65.445 -110.325 -65.115 -109.995 ;
        RECT -65.445 -111.685 -65.115 -111.355 ;
        RECT -65.445 -113.045 -65.115 -112.715 ;
        RECT -65.445 -114.405 -65.115 -114.075 ;
        RECT -65.445 -115.765 -65.115 -115.435 ;
        RECT -65.445 -117.125 -65.115 -116.795 ;
        RECT -65.445 -118.485 -65.115 -118.155 ;
        RECT -65.445 -119.845 -65.115 -119.515 ;
        RECT -65.445 -121.205 -65.115 -120.875 ;
        RECT -65.445 -122.565 -65.115 -122.235 ;
        RECT -65.445 -123.925 -65.115 -123.595 ;
        RECT -65.445 -125.285 -65.115 -124.955 ;
        RECT -65.445 -126.645 -65.115 -126.315 ;
        RECT -65.445 -128.005 -65.115 -127.675 ;
        RECT -65.445 -129.365 -65.115 -129.035 ;
        RECT -65.445 -130.725 -65.115 -130.395 ;
        RECT -65.445 -132.085 -65.115 -131.755 ;
        RECT -65.445 -133.445 -65.115 -133.115 ;
        RECT -65.445 -134.805 -65.115 -134.475 ;
        RECT -65.445 -136.165 -65.115 -135.835 ;
        RECT -65.445 -137.525 -65.115 -137.195 ;
        RECT -65.445 -138.885 -65.115 -138.555 ;
        RECT -65.445 -140.245 -65.115 -139.915 ;
        RECT -65.445 -141.605 -65.115 -141.275 ;
        RECT -65.445 -142.965 -65.115 -142.635 ;
        RECT -65.445 -144.325 -65.115 -143.995 ;
        RECT -65.445 -145.685 -65.115 -145.355 ;
        RECT -65.445 -147.045 -65.115 -146.715 ;
        RECT -65.445 -149.765 -65.115 -149.435 ;
        RECT -65.445 -151.125 -65.115 -150.795 ;
        RECT -65.445 -152.485 -65.115 -152.155 ;
        RECT -65.445 -153.845 -65.115 -153.515 ;
        RECT -65.445 -156.565 -65.115 -156.235 ;
        RECT -65.445 -157.925 -65.115 -157.595 ;
        RECT -65.445 -160.17 -65.115 -159.04 ;
        RECT -65.44 -160.285 -65.12 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.085 127.225 -63.755 128.355 ;
        RECT -64.085 124.955 -63.755 125.285 ;
        RECT -64.085 123.595 -63.755 123.925 ;
        RECT -64.085 122.235 -63.755 122.565 ;
        RECT -64.085 120.875 -63.755 121.205 ;
        RECT -64.085 119.515 -63.755 119.845 ;
        RECT -64.085 118.155 -63.755 118.485 ;
        RECT -64.085 116.795 -63.755 117.125 ;
        RECT -64.085 115.435 -63.755 115.765 ;
        RECT -64.085 114.075 -63.755 114.405 ;
        RECT -64.085 112.715 -63.755 113.045 ;
        RECT -64.085 111.355 -63.755 111.685 ;
        RECT -64.085 109.995 -63.755 110.325 ;
        RECT -64.085 108.635 -63.755 108.965 ;
        RECT -64.085 107.275 -63.755 107.605 ;
        RECT -64.085 105.915 -63.755 106.245 ;
        RECT -64.085 104.555 -63.755 104.885 ;
        RECT -64.085 103.195 -63.755 103.525 ;
        RECT -64.085 101.835 -63.755 102.165 ;
        RECT -64.085 100.475 -63.755 100.805 ;
        RECT -64.085 99.115 -63.755 99.445 ;
        RECT -64.085 97.755 -63.755 98.085 ;
        RECT -64.085 96.395 -63.755 96.725 ;
        RECT -64.085 95.035 -63.755 95.365 ;
        RECT -64.085 93.675 -63.755 94.005 ;
        RECT -64.085 92.315 -63.755 92.645 ;
        RECT -64.085 90.955 -63.755 91.285 ;
        RECT -64.085 89.595 -63.755 89.925 ;
        RECT -64.085 88.235 -63.755 88.565 ;
        RECT -64.085 86.875 -63.755 87.205 ;
        RECT -64.085 85.515 -63.755 85.845 ;
        RECT -64.085 84.155 -63.755 84.485 ;
        RECT -64.085 82.795 -63.755 83.125 ;
        RECT -64.085 81.435 -63.755 81.765 ;
        RECT -64.085 80.075 -63.755 80.405 ;
        RECT -64.085 78.715 -63.755 79.045 ;
        RECT -64.085 77.355 -63.755 77.685 ;
        RECT -64.085 75.995 -63.755 76.325 ;
        RECT -64.085 74.635 -63.755 74.965 ;
        RECT -64.085 73.275 -63.755 73.605 ;
        RECT -64.085 71.915 -63.755 72.245 ;
        RECT -64.085 70.555 -63.755 70.885 ;
        RECT -64.085 69.195 -63.755 69.525 ;
        RECT -64.085 67.835 -63.755 68.165 ;
        RECT -64.085 66.475 -63.755 66.805 ;
        RECT -64.085 65.115 -63.755 65.445 ;
        RECT -64.085 63.755 -63.755 64.085 ;
        RECT -64.085 62.395 -63.755 62.725 ;
        RECT -64.085 61.035 -63.755 61.365 ;
        RECT -64.085 59.675 -63.755 60.005 ;
        RECT -64.085 58.315 -63.755 58.645 ;
        RECT -64.085 56.955 -63.755 57.285 ;
        RECT -64.085 55.595 -63.755 55.925 ;
        RECT -64.085 54.235 -63.755 54.565 ;
        RECT -64.085 52.875 -63.755 53.205 ;
        RECT -64.085 51.515 -63.755 51.845 ;
        RECT -64.085 50.155 -63.755 50.485 ;
        RECT -64.085 48.795 -63.755 49.125 ;
        RECT -64.085 47.435 -63.755 47.765 ;
        RECT -64.085 46.075 -63.755 46.405 ;
        RECT -64.085 44.715 -63.755 45.045 ;
        RECT -64.085 43.355 -63.755 43.685 ;
        RECT -64.085 41.995 -63.755 42.325 ;
        RECT -64.085 40.635 -63.755 40.965 ;
        RECT -64.085 39.275 -63.755 39.605 ;
        RECT -64.085 37.915 -63.755 38.245 ;
        RECT -64.085 36.555 -63.755 36.885 ;
        RECT -64.085 35.195 -63.755 35.525 ;
        RECT -64.085 33.835 -63.755 34.165 ;
        RECT -64.085 32.475 -63.755 32.805 ;
        RECT -64.085 31.115 -63.755 31.445 ;
        RECT -64.085 29.755 -63.755 30.085 ;
        RECT -64.085 28.395 -63.755 28.725 ;
        RECT -64.085 27.035 -63.755 27.365 ;
        RECT -64.085 25.675 -63.755 26.005 ;
        RECT -64.085 24.315 -63.755 24.645 ;
        RECT -64.085 22.955 -63.755 23.285 ;
        RECT -64.085 21.595 -63.755 21.925 ;
        RECT -64.085 20.235 -63.755 20.565 ;
        RECT -64.085 18.875 -63.755 19.205 ;
        RECT -64.085 17.515 -63.755 17.845 ;
        RECT -64.085 16.155 -63.755 16.485 ;
        RECT -64.085 14.795 -63.755 15.125 ;
        RECT -64.085 13.435 -63.755 13.765 ;
        RECT -64.085 12.075 -63.755 12.405 ;
        RECT -64.085 10.715 -63.755 11.045 ;
        RECT -64.085 9.355 -63.755 9.685 ;
        RECT -64.085 7.995 -63.755 8.325 ;
        RECT -64.085 6.635 -63.755 6.965 ;
        RECT -64.085 5.275 -63.755 5.605 ;
        RECT -64.085 3.915 -63.755 4.245 ;
        RECT -64.085 2.555 -63.755 2.885 ;
        RECT -64.085 1.195 -63.755 1.525 ;
        RECT -64.085 -0.165 -63.755 0.165 ;
        RECT -64.085 -1.525 -63.755 -1.195 ;
        RECT -64.085 -2.885 -63.755 -2.555 ;
        RECT -64.085 -4.245 -63.755 -3.915 ;
        RECT -64.085 -5.605 -63.755 -5.275 ;
        RECT -64.085 -6.965 -63.755 -6.635 ;
        RECT -64.085 -8.325 -63.755 -7.995 ;
        RECT -64.085 -9.685 -63.755 -9.355 ;
        RECT -64.085 -11.045 -63.755 -10.715 ;
        RECT -64.085 -12.405 -63.755 -12.075 ;
        RECT -64.085 -13.765 -63.755 -13.435 ;
        RECT -64.085 -15.125 -63.755 -14.795 ;
        RECT -64.085 -16.485 -63.755 -16.155 ;
        RECT -64.085 -17.845 -63.755 -17.515 ;
        RECT -64.085 -19.205 -63.755 -18.875 ;
        RECT -64.085 -20.565 -63.755 -20.235 ;
        RECT -64.085 -21.925 -63.755 -21.595 ;
        RECT -64.085 -23.285 -63.755 -22.955 ;
        RECT -64.085 -24.645 -63.755 -24.315 ;
        RECT -64.085 -26.005 -63.755 -25.675 ;
        RECT -64.085 -27.365 -63.755 -27.035 ;
        RECT -64.085 -28.725 -63.755 -28.395 ;
        RECT -64.085 -30.085 -63.755 -29.755 ;
        RECT -64.085 -31.445 -63.755 -31.115 ;
        RECT -64.085 -32.805 -63.755 -32.475 ;
        RECT -64.085 -34.165 -63.755 -33.835 ;
        RECT -64.085 -35.525 -63.755 -35.195 ;
        RECT -64.085 -36.885 -63.755 -36.555 ;
        RECT -64.085 -38.245 -63.755 -37.915 ;
        RECT -64.085 -39.605 -63.755 -39.275 ;
        RECT -64.085 -40.965 -63.755 -40.635 ;
        RECT -64.085 -42.325 -63.755 -41.995 ;
        RECT -64.085 -43.685 -63.755 -43.355 ;
        RECT -64.085 -45.045 -63.755 -44.715 ;
        RECT -64.085 -46.405 -63.755 -46.075 ;
        RECT -64.085 -47.765 -63.755 -47.435 ;
        RECT -64.085 -49.125 -63.755 -48.795 ;
        RECT -64.085 -50.485 -63.755 -50.155 ;
        RECT -64.085 -51.845 -63.755 -51.515 ;
        RECT -64.085 -53.205 -63.755 -52.875 ;
        RECT -64.085 -54.565 -63.755 -54.235 ;
        RECT -64.085 -55.925 -63.755 -55.595 ;
        RECT -64.085 -57.285 -63.755 -56.955 ;
        RECT -64.085 -58.645 -63.755 -58.315 ;
        RECT -64.085 -60.005 -63.755 -59.675 ;
        RECT -64.085 -61.365 -63.755 -61.035 ;
        RECT -64.085 -62.725 -63.755 -62.395 ;
        RECT -64.085 -64.085 -63.755 -63.755 ;
        RECT -64.085 -65.445 -63.755 -65.115 ;
        RECT -64.085 -66.805 -63.755 -66.475 ;
        RECT -64.085 -68.165 -63.755 -67.835 ;
        RECT -64.085 -69.525 -63.755 -69.195 ;
        RECT -64.085 -70.885 -63.755 -70.555 ;
        RECT -64.085 -72.245 -63.755 -71.915 ;
        RECT -64.085 -73.605 -63.755 -73.275 ;
        RECT -64.085 -74.965 -63.755 -74.635 ;
        RECT -64.085 -76.325 -63.755 -75.995 ;
        RECT -64.085 -77.685 -63.755 -77.355 ;
        RECT -64.085 -79.045 -63.755 -78.715 ;
        RECT -64.085 -80.405 -63.755 -80.075 ;
        RECT -64.085 -81.765 -63.755 -81.435 ;
        RECT -64.085 -83.125 -63.755 -82.795 ;
        RECT -64.085 -84.485 -63.755 -84.155 ;
        RECT -64.085 -85.845 -63.755 -85.515 ;
        RECT -64.085 -87.205 -63.755 -86.875 ;
        RECT -64.085 -88.565 -63.755 -88.235 ;
        RECT -64.085 -89.925 -63.755 -89.595 ;
        RECT -64.085 -91.285 -63.755 -90.955 ;
        RECT -64.085 -92.645 -63.755 -92.315 ;
        RECT -64.085 -94.005 -63.755 -93.675 ;
        RECT -64.085 -95.365 -63.755 -95.035 ;
        RECT -64.085 -96.725 -63.755 -96.395 ;
        RECT -64.085 -98.085 -63.755 -97.755 ;
        RECT -64.085 -99.445 -63.755 -99.115 ;
        RECT -64.085 -100.805 -63.755 -100.475 ;
        RECT -64.085 -102.165 -63.755 -101.835 ;
        RECT -64.085 -103.525 -63.755 -103.195 ;
        RECT -64.085 -104.885 -63.755 -104.555 ;
        RECT -64.085 -106.245 -63.755 -105.915 ;
        RECT -64.085 -107.605 -63.755 -107.275 ;
        RECT -64.085 -108.965 -63.755 -108.635 ;
        RECT -64.085 -110.325 -63.755 -109.995 ;
        RECT -64.085 -111.685 -63.755 -111.355 ;
        RECT -64.085 -113.045 -63.755 -112.715 ;
        RECT -64.085 -114.405 -63.755 -114.075 ;
        RECT -64.085 -115.765 -63.755 -115.435 ;
        RECT -64.085 -117.125 -63.755 -116.795 ;
        RECT -64.085 -118.485 -63.755 -118.155 ;
        RECT -64.085 -119.845 -63.755 -119.515 ;
        RECT -64.085 -121.205 -63.755 -120.875 ;
        RECT -64.085 -122.565 -63.755 -122.235 ;
        RECT -64.085 -123.925 -63.755 -123.595 ;
        RECT -64.085 -125.285 -63.755 -124.955 ;
        RECT -64.085 -126.645 -63.755 -126.315 ;
        RECT -64.085 -128.005 -63.755 -127.675 ;
        RECT -64.085 -129.365 -63.755 -129.035 ;
        RECT -64.085 -130.725 -63.755 -130.395 ;
        RECT -64.085 -132.085 -63.755 -131.755 ;
        RECT -64.085 -133.445 -63.755 -133.115 ;
        RECT -64.085 -134.805 -63.755 -134.475 ;
        RECT -64.085 -136.165 -63.755 -135.835 ;
        RECT -64.085 -137.525 -63.755 -137.195 ;
        RECT -64.085 -138.885 -63.755 -138.555 ;
        RECT -64.085 -140.245 -63.755 -139.915 ;
        RECT -64.085 -141.605 -63.755 -141.275 ;
        RECT -64.085 -142.965 -63.755 -142.635 ;
        RECT -64.085 -144.325 -63.755 -143.995 ;
        RECT -64.085 -145.685 -63.755 -145.355 ;
        RECT -64.085 -147.045 -63.755 -146.715 ;
        RECT -64.085 -149.765 -63.755 -149.435 ;
        RECT -64.085 -153.845 -63.755 -153.515 ;
        RECT -64.085 -155.285 -63.755 -154.955 ;
        RECT -64.085 -156.565 -63.755 -156.235 ;
        RECT -64.085 -157.925 -63.755 -157.595 ;
        RECT -64.085 -160.17 -63.755 -159.04 ;
        RECT -64.08 -160.285 -63.76 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.725 127.225 -62.395 128.355 ;
        RECT -62.725 124.955 -62.395 125.285 ;
        RECT -62.725 123.595 -62.395 123.925 ;
        RECT -62.725 122.235 -62.395 122.565 ;
        RECT -62.725 120.875 -62.395 121.205 ;
        RECT -62.725 119.515 -62.395 119.845 ;
        RECT -62.725 118.155 -62.395 118.485 ;
        RECT -62.725 116.795 -62.395 117.125 ;
        RECT -62.725 115.435 -62.395 115.765 ;
        RECT -62.725 114.075 -62.395 114.405 ;
        RECT -62.725 112.715 -62.395 113.045 ;
        RECT -62.725 111.355 -62.395 111.685 ;
        RECT -62.725 109.995 -62.395 110.325 ;
        RECT -62.725 108.635 -62.395 108.965 ;
        RECT -62.725 107.275 -62.395 107.605 ;
        RECT -62.725 105.915 -62.395 106.245 ;
        RECT -62.725 104.555 -62.395 104.885 ;
        RECT -62.725 103.195 -62.395 103.525 ;
        RECT -62.725 101.835 -62.395 102.165 ;
        RECT -62.725 100.475 -62.395 100.805 ;
        RECT -62.725 99.115 -62.395 99.445 ;
        RECT -62.725 97.755 -62.395 98.085 ;
        RECT -62.725 96.395 -62.395 96.725 ;
        RECT -62.725 95.035 -62.395 95.365 ;
        RECT -62.725 93.675 -62.395 94.005 ;
        RECT -62.725 92.315 -62.395 92.645 ;
        RECT -62.725 90.955 -62.395 91.285 ;
        RECT -62.725 89.595 -62.395 89.925 ;
        RECT -62.725 88.235 -62.395 88.565 ;
        RECT -62.725 86.875 -62.395 87.205 ;
        RECT -62.725 85.515 -62.395 85.845 ;
        RECT -62.725 84.155 -62.395 84.485 ;
        RECT -62.725 82.795 -62.395 83.125 ;
        RECT -62.725 81.435 -62.395 81.765 ;
        RECT -62.725 80.075 -62.395 80.405 ;
        RECT -62.725 78.715 -62.395 79.045 ;
        RECT -62.725 77.355 -62.395 77.685 ;
        RECT -62.725 75.995 -62.395 76.325 ;
        RECT -62.725 74.635 -62.395 74.965 ;
        RECT -62.725 73.275 -62.395 73.605 ;
        RECT -62.725 71.915 -62.395 72.245 ;
        RECT -62.725 70.555 -62.395 70.885 ;
        RECT -62.725 69.195 -62.395 69.525 ;
        RECT -62.725 67.835 -62.395 68.165 ;
        RECT -62.725 66.475 -62.395 66.805 ;
        RECT -62.725 65.115 -62.395 65.445 ;
        RECT -62.725 63.755 -62.395 64.085 ;
        RECT -62.725 62.395 -62.395 62.725 ;
        RECT -62.725 61.035 -62.395 61.365 ;
        RECT -62.725 59.675 -62.395 60.005 ;
        RECT -62.725 58.315 -62.395 58.645 ;
        RECT -62.725 56.955 -62.395 57.285 ;
        RECT -62.725 55.595 -62.395 55.925 ;
        RECT -62.725 54.235 -62.395 54.565 ;
        RECT -62.725 52.875 -62.395 53.205 ;
        RECT -62.725 51.515 -62.395 51.845 ;
        RECT -62.725 50.155 -62.395 50.485 ;
        RECT -62.725 48.795 -62.395 49.125 ;
        RECT -62.725 47.435 -62.395 47.765 ;
        RECT -62.725 46.075 -62.395 46.405 ;
        RECT -62.725 44.715 -62.395 45.045 ;
        RECT -62.725 43.355 -62.395 43.685 ;
        RECT -62.725 41.995 -62.395 42.325 ;
        RECT -62.725 40.635 -62.395 40.965 ;
        RECT -62.725 39.275 -62.395 39.605 ;
        RECT -62.725 37.915 -62.395 38.245 ;
        RECT -62.725 36.555 -62.395 36.885 ;
        RECT -62.725 35.195 -62.395 35.525 ;
        RECT -62.725 33.835 -62.395 34.165 ;
        RECT -62.725 32.475 -62.395 32.805 ;
        RECT -62.725 31.115 -62.395 31.445 ;
        RECT -62.725 29.755 -62.395 30.085 ;
        RECT -62.725 28.395 -62.395 28.725 ;
        RECT -62.725 27.035 -62.395 27.365 ;
        RECT -62.725 25.675 -62.395 26.005 ;
        RECT -62.725 24.315 -62.395 24.645 ;
        RECT -62.725 22.955 -62.395 23.285 ;
        RECT -62.725 21.595 -62.395 21.925 ;
        RECT -62.725 20.235 -62.395 20.565 ;
        RECT -62.725 18.875 -62.395 19.205 ;
        RECT -62.725 17.515 -62.395 17.845 ;
        RECT -62.725 16.155 -62.395 16.485 ;
        RECT -62.725 14.795 -62.395 15.125 ;
        RECT -62.725 13.435 -62.395 13.765 ;
        RECT -62.725 12.075 -62.395 12.405 ;
        RECT -62.725 10.715 -62.395 11.045 ;
        RECT -62.725 9.355 -62.395 9.685 ;
        RECT -62.725 7.995 -62.395 8.325 ;
        RECT -62.725 6.635 -62.395 6.965 ;
        RECT -62.725 5.275 -62.395 5.605 ;
        RECT -62.725 3.915 -62.395 4.245 ;
        RECT -62.725 2.555 -62.395 2.885 ;
        RECT -62.725 1.195 -62.395 1.525 ;
        RECT -62.725 -0.165 -62.395 0.165 ;
        RECT -62.725 -1.525 -62.395 -1.195 ;
        RECT -62.725 -2.885 -62.395 -2.555 ;
        RECT -62.725 -4.245 -62.395 -3.915 ;
        RECT -62.725 -5.605 -62.395 -5.275 ;
        RECT -62.725 -6.965 -62.395 -6.635 ;
        RECT -62.725 -8.325 -62.395 -7.995 ;
        RECT -62.725 -9.685 -62.395 -9.355 ;
        RECT -62.725 -11.045 -62.395 -10.715 ;
        RECT -62.725 -12.405 -62.395 -12.075 ;
        RECT -62.725 -13.765 -62.395 -13.435 ;
        RECT -62.725 -15.125 -62.395 -14.795 ;
        RECT -62.725 -16.485 -62.395 -16.155 ;
        RECT -62.725 -17.845 -62.395 -17.515 ;
        RECT -62.725 -19.205 -62.395 -18.875 ;
        RECT -62.725 -20.565 -62.395 -20.235 ;
        RECT -62.725 -21.925 -62.395 -21.595 ;
        RECT -62.725 -23.285 -62.395 -22.955 ;
        RECT -62.725 -24.645 -62.395 -24.315 ;
        RECT -62.725 -26.005 -62.395 -25.675 ;
        RECT -62.725 -27.365 -62.395 -27.035 ;
        RECT -62.725 -28.725 -62.395 -28.395 ;
        RECT -62.725 -30.085 -62.395 -29.755 ;
        RECT -62.725 -31.445 -62.395 -31.115 ;
        RECT -62.725 -32.805 -62.395 -32.475 ;
        RECT -62.725 -34.165 -62.395 -33.835 ;
        RECT -62.725 -35.525 -62.395 -35.195 ;
        RECT -62.725 -36.885 -62.395 -36.555 ;
        RECT -62.725 -38.245 -62.395 -37.915 ;
        RECT -62.725 -39.605 -62.395 -39.275 ;
        RECT -62.725 -40.965 -62.395 -40.635 ;
        RECT -62.725 -42.325 -62.395 -41.995 ;
        RECT -62.725 -43.685 -62.395 -43.355 ;
        RECT -62.725 -45.045 -62.395 -44.715 ;
        RECT -62.725 -46.405 -62.395 -46.075 ;
        RECT -62.725 -47.765 -62.395 -47.435 ;
        RECT -62.725 -49.125 -62.395 -48.795 ;
        RECT -62.725 -50.485 -62.395 -50.155 ;
        RECT -62.725 -51.845 -62.395 -51.515 ;
        RECT -62.725 -53.205 -62.395 -52.875 ;
        RECT -62.725 -54.565 -62.395 -54.235 ;
        RECT -62.725 -55.925 -62.395 -55.595 ;
        RECT -62.725 -57.285 -62.395 -56.955 ;
        RECT -62.725 -58.645 -62.395 -58.315 ;
        RECT -62.725 -60.005 -62.395 -59.675 ;
        RECT -62.725 -61.365 -62.395 -61.035 ;
        RECT -62.725 -62.725 -62.395 -62.395 ;
        RECT -62.725 -64.085 -62.395 -63.755 ;
        RECT -62.725 -65.445 -62.395 -65.115 ;
        RECT -62.725 -66.805 -62.395 -66.475 ;
        RECT -62.725 -68.165 -62.395 -67.835 ;
        RECT -62.725 -69.525 -62.395 -69.195 ;
        RECT -62.725 -70.885 -62.395 -70.555 ;
        RECT -62.725 -72.245 -62.395 -71.915 ;
        RECT -62.725 -73.605 -62.395 -73.275 ;
        RECT -62.725 -74.965 -62.395 -74.635 ;
        RECT -62.725 -76.325 -62.395 -75.995 ;
        RECT -62.725 -77.685 -62.395 -77.355 ;
        RECT -62.725 -79.045 -62.395 -78.715 ;
        RECT -62.725 -80.405 -62.395 -80.075 ;
        RECT -62.725 -81.765 -62.395 -81.435 ;
        RECT -62.725 -83.125 -62.395 -82.795 ;
        RECT -62.725 -84.485 -62.395 -84.155 ;
        RECT -62.725 -85.845 -62.395 -85.515 ;
        RECT -62.725 -87.205 -62.395 -86.875 ;
        RECT -62.725 -88.565 -62.395 -88.235 ;
        RECT -62.725 -89.925 -62.395 -89.595 ;
        RECT -62.725 -91.285 -62.395 -90.955 ;
        RECT -62.725 -92.645 -62.395 -92.315 ;
        RECT -62.725 -94.005 -62.395 -93.675 ;
        RECT -62.725 -95.365 -62.395 -95.035 ;
        RECT -62.725 -96.725 -62.395 -96.395 ;
        RECT -62.725 -98.085 -62.395 -97.755 ;
        RECT -62.725 -99.445 -62.395 -99.115 ;
        RECT -62.725 -100.805 -62.395 -100.475 ;
        RECT -62.725 -102.165 -62.395 -101.835 ;
        RECT -62.725 -103.525 -62.395 -103.195 ;
        RECT -62.725 -104.885 -62.395 -104.555 ;
        RECT -62.725 -106.245 -62.395 -105.915 ;
        RECT -62.725 -107.605 -62.395 -107.275 ;
        RECT -62.725 -108.965 -62.395 -108.635 ;
        RECT -62.725 -110.325 -62.395 -109.995 ;
        RECT -62.725 -111.685 -62.395 -111.355 ;
        RECT -62.725 -113.045 -62.395 -112.715 ;
        RECT -62.725 -114.405 -62.395 -114.075 ;
        RECT -62.725 -115.765 -62.395 -115.435 ;
        RECT -62.725 -117.125 -62.395 -116.795 ;
        RECT -62.725 -118.485 -62.395 -118.155 ;
        RECT -62.725 -119.845 -62.395 -119.515 ;
        RECT -62.725 -121.205 -62.395 -120.875 ;
        RECT -62.725 -122.565 -62.395 -122.235 ;
        RECT -62.725 -123.925 -62.395 -123.595 ;
        RECT -62.725 -125.285 -62.395 -124.955 ;
        RECT -62.725 -126.645 -62.395 -126.315 ;
        RECT -62.725 -128.005 -62.395 -127.675 ;
        RECT -62.725 -129.365 -62.395 -129.035 ;
        RECT -62.725 -130.725 -62.395 -130.395 ;
        RECT -62.725 -132.085 -62.395 -131.755 ;
        RECT -62.725 -133.445 -62.395 -133.115 ;
        RECT -62.725 -134.805 -62.395 -134.475 ;
        RECT -62.725 -136.165 -62.395 -135.835 ;
        RECT -62.725 -137.525 -62.395 -137.195 ;
        RECT -62.725 -138.885 -62.395 -138.555 ;
        RECT -62.725 -140.245 -62.395 -139.915 ;
        RECT -62.725 -141.605 -62.395 -141.275 ;
        RECT -62.725 -142.965 -62.395 -142.635 ;
        RECT -62.725 -144.325 -62.395 -143.995 ;
        RECT -62.725 -145.685 -62.395 -145.355 ;
        RECT -62.725 -147.045 -62.395 -146.715 ;
        RECT -62.725 -149.765 -62.395 -149.435 ;
        RECT -62.725 -152.485 -62.395 -152.155 ;
        RECT -62.725 -153.845 -62.395 -153.515 ;
        RECT -62.725 -155.285 -62.395 -154.955 ;
        RECT -62.725 -156.565 -62.395 -156.235 ;
        RECT -62.725 -157.925 -62.395 -157.595 ;
        RECT -62.725 -160.17 -62.395 -159.04 ;
        RECT -62.72 -160.285 -62.4 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.365 127.225 -61.035 128.355 ;
        RECT -61.365 124.955 -61.035 125.285 ;
        RECT -61.365 123.595 -61.035 123.925 ;
        RECT -61.365 122.235 -61.035 122.565 ;
        RECT -61.365 120.875 -61.035 121.205 ;
        RECT -61.365 119.515 -61.035 119.845 ;
        RECT -61.365 118.155 -61.035 118.485 ;
        RECT -61.365 116.795 -61.035 117.125 ;
        RECT -61.365 115.435 -61.035 115.765 ;
        RECT -61.365 114.075 -61.035 114.405 ;
        RECT -61.365 112.715 -61.035 113.045 ;
        RECT -61.365 111.355 -61.035 111.685 ;
        RECT -61.365 109.995 -61.035 110.325 ;
        RECT -61.365 108.635 -61.035 108.965 ;
        RECT -61.365 107.275 -61.035 107.605 ;
        RECT -61.365 105.915 -61.035 106.245 ;
        RECT -61.365 104.555 -61.035 104.885 ;
        RECT -61.365 103.195 -61.035 103.525 ;
        RECT -61.365 101.835 -61.035 102.165 ;
        RECT -61.365 100.475 -61.035 100.805 ;
        RECT -61.365 99.115 -61.035 99.445 ;
        RECT -61.365 97.755 -61.035 98.085 ;
        RECT -61.365 96.395 -61.035 96.725 ;
        RECT -61.365 95.035 -61.035 95.365 ;
        RECT -61.365 93.675 -61.035 94.005 ;
        RECT -61.365 92.315 -61.035 92.645 ;
        RECT -61.365 90.955 -61.035 91.285 ;
        RECT -61.365 89.595 -61.035 89.925 ;
        RECT -61.365 88.235 -61.035 88.565 ;
        RECT -61.365 86.875 -61.035 87.205 ;
        RECT -61.365 85.515 -61.035 85.845 ;
        RECT -61.365 84.155 -61.035 84.485 ;
        RECT -61.365 82.795 -61.035 83.125 ;
        RECT -61.365 81.435 -61.035 81.765 ;
        RECT -61.365 80.075 -61.035 80.405 ;
        RECT -61.365 78.715 -61.035 79.045 ;
        RECT -61.365 77.355 -61.035 77.685 ;
        RECT -61.365 75.995 -61.035 76.325 ;
        RECT -61.365 74.635 -61.035 74.965 ;
        RECT -61.365 73.275 -61.035 73.605 ;
        RECT -61.365 71.915 -61.035 72.245 ;
        RECT -61.365 70.555 -61.035 70.885 ;
        RECT -61.365 69.195 -61.035 69.525 ;
        RECT -61.365 67.835 -61.035 68.165 ;
        RECT -61.365 66.475 -61.035 66.805 ;
        RECT -61.365 65.115 -61.035 65.445 ;
        RECT -61.365 63.755 -61.035 64.085 ;
        RECT -61.365 62.395 -61.035 62.725 ;
        RECT -61.365 61.035 -61.035 61.365 ;
        RECT -61.365 59.675 -61.035 60.005 ;
        RECT -61.365 58.315 -61.035 58.645 ;
        RECT -61.365 56.955 -61.035 57.285 ;
        RECT -61.365 55.595 -61.035 55.925 ;
        RECT -61.365 54.235 -61.035 54.565 ;
        RECT -61.365 52.875 -61.035 53.205 ;
        RECT -61.365 51.515 -61.035 51.845 ;
        RECT -61.365 50.155 -61.035 50.485 ;
        RECT -61.365 48.795 -61.035 49.125 ;
        RECT -61.365 47.435 -61.035 47.765 ;
        RECT -61.365 46.075 -61.035 46.405 ;
        RECT -61.365 44.715 -61.035 45.045 ;
        RECT -61.365 43.355 -61.035 43.685 ;
        RECT -61.365 41.995 -61.035 42.325 ;
        RECT -61.365 40.635 -61.035 40.965 ;
        RECT -61.365 39.275 -61.035 39.605 ;
        RECT -61.365 37.915 -61.035 38.245 ;
        RECT -61.365 36.555 -61.035 36.885 ;
        RECT -61.365 35.195 -61.035 35.525 ;
        RECT -61.365 33.835 -61.035 34.165 ;
        RECT -61.365 32.475 -61.035 32.805 ;
        RECT -61.365 31.115 -61.035 31.445 ;
        RECT -61.365 29.755 -61.035 30.085 ;
        RECT -61.365 28.395 -61.035 28.725 ;
        RECT -61.365 27.035 -61.035 27.365 ;
        RECT -61.365 25.675 -61.035 26.005 ;
        RECT -61.365 24.315 -61.035 24.645 ;
        RECT -61.365 22.955 -61.035 23.285 ;
        RECT -61.365 21.595 -61.035 21.925 ;
        RECT -61.365 20.235 -61.035 20.565 ;
        RECT -61.365 18.875 -61.035 19.205 ;
        RECT -61.365 17.515 -61.035 17.845 ;
        RECT -61.365 16.155 -61.035 16.485 ;
        RECT -61.365 14.795 -61.035 15.125 ;
        RECT -61.365 13.435 -61.035 13.765 ;
        RECT -61.365 12.075 -61.035 12.405 ;
        RECT -61.365 10.715 -61.035 11.045 ;
        RECT -61.365 9.355 -61.035 9.685 ;
        RECT -61.365 7.995 -61.035 8.325 ;
        RECT -61.365 6.635 -61.035 6.965 ;
        RECT -61.365 5.275 -61.035 5.605 ;
        RECT -61.365 3.915 -61.035 4.245 ;
        RECT -61.365 2.555 -61.035 2.885 ;
        RECT -61.365 1.195 -61.035 1.525 ;
        RECT -61.365 -0.165 -61.035 0.165 ;
        RECT -61.365 -1.525 -61.035 -1.195 ;
        RECT -61.365 -2.885 -61.035 -2.555 ;
        RECT -61.365 -4.245 -61.035 -3.915 ;
        RECT -61.365 -5.605 -61.035 -5.275 ;
        RECT -61.365 -6.965 -61.035 -6.635 ;
        RECT -61.365 -8.325 -61.035 -7.995 ;
        RECT -61.365 -9.685 -61.035 -9.355 ;
        RECT -61.365 -11.045 -61.035 -10.715 ;
        RECT -61.365 -12.405 -61.035 -12.075 ;
        RECT -61.365 -13.765 -61.035 -13.435 ;
        RECT -61.365 -15.125 -61.035 -14.795 ;
        RECT -61.365 -16.485 -61.035 -16.155 ;
        RECT -61.365 -17.845 -61.035 -17.515 ;
        RECT -61.365 -19.205 -61.035 -18.875 ;
        RECT -61.365 -20.565 -61.035 -20.235 ;
        RECT -61.365 -21.925 -61.035 -21.595 ;
        RECT -61.365 -23.285 -61.035 -22.955 ;
        RECT -61.365 -24.645 -61.035 -24.315 ;
        RECT -61.365 -26.005 -61.035 -25.675 ;
        RECT -61.365 -27.365 -61.035 -27.035 ;
        RECT -61.365 -28.725 -61.035 -28.395 ;
        RECT -61.365 -30.085 -61.035 -29.755 ;
        RECT -61.365 -31.445 -61.035 -31.115 ;
        RECT -61.365 -32.805 -61.035 -32.475 ;
        RECT -61.365 -34.165 -61.035 -33.835 ;
        RECT -61.365 -35.525 -61.035 -35.195 ;
        RECT -61.365 -36.885 -61.035 -36.555 ;
        RECT -61.365 -38.245 -61.035 -37.915 ;
        RECT -61.365 -39.605 -61.035 -39.275 ;
        RECT -61.365 -40.965 -61.035 -40.635 ;
        RECT -61.365 -42.325 -61.035 -41.995 ;
        RECT -61.365 -43.685 -61.035 -43.355 ;
        RECT -61.365 -45.045 -61.035 -44.715 ;
        RECT -61.365 -46.405 -61.035 -46.075 ;
        RECT -61.365 -47.765 -61.035 -47.435 ;
        RECT -61.365 -49.125 -61.035 -48.795 ;
        RECT -61.365 -50.485 -61.035 -50.155 ;
        RECT -61.365 -51.845 -61.035 -51.515 ;
        RECT -61.365 -53.205 -61.035 -52.875 ;
        RECT -61.365 -54.565 -61.035 -54.235 ;
        RECT -61.365 -55.925 -61.035 -55.595 ;
        RECT -61.365 -57.285 -61.035 -56.955 ;
        RECT -61.365 -58.645 -61.035 -58.315 ;
        RECT -61.365 -60.005 -61.035 -59.675 ;
        RECT -61.365 -61.365 -61.035 -61.035 ;
        RECT -61.365 -62.725 -61.035 -62.395 ;
        RECT -61.365 -64.085 -61.035 -63.755 ;
        RECT -61.365 -65.445 -61.035 -65.115 ;
        RECT -61.365 -66.805 -61.035 -66.475 ;
        RECT -61.365 -68.165 -61.035 -67.835 ;
        RECT -61.365 -69.525 -61.035 -69.195 ;
        RECT -61.365 -70.885 -61.035 -70.555 ;
        RECT -61.365 -72.245 -61.035 -71.915 ;
        RECT -61.365 -73.605 -61.035 -73.275 ;
        RECT -61.365 -74.965 -61.035 -74.635 ;
        RECT -61.365 -76.325 -61.035 -75.995 ;
        RECT -61.365 -77.685 -61.035 -77.355 ;
        RECT -61.365 -79.045 -61.035 -78.715 ;
        RECT -61.365 -80.405 -61.035 -80.075 ;
        RECT -61.365 -81.765 -61.035 -81.435 ;
        RECT -61.365 -83.125 -61.035 -82.795 ;
        RECT -61.365 -84.485 -61.035 -84.155 ;
        RECT -61.365 -85.845 -61.035 -85.515 ;
        RECT -61.365 -87.205 -61.035 -86.875 ;
        RECT -61.365 -88.565 -61.035 -88.235 ;
        RECT -61.365 -89.925 -61.035 -89.595 ;
        RECT -61.365 -91.285 -61.035 -90.955 ;
        RECT -61.365 -92.645 -61.035 -92.315 ;
        RECT -61.365 -94.005 -61.035 -93.675 ;
        RECT -61.365 -95.365 -61.035 -95.035 ;
        RECT -61.365 -96.725 -61.035 -96.395 ;
        RECT -61.365 -98.085 -61.035 -97.755 ;
        RECT -61.365 -99.445 -61.035 -99.115 ;
        RECT -61.365 -100.805 -61.035 -100.475 ;
        RECT -61.365 -102.165 -61.035 -101.835 ;
        RECT -61.365 -103.525 -61.035 -103.195 ;
        RECT -61.365 -104.885 -61.035 -104.555 ;
        RECT -61.365 -106.245 -61.035 -105.915 ;
        RECT -61.365 -107.605 -61.035 -107.275 ;
        RECT -61.365 -108.965 -61.035 -108.635 ;
        RECT -61.365 -110.325 -61.035 -109.995 ;
        RECT -61.365 -111.685 -61.035 -111.355 ;
        RECT -61.365 -113.045 -61.035 -112.715 ;
        RECT -61.365 -114.405 -61.035 -114.075 ;
        RECT -61.365 -115.765 -61.035 -115.435 ;
        RECT -61.365 -117.125 -61.035 -116.795 ;
        RECT -61.365 -118.485 -61.035 -118.155 ;
        RECT -61.365 -119.845 -61.035 -119.515 ;
        RECT -61.365 -121.205 -61.035 -120.875 ;
        RECT -61.365 -122.565 -61.035 -122.235 ;
        RECT -61.365 -123.925 -61.035 -123.595 ;
        RECT -61.365 -125.285 -61.035 -124.955 ;
        RECT -61.365 -126.645 -61.035 -126.315 ;
        RECT -61.365 -128.005 -61.035 -127.675 ;
        RECT -61.365 -129.365 -61.035 -129.035 ;
        RECT -61.365 -130.725 -61.035 -130.395 ;
        RECT -61.365 -132.085 -61.035 -131.755 ;
        RECT -61.365 -133.445 -61.035 -133.115 ;
        RECT -61.365 -134.805 -61.035 -134.475 ;
        RECT -61.365 -136.165 -61.035 -135.835 ;
        RECT -61.365 -137.525 -61.035 -137.195 ;
        RECT -61.365 -138.885 -61.035 -138.555 ;
        RECT -61.365 -140.245 -61.035 -139.915 ;
        RECT -61.365 -141.605 -61.035 -141.275 ;
        RECT -61.365 -142.965 -61.035 -142.635 ;
        RECT -61.365 -144.325 -61.035 -143.995 ;
        RECT -61.365 -145.685 -61.035 -145.355 ;
        RECT -61.365 -147.045 -61.035 -146.715 ;
        RECT -61.365 -149.765 -61.035 -149.435 ;
        RECT -61.365 -152.485 -61.035 -152.155 ;
        RECT -61.365 -153.845 -61.035 -153.515 ;
        RECT -61.365 -155.285 -61.035 -154.955 ;
        RECT -61.365 -156.565 -61.035 -156.235 ;
        RECT -61.365 -157.925 -61.035 -157.595 ;
        RECT -61.365 -160.17 -61.035 -159.04 ;
        RECT -61.36 -160.285 -61.04 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 -88.565 -59.675 -88.235 ;
        RECT -60.005 -89.925 -59.675 -89.595 ;
        RECT -60.005 -91.285 -59.675 -90.955 ;
        RECT -60 -91.285 -59.68 128.47 ;
        RECT -60.005 127.225 -59.675 128.355 ;
        RECT -60.005 124.955 -59.675 125.285 ;
        RECT -60.005 123.595 -59.675 123.925 ;
        RECT -60.005 122.235 -59.675 122.565 ;
        RECT -60.005 120.875 -59.675 121.205 ;
        RECT -60.005 119.515 -59.675 119.845 ;
        RECT -60.005 118.155 -59.675 118.485 ;
        RECT -60.005 116.795 -59.675 117.125 ;
        RECT -60.005 115.435 -59.675 115.765 ;
        RECT -60.005 114.075 -59.675 114.405 ;
        RECT -60.005 112.715 -59.675 113.045 ;
        RECT -60.005 111.355 -59.675 111.685 ;
        RECT -60.005 109.995 -59.675 110.325 ;
        RECT -60.005 108.635 -59.675 108.965 ;
        RECT -60.005 107.275 -59.675 107.605 ;
        RECT -60.005 105.915 -59.675 106.245 ;
        RECT -60.005 104.555 -59.675 104.885 ;
        RECT -60.005 103.195 -59.675 103.525 ;
        RECT -60.005 101.835 -59.675 102.165 ;
        RECT -60.005 100.475 -59.675 100.805 ;
        RECT -60.005 99.115 -59.675 99.445 ;
        RECT -60.005 97.755 -59.675 98.085 ;
        RECT -60.005 96.395 -59.675 96.725 ;
        RECT -60.005 95.035 -59.675 95.365 ;
        RECT -60.005 93.675 -59.675 94.005 ;
        RECT -60.005 92.315 -59.675 92.645 ;
        RECT -60.005 90.955 -59.675 91.285 ;
        RECT -60.005 89.595 -59.675 89.925 ;
        RECT -60.005 88.235 -59.675 88.565 ;
        RECT -60.005 86.875 -59.675 87.205 ;
        RECT -60.005 85.515 -59.675 85.845 ;
        RECT -60.005 84.155 -59.675 84.485 ;
        RECT -60.005 82.795 -59.675 83.125 ;
        RECT -60.005 81.435 -59.675 81.765 ;
        RECT -60.005 80.075 -59.675 80.405 ;
        RECT -60.005 78.715 -59.675 79.045 ;
        RECT -60.005 77.355 -59.675 77.685 ;
        RECT -60.005 75.995 -59.675 76.325 ;
        RECT -60.005 74.635 -59.675 74.965 ;
        RECT -60.005 73.275 -59.675 73.605 ;
        RECT -60.005 72.445 -59.675 72.775 ;
        RECT -60.005 70.395 -59.675 70.725 ;
        RECT -60.005 68.035 -59.675 68.365 ;
        RECT -60.005 66.885 -59.675 67.215 ;
        RECT -60.005 64.875 -59.675 65.205 ;
        RECT -60.005 63.725 -59.675 64.055 ;
        RECT -60.005 61.715 -59.675 62.045 ;
        RECT -60.005 60.395 -59.675 60.725 ;
        RECT -60.005 58.555 -59.675 58.885 ;
        RECT -60.005 57.405 -59.675 57.735 ;
        RECT -60.005 55.395 -59.675 55.725 ;
        RECT -60.005 54.245 -59.675 54.575 ;
        RECT -60.005 51.885 -59.675 52.215 ;
        RECT -60.005 49.83 -59.675 50.16 ;
        RECT -60.005 48.795 -59.675 49.125 ;
        RECT -60.005 47.435 -59.675 47.765 ;
        RECT -60.005 46.075 -59.675 46.405 ;
        RECT -60.005 44.715 -59.675 45.045 ;
        RECT -60.005 43.355 -59.675 43.685 ;
        RECT -60.005 41.995 -59.675 42.325 ;
        RECT -60.005 40.635 -59.675 40.965 ;
        RECT -60.005 39.275 -59.675 39.605 ;
        RECT -60.005 37.915 -59.675 38.245 ;
        RECT -60.005 36.555 -59.675 36.885 ;
        RECT -60.005 35.195 -59.675 35.525 ;
        RECT -60.005 33.835 -59.675 34.165 ;
        RECT -60.005 32.475 -59.675 32.805 ;
        RECT -60.005 31.115 -59.675 31.445 ;
        RECT -60.005 29.755 -59.675 30.085 ;
        RECT -60.005 28.395 -59.675 28.725 ;
        RECT -60.005 27.035 -59.675 27.365 ;
        RECT -60.005 25.675 -59.675 26.005 ;
        RECT -60.005 24.315 -59.675 24.645 ;
        RECT -60.005 22.955 -59.675 23.285 ;
        RECT -60.005 21.595 -59.675 21.925 ;
        RECT -60.005 20.235 -59.675 20.565 ;
        RECT -60.005 18.875 -59.675 19.205 ;
        RECT -60.005 17.515 -59.675 17.845 ;
        RECT -60.005 16.155 -59.675 16.485 ;
        RECT -60.005 14.795 -59.675 15.125 ;
        RECT -60.005 13.435 -59.675 13.765 ;
        RECT -60.005 12.075 -59.675 12.405 ;
        RECT -60.005 10.715 -59.675 11.045 ;
        RECT -60.005 9.355 -59.675 9.685 ;
        RECT -60.005 7.995 -59.675 8.325 ;
        RECT -60.005 6.635 -59.675 6.965 ;
        RECT -60.005 5.275 -59.675 5.605 ;
        RECT -60.005 3.915 -59.675 4.245 ;
        RECT -60.005 2.555 -59.675 2.885 ;
        RECT -60.005 1.195 -59.675 1.525 ;
        RECT -60.005 -0.165 -59.675 0.165 ;
        RECT -60.005 -1.525 -59.675 -1.195 ;
        RECT -60.005 -2.885 -59.675 -2.555 ;
        RECT -60.005 -4.245 -59.675 -3.915 ;
        RECT -60.005 -5.605 -59.675 -5.275 ;
        RECT -60.005 -6.965 -59.675 -6.635 ;
        RECT -60.005 -8.325 -59.675 -7.995 ;
        RECT -60.005 -9.685 -59.675 -9.355 ;
        RECT -60.005 -11.045 -59.675 -10.715 ;
        RECT -60.005 -12.405 -59.675 -12.075 ;
        RECT -60.005 -13.765 -59.675 -13.435 ;
        RECT -60.005 -15.125 -59.675 -14.795 ;
        RECT -60.005 -16.485 -59.675 -16.155 ;
        RECT -60.005 -17.845 -59.675 -17.515 ;
        RECT -60.005 -19.205 -59.675 -18.875 ;
        RECT -60.005 -20.565 -59.675 -20.235 ;
        RECT -60.005 -21.925 -59.675 -21.595 ;
        RECT -60.005 -23.285 -59.675 -22.955 ;
        RECT -60.005 -24.645 -59.675 -24.315 ;
        RECT -60.005 -26.005 -59.675 -25.675 ;
        RECT -60.005 -27.365 -59.675 -27.035 ;
        RECT -60.005 -28.725 -59.675 -28.395 ;
        RECT -60.005 -30.085 -59.675 -29.755 ;
        RECT -60.005 -31.445 -59.675 -31.115 ;
        RECT -60.005 -32.805 -59.675 -32.475 ;
        RECT -60.005 -34.165 -59.675 -33.835 ;
        RECT -60.005 -35.525 -59.675 -35.195 ;
        RECT -60.005 -36.885 -59.675 -36.555 ;
        RECT -60.005 -38.245 -59.675 -37.915 ;
        RECT -60.005 -39.605 -59.675 -39.275 ;
        RECT -60.005 -40.965 -59.675 -40.635 ;
        RECT -60.005 -42.325 -59.675 -41.995 ;
        RECT -60.005 -43.685 -59.675 -43.355 ;
        RECT -60.005 -45.045 -59.675 -44.715 ;
        RECT -60.005 -46.405 -59.675 -46.075 ;
        RECT -60.005 -47.765 -59.675 -47.435 ;
        RECT -60.005 -49.125 -59.675 -48.795 ;
        RECT -60.005 -50.485 -59.675 -50.155 ;
        RECT -60.005 -51.845 -59.675 -51.515 ;
        RECT -60.005 -53.205 -59.675 -52.875 ;
        RECT -60.005 -54.565 -59.675 -54.235 ;
        RECT -60.005 -55.925 -59.675 -55.595 ;
        RECT -60.005 -57.285 -59.675 -56.955 ;
        RECT -60.005 -58.645 -59.675 -58.315 ;
        RECT -60.005 -60.005 -59.675 -59.675 ;
        RECT -60.005 -61.365 -59.675 -61.035 ;
        RECT -60.005 -62.725 -59.675 -62.395 ;
        RECT -60.005 -64.085 -59.675 -63.755 ;
        RECT -60.005 -65.445 -59.675 -65.115 ;
        RECT -60.005 -66.805 -59.675 -66.475 ;
        RECT -60.005 -68.165 -59.675 -67.835 ;
        RECT -60.005 -69.525 -59.675 -69.195 ;
        RECT -60.005 -70.885 -59.675 -70.555 ;
        RECT -60.005 -72.245 -59.675 -71.915 ;
        RECT -60.005 -73.605 -59.675 -73.275 ;
        RECT -60.005 -74.965 -59.675 -74.635 ;
        RECT -60.005 -76.325 -59.675 -75.995 ;
        RECT -60.005 -77.685 -59.675 -77.355 ;
        RECT -60.005 -79.045 -59.675 -78.715 ;
        RECT -60.005 -80.405 -59.675 -80.075 ;
        RECT -60.005 -81.765 -59.675 -81.435 ;
        RECT -60.005 -83.125 -59.675 -82.795 ;
        RECT -60.005 -84.485 -59.675 -84.155 ;
        RECT -60.005 -85.845 -59.675 -85.515 ;
        RECT -60.005 -87.205 -59.675 -86.875 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.165 127.225 -67.835 128.355 ;
        RECT -68.165 124.955 -67.835 125.285 ;
        RECT -68.165 123.595 -67.835 123.925 ;
        RECT -68.165 122.235 -67.835 122.565 ;
        RECT -68.165 120.875 -67.835 121.205 ;
        RECT -68.165 119.515 -67.835 119.845 ;
        RECT -68.165 118.155 -67.835 118.485 ;
        RECT -68.165 116.795 -67.835 117.125 ;
        RECT -68.165 115.435 -67.835 115.765 ;
        RECT -68.165 114.075 -67.835 114.405 ;
        RECT -68.165 112.715 -67.835 113.045 ;
        RECT -68.165 111.355 -67.835 111.685 ;
        RECT -68.165 109.995 -67.835 110.325 ;
        RECT -68.165 108.635 -67.835 108.965 ;
        RECT -68.165 107.275 -67.835 107.605 ;
        RECT -68.165 105.915 -67.835 106.245 ;
        RECT -68.165 104.555 -67.835 104.885 ;
        RECT -68.165 103.195 -67.835 103.525 ;
        RECT -68.165 101.835 -67.835 102.165 ;
        RECT -68.165 100.475 -67.835 100.805 ;
        RECT -68.165 99.115 -67.835 99.445 ;
        RECT -68.165 97.755 -67.835 98.085 ;
        RECT -68.165 96.395 -67.835 96.725 ;
        RECT -68.165 95.035 -67.835 95.365 ;
        RECT -68.165 93.675 -67.835 94.005 ;
        RECT -68.165 92.315 -67.835 92.645 ;
        RECT -68.165 90.955 -67.835 91.285 ;
        RECT -68.165 89.595 -67.835 89.925 ;
        RECT -68.165 88.235 -67.835 88.565 ;
        RECT -68.165 86.875 -67.835 87.205 ;
        RECT -68.165 85.515 -67.835 85.845 ;
        RECT -68.165 84.155 -67.835 84.485 ;
        RECT -68.165 82.795 -67.835 83.125 ;
        RECT -68.165 81.435 -67.835 81.765 ;
        RECT -68.165 80.075 -67.835 80.405 ;
        RECT -68.165 78.715 -67.835 79.045 ;
        RECT -68.165 77.355 -67.835 77.685 ;
        RECT -68.165 75.995 -67.835 76.325 ;
        RECT -68.165 74.635 -67.835 74.965 ;
        RECT -68.165 73.275 -67.835 73.605 ;
        RECT -68.165 71.915 -67.835 72.245 ;
        RECT -68.165 70.555 -67.835 70.885 ;
        RECT -68.165 69.195 -67.835 69.525 ;
        RECT -68.165 67.835 -67.835 68.165 ;
        RECT -68.165 66.475 -67.835 66.805 ;
        RECT -68.165 65.115 -67.835 65.445 ;
        RECT -68.165 63.755 -67.835 64.085 ;
        RECT -68.165 62.395 -67.835 62.725 ;
        RECT -68.165 61.035 -67.835 61.365 ;
        RECT -68.165 59.675 -67.835 60.005 ;
        RECT -68.165 58.315 -67.835 58.645 ;
        RECT -68.165 56.955 -67.835 57.285 ;
        RECT -68.165 55.595 -67.835 55.925 ;
        RECT -68.165 54.235 -67.835 54.565 ;
        RECT -68.165 52.875 -67.835 53.205 ;
        RECT -68.165 51.515 -67.835 51.845 ;
        RECT -68.165 50.155 -67.835 50.485 ;
        RECT -68.165 48.795 -67.835 49.125 ;
        RECT -68.165 47.435 -67.835 47.765 ;
        RECT -68.165 46.075 -67.835 46.405 ;
        RECT -68.165 44.715 -67.835 45.045 ;
        RECT -68.165 43.355 -67.835 43.685 ;
        RECT -68.165 41.995 -67.835 42.325 ;
        RECT -68.165 40.635 -67.835 40.965 ;
        RECT -68.165 39.275 -67.835 39.605 ;
        RECT -68.165 37.915 -67.835 38.245 ;
        RECT -68.165 36.555 -67.835 36.885 ;
        RECT -68.165 35.195 -67.835 35.525 ;
        RECT -68.165 33.835 -67.835 34.165 ;
        RECT -68.165 32.475 -67.835 32.805 ;
        RECT -68.165 31.115 -67.835 31.445 ;
        RECT -68.165 29.755 -67.835 30.085 ;
        RECT -68.165 28.395 -67.835 28.725 ;
        RECT -68.165 27.035 -67.835 27.365 ;
        RECT -68.165 25.675 -67.835 26.005 ;
        RECT -68.165 24.315 -67.835 24.645 ;
        RECT -68.165 22.955 -67.835 23.285 ;
        RECT -68.165 21.595 -67.835 21.925 ;
        RECT -68.165 20.235 -67.835 20.565 ;
        RECT -68.165 18.875 -67.835 19.205 ;
        RECT -68.165 17.515 -67.835 17.845 ;
        RECT -68.165 16.155 -67.835 16.485 ;
        RECT -68.165 14.795 -67.835 15.125 ;
        RECT -68.165 13.435 -67.835 13.765 ;
        RECT -68.165 12.075 -67.835 12.405 ;
        RECT -68.165 10.715 -67.835 11.045 ;
        RECT -68.165 9.355 -67.835 9.685 ;
        RECT -68.165 7.995 -67.835 8.325 ;
        RECT -68.165 6.635 -67.835 6.965 ;
        RECT -68.165 5.275 -67.835 5.605 ;
        RECT -68.165 3.915 -67.835 4.245 ;
        RECT -68.165 2.555 -67.835 2.885 ;
        RECT -68.165 1.195 -67.835 1.525 ;
        RECT -68.165 -0.165 -67.835 0.165 ;
        RECT -68.165 -1.525 -67.835 -1.195 ;
        RECT -68.165 -2.885 -67.835 -2.555 ;
        RECT -68.165 -4.245 -67.835 -3.915 ;
        RECT -68.165 -5.605 -67.835 -5.275 ;
        RECT -68.165 -6.965 -67.835 -6.635 ;
        RECT -68.165 -8.325 -67.835 -7.995 ;
        RECT -68.165 -9.685 -67.835 -9.355 ;
        RECT -68.165 -11.045 -67.835 -10.715 ;
        RECT -68.165 -12.405 -67.835 -12.075 ;
        RECT -68.165 -13.765 -67.835 -13.435 ;
        RECT -68.165 -15.125 -67.835 -14.795 ;
        RECT -68.165 -16.485 -67.835 -16.155 ;
        RECT -68.165 -17.845 -67.835 -17.515 ;
        RECT -68.165 -19.205 -67.835 -18.875 ;
        RECT -68.165 -20.565 -67.835 -20.235 ;
        RECT -68.165 -21.925 -67.835 -21.595 ;
        RECT -68.165 -23.285 -67.835 -22.955 ;
        RECT -68.165 -24.645 -67.835 -24.315 ;
        RECT -68.165 -26.005 -67.835 -25.675 ;
        RECT -68.165 -27.365 -67.835 -27.035 ;
        RECT -68.165 -28.725 -67.835 -28.395 ;
        RECT -68.165 -30.085 -67.835 -29.755 ;
        RECT -68.165 -31.445 -67.835 -31.115 ;
        RECT -68.165 -32.805 -67.835 -32.475 ;
        RECT -68.165 -34.165 -67.835 -33.835 ;
        RECT -68.165 -35.525 -67.835 -35.195 ;
        RECT -68.165 -36.885 -67.835 -36.555 ;
        RECT -68.165 -38.245 -67.835 -37.915 ;
        RECT -68.165 -39.605 -67.835 -39.275 ;
        RECT -68.165 -40.965 -67.835 -40.635 ;
        RECT -68.165 -42.325 -67.835 -41.995 ;
        RECT -68.165 -43.685 -67.835 -43.355 ;
        RECT -68.165 -45.045 -67.835 -44.715 ;
        RECT -68.165 -46.405 -67.835 -46.075 ;
        RECT -68.165 -47.765 -67.835 -47.435 ;
        RECT -68.165 -49.125 -67.835 -48.795 ;
        RECT -68.165 -50.485 -67.835 -50.155 ;
        RECT -68.165 -51.845 -67.835 -51.515 ;
        RECT -68.165 -53.205 -67.835 -52.875 ;
        RECT -68.165 -54.565 -67.835 -54.235 ;
        RECT -68.165 -55.925 -67.835 -55.595 ;
        RECT -68.165 -57.285 -67.835 -56.955 ;
        RECT -68.165 -58.645 -67.835 -58.315 ;
        RECT -68.165 -60.005 -67.835 -59.675 ;
        RECT -68.165 -61.365 -67.835 -61.035 ;
        RECT -68.165 -62.725 -67.835 -62.395 ;
        RECT -68.165 -64.085 -67.835 -63.755 ;
        RECT -68.165 -65.445 -67.835 -65.115 ;
        RECT -68.165 -66.805 -67.835 -66.475 ;
        RECT -68.165 -68.165 -67.835 -67.835 ;
        RECT -68.165 -69.525 -67.835 -69.195 ;
        RECT -68.165 -70.885 -67.835 -70.555 ;
        RECT -68.165 -72.245 -67.835 -71.915 ;
        RECT -68.165 -73.605 -67.835 -73.275 ;
        RECT -68.165 -74.965 -67.835 -74.635 ;
        RECT -68.165 -76.325 -67.835 -75.995 ;
        RECT -68.165 -77.685 -67.835 -77.355 ;
        RECT -68.165 -79.045 -67.835 -78.715 ;
        RECT -68.165 -80.405 -67.835 -80.075 ;
        RECT -68.165 -81.765 -67.835 -81.435 ;
        RECT -68.165 -83.125 -67.835 -82.795 ;
        RECT -68.165 -84.485 -67.835 -84.155 ;
        RECT -68.165 -85.845 -67.835 -85.515 ;
        RECT -68.165 -87.205 -67.835 -86.875 ;
        RECT -68.165 -88.565 -67.835 -88.235 ;
        RECT -68.165 -89.925 -67.835 -89.595 ;
        RECT -68.165 -91.285 -67.835 -90.955 ;
        RECT -68.165 -92.645 -67.835 -92.315 ;
        RECT -68.165 -94.005 -67.835 -93.675 ;
        RECT -68.165 -95.365 -67.835 -95.035 ;
        RECT -68.165 -96.725 -67.835 -96.395 ;
        RECT -68.165 -98.085 -67.835 -97.755 ;
        RECT -68.165 -99.445 -67.835 -99.115 ;
        RECT -68.165 -100.805 -67.835 -100.475 ;
        RECT -68.165 -102.165 -67.835 -101.835 ;
        RECT -68.165 -103.525 -67.835 -103.195 ;
        RECT -68.165 -104.885 -67.835 -104.555 ;
        RECT -68.165 -106.245 -67.835 -105.915 ;
        RECT -68.165 -107.605 -67.835 -107.275 ;
        RECT -68.165 -108.965 -67.835 -108.635 ;
        RECT -68.165 -110.325 -67.835 -109.995 ;
        RECT -68.165 -111.685 -67.835 -111.355 ;
        RECT -68.165 -113.045 -67.835 -112.715 ;
        RECT -68.165 -114.405 -67.835 -114.075 ;
        RECT -68.165 -115.765 -67.835 -115.435 ;
        RECT -68.165 -117.125 -67.835 -116.795 ;
        RECT -68.165 -118.485 -67.835 -118.155 ;
        RECT -68.165 -119.845 -67.835 -119.515 ;
        RECT -68.165 -121.205 -67.835 -120.875 ;
        RECT -68.165 -122.565 -67.835 -122.235 ;
        RECT -68.165 -123.925 -67.835 -123.595 ;
        RECT -68.165 -125.285 -67.835 -124.955 ;
        RECT -68.165 -126.645 -67.835 -126.315 ;
        RECT -68.165 -128.005 -67.835 -127.675 ;
        RECT -68.165 -129.365 -67.835 -129.035 ;
        RECT -68.165 -130.725 -67.835 -130.395 ;
        RECT -68.165 -132.085 -67.835 -131.755 ;
        RECT -68.165 -133.445 -67.835 -133.115 ;
        RECT -68.165 -134.805 -67.835 -134.475 ;
        RECT -68.165 -136.165 -67.835 -135.835 ;
        RECT -68.165 -137.525 -67.835 -137.195 ;
        RECT -68.165 -138.885 -67.835 -138.555 ;
        RECT -68.165 -140.245 -67.835 -139.915 ;
        RECT -68.165 -141.605 -67.835 -141.275 ;
        RECT -68.165 -142.965 -67.835 -142.635 ;
        RECT -68.165 -144.325 -67.835 -143.995 ;
        RECT -68.165 -145.685 -67.835 -145.355 ;
        RECT -68.165 -147.045 -67.835 -146.715 ;
        RECT -68.165 -148.405 -67.835 -148.075 ;
        RECT -68.165 -149.765 -67.835 -149.435 ;
        RECT -68.165 -151.125 -67.835 -150.795 ;
        RECT -68.165 -152.485 -67.835 -152.155 ;
        RECT -68.165 -153.845 -67.835 -153.515 ;
        RECT -68.165 -155.205 -67.835 -154.875 ;
        RECT -68.165 -156.565 -67.835 -156.235 ;
        RECT -68.165 -157.925 -67.835 -157.595 ;
        RECT -68.165 -160.17 -67.835 -159.04 ;
        RECT -68.16 -160.285 -67.84 128.47 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.805 -87.205 -66.475 -86.875 ;
        RECT -66.805 -88.565 -66.475 -88.235 ;
        RECT -66.805 -89.925 -66.475 -89.595 ;
        RECT -66.805 -91.285 -66.475 -90.955 ;
        RECT -66.805 -92.645 -66.475 -92.315 ;
        RECT -66.805 -94.005 -66.475 -93.675 ;
        RECT -66.805 -95.365 -66.475 -95.035 ;
        RECT -66.805 -96.725 -66.475 -96.395 ;
        RECT -66.805 -98.085 -66.475 -97.755 ;
        RECT -66.805 -99.445 -66.475 -99.115 ;
        RECT -66.805 -100.805 -66.475 -100.475 ;
        RECT -66.805 -102.165 -66.475 -101.835 ;
        RECT -66.805 -103.525 -66.475 -103.195 ;
        RECT -66.805 -104.885 -66.475 -104.555 ;
        RECT -66.805 -106.245 -66.475 -105.915 ;
        RECT -66.805 -107.605 -66.475 -107.275 ;
        RECT -66.805 -108.965 -66.475 -108.635 ;
        RECT -66.805 -110.325 -66.475 -109.995 ;
        RECT -66.805 -111.685 -66.475 -111.355 ;
        RECT -66.805 -113.045 -66.475 -112.715 ;
        RECT -66.805 -114.405 -66.475 -114.075 ;
        RECT -66.805 -115.765 -66.475 -115.435 ;
        RECT -66.805 -117.125 -66.475 -116.795 ;
        RECT -66.805 -118.485 -66.475 -118.155 ;
        RECT -66.805 -119.845 -66.475 -119.515 ;
        RECT -66.805 -121.205 -66.475 -120.875 ;
        RECT -66.805 -122.565 -66.475 -122.235 ;
        RECT -66.805 -123.925 -66.475 -123.595 ;
        RECT -66.805 -125.285 -66.475 -124.955 ;
        RECT -66.805 -126.645 -66.475 -126.315 ;
        RECT -66.805 -128.005 -66.475 -127.675 ;
        RECT -66.805 -129.365 -66.475 -129.035 ;
        RECT -66.805 -130.725 -66.475 -130.395 ;
        RECT -66.805 -132.085 -66.475 -131.755 ;
        RECT -66.805 -133.445 -66.475 -133.115 ;
        RECT -66.805 -134.805 -66.475 -134.475 ;
        RECT -66.805 -136.165 -66.475 -135.835 ;
        RECT -66.805 -137.525 -66.475 -137.195 ;
        RECT -66.805 -138.885 -66.475 -138.555 ;
        RECT -66.805 -140.245 -66.475 -139.915 ;
        RECT -66.805 -141.605 -66.475 -141.275 ;
        RECT -66.805 -142.965 -66.475 -142.635 ;
        RECT -66.805 -144.325 -66.475 -143.995 ;
        RECT -66.805 -145.685 -66.475 -145.355 ;
        RECT -66.805 -147.045 -66.475 -146.715 ;
        RECT -66.805 -148.405 -66.475 -148.075 ;
        RECT -66.805 -149.765 -66.475 -149.435 ;
        RECT -66.805 -151.125 -66.475 -150.795 ;
        RECT -66.805 -152.485 -66.475 -152.155 ;
        RECT -66.805 -153.845 -66.475 -153.515 ;
        RECT -66.805 -155.205 -66.475 -154.875 ;
        RECT -66.805 -156.565 -66.475 -156.235 ;
        RECT -66.805 -157.925 -66.475 -157.595 ;
        RECT -66.805 -160.17 -66.475 -159.04 ;
        RECT -66.8 -160.285 -66.48 128.47 ;
        RECT -66.805 127.225 -66.475 128.355 ;
        RECT -66.805 124.955 -66.475 125.285 ;
        RECT -66.805 123.595 -66.475 123.925 ;
        RECT -66.805 122.235 -66.475 122.565 ;
        RECT -66.805 120.875 -66.475 121.205 ;
        RECT -66.805 119.515 -66.475 119.845 ;
        RECT -66.805 118.155 -66.475 118.485 ;
        RECT -66.805 116.795 -66.475 117.125 ;
        RECT -66.805 115.435 -66.475 115.765 ;
        RECT -66.805 114.075 -66.475 114.405 ;
        RECT -66.805 112.715 -66.475 113.045 ;
        RECT -66.805 111.355 -66.475 111.685 ;
        RECT -66.805 109.995 -66.475 110.325 ;
        RECT -66.805 108.635 -66.475 108.965 ;
        RECT -66.805 107.275 -66.475 107.605 ;
        RECT -66.805 105.915 -66.475 106.245 ;
        RECT -66.805 104.555 -66.475 104.885 ;
        RECT -66.805 103.195 -66.475 103.525 ;
        RECT -66.805 101.835 -66.475 102.165 ;
        RECT -66.805 100.475 -66.475 100.805 ;
        RECT -66.805 99.115 -66.475 99.445 ;
        RECT -66.805 97.755 -66.475 98.085 ;
        RECT -66.805 96.395 -66.475 96.725 ;
        RECT -66.805 95.035 -66.475 95.365 ;
        RECT -66.805 93.675 -66.475 94.005 ;
        RECT -66.805 92.315 -66.475 92.645 ;
        RECT -66.805 90.955 -66.475 91.285 ;
        RECT -66.805 89.595 -66.475 89.925 ;
        RECT -66.805 88.235 -66.475 88.565 ;
        RECT -66.805 86.875 -66.475 87.205 ;
        RECT -66.805 85.515 -66.475 85.845 ;
        RECT -66.805 84.155 -66.475 84.485 ;
        RECT -66.805 82.795 -66.475 83.125 ;
        RECT -66.805 81.435 -66.475 81.765 ;
        RECT -66.805 80.075 -66.475 80.405 ;
        RECT -66.805 78.715 -66.475 79.045 ;
        RECT -66.805 77.355 -66.475 77.685 ;
        RECT -66.805 75.995 -66.475 76.325 ;
        RECT -66.805 74.635 -66.475 74.965 ;
        RECT -66.805 73.275 -66.475 73.605 ;
        RECT -66.805 71.915 -66.475 72.245 ;
        RECT -66.805 70.555 -66.475 70.885 ;
        RECT -66.805 69.195 -66.475 69.525 ;
        RECT -66.805 67.835 -66.475 68.165 ;
        RECT -66.805 66.475 -66.475 66.805 ;
        RECT -66.805 65.115 -66.475 65.445 ;
        RECT -66.805 63.755 -66.475 64.085 ;
        RECT -66.805 62.395 -66.475 62.725 ;
        RECT -66.805 61.035 -66.475 61.365 ;
        RECT -66.805 59.675 -66.475 60.005 ;
        RECT -66.805 58.315 -66.475 58.645 ;
        RECT -66.805 56.955 -66.475 57.285 ;
        RECT -66.805 55.595 -66.475 55.925 ;
        RECT -66.805 54.235 -66.475 54.565 ;
        RECT -66.805 52.875 -66.475 53.205 ;
        RECT -66.805 51.515 -66.475 51.845 ;
        RECT -66.805 50.155 -66.475 50.485 ;
        RECT -66.805 48.795 -66.475 49.125 ;
        RECT -66.805 47.435 -66.475 47.765 ;
        RECT -66.805 46.075 -66.475 46.405 ;
        RECT -66.805 44.715 -66.475 45.045 ;
        RECT -66.805 43.355 -66.475 43.685 ;
        RECT -66.805 41.995 -66.475 42.325 ;
        RECT -66.805 40.635 -66.475 40.965 ;
        RECT -66.805 39.275 -66.475 39.605 ;
        RECT -66.805 37.915 -66.475 38.245 ;
        RECT -66.805 36.555 -66.475 36.885 ;
        RECT -66.805 35.195 -66.475 35.525 ;
        RECT -66.805 33.835 -66.475 34.165 ;
        RECT -66.805 32.475 -66.475 32.805 ;
        RECT -66.805 31.115 -66.475 31.445 ;
        RECT -66.805 29.755 -66.475 30.085 ;
        RECT -66.805 28.395 -66.475 28.725 ;
        RECT -66.805 27.035 -66.475 27.365 ;
        RECT -66.805 25.675 -66.475 26.005 ;
        RECT -66.805 24.315 -66.475 24.645 ;
        RECT -66.805 22.955 -66.475 23.285 ;
        RECT -66.805 21.595 -66.475 21.925 ;
        RECT -66.805 20.235 -66.475 20.565 ;
        RECT -66.805 18.875 -66.475 19.205 ;
        RECT -66.805 17.515 -66.475 17.845 ;
        RECT -66.805 16.155 -66.475 16.485 ;
        RECT -66.805 14.795 -66.475 15.125 ;
        RECT -66.805 13.435 -66.475 13.765 ;
        RECT -66.805 12.075 -66.475 12.405 ;
        RECT -66.805 10.715 -66.475 11.045 ;
        RECT -66.805 9.355 -66.475 9.685 ;
        RECT -66.805 7.995 -66.475 8.325 ;
        RECT -66.805 6.635 -66.475 6.965 ;
        RECT -66.805 5.275 -66.475 5.605 ;
        RECT -66.805 3.915 -66.475 4.245 ;
        RECT -66.805 2.555 -66.475 2.885 ;
        RECT -66.805 1.195 -66.475 1.525 ;
        RECT -66.805 -0.165 -66.475 0.165 ;
        RECT -66.805 -1.525 -66.475 -1.195 ;
        RECT -66.805 -2.885 -66.475 -2.555 ;
        RECT -66.805 -4.245 -66.475 -3.915 ;
        RECT -66.805 -5.605 -66.475 -5.275 ;
        RECT -66.805 -6.965 -66.475 -6.635 ;
        RECT -66.805 -8.325 -66.475 -7.995 ;
        RECT -66.805 -9.685 -66.475 -9.355 ;
        RECT -66.805 -11.045 -66.475 -10.715 ;
        RECT -66.805 -12.405 -66.475 -12.075 ;
        RECT -66.805 -13.765 -66.475 -13.435 ;
        RECT -66.805 -15.125 -66.475 -14.795 ;
        RECT -66.805 -16.485 -66.475 -16.155 ;
        RECT -66.805 -17.845 -66.475 -17.515 ;
        RECT -66.805 -19.205 -66.475 -18.875 ;
        RECT -66.805 -20.565 -66.475 -20.235 ;
        RECT -66.805 -21.925 -66.475 -21.595 ;
        RECT -66.805 -23.285 -66.475 -22.955 ;
        RECT -66.805 -24.645 -66.475 -24.315 ;
        RECT -66.805 -26.005 -66.475 -25.675 ;
        RECT -66.805 -27.365 -66.475 -27.035 ;
        RECT -66.805 -28.725 -66.475 -28.395 ;
        RECT -66.805 -30.085 -66.475 -29.755 ;
        RECT -66.805 -31.445 -66.475 -31.115 ;
        RECT -66.805 -32.805 -66.475 -32.475 ;
        RECT -66.805 -34.165 -66.475 -33.835 ;
        RECT -66.805 -35.525 -66.475 -35.195 ;
        RECT -66.805 -36.885 -66.475 -36.555 ;
        RECT -66.805 -38.245 -66.475 -37.915 ;
        RECT -66.805 -39.605 -66.475 -39.275 ;
        RECT -66.805 -40.965 -66.475 -40.635 ;
        RECT -66.805 -42.325 -66.475 -41.995 ;
        RECT -66.805 -43.685 -66.475 -43.355 ;
        RECT -66.805 -45.045 -66.475 -44.715 ;
        RECT -66.805 -46.405 -66.475 -46.075 ;
        RECT -66.805 -47.765 -66.475 -47.435 ;
        RECT -66.805 -49.125 -66.475 -48.795 ;
        RECT -66.805 -50.485 -66.475 -50.155 ;
        RECT -66.805 -51.845 -66.475 -51.515 ;
        RECT -66.805 -53.205 -66.475 -52.875 ;
        RECT -66.805 -54.565 -66.475 -54.235 ;
        RECT -66.805 -55.925 -66.475 -55.595 ;
        RECT -66.805 -57.285 -66.475 -56.955 ;
        RECT -66.805 -58.645 -66.475 -58.315 ;
        RECT -66.805 -60.005 -66.475 -59.675 ;
        RECT -66.805 -61.365 -66.475 -61.035 ;
        RECT -66.805 -62.725 -66.475 -62.395 ;
        RECT -66.805 -64.085 -66.475 -63.755 ;
        RECT -66.805 -65.445 -66.475 -65.115 ;
        RECT -66.805 -66.805 -66.475 -66.475 ;
        RECT -66.805 -68.165 -66.475 -67.835 ;
        RECT -66.805 -69.525 -66.475 -69.195 ;
        RECT -66.805 -70.885 -66.475 -70.555 ;
        RECT -66.805 -72.245 -66.475 -71.915 ;
        RECT -66.805 -73.605 -66.475 -73.275 ;
        RECT -66.805 -74.965 -66.475 -74.635 ;
        RECT -66.805 -76.325 -66.475 -75.995 ;
        RECT -66.805 -77.685 -66.475 -77.355 ;
        RECT -66.805 -79.045 -66.475 -78.715 ;
        RECT -66.805 -80.405 -66.475 -80.075 ;
        RECT -66.805 -81.765 -66.475 -81.435 ;
        RECT -66.805 -83.125 -66.475 -82.795 ;
        RECT -66.805 -84.485 -66.475 -84.155 ;
        RECT -66.805 -85.845 -66.475 -85.515 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -21.24 -163.165 -20.92 -162.845 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -27.36 -163.165 -27.04 -162.845 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -33.48 -163.165 -33.16 -162.845 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -39.6 -163.165 -39.28 -162.845 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -46.4 -163.165 -46.08 -162.845 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -52.52 -163.165 -52.2 -162.845 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -58.64 -163.165 -58.32 -162.845 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -64.76 -163.165 -64.44 -162.845 ;
    END
  END addr[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -9.68 -163.165 -9.36 -162.845 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.6 -163.165 6 -162.765 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.6 -163.165 67 -162.765 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.7 -163.165 73.1 -162.765 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.8 -163.165 79.2 -162.765 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.9 -163.165 85.3 -162.765 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91 -163.165 91.4 -162.765 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 97.1 -163.165 97.5 -162.765 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.2 -163.165 103.6 -162.765 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.3 -163.165 109.7 -162.765 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.4 -163.165 115.8 -162.765 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.5 -163.165 121.9 -162.765 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 11.7 -163.165 12.1 -162.765 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 127.6 -163.165 128 -162.765 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.7 -163.165 134.1 -162.765 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 139.8 -163.165 140.2 -162.765 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 145.9 -163.165 146.3 -162.765 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152 -163.165 152.4 -162.765 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.1 -163.165 158.5 -162.765 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 164.2 -163.165 164.6 -162.765 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 170.3 -163.165 170.7 -162.765 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.4 -163.165 176.8 -162.765 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.5 -163.165 182.9 -162.765 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.8 -163.165 18.2 -162.765 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 188.6 -163.165 189 -162.765 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.7 -163.165 195.1 -162.765 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 23.9 -163.165 24.3 -162.765 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30 -163.165 30.4 -162.765 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.1 -163.165 36.5 -162.765 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 42.2 -163.165 42.6 -162.765 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.3 -163.165 48.7 -162.765 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 54.4 -163.165 54.8 -162.765 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.5 -163.165 60.9 -162.765 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4 -163.165 4.4 -162.765 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65 -163.165 65.4 -162.765 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.1 -163.165 71.5 -162.765 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.2 -163.165 77.6 -162.765 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.3 -163.165 83.7 -162.765 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.4 -163.165 89.8 -162.765 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.5 -163.165 95.9 -162.765 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.6 -163.165 102 -162.765 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.7 -163.165 108.1 -162.765 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.8 -163.165 114.2 -162.765 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.9 -163.165 120.3 -162.765 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 10.1 -163.165 10.5 -162.765 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126 -163.165 126.4 -162.765 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.1 -163.165 132.5 -162.765 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.2 -163.165 138.6 -162.765 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 144.3 -163.165 144.7 -162.765 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 150.4 -163.165 150.8 -162.765 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.5 -163.165 156.9 -162.765 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 162.6 -163.165 163 -162.765 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 168.7 -163.165 169.1 -162.765 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 174.8 -163.165 175.2 -162.765 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 180.9 -163.165 181.3 -162.765 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.2 -163.165 16.6 -162.765 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 187 -163.165 187.4 -162.765 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.1 -163.165 193.5 -162.765 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.3 -163.165 22.7 -162.765 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.4 -163.165 28.8 -162.765 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 34.5 -163.165 34.9 -162.765 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 40.6 -163.165 41 -162.765 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.7 -163.165 47.1 -162.765 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.8 -163.165 53.2 -162.765 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.9 -163.165 59.3 -162.765 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -15.12 -163.165 -14.8 -162.845 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.4 -163.165 6.8 -162.765 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.2 -163.165 55.6 -162.765 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 104 -163.165 104.4 -162.765 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.8 -163.165 153.2 -162.765 ;
    END
  END wmask[3]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -73.425 -163.165 212.825 131.35 ;
    LAYER met2 SPACING 0.14 ;
      RECT -73.425 -163.165 212.825 131.35 ;
    LAYER met3 SPACING 0.3 ;
      RECT 0.515 -35.525 0.845 -35.195 ;
      RECT 0.52 -47.085 0.84 -35.195 ;
      RECT 0.515 -47.085 0.845 -46.755 ;
      RECT -0.165 -34.165 0.165 -33.835 ;
      RECT -0.16 -47.765 0.16 -33.835 ;
      RECT -0.165 -47.765 0.165 -47.435 ;
      RECT -8.325 -39.605 -7.995 -39.275 ;
      RECT -8.32 -100.125 -8 -39.275 ;
      RECT -8.325 -100.125 -7.995 -99.795 ;
      RECT -9.005 -86.525 -8.675 -86.195 ;
      RECT -9 -137.525 -8.68 -86.195 ;
      RECT -9.005 -137.525 -8.675 -137.195 ;
      RECT -9.005 -20.565 -8.675 -20.235 ;
      RECT -9 -81.085 -8.68 -20.235 ;
      RECT -9.005 -81.085 -8.675 -80.755 ;
      RECT -9.685 -137.525 -9.355 -137.195 ;
      RECT -9.68 -162.355 -9.36 -137.195 ;
      RECT -9.685 -151.125 -9.355 -150.795 ;
      RECT -10.365 -147.045 -10.035 -146.715 ;
      RECT -10.36 -151.805 -10.04 -146.715 ;
      RECT -10.365 -151.805 -10.035 -151.475 ;
      RECT -11.045 -11.045 -10.715 -10.715 ;
      RECT -11.04 -100.805 -10.72 -10.715 ;
      RECT -11.045 -100.805 -10.715 -100.475 ;
      RECT -11.725 -18.525 -11.395 -18.195 ;
      RECT -11.72 -87.885 -11.4 -18.195 ;
      RECT -11.725 -87.885 -11.395 -87.555 ;
      RECT -12.405 -10.365 -12.075 -10.035 ;
      RECT -12.4 -23.285 -12.08 -10.035 ;
      RECT -12.405 -23.285 -12.075 -22.955 ;
      RECT -13.085 -19.205 -12.755 -18.875 ;
      RECT -13.08 -80.405 -12.76 -18.875 ;
      RECT -13.085 -80.405 -12.755 -80.075 ;
      RECT -13.765 -89.69 -13.435 -89.36 ;
      RECT -13.76 -91.965 -13.44 -89.36 ;
      RECT -13.765 -91.965 -13.435 -91.635 ;
      RECT -14.445 -90.17 -14.115 -89.84 ;
      RECT -14.44 -92.645 -14.12 -89.84 ;
      RECT -14.445 -92.645 -14.115 -92.315 ;
      RECT -15.125 -152.485 -14.795 -152.155 ;
      RECT -15.12 -162.355 -14.8 -152.155 ;
      RECT -15.125 -90.65 -14.795 -90.32 ;
      RECT -15.12 -151.805 -14.8 -90.32 ;
      RECT -15.125 -151.805 -14.795 -151.475 ;
      RECT -15.805 -91.13 -15.475 -90.8 ;
      RECT -15.8 -93.325 -15.48 -90.8 ;
      RECT -15.805 -93.325 -15.475 -92.995 ;
      RECT -16.485 -32.805 -16.155 -32.475 ;
      RECT -16.48 -98.085 -16.16 -32.475 ;
      RECT -16.485 -98.085 -16.155 -97.755 ;
      RECT -16.485 -9.685 -16.155 -9.355 ;
      RECT -16.48 -23.285 -16.16 -9.355 ;
      RECT -16.485 -23.285 -16.155 -22.955 ;
      RECT -17.165 -93.325 -16.835 -92.995 ;
      RECT -17.16 -153.165 -16.84 -92.995 ;
      RECT -17.165 -153.165 -16.835 -152.835 ;
      RECT -17.165 -9.005 -16.835 -8.675 ;
      RECT -17.16 -23.285 -16.84 -8.675 ;
      RECT -17.165 -23.285 -16.835 -22.955 ;
      RECT -17.845 -42.93 -17.515 -42.6 ;
      RECT -17.84 -46.405 -17.52 -42.6 ;
      RECT -17.845 -46.405 -17.515 -46.075 ;
      RECT -17.845 -19.95 -17.515 -19.62 ;
      RECT -17.84 -23.285 -17.52 -19.62 ;
      RECT -17.845 -23.285 -17.515 -22.955 ;
      RECT -18.525 -43.41 -18.195 -43.08 ;
      RECT -18.52 -47.085 -18.2 -43.08 ;
      RECT -18.525 -47.085 -18.195 -46.755 ;
      RECT -18.525 -20.43 -18.195 -20.1 ;
      RECT -18.52 -23.965 -18.2 -20.1 ;
      RECT -18.525 -23.965 -18.195 -23.635 ;
      RECT -19.205 -43.89 -18.875 -43.56 ;
      RECT -19.2 -47.765 -18.88 -43.56 ;
      RECT -19.205 -47.765 -18.875 -47.435 ;
      RECT -19.205 -20.91 -18.875 -20.58 ;
      RECT -19.2 -24.645 -18.88 -20.58 ;
      RECT -19.205 -24.645 -18.875 -24.315 ;
      RECT -19.885 -44.37 -19.555 -44.04 ;
      RECT -19.88 -48.445 -19.56 -44.04 ;
      RECT -19.885 -48.445 -19.555 -48.115 ;
      RECT -19.885 -21.39 -19.555 -21.06 ;
      RECT -19.88 -25.325 -19.56 -21.06 ;
      RECT -19.885 -25.325 -19.555 -24.995 ;
      RECT -20.565 -68.165 -20.235 -67.835 ;
      RECT -20.56 -98.765 -20.24 -67.835 ;
      RECT -20.565 -98.765 -20.235 -98.435 ;
      RECT -20.565 -44.85 -20.235 -44.52 ;
      RECT -20.56 -49.125 -20.24 -44.52 ;
      RECT -20.565 -49.125 -20.235 -48.795 ;
      RECT -20.565 -21.87 -20.235 -21.54 ;
      RECT -20.56 -26.005 -20.24 -21.54 ;
      RECT -20.565 -26.005 -20.235 -25.675 ;
      RECT -21.245 -152.485 -20.915 -152.155 ;
      RECT -21.24 -162.355 -20.92 -152.155 ;
      RECT -21.245 -91.965 -20.915 -91.635 ;
      RECT -21.24 -151.805 -20.92 -91.635 ;
      RECT -21.245 -151.805 -20.915 -151.475 ;
      RECT -21.245 -45.33 -20.915 -45 ;
      RECT -21.24 -49.805 -20.92 -45 ;
      RECT -21.245 -49.805 -20.915 -49.475 ;
      RECT -21.245 -22.35 -20.915 -22.02 ;
      RECT -21.24 -26.685 -20.92 -22.02 ;
      RECT -21.245 -26.685 -20.915 -26.355 ;
      RECT -21.925 -6.965 -21.595 -6.635 ;
      RECT -21.92 -27.365 -21.6 -6.635 ;
      RECT -21.925 -27.365 -21.595 -27.035 ;
      RECT -23.285 -92.645 -22.955 -92.315 ;
      RECT -23.28 -153.165 -22.96 -92.315 ;
      RECT -23.285 -153.165 -22.955 -152.835 ;
      RECT -26.685 -6.285 -26.355 -5.955 ;
      RECT -26.68 -27.365 -26.36 -5.955 ;
      RECT -26.685 -27.365 -26.355 -27.035 ;
      RECT -27.365 -152.485 -27.035 -152.155 ;
      RECT -27.36 -162.355 -27.04 -152.155 ;
      RECT -28.725 -91.965 -28.395 -91.635 ;
      RECT -28.72 -151.805 -28.4 -91.635 ;
      RECT -28.725 -151.805 -28.395 -151.475 ;
      RECT -29.405 -92.645 -29.075 -92.315 ;
      RECT -29.4 -153.165 -29.08 -92.315 ;
      RECT -29.405 -153.165 -29.075 -152.835 ;
      RECT -33.485 -152.485 -33.155 -152.155 ;
      RECT -33.48 -162.355 -33.16 -152.155 ;
      RECT -34.165 -91.965 -33.835 -91.635 ;
      RECT -34.16 -153.165 -33.84 -91.635 ;
      RECT -34.165 -153.165 -33.835 -152.835 ;
      RECT -35.525 -91.965 -35.195 -91.635 ;
      RECT -35.52 -151.805 -35.2 -91.635 ;
      RECT -35.525 -151.805 -35.195 -151.475 ;
      RECT -38.925 -91.965 -38.595 -91.635 ;
      RECT -38.92 -153.165 -38.6 -91.635 ;
      RECT -38.925 -153.165 -38.595 -152.835 ;
      RECT -39.605 -152.485 -39.275 -152.155 ;
      RECT -39.6 -162.355 -39.28 -152.155 ;
      RECT -41.645 -91.965 -41.315 -91.635 ;
      RECT -41.64 -151.805 -41.32 -91.635 ;
      RECT -41.645 -151.805 -41.315 -151.475 ;
      RECT -43.685 -91.965 -43.355 -91.635 ;
      RECT -43.68 -153.165 -43.36 -91.635 ;
      RECT -43.685 -153.165 -43.355 -152.835 ;
      RECT -46.405 -152.485 -46.075 -152.155 ;
      RECT -46.4 -162.355 -46.08 -152.155 ;
      RECT -47.765 -91.965 -47.435 -91.635 ;
      RECT -47.76 -151.805 -47.44 -91.635 ;
      RECT -47.765 -151.805 -47.435 -151.475 ;
      RECT -49.4 60.84 -48.12 61.43 ;
      RECT -48.44 -97.405 -48.12 61.43 ;
      RECT -48.445 -97.405 -48.115 -97.075 ;
      RECT -49.125 -91.965 -48.795 -91.635 ;
      RECT -49.12 -153.165 -48.8 -91.635 ;
      RECT -49.125 -153.165 -48.795 -152.835 ;
      RECT -52.525 -152.485 -52.195 -152.155 ;
      RECT -52.52 -162.355 -52.2 -152.155 ;
      RECT -53.885 -93.325 -53.555 -92.995 ;
      RECT -53.88 -151.805 -53.56 -92.995 ;
      RECT -53.885 -151.805 -53.555 -151.475 ;
      RECT -55.245 37.915 -54.915 38.245 ;
      RECT -55.24 -11.045 -54.92 38.245 ;
      RECT -55.245 -11.045 -54.915 -10.715 ;
      RECT -55.925 37.235 -55.595 37.565 ;
      RECT -55.92 -100.805 -55.6 37.565 ;
      RECT -55.925 -100.805 -55.595 -100.475 ;
      RECT -56.605 -91.285 -56.275 -90.955 ;
      RECT -56.6 -99.445 -56.28 -90.955 ;
      RECT -56.605 -99.445 -56.275 -99.115 ;
      RECT -58.645 -152.485 -58.315 -152.155 ;
      RECT -58.64 -162.355 -58.32 -152.155 ;
      RECT -60.005 -91.965 -59.675 -91.635 ;
      RECT -60 -151.805 -59.68 -91.635 ;
      RECT -60.005 -151.805 -59.675 -151.475 ;
      RECT -60.685 -92.645 -60.355 -92.315 ;
      RECT -60.68 -153.165 -60.36 -92.315 ;
      RECT -60.685 -153.165 -60.355 -152.835 ;
      RECT -64.765 -152.485 -64.435 -152.155 ;
      RECT -64.76 -162.355 -64.44 -152.155 ;
      RECT 196.3 -80.215 196.7 -20.12 ;
      RECT 195.5 -79.355 195.9 -20.12 ;
      RECT 194.7 -162.275 195.1 -79.445 ;
      RECT 193.9 -63.5 194.3 -48.905 ;
      RECT 193.9 -45.08 194.3 -15.74 ;
      RECT 193.1 -162.275 193.5 -73.605 ;
      RECT 193.1 -64 193.5 -49.36 ;
      RECT 193.1 -45.51 193.5 -12.47 ;
      RECT 190.2 -80.215 190.6 -20.12 ;
      RECT 189.4 -79.355 189.8 -20.12 ;
      RECT 188.6 -162.275 189 -79.445 ;
      RECT 187.8 -63.5 188.2 -48.905 ;
      RECT 187.8 -45.08 188.2 -15.74 ;
      RECT 187 -162.275 187.4 -73.605 ;
      RECT 187 -64 187.4 -49.36 ;
      RECT 187 -45.51 187.4 -12.47 ;
      RECT 184.1 -80.215 184.5 -20.12 ;
      RECT 183.3 -79.355 183.7 -20.12 ;
      RECT 182.5 -162.275 182.9 -79.445 ;
      RECT 181.7 -63.5 182.1 -48.905 ;
      RECT 181.7 -45.08 182.1 -15.74 ;
      RECT 180.9 -162.275 181.3 -73.605 ;
      RECT 180.9 -64 181.3 -49.36 ;
      RECT 180.9 -45.51 181.3 -12.47 ;
      RECT 178 -80.215 178.4 -20.12 ;
      RECT 177.2 -79.355 177.6 -20.12 ;
      RECT 176.4 -162.275 176.8 -79.445 ;
      RECT 175.6 -63.5 176 -48.905 ;
      RECT 175.6 -45.08 176 -15.74 ;
      RECT 174.8 -162.275 175.2 -73.605 ;
      RECT 174.8 -64 175.2 -49.36 ;
      RECT 174.8 -45.51 175.2 -12.47 ;
      RECT 171.9 -80.215 172.3 -20.12 ;
      RECT 171.1 -79.355 171.5 -20.12 ;
      RECT 170.3 -162.275 170.7 -79.445 ;
      RECT 169.5 -63.5 169.9 -48.905 ;
      RECT 169.5 -45.08 169.9 -15.74 ;
      RECT 168.7 -162.275 169.1 -73.605 ;
      RECT 168.7 -64 169.1 -49.36 ;
      RECT 168.7 -45.51 169.1 -12.47 ;
      RECT 165.8 -80.215 166.2 -20.12 ;
      RECT 165 -79.355 165.4 -20.12 ;
      RECT 164.2 -162.275 164.6 -79.445 ;
      RECT 163.4 -63.5 163.8 -48.905 ;
      RECT 163.4 -45.08 163.8 -15.74 ;
      RECT 162.6 -162.275 163 -73.605 ;
      RECT 162.6 -64 163 -49.36 ;
      RECT 162.6 -45.51 163 -12.47 ;
      RECT 159.7 -80.215 160.1 -20.12 ;
      RECT 158.9 -79.355 159.3 -20.12 ;
      RECT 158.1 -162.275 158.5 -79.445 ;
      RECT 157.3 -63.5 157.7 -48.905 ;
      RECT 157.3 -45.08 157.7 -15.74 ;
      RECT 156.5 -162.275 156.9 -73.605 ;
      RECT 156.5 -64 156.9 -49.36 ;
      RECT 156.5 -45.51 156.9 -12.47 ;
      RECT 154.4 -87.06 154.8 -20.12 ;
      RECT 153.6 -80.215 154 -20.12 ;
      RECT 152.8 -162.275 153.2 -87.15 ;
      RECT 152.8 -79.355 153.2 -20.12 ;
      RECT 152 -162.275 152.4 -79.445 ;
      RECT 151.2 -63.5 151.6 -48.905 ;
      RECT 151.2 -45.08 151.6 -15.74 ;
      RECT 150.4 -162.275 150.8 -73.605 ;
      RECT 150.4 -64 150.8 -49.36 ;
      RECT 150.4 -45.51 150.8 -12.47 ;
      RECT 147.5 -80.215 147.9 -20.12 ;
      RECT 146.7 -79.355 147.1 -20.12 ;
      RECT 145.9 -162.275 146.3 -79.445 ;
      RECT 145.1 -63.5 145.5 -48.905 ;
      RECT 145.1 -45.08 145.5 -15.74 ;
      RECT 144.3 -162.275 144.7 -73.605 ;
      RECT 144.3 -64 144.7 -49.36 ;
      RECT 144.3 -45.51 144.7 -12.47 ;
      RECT 141.4 -80.215 141.8 -20.12 ;
      RECT 140.6 -79.355 141 -20.12 ;
      RECT 139.8 -162.275 140.2 -79.445 ;
      RECT 139 -63.5 139.4 -48.905 ;
      RECT 139 -45.08 139.4 -15.74 ;
      RECT 138.2 -162.275 138.6 -73.605 ;
      RECT 138.2 -64 138.6 -49.36 ;
      RECT 138.2 -45.51 138.6 -12.47 ;
      RECT 135.3 -80.215 135.7 -20.12 ;
      RECT 134.5 -79.355 134.9 -20.12 ;
      RECT 133.7 -162.275 134.1 -79.445 ;
      RECT 132.9 -63.5 133.3 -48.905 ;
      RECT 132.9 -45.08 133.3 -15.74 ;
      RECT 132.1 -162.275 132.5 -73.605 ;
      RECT 132.1 -64 132.5 -49.36 ;
      RECT 132.1 -45.51 132.5 -12.47 ;
      RECT 129.2 -80.215 129.6 -20.12 ;
      RECT 128.4 -79.355 128.8 -20.12 ;
      RECT 127.6 -162.275 128 -79.445 ;
      RECT 126.8 -63.5 127.2 -48.905 ;
      RECT 126.8 -45.08 127.2 -15.74 ;
      RECT 126 -162.275 126.4 -73.605 ;
      RECT 126 -64 126.4 -49.36 ;
      RECT 126 -45.51 126.4 -12.47 ;
      RECT 123.1 -80.215 123.5 -20.12 ;
      RECT 122.3 -79.355 122.7 -20.12 ;
      RECT 121.5 -162.275 121.9 -79.445 ;
      RECT 120.7 -63.5 121.1 -48.905 ;
      RECT 120.7 -45.08 121.1 -15.74 ;
      RECT 119.9 -162.275 120.3 -73.605 ;
      RECT 119.9 -64 120.3 -49.36 ;
      RECT 119.9 -45.51 120.3 -12.47 ;
      RECT 117 -80.215 117.4 -20.12 ;
      RECT 116.2 -79.355 116.6 -20.12 ;
      RECT 115.4 -162.275 115.8 -79.445 ;
      RECT 114.6 -63.5 115 -48.905 ;
      RECT 114.6 -45.08 115 -15.74 ;
      RECT 113.8 -162.275 114.2 -73.605 ;
      RECT 113.8 -64 114.2 -49.36 ;
      RECT 113.8 -45.51 114.2 -12.47 ;
      RECT 110.9 -80.215 111.3 -20.12 ;
      RECT 110.1 -79.355 110.5 -20.12 ;
      RECT 109.3 -162.275 109.7 -79.445 ;
      RECT 108.5 -63.5 108.9 -48.905 ;
      RECT 108.5 -45.08 108.9 -15.74 ;
      RECT 107.7 -162.275 108.1 -73.605 ;
      RECT 107.7 -64 108.1 -49.36 ;
      RECT 107.7 -45.51 108.1 -12.47 ;
      RECT 105.6 -87.06 106 -20.12 ;
      RECT 104.8 -80.215 105.2 -20.12 ;
      RECT 104 -162.275 104.4 -87.15 ;
      RECT 104 -79.355 104.4 -20.12 ;
      RECT 103.2 -162.275 103.6 -79.445 ;
      RECT 102.4 -63.5 102.8 -48.905 ;
      RECT 102.4 -45.08 102.8 -15.74 ;
      RECT 101.6 -162.275 102 -73.605 ;
      RECT 101.6 -64 102 -49.36 ;
      RECT 101.6 -45.51 102 -12.47 ;
      RECT 98.7 -80.215 99.1 -20.12 ;
      RECT 97.9 -79.355 98.3 -20.12 ;
      RECT 97.1 -162.275 97.5 -79.445 ;
      RECT 96.3 -63.5 96.7 -48.905 ;
      RECT 96.3 -45.08 96.7 -15.74 ;
      RECT 95.5 -162.275 95.9 -73.605 ;
      RECT 95.5 -64 95.9 -49.36 ;
      RECT 95.5 -45.51 95.9 -12.47 ;
      RECT 92.6 -80.215 93 -20.12 ;
      RECT 91.8 -79.355 92.2 -20.12 ;
      RECT 91 -162.275 91.4 -79.445 ;
      RECT 90.2 -63.5 90.6 -48.905 ;
      RECT 90.2 -45.08 90.6 -15.74 ;
      RECT 89.4 -162.275 89.8 -73.605 ;
      RECT 89.4 -64 89.8 -49.36 ;
      RECT 89.4 -45.51 89.8 -12.47 ;
      RECT 86.5 -80.215 86.9 -20.12 ;
      RECT 85.7 -79.355 86.1 -20.12 ;
      RECT 84.9 -162.275 85.3 -79.445 ;
      RECT 84.1 -63.5 84.5 -48.905 ;
      RECT 84.1 -45.08 84.5 -15.74 ;
      RECT 83.3 -162.275 83.7 -73.605 ;
      RECT 83.3 -64 83.7 -49.36 ;
      RECT 83.3 -45.51 83.7 -12.47 ;
      RECT 80.4 -80.215 80.8 -20.12 ;
      RECT 79.6 -79.355 80 -20.12 ;
      RECT 78.8 -162.275 79.2 -79.445 ;
      RECT 78 -63.5 78.4 -48.905 ;
      RECT 78 -45.08 78.4 -15.74 ;
      RECT 77.2 -162.275 77.6 -73.605 ;
      RECT 77.2 -64 77.6 -49.36 ;
      RECT 77.2 -45.51 77.6 -12.47 ;
      RECT 74.3 -80.215 74.7 -20.12 ;
      RECT 73.5 -79.355 73.9 -20.12 ;
      RECT 72.7 -162.275 73.1 -79.445 ;
      RECT 71.9 -63.5 72.3 -48.905 ;
      RECT 71.9 -45.08 72.3 -15.74 ;
      RECT 71.1 -162.275 71.5 -73.605 ;
      RECT 71.1 -64 71.5 -49.36 ;
      RECT 71.1 -45.51 71.5 -12.47 ;
      RECT 68.2 -80.215 68.6 -20.12 ;
      RECT 67.4 -79.355 67.8 -20.12 ;
      RECT 66.6 -162.275 67 -79.445 ;
      RECT 65.8 -63.5 66.2 -48.905 ;
      RECT 65.8 -45.08 66.2 -15.74 ;
      RECT 65 -162.275 65.4 -73.605 ;
      RECT 65 -64 65.4 -49.36 ;
      RECT 65 -45.51 65.4 -12.47 ;
      RECT 62.1 -80.215 62.5 -20.12 ;
      RECT 61.3 -79.355 61.7 -20.12 ;
      RECT 60.5 -162.275 60.9 -79.445 ;
      RECT 59.7 -63.5 60.1 -48.905 ;
      RECT 59.7 -45.08 60.1 -15.74 ;
      RECT 58.9 -162.275 59.3 -73.605 ;
      RECT 58.9 -64 59.3 -49.36 ;
      RECT 58.9 -45.51 59.3 -12.47 ;
      RECT 56.8 -87.06 57.2 -20.12 ;
      RECT 56 -80.215 56.4 -20.12 ;
      RECT 55.2 -162.275 55.6 -87.15 ;
      RECT 55.2 -79.355 55.6 -20.12 ;
      RECT 54.4 -162.275 54.8 -79.445 ;
      RECT 53.6 -63.5 54 -48.905 ;
      RECT 53.6 -45.08 54 -15.74 ;
      RECT 52.8 -162.275 53.2 -73.605 ;
      RECT 52.8 -64 53.2 -49.36 ;
      RECT 52.8 -45.51 53.2 -12.47 ;
      RECT 49.9 -80.215 50.3 -20.12 ;
      RECT 49.1 -79.355 49.5 -20.12 ;
      RECT 48.3 -162.275 48.7 -79.445 ;
      RECT 47.5 -63.5 47.9 -48.905 ;
      RECT 47.5 -45.08 47.9 -15.74 ;
      RECT 46.7 -162.275 47.1 -73.605 ;
      RECT 46.7 -64 47.1 -49.36 ;
      RECT 46.7 -45.51 47.1 -12.47 ;
      RECT 43.8 -80.215 44.2 -20.12 ;
      RECT 43 -79.355 43.4 -20.12 ;
      RECT 42.2 -162.275 42.6 -79.445 ;
      RECT 41.4 -63.5 41.8 -48.905 ;
      RECT 41.4 -45.08 41.8 -15.74 ;
      RECT 40.6 -162.275 41 -73.605 ;
      RECT 40.6 -64 41 -49.36 ;
      RECT 40.6 -45.51 41 -12.47 ;
      RECT 37.7 -80.215 38.1 -20.12 ;
      RECT 36.9 -79.355 37.3 -20.12 ;
      RECT 36.1 -162.275 36.5 -79.445 ;
      RECT 35.3 -63.5 35.7 -48.905 ;
      RECT 35.3 -45.08 35.7 -15.74 ;
      RECT 34.5 -162.275 34.9 -73.605 ;
      RECT 34.5 -64 34.9 -49.36 ;
      RECT 34.5 -45.51 34.9 -12.47 ;
      RECT 31.6 -80.215 32 -20.12 ;
      RECT 30.8 -79.355 31.2 -20.12 ;
      RECT 30 -162.275 30.4 -79.445 ;
      RECT 29.2 -63.5 29.6 -48.905 ;
      RECT 29.2 -45.08 29.6 -15.74 ;
      RECT 28.4 -162.275 28.8 -73.605 ;
      RECT 28.4 -64 28.8 -49.36 ;
      RECT 28.4 -45.51 28.8 -12.47 ;
      RECT 25.5 -80.215 25.9 -20.12 ;
      RECT 24.7 -79.355 25.1 -20.12 ;
      RECT 23.9 -162.275 24.3 -79.445 ;
      RECT 23.1 -63.5 23.5 -48.905 ;
      RECT 23.1 -45.08 23.5 -15.74 ;
      RECT 22.3 -162.275 22.7 -73.605 ;
      RECT 22.3 -64 22.7 -49.36 ;
      RECT 22.3 -45.51 22.7 -12.47 ;
      RECT 19.4 -80.215 19.8 -20.12 ;
      RECT 18.6 -79.355 19 -20.12 ;
      RECT 17.8 -162.275 18.2 -79.445 ;
      RECT 17 -63.5 17.4 -48.905 ;
      RECT 17 -45.08 17.4 -15.74 ;
      RECT 16.2 -162.275 16.6 -73.605 ;
      RECT 16.2 -64 16.6 -49.36 ;
      RECT 16.2 -45.51 16.6 -12.47 ;
      RECT 13.3 -80.215 13.7 -20.12 ;
      RECT 12.5 -79.355 12.9 -20.12 ;
      RECT 11.7 -162.275 12.1 -79.445 ;
      RECT 10.9 -63.5 11.3 -48.905 ;
      RECT 10.9 -45.08 11.3 -15.74 ;
      RECT 10.1 -162.275 10.5 -73.605 ;
      RECT 10.1 -64 10.5 -49.36 ;
      RECT 10.1 -45.51 10.5 -12.47 ;
      RECT 8 -87.06 8.4 -20.12 ;
      RECT 7.2 -80.215 7.6 -20.12 ;
      RECT 6.4 -162.275 6.8 -87.15 ;
      RECT 6.4 -79.355 6.8 -20.12 ;
      RECT 5.6 -162.275 6 -79.445 ;
      RECT 4.8 -63.5 5.2 -48.905 ;
      RECT 4.8 -45.08 5.2 -15.74 ;
      RECT 4 -162.275 4.4 -73.605 ;
      RECT 4 -64 4.4 -49.36 ;
      RECT 4 -45.51 4.4 -12.47 ;
  END
END sram22_256x32m4w8

END LIBRARY
