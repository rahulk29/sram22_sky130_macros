VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_512x128m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_512x128m4w8   ;
    SIZE 1206.240 BY 467.760 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 412.510 0.000 412.650 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 418.610 0.000 418.750 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 424.710 0.000 424.850 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 430.810 0.000 430.950 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 436.910 0.000 437.050 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 443.010 0.000 443.150 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 449.110 0.000 449.250 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 455.210 0.000 455.350 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 461.310 0.000 461.450 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 467.410 0.000 467.550 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 473.510 0.000 473.650 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 479.610 0.000 479.750 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 485.710 0.000 485.850 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 491.810 0.000 491.950 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 497.910 0.000 498.050 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 504.010 0.000 504.150 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 510.110 0.000 510.250 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 516.210 0.000 516.350 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 522.310 0.000 522.450 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 528.410 0.000 528.550 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 534.510 0.000 534.650 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 540.610 0.000 540.750 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 546.710 0.000 546.850 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 552.810 0.000 552.950 0.140 ; 
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 558.910 0.000 559.050 0.140 ; 
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 565.010 0.000 565.150 0.140 ; 
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 571.110 0.000 571.250 0.140 ; 
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 577.210 0.000 577.350 0.140 ; 
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 583.310 0.000 583.450 0.140 ; 
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 589.410 0.000 589.550 0.140 ; 
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 595.510 0.000 595.650 0.140 ; 
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 601.610 0.000 601.750 0.140 ; 
        END 
    END dout[31] 
    PIN dout[32] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 607.710 0.000 607.850 0.140 ; 
        END 
    END dout[32] 
    PIN dout[33] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 613.810 0.000 613.950 0.140 ; 
        END 
    END dout[33] 
    PIN dout[34] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 619.910 0.000 620.050 0.140 ; 
        END 
    END dout[34] 
    PIN dout[35] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 626.010 0.000 626.150 0.140 ; 
        END 
    END dout[35] 
    PIN dout[36] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 632.110 0.000 632.250 0.140 ; 
        END 
    END dout[36] 
    PIN dout[37] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 638.210 0.000 638.350 0.140 ; 
        END 
    END dout[37] 
    PIN dout[38] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 644.310 0.000 644.450 0.140 ; 
        END 
    END dout[38] 
    PIN dout[39] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 650.410 0.000 650.550 0.140 ; 
        END 
    END dout[39] 
    PIN dout[40] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 656.510 0.000 656.650 0.140 ; 
        END 
    END dout[40] 
    PIN dout[41] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 662.610 0.000 662.750 0.140 ; 
        END 
    END dout[41] 
    PIN dout[42] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 668.710 0.000 668.850 0.140 ; 
        END 
    END dout[42] 
    PIN dout[43] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 674.810 0.000 674.950 0.140 ; 
        END 
    END dout[43] 
    PIN dout[44] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 680.910 0.000 681.050 0.140 ; 
        END 
    END dout[44] 
    PIN dout[45] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 687.010 0.000 687.150 0.140 ; 
        END 
    END dout[45] 
    PIN dout[46] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 693.110 0.000 693.250 0.140 ; 
        END 
    END dout[46] 
    PIN dout[47] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 699.210 0.000 699.350 0.140 ; 
        END 
    END dout[47] 
    PIN dout[48] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 705.310 0.000 705.450 0.140 ; 
        END 
    END dout[48] 
    PIN dout[49] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 711.410 0.000 711.550 0.140 ; 
        END 
    END dout[49] 
    PIN dout[50] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 717.510 0.000 717.650 0.140 ; 
        END 
    END dout[50] 
    PIN dout[51] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 723.610 0.000 723.750 0.140 ; 
        END 
    END dout[51] 
    PIN dout[52] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 729.710 0.000 729.850 0.140 ; 
        END 
    END dout[52] 
    PIN dout[53] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 735.810 0.000 735.950 0.140 ; 
        END 
    END dout[53] 
    PIN dout[54] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 741.910 0.000 742.050 0.140 ; 
        END 
    END dout[54] 
    PIN dout[55] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 748.010 0.000 748.150 0.140 ; 
        END 
    END dout[55] 
    PIN dout[56] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 754.110 0.000 754.250 0.140 ; 
        END 
    END dout[56] 
    PIN dout[57] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 760.210 0.000 760.350 0.140 ; 
        END 
    END dout[57] 
    PIN dout[58] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 766.310 0.000 766.450 0.140 ; 
        END 
    END dout[58] 
    PIN dout[59] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 772.410 0.000 772.550 0.140 ; 
        END 
    END dout[59] 
    PIN dout[60] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 778.510 0.000 778.650 0.140 ; 
        END 
    END dout[60] 
    PIN dout[61] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 784.610 0.000 784.750 0.140 ; 
        END 
    END dout[61] 
    PIN dout[62] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 790.710 0.000 790.850 0.140 ; 
        END 
    END dout[62] 
    PIN dout[63] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 796.810 0.000 796.950 0.140 ; 
        END 
    END dout[63] 
    PIN dout[64] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 802.910 0.000 803.050 0.140 ; 
        END 
    END dout[64] 
    PIN dout[65] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 809.010 0.000 809.150 0.140 ; 
        END 
    END dout[65] 
    PIN dout[66] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 815.110 0.000 815.250 0.140 ; 
        END 
    END dout[66] 
    PIN dout[67] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 821.210 0.000 821.350 0.140 ; 
        END 
    END dout[67] 
    PIN dout[68] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 827.310 0.000 827.450 0.140 ; 
        END 
    END dout[68] 
    PIN dout[69] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 833.410 0.000 833.550 0.140 ; 
        END 
    END dout[69] 
    PIN dout[70] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 839.510 0.000 839.650 0.140 ; 
        END 
    END dout[70] 
    PIN dout[71] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 845.610 0.000 845.750 0.140 ; 
        END 
    END dout[71] 
    PIN dout[72] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 851.710 0.000 851.850 0.140 ; 
        END 
    END dout[72] 
    PIN dout[73] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 857.810 0.000 857.950 0.140 ; 
        END 
    END dout[73] 
    PIN dout[74] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 863.910 0.000 864.050 0.140 ; 
        END 
    END dout[74] 
    PIN dout[75] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 870.010 0.000 870.150 0.140 ; 
        END 
    END dout[75] 
    PIN dout[76] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 876.110 0.000 876.250 0.140 ; 
        END 
    END dout[76] 
    PIN dout[77] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 882.210 0.000 882.350 0.140 ; 
        END 
    END dout[77] 
    PIN dout[78] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 888.310 0.000 888.450 0.140 ; 
        END 
    END dout[78] 
    PIN dout[79] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 894.410 0.000 894.550 0.140 ; 
        END 
    END dout[79] 
    PIN dout[80] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 900.510 0.000 900.650 0.140 ; 
        END 
    END dout[80] 
    PIN dout[81] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 906.610 0.000 906.750 0.140 ; 
        END 
    END dout[81] 
    PIN dout[82] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 912.710 0.000 912.850 0.140 ; 
        END 
    END dout[82] 
    PIN dout[83] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 918.810 0.000 918.950 0.140 ; 
        END 
    END dout[83] 
    PIN dout[84] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 924.910 0.000 925.050 0.140 ; 
        END 
    END dout[84] 
    PIN dout[85] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 931.010 0.000 931.150 0.140 ; 
        END 
    END dout[85] 
    PIN dout[86] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 937.110 0.000 937.250 0.140 ; 
        END 
    END dout[86] 
    PIN dout[87] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 943.210 0.000 943.350 0.140 ; 
        END 
    END dout[87] 
    PIN dout[88] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 949.310 0.000 949.450 0.140 ; 
        END 
    END dout[88] 
    PIN dout[89] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 955.410 0.000 955.550 0.140 ; 
        END 
    END dout[89] 
    PIN dout[90] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 961.510 0.000 961.650 0.140 ; 
        END 
    END dout[90] 
    PIN dout[91] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 967.610 0.000 967.750 0.140 ; 
        END 
    END dout[91] 
    PIN dout[92] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 973.710 0.000 973.850 0.140 ; 
        END 
    END dout[92] 
    PIN dout[93] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 979.810 0.000 979.950 0.140 ; 
        END 
    END dout[93] 
    PIN dout[94] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 985.910 0.000 986.050 0.140 ; 
        END 
    END dout[94] 
    PIN dout[95] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 992.010 0.000 992.150 0.140 ; 
        END 
    END dout[95] 
    PIN dout[96] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 998.110 0.000 998.250 0.140 ; 
        END 
    END dout[96] 
    PIN dout[97] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1004.210 0.000 1004.350 0.140 ; 
        END 
    END dout[97] 
    PIN dout[98] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1010.310 0.000 1010.450 0.140 ; 
        END 
    END dout[98] 
    PIN dout[99] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1016.410 0.000 1016.550 0.140 ; 
        END 
    END dout[99] 
    PIN dout[100] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1022.510 0.000 1022.650 0.140 ; 
        END 
    END dout[100] 
    PIN dout[101] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1028.610 0.000 1028.750 0.140 ; 
        END 
    END dout[101] 
    PIN dout[102] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1034.710 0.000 1034.850 0.140 ; 
        END 
    END dout[102] 
    PIN dout[103] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1040.810 0.000 1040.950 0.140 ; 
        END 
    END dout[103] 
    PIN dout[104] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1046.910 0.000 1047.050 0.140 ; 
        END 
    END dout[104] 
    PIN dout[105] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1053.010 0.000 1053.150 0.140 ; 
        END 
    END dout[105] 
    PIN dout[106] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1059.110 0.000 1059.250 0.140 ; 
        END 
    END dout[106] 
    PIN dout[107] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1065.210 0.000 1065.350 0.140 ; 
        END 
    END dout[107] 
    PIN dout[108] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1071.310 0.000 1071.450 0.140 ; 
        END 
    END dout[108] 
    PIN dout[109] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1077.410 0.000 1077.550 0.140 ; 
        END 
    END dout[109] 
    PIN dout[110] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1083.510 0.000 1083.650 0.140 ; 
        END 
    END dout[110] 
    PIN dout[111] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1089.610 0.000 1089.750 0.140 ; 
        END 
    END dout[111] 
    PIN dout[112] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1095.710 0.000 1095.850 0.140 ; 
        END 
    END dout[112] 
    PIN dout[113] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1101.810 0.000 1101.950 0.140 ; 
        END 
    END dout[113] 
    PIN dout[114] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1107.910 0.000 1108.050 0.140 ; 
        END 
    END dout[114] 
    PIN dout[115] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1114.010 0.000 1114.150 0.140 ; 
        END 
    END dout[115] 
    PIN dout[116] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1120.110 0.000 1120.250 0.140 ; 
        END 
    END dout[116] 
    PIN dout[117] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1126.210 0.000 1126.350 0.140 ; 
        END 
    END dout[117] 
    PIN dout[118] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1132.310 0.000 1132.450 0.140 ; 
        END 
    END dout[118] 
    PIN dout[119] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1138.410 0.000 1138.550 0.140 ; 
        END 
    END dout[119] 
    PIN dout[120] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1144.510 0.000 1144.650 0.140 ; 
        END 
    END dout[120] 
    PIN dout[121] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1150.610 0.000 1150.750 0.140 ; 
        END 
    END dout[121] 
    PIN dout[122] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1156.710 0.000 1156.850 0.140 ; 
        END 
    END dout[122] 
    PIN dout[123] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1162.810 0.000 1162.950 0.140 ; 
        END 
    END dout[123] 
    PIN dout[124] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1168.910 0.000 1169.050 0.140 ; 
        END 
    END dout[124] 
    PIN dout[125] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1175.010 0.000 1175.150 0.140 ; 
        END 
    END dout[125] 
    PIN dout[126] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1181.110 0.000 1181.250 0.140 ; 
        END 
    END dout[126] 
    PIN dout[127] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1187.210 0.000 1187.350 0.140 ; 
        END 
    END dout[127] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 412.090 0.000 412.230 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 418.190 0.000 418.330 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 424.290 0.000 424.430 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 430.390 0.000 430.530 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 436.490 0.000 436.630 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 442.590 0.000 442.730 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 448.690 0.000 448.830 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 454.790 0.000 454.930 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 460.890 0.000 461.030 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 466.990 0.000 467.130 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 473.090 0.000 473.230 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 479.190 0.000 479.330 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 485.290 0.000 485.430 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 491.390 0.000 491.530 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 497.490 0.000 497.630 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 503.590 0.000 503.730 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 509.690 0.000 509.830 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 515.790 0.000 515.930 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 521.890 0.000 522.030 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 527.990 0.000 528.130 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 534.090 0.000 534.230 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 540.190 0.000 540.330 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 546.290 0.000 546.430 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 552.390 0.000 552.530 0.140 ; 
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 558.490 0.000 558.630 0.140 ; 
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 564.590 0.000 564.730 0.140 ; 
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 570.690 0.000 570.830 0.140 ; 
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 576.790 0.000 576.930 0.140 ; 
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 582.890 0.000 583.030 0.140 ; 
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 588.990 0.000 589.130 0.140 ; 
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 595.090 0.000 595.230 0.140 ; 
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 601.190 0.000 601.330 0.140 ; 
        END 
    END din[31] 
    PIN din[32] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 607.290 0.000 607.430 0.140 ; 
        END 
    END din[32] 
    PIN din[33] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 613.390 0.000 613.530 0.140 ; 
        END 
    END din[33] 
    PIN din[34] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 619.490 0.000 619.630 0.140 ; 
        END 
    END din[34] 
    PIN din[35] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 625.590 0.000 625.730 0.140 ; 
        END 
    END din[35] 
    PIN din[36] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 631.690 0.000 631.830 0.140 ; 
        END 
    END din[36] 
    PIN din[37] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 637.790 0.000 637.930 0.140 ; 
        END 
    END din[37] 
    PIN din[38] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 643.890 0.000 644.030 0.140 ; 
        END 
    END din[38] 
    PIN din[39] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 649.990 0.000 650.130 0.140 ; 
        END 
    END din[39] 
    PIN din[40] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 656.090 0.000 656.230 0.140 ; 
        END 
    END din[40] 
    PIN din[41] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 662.190 0.000 662.330 0.140 ; 
        END 
    END din[41] 
    PIN din[42] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 668.290 0.000 668.430 0.140 ; 
        END 
    END din[42] 
    PIN din[43] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 674.390 0.000 674.530 0.140 ; 
        END 
    END din[43] 
    PIN din[44] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 680.490 0.000 680.630 0.140 ; 
        END 
    END din[44] 
    PIN din[45] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 686.590 0.000 686.730 0.140 ; 
        END 
    END din[45] 
    PIN din[46] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 692.690 0.000 692.830 0.140 ; 
        END 
    END din[46] 
    PIN din[47] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 698.790 0.000 698.930 0.140 ; 
        END 
    END din[47] 
    PIN din[48] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 704.890 0.000 705.030 0.140 ; 
        END 
    END din[48] 
    PIN din[49] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 710.990 0.000 711.130 0.140 ; 
        END 
    END din[49] 
    PIN din[50] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 717.090 0.000 717.230 0.140 ; 
        END 
    END din[50] 
    PIN din[51] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 723.190 0.000 723.330 0.140 ; 
        END 
    END din[51] 
    PIN din[52] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 729.290 0.000 729.430 0.140 ; 
        END 
    END din[52] 
    PIN din[53] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 735.390 0.000 735.530 0.140 ; 
        END 
    END din[53] 
    PIN din[54] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 741.490 0.000 741.630 0.140 ; 
        END 
    END din[54] 
    PIN din[55] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 747.590 0.000 747.730 0.140 ; 
        END 
    END din[55] 
    PIN din[56] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 753.690 0.000 753.830 0.140 ; 
        END 
    END din[56] 
    PIN din[57] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 759.790 0.000 759.930 0.140 ; 
        END 
    END din[57] 
    PIN din[58] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 765.890 0.000 766.030 0.140 ; 
        END 
    END din[58] 
    PIN din[59] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 771.990 0.000 772.130 0.140 ; 
        END 
    END din[59] 
    PIN din[60] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 778.090 0.000 778.230 0.140 ; 
        END 
    END din[60] 
    PIN din[61] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 784.190 0.000 784.330 0.140 ; 
        END 
    END din[61] 
    PIN din[62] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 790.290 0.000 790.430 0.140 ; 
        END 
    END din[62] 
    PIN din[63] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 796.390 0.000 796.530 0.140 ; 
        END 
    END din[63] 
    PIN din[64] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 802.490 0.000 802.630 0.140 ; 
        END 
    END din[64] 
    PIN din[65] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 808.590 0.000 808.730 0.140 ; 
        END 
    END din[65] 
    PIN din[66] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 814.690 0.000 814.830 0.140 ; 
        END 
    END din[66] 
    PIN din[67] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 820.790 0.000 820.930 0.140 ; 
        END 
    END din[67] 
    PIN din[68] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 826.890 0.000 827.030 0.140 ; 
        END 
    END din[68] 
    PIN din[69] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 832.990 0.000 833.130 0.140 ; 
        END 
    END din[69] 
    PIN din[70] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 839.090 0.000 839.230 0.140 ; 
        END 
    END din[70] 
    PIN din[71] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 845.190 0.000 845.330 0.140 ; 
        END 
    END din[71] 
    PIN din[72] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 851.290 0.000 851.430 0.140 ; 
        END 
    END din[72] 
    PIN din[73] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 857.390 0.000 857.530 0.140 ; 
        END 
    END din[73] 
    PIN din[74] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 863.490 0.000 863.630 0.140 ; 
        END 
    END din[74] 
    PIN din[75] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 869.590 0.000 869.730 0.140 ; 
        END 
    END din[75] 
    PIN din[76] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 875.690 0.000 875.830 0.140 ; 
        END 
    END din[76] 
    PIN din[77] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 881.790 0.000 881.930 0.140 ; 
        END 
    END din[77] 
    PIN din[78] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 887.890 0.000 888.030 0.140 ; 
        END 
    END din[78] 
    PIN din[79] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 893.990 0.000 894.130 0.140 ; 
        END 
    END din[79] 
    PIN din[80] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 900.090 0.000 900.230 0.140 ; 
        END 
    END din[80] 
    PIN din[81] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 906.190 0.000 906.330 0.140 ; 
        END 
    END din[81] 
    PIN din[82] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 912.290 0.000 912.430 0.140 ; 
        END 
    END din[82] 
    PIN din[83] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 918.390 0.000 918.530 0.140 ; 
        END 
    END din[83] 
    PIN din[84] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 924.490 0.000 924.630 0.140 ; 
        END 
    END din[84] 
    PIN din[85] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 930.590 0.000 930.730 0.140 ; 
        END 
    END din[85] 
    PIN din[86] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 936.690 0.000 936.830 0.140 ; 
        END 
    END din[86] 
    PIN din[87] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 942.790 0.000 942.930 0.140 ; 
        END 
    END din[87] 
    PIN din[88] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 948.890 0.000 949.030 0.140 ; 
        END 
    END din[88] 
    PIN din[89] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 954.990 0.000 955.130 0.140 ; 
        END 
    END din[89] 
    PIN din[90] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 961.090 0.000 961.230 0.140 ; 
        END 
    END din[90] 
    PIN din[91] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 967.190 0.000 967.330 0.140 ; 
        END 
    END din[91] 
    PIN din[92] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 973.290 0.000 973.430 0.140 ; 
        END 
    END din[92] 
    PIN din[93] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 979.390 0.000 979.530 0.140 ; 
        END 
    END din[93] 
    PIN din[94] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 985.490 0.000 985.630 0.140 ; 
        END 
    END din[94] 
    PIN din[95] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 991.590 0.000 991.730 0.140 ; 
        END 
    END din[95] 
    PIN din[96] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 997.690 0.000 997.830 0.140 ; 
        END 
    END din[96] 
    PIN din[97] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1003.790 0.000 1003.930 0.140 ; 
        END 
    END din[97] 
    PIN din[98] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1009.890 0.000 1010.030 0.140 ; 
        END 
    END din[98] 
    PIN din[99] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1015.990 0.000 1016.130 0.140 ; 
        END 
    END din[99] 
    PIN din[100] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1022.090 0.000 1022.230 0.140 ; 
        END 
    END din[100] 
    PIN din[101] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1028.190 0.000 1028.330 0.140 ; 
        END 
    END din[101] 
    PIN din[102] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1034.290 0.000 1034.430 0.140 ; 
        END 
    END din[102] 
    PIN din[103] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1040.390 0.000 1040.530 0.140 ; 
        END 
    END din[103] 
    PIN din[104] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1046.490 0.000 1046.630 0.140 ; 
        END 
    END din[104] 
    PIN din[105] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1052.590 0.000 1052.730 0.140 ; 
        END 
    END din[105] 
    PIN din[106] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1058.690 0.000 1058.830 0.140 ; 
        END 
    END din[106] 
    PIN din[107] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1064.790 0.000 1064.930 0.140 ; 
        END 
    END din[107] 
    PIN din[108] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1070.890 0.000 1071.030 0.140 ; 
        END 
    END din[108] 
    PIN din[109] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1076.990 0.000 1077.130 0.140 ; 
        END 
    END din[109] 
    PIN din[110] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1083.090 0.000 1083.230 0.140 ; 
        END 
    END din[110] 
    PIN din[111] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1089.190 0.000 1089.330 0.140 ; 
        END 
    END din[111] 
    PIN din[112] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1095.290 0.000 1095.430 0.140 ; 
        END 
    END din[112] 
    PIN din[113] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1101.390 0.000 1101.530 0.140 ; 
        END 
    END din[113] 
    PIN din[114] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1107.490 0.000 1107.630 0.140 ; 
        END 
    END din[114] 
    PIN din[115] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1113.590 0.000 1113.730 0.140 ; 
        END 
    END din[115] 
    PIN din[116] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1119.690 0.000 1119.830 0.140 ; 
        END 
    END din[116] 
    PIN din[117] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1125.790 0.000 1125.930 0.140 ; 
        END 
    END din[117] 
    PIN din[118] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1131.890 0.000 1132.030 0.140 ; 
        END 
    END din[118] 
    PIN din[119] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1137.990 0.000 1138.130 0.140 ; 
        END 
    END din[119] 
    PIN din[120] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1144.090 0.000 1144.230 0.140 ; 
        END 
    END din[120] 
    PIN din[121] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1150.190 0.000 1150.330 0.140 ; 
        END 
    END din[121] 
    PIN din[122] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1156.290 0.000 1156.430 0.140 ; 
        END 
    END din[122] 
    PIN din[123] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1162.390 0.000 1162.530 0.140 ; 
        END 
    END din[123] 
    PIN din[124] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1168.490 0.000 1168.630 0.140 ; 
        END 
    END din[124] 
    PIN din[125] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1174.590 0.000 1174.730 0.140 ; 
        END 
    END din[125] 
    PIN din[126] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1180.690 0.000 1180.830 0.140 ; 
        END 
    END din[126] 
    PIN din[127] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.815400 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1186.790 0.000 1186.930 0.140 ; 
        END 
    END din[127] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 411.740 0.000 411.880 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 460.540 0.000 460.680 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 509.340 0.000 509.480 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 558.140 0.000 558.280 0.140 ; 
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 606.940 0.000 607.080 0.140 ; 
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 655.740 0.000 655.880 0.140 ; 
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 704.540 0.000 704.680 0.140 ; 
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 753.340 0.000 753.480 0.140 ; 
        END 
    END wmask[7] 
    PIN wmask[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 802.140 0.000 802.280 0.140 ; 
        END 
    END wmask[8] 
    PIN wmask[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 850.940 0.000 851.080 0.140 ; 
        END 
    END wmask[9] 
    PIN wmask[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 899.740 0.000 899.880 0.140 ; 
        END 
    END wmask[10] 
    PIN wmask[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 948.540 0.000 948.680 0.140 ; 
        END 
    END wmask[11] 
    PIN wmask[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 997.340 0.000 997.480 0.140 ; 
        END 
    END wmask[12] 
    PIN wmask[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1046.140 0.000 1046.280 0.140 ; 
        END 
    END wmask[13] 
    PIN wmask[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1094.940 0.000 1095.080 0.140 ; 
        END 
    END wmask[14] 
    PIN wmask[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.625800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1143.740 0.000 1143.880 0.140 ; 
        END 
    END wmask[15] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 354.760 0.000 355.080 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 348.640 0.000 348.960 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 342.520 0.000 342.840 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 336.400 0.000 336.720 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 330.280 0.000 330.600 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 324.160 0.000 324.480 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 318.040 0.000 318.360 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 311.920 0.000 312.240 0.320 ; 
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 305.800 0.000 306.120 0.320 ; 
        END 
    END addr[8] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 367.000 0.000 367.320 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.027900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 360.880 0.000 361.200 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 79.515000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 370.400 0.000 370.720 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 83.421000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 371.080 0.000 371.400 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 411.520 6.240 ; 
                RECT 1187.760 5.920 1206.080 6.240 ; 
                RECT 0.160 7.280 1206.080 7.600 ; 
                RECT 0.160 8.640 1206.080 8.960 ; 
                RECT 0.160 10.000 370.040 10.320 ; 
                RECT 1196.600 10.000 1206.080 10.320 ; 
                RECT 0.160 11.360 401.320 11.680 ; 
                RECT 1196.600 11.360 1206.080 11.680 ; 
                RECT 0.160 12.720 401.320 13.040 ; 
                RECT 1196.600 12.720 1206.080 13.040 ; 
                RECT 0.160 14.080 401.320 14.400 ; 
                RECT 1196.600 14.080 1206.080 14.400 ; 
                RECT 0.160 15.440 401.320 15.760 ; 
                RECT 1196.600 15.440 1206.080 15.760 ; 
                RECT 0.160 16.800 401.320 17.120 ; 
                RECT 1196.600 16.800 1206.080 17.120 ; 
                RECT 0.160 18.160 401.320 18.480 ; 
                RECT 1196.600 18.160 1206.080 18.480 ; 
                RECT 0.160 19.520 401.320 19.840 ; 
                RECT 1196.600 19.520 1206.080 19.840 ; 
                RECT 0.160 20.880 302.040 21.200 ; 
                RECT 371.760 20.880 401.320 21.200 ; 
                RECT 1196.600 20.880 1206.080 21.200 ; 
                RECT 0.160 22.240 401.320 22.560 ; 
                RECT 1196.600 22.240 1206.080 22.560 ; 
                RECT 0.160 23.600 401.320 23.920 ; 
                RECT 1196.600 23.600 1206.080 23.920 ; 
                RECT 0.160 24.960 302.040 25.280 ; 
                RECT 371.080 24.960 401.320 25.280 ; 
                RECT 1196.600 24.960 1206.080 25.280 ; 
                RECT 0.160 26.320 401.320 26.640 ; 
                RECT 1196.600 26.320 1206.080 26.640 ; 
                RECT 0.160 27.680 400.640 28.000 ; 
                RECT 1196.600 27.680 1206.080 28.000 ; 
                RECT 0.160 29.040 401.320 29.360 ; 
                RECT 1196.600 29.040 1206.080 29.360 ; 
                RECT 0.160 30.400 401.320 30.720 ; 
                RECT 1196.600 30.400 1206.080 30.720 ; 
                RECT 0.160 31.760 401.320 32.080 ; 
                RECT 1196.600 31.760 1206.080 32.080 ; 
                RECT 0.160 33.120 401.320 33.440 ; 
                RECT 1196.600 33.120 1206.080 33.440 ; 
                RECT 0.160 34.480 401.320 34.800 ; 
                RECT 1196.600 34.480 1206.080 34.800 ; 
                RECT 0.160 35.840 401.320 36.160 ; 
                RECT 1196.600 35.840 1206.080 36.160 ; 
                RECT 0.160 37.200 401.320 37.520 ; 
                RECT 1196.600 37.200 1206.080 37.520 ; 
                RECT 0.160 38.560 401.320 38.880 ; 
                RECT 1196.600 38.560 1206.080 38.880 ; 
                RECT 0.160 39.920 401.320 40.240 ; 
                RECT 1196.600 39.920 1206.080 40.240 ; 
                RECT 0.160 41.280 401.320 41.600 ; 
                RECT 1196.600 41.280 1206.080 41.600 ; 
                RECT 0.160 42.640 200.040 42.960 ; 
                RECT 348.640 42.640 401.320 42.960 ; 
                RECT 1196.600 42.640 1206.080 42.960 ; 
                RECT 0.160 44.000 198.680 44.320 ; 
                RECT 354.760 44.000 401.320 44.320 ; 
                RECT 1196.600 44.000 1206.080 44.320 ; 
                RECT 0.160 45.360 178.960 45.680 ; 
                RECT 371.760 45.360 401.320 45.680 ; 
                RECT 1196.600 45.360 1206.080 45.680 ; 
                RECT 0.160 46.720 178.280 47.040 ; 
                RECT 367.000 46.720 401.320 47.040 ; 
                RECT 1196.600 46.720 1206.080 47.040 ; 
                RECT 0.160 48.080 401.320 48.400 ; 
                RECT 1196.600 48.080 1206.080 48.400 ; 
                RECT 0.160 49.440 338.080 49.760 ; 
                RECT 367.680 49.440 401.320 49.760 ; 
                RECT 1196.600 49.440 1206.080 49.760 ; 
                RECT 0.160 50.800 338.080 51.120 ; 
                RECT 367.680 50.800 401.320 51.120 ; 
                RECT 1196.600 50.800 1206.080 51.120 ; 
                RECT 0.160 52.160 338.080 52.480 ; 
                RECT 1196.600 52.160 1206.080 52.480 ; 
                RECT 0.160 53.520 338.080 53.840 ; 
                RECT 1196.600 53.520 1206.080 53.840 ; 
                RECT 0.160 54.880 197.320 55.200 ; 
                RECT 335.720 54.880 338.080 55.200 ; 
                RECT 367.680 54.880 401.320 55.200 ; 
                RECT 1196.600 54.880 1206.080 55.200 ; 
                RECT 0.160 56.240 401.320 56.560 ; 
                RECT 1196.600 56.240 1206.080 56.560 ; 
                RECT 0.160 57.600 401.320 57.920 ; 
                RECT 1196.600 57.600 1206.080 57.920 ; 
                RECT 0.160 58.960 401.320 59.280 ; 
                RECT 1196.600 58.960 1206.080 59.280 ; 
                RECT 0.160 60.320 401.320 60.640 ; 
                RECT 1196.600 60.320 1206.080 60.640 ; 
                RECT 0.160 61.680 198.680 62.000 ; 
                RECT 204.480 61.680 210.240 62.000 ; 
                RECT 368.360 61.680 401.320 62.000 ; 
                RECT 1196.600 61.680 1206.080 62.000 ; 
                RECT 0.160 63.040 200.040 63.360 ; 
                RECT 203.800 63.040 210.240 63.360 ; 
                RECT 385.360 63.040 401.320 63.360 ; 
                RECT 1196.600 63.040 1206.080 63.360 ; 
                RECT 0.160 64.400 210.240 64.720 ; 
                RECT 385.360 64.400 401.320 64.720 ; 
                RECT 1196.600 64.400 1206.080 64.720 ; 
                RECT 0.160 65.760 210.240 66.080 ; 
                RECT 382.640 65.760 401.320 66.080 ; 
                RECT 1196.600 65.760 1206.080 66.080 ; 
                RECT 0.160 67.120 210.240 67.440 ; 
                RECT 385.360 67.120 401.320 67.440 ; 
                RECT 1196.600 67.120 1206.080 67.440 ; 
                RECT 0.160 68.480 210.240 68.800 ; 
                RECT 385.360 68.480 401.320 68.800 ; 
                RECT 1196.600 68.480 1206.080 68.800 ; 
                RECT 0.160 69.840 210.240 70.160 ; 
                RECT 382.640 69.840 401.320 70.160 ; 
                RECT 1196.600 69.840 1206.080 70.160 ; 
                RECT 0.160 71.200 210.240 71.520 ; 
                RECT 385.360 71.200 401.320 71.520 ; 
                RECT 1196.600 71.200 1206.080 71.520 ; 
                RECT 0.160 72.560 210.240 72.880 ; 
                RECT 382.640 72.560 401.320 72.880 ; 
                RECT 1196.600 72.560 1206.080 72.880 ; 
                RECT 0.160 73.920 210.240 74.240 ; 
                RECT 385.360 73.920 401.320 74.240 ; 
                RECT 1196.600 73.920 1206.080 74.240 ; 
                RECT 0.160 75.280 174.880 75.600 ; 
                RECT 185.440 75.280 210.240 75.600 ; 
                RECT 390.800 75.280 401.320 75.600 ; 
                RECT 1196.600 75.280 1206.080 75.600 ; 
                RECT 0.160 76.640 176.240 76.960 ; 
                RECT 179.320 76.640 210.240 76.960 ; 
                RECT 368.360 76.640 401.320 76.960 ; 
                RECT 1196.600 76.640 1206.080 76.960 ; 
                RECT 0.160 78.000 177.600 78.320 ; 
                RECT 182.040 78.000 189.160 78.320 ; 
                RECT 192.240 78.000 210.240 78.320 ; 
                RECT 388.080 78.000 401.320 78.320 ; 
                RECT 1196.600 78.000 1206.080 78.320 ; 
                RECT 0.160 79.360 210.240 79.680 ; 
                RECT 368.360 79.360 401.320 79.680 ; 
                RECT 1196.600 79.360 1206.080 79.680 ; 
                RECT 0.160 80.720 183.720 81.040 ; 
                RECT 192.240 80.720 210.240 81.040 ; 
                RECT 390.800 80.720 401.320 81.040 ; 
                RECT 1196.600 80.720 1206.080 81.040 ; 
                RECT 0.160 82.080 176.240 82.400 ; 
                RECT 185.440 82.080 210.240 82.400 ; 
                RECT 390.800 82.080 401.320 82.400 ; 
                RECT 1196.600 82.080 1206.080 82.400 ; 
                RECT 0.160 83.440 180.320 83.760 ; 
                RECT 185.440 83.440 210.240 83.760 ; 
                RECT 390.800 83.440 401.320 83.760 ; 
                RECT 1196.600 83.440 1206.080 83.760 ; 
                RECT 0.160 84.800 210.240 85.120 ; 
                RECT 388.080 84.800 401.320 85.120 ; 
                RECT 1196.600 84.800 1206.080 85.120 ; 
                RECT 0.160 86.160 176.240 86.480 ; 
                RECT 178.640 86.160 183.720 86.480 ; 
                RECT 192.920 86.160 210.240 86.480 ; 
                RECT 390.800 86.160 401.320 86.480 ; 
                RECT 1196.600 86.160 1206.080 86.480 ; 
                RECT 0.160 87.520 183.720 87.840 ; 
                RECT 191.560 87.520 210.240 87.840 ; 
                RECT 368.360 87.520 401.320 87.840 ; 
                RECT 1196.600 87.520 1206.080 87.840 ; 
                RECT 0.160 88.880 183.040 89.200 ; 
                RECT 185.440 88.880 210.240 89.200 ; 
                RECT 396.240 88.880 401.320 89.200 ; 
                RECT 1196.600 88.880 1206.080 89.200 ; 
                RECT 0.160 90.240 210.240 90.560 ; 
                RECT 396.240 90.240 401.320 90.560 ; 
                RECT 1196.600 90.240 1206.080 90.560 ; 
                RECT 0.160 91.600 183.720 91.920 ; 
                RECT 192.240 91.600 210.240 91.920 ; 
                RECT 393.520 91.600 401.320 91.920 ; 
                RECT 1196.600 91.600 1206.080 91.920 ; 
                RECT 0.160 92.960 181.000 93.280 ; 
                RECT 185.440 92.960 210.240 93.280 ; 
                RECT 396.240 92.960 401.320 93.280 ; 
                RECT 1196.600 92.960 1206.080 93.280 ; 
                RECT 0.160 94.320 183.040 94.640 ; 
                RECT 185.440 94.320 210.240 94.640 ; 
                RECT 396.240 94.320 401.320 94.640 ; 
                RECT 1196.600 94.320 1206.080 94.640 ; 
                RECT 0.160 95.680 186.440 96.000 ; 
                RECT 197.000 95.680 210.240 96.000 ; 
                RECT 393.520 95.680 401.320 96.000 ; 
                RECT 1196.600 95.680 1206.080 96.000 ; 
                RECT 0.160 97.040 174.200 97.360 ; 
                RECT 192.240 97.040 210.240 97.360 ; 
                RECT 396.240 97.040 401.320 97.360 ; 
                RECT 1196.600 97.040 1206.080 97.360 ; 
                RECT 0.160 98.400 183.040 98.720 ; 
                RECT 185.440 98.400 192.560 98.720 ; 
                RECT 198.360 98.400 210.240 98.720 ; 
                RECT 393.520 98.400 401.320 98.720 ; 
                RECT 1196.600 98.400 1206.080 98.720 ; 
                RECT 0.160 99.760 195.280 100.080 ; 
                RECT 199.040 99.760 210.240 100.080 ; 
                RECT 396.240 99.760 401.320 100.080 ; 
                RECT 1196.600 99.760 1206.080 100.080 ; 
                RECT 0.160 101.120 174.880 101.440 ; 
                RECT 188.160 101.120 210.240 101.440 ; 
                RECT 1196.600 101.120 1206.080 101.440 ; 
                RECT 0.160 102.480 183.720 102.800 ; 
                RECT 192.920 102.480 210.240 102.800 ; 
                RECT 368.360 102.480 401.320 102.800 ; 
                RECT 1196.600 102.480 1206.080 102.800 ; 
                RECT 0.160 103.840 181.000 104.160 ; 
                RECT 192.240 103.840 210.240 104.160 ; 
                RECT 1196.600 103.840 1206.080 104.160 ; 
                RECT 0.160 105.200 210.240 105.520 ; 
                RECT 368.360 105.200 401.320 105.520 ; 
                RECT 1196.600 105.200 1206.080 105.520 ; 
                RECT 0.160 106.560 176.920 106.880 ; 
                RECT 179.320 106.560 210.240 106.880 ; 
                RECT 1196.600 106.560 1206.080 106.880 ; 
                RECT 0.160 107.920 176.240 108.240 ; 
                RECT 185.440 107.920 210.240 108.240 ; 
                RECT 1196.600 107.920 1206.080 108.240 ; 
                RECT 0.160 109.280 210.240 109.600 ; 
                RECT 1196.600 109.280 1206.080 109.600 ; 
                RECT 0.160 110.640 210.240 110.960 ; 
                RECT 1196.600 110.640 1206.080 110.960 ; 
                RECT 0.160 112.000 183.040 112.320 ; 
                RECT 185.440 112.000 210.240 112.320 ; 
                RECT 1196.600 112.000 1206.080 112.320 ; 
                RECT 0.160 113.360 183.720 113.680 ; 
                RECT 186.120 113.360 210.240 113.680 ; 
                RECT 368.360 113.360 401.320 113.680 ; 
                RECT 1196.600 113.360 1206.080 113.680 ; 
                RECT 0.160 114.720 183.040 115.040 ; 
                RECT 185.440 114.720 401.320 115.040 ; 
                RECT 1196.600 114.720 1206.080 115.040 ; 
                RECT 0.160 116.080 401.320 116.400 ; 
                RECT 1196.600 116.080 1206.080 116.400 ; 
                RECT 0.160 117.440 173.520 117.760 ; 
                RECT 185.440 117.440 375.480 117.760 ; 
                RECT 1196.600 117.440 1206.080 117.760 ; 
                RECT 0.160 118.800 183.720 119.120 ; 
                RECT 186.120 118.800 395.880 119.120 ; 
                RECT 1196.600 118.800 1206.080 119.120 ; 
                RECT 0.160 120.160 395.880 120.480 ; 
                RECT 1196.600 120.160 1206.080 120.480 ; 
                RECT 0.160 121.520 390.440 121.840 ; 
                RECT 1196.600 121.520 1206.080 121.840 ; 
                RECT 0.160 122.880 170.800 123.200 ; 
                RECT 184.760 122.880 390.440 123.200 ; 
                RECT 1196.600 122.880 1206.080 123.200 ; 
                RECT 0.160 124.240 176.240 124.560 ; 
                RECT 192.240 124.240 385.000 124.560 ; 
                RECT 1196.600 124.240 1206.080 124.560 ; 
                RECT 0.160 125.600 189.840 125.920 ; 
                RECT 192.240 125.600 385.000 125.920 ; 
                RECT 1196.600 125.600 1206.080 125.920 ; 
                RECT 0.160 126.960 379.560 127.280 ; 
                RECT 1196.600 126.960 1206.080 127.280 ; 
                RECT 0.160 128.320 176.240 128.640 ; 
                RECT 194.280 128.320 379.560 128.640 ; 
                RECT 1196.600 128.320 1206.080 128.640 ; 
                RECT 0.160 129.680 379.560 130.000 ; 
                RECT 1196.600 129.680 1206.080 130.000 ; 
                RECT 0.160 131.040 401.320 131.360 ; 
                RECT 1196.600 131.040 1206.080 131.360 ; 
                RECT 0.160 132.400 401.320 132.720 ; 
                RECT 1196.600 132.400 1206.080 132.720 ; 
                RECT 0.160 133.760 174.200 134.080 ; 
                RECT 177.960 133.760 401.320 134.080 ; 
                RECT 1196.600 133.760 1206.080 134.080 ; 
                RECT 0.160 135.120 174.880 135.440 ; 
                RECT 182.040 135.120 401.320 135.440 ; 
                RECT 1196.600 135.120 1206.080 135.440 ; 
                RECT 0.160 136.480 179.640 136.800 ; 
                RECT 192.240 136.480 401.320 136.800 ; 
                RECT 1196.600 136.480 1206.080 136.800 ; 
                RECT 0.160 137.840 401.320 138.160 ; 
                RECT 1196.600 137.840 1206.080 138.160 ; 
                RECT 0.160 139.200 401.320 139.520 ; 
                RECT 1196.600 139.200 1206.080 139.520 ; 
                RECT 0.160 140.560 153.120 140.880 ; 
                RECT 171.160 140.560 401.320 140.880 ; 
                RECT 1196.600 140.560 1206.080 140.880 ; 
                RECT 0.160 141.920 153.120 142.240 ; 
                RECT 171.160 141.920 176.240 142.240 ; 
                RECT 181.360 141.920 401.320 142.240 ; 
                RECT 1196.600 141.920 1206.080 142.240 ; 
                RECT 0.160 143.280 153.120 143.600 ; 
                RECT 171.160 143.280 401.320 143.600 ; 
                RECT 1196.600 143.280 1206.080 143.600 ; 
                RECT 0.160 144.640 153.120 144.960 ; 
                RECT 171.160 144.640 189.840 144.960 ; 
                RECT 192.240 144.640 401.320 144.960 ; 
                RECT 1196.600 144.640 1206.080 144.960 ; 
                RECT 0.160 146.000 153.120 146.320 ; 
                RECT 171.160 146.000 401.320 146.320 ; 
                RECT 1196.600 146.000 1206.080 146.320 ; 
                RECT 0.160 147.360 153.120 147.680 ; 
                RECT 171.160 147.360 263.280 147.680 ; 
                RECT 368.360 147.360 401.320 147.680 ; 
                RECT 1196.600 147.360 1206.080 147.680 ; 
                RECT 0.160 148.720 153.120 149.040 ; 
                RECT 171.160 148.720 177.600 149.040 ; 
                RECT 179.320 148.720 263.280 149.040 ; 
                RECT 368.360 148.720 401.320 149.040 ; 
                RECT 1196.600 148.720 1206.080 149.040 ; 
                RECT 0.160 150.080 153.120 150.400 ; 
                RECT 171.160 150.080 263.280 150.400 ; 
                RECT 368.360 150.080 401.320 150.400 ; 
                RECT 1196.600 150.080 1206.080 150.400 ; 
                RECT 0.160 151.440 153.120 151.760 ; 
                RECT 171.160 151.440 263.280 151.760 ; 
                RECT 368.360 151.440 401.320 151.760 ; 
                RECT 1196.600 151.440 1206.080 151.760 ; 
                RECT 0.160 152.800 153.120 153.120 ; 
                RECT 171.160 152.800 263.280 153.120 ; 
                RECT 368.360 152.800 401.320 153.120 ; 
                RECT 1196.600 152.800 1206.080 153.120 ; 
                RECT 0.160 154.160 153.120 154.480 ; 
                RECT 171.160 154.160 183.040 154.480 ; 
                RECT 191.560 154.160 263.280 154.480 ; 
                RECT 368.360 154.160 401.320 154.480 ; 
                RECT 1196.600 154.160 1206.080 154.480 ; 
                RECT 0.160 155.520 153.120 155.840 ; 
                RECT 171.160 155.520 263.280 155.840 ; 
                RECT 368.360 155.520 382.280 155.840 ; 
                RECT 1196.600 155.520 1206.080 155.840 ; 
                RECT 0.160 156.880 153.120 157.200 ; 
                RECT 171.160 156.880 263.280 157.200 ; 
                RECT 368.360 156.880 382.280 157.200 ; 
                RECT 1196.600 156.880 1206.080 157.200 ; 
                RECT 0.160 158.240 153.120 158.560 ; 
                RECT 171.160 158.240 263.280 158.560 ; 
                RECT 368.360 158.240 387.720 158.560 ; 
                RECT 1196.600 158.240 1206.080 158.560 ; 
                RECT 0.160 159.600 153.120 159.920 ; 
                RECT 171.840 159.600 387.720 159.920 ; 
                RECT 1196.600 159.600 1206.080 159.920 ; 
                RECT 0.160 160.960 153.120 161.280 ; 
                RECT 171.160 160.960 387.720 161.280 ; 
                RECT 1196.600 160.960 1206.080 161.280 ; 
                RECT 0.160 162.320 153.120 162.640 ; 
                RECT 171.160 162.320 393.160 162.640 ; 
                RECT 1196.600 162.320 1206.080 162.640 ; 
                RECT 0.160 163.680 153.120 164.000 ; 
                RECT 171.160 163.680 263.960 164.000 ; 
                RECT 368.360 163.680 393.160 164.000 ; 
                RECT 1196.600 163.680 1206.080 164.000 ; 
                RECT 0.160 165.040 153.120 165.360 ; 
                RECT 171.160 165.040 263.960 165.360 ; 
                RECT 368.360 165.040 398.600 165.360 ; 
                RECT 1196.600 165.040 1206.080 165.360 ; 
                RECT 0.160 166.400 153.120 166.720 ; 
                RECT 171.160 166.400 263.960 166.720 ; 
                RECT 368.360 166.400 398.600 166.720 ; 
                RECT 1196.600 166.400 1206.080 166.720 ; 
                RECT 0.160 167.760 153.120 168.080 ; 
                RECT 171.160 167.760 263.960 168.080 ; 
                RECT 1196.600 167.760 1206.080 168.080 ; 
                RECT 0.160 169.120 153.120 169.440 ; 
                RECT 171.160 169.120 178.960 169.440 ; 
                RECT 182.040 169.120 263.960 169.440 ; 
                RECT 1196.600 169.120 1206.080 169.440 ; 
                RECT 0.160 170.480 153.120 170.800 ; 
                RECT 171.160 170.480 263.960 170.800 ; 
                RECT 1196.600 170.480 1206.080 170.800 ; 
                RECT 0.160 171.840 153.120 172.160 ; 
                RECT 171.160 171.840 263.960 172.160 ; 
                RECT 1196.600 171.840 1206.080 172.160 ; 
                RECT 0.160 173.200 153.120 173.520 ; 
                RECT 171.160 173.200 263.960 173.520 ; 
                RECT 368.360 173.200 401.320 173.520 ; 
                RECT 1196.600 173.200 1206.080 173.520 ; 
                RECT 0.160 174.560 153.120 174.880 ; 
                RECT 171.160 174.560 263.960 174.880 ; 
                RECT 368.360 174.560 401.320 174.880 ; 
                RECT 1196.600 174.560 1206.080 174.880 ; 
                RECT 0.160 175.920 153.120 176.240 ; 
                RECT 171.160 175.920 263.960 176.240 ; 
                RECT 368.360 175.920 401.320 176.240 ; 
                RECT 1196.600 175.920 1206.080 176.240 ; 
                RECT 0.160 177.280 153.120 177.600 ; 
                RECT 171.160 177.280 263.960 177.600 ; 
                RECT 368.360 177.280 401.320 177.600 ; 
                RECT 1196.600 177.280 1206.080 177.600 ; 
                RECT 0.160 178.640 153.120 178.960 ; 
                RECT 171.160 178.640 263.960 178.960 ; 
                RECT 368.360 178.640 401.320 178.960 ; 
                RECT 1196.600 178.640 1206.080 178.960 ; 
                RECT 0.160 180.000 153.120 180.320 ; 
                RECT 171.160 180.000 176.240 180.320 ; 
                RECT 182.040 180.000 263.960 180.320 ; 
                RECT 368.360 180.000 401.320 180.320 ; 
                RECT 1196.600 180.000 1206.080 180.320 ; 
                RECT 0.160 181.360 263.960 181.680 ; 
                RECT 368.360 181.360 401.320 181.680 ; 
                RECT 1196.600 181.360 1206.080 181.680 ; 
                RECT 0.160 182.720 263.960 183.040 ; 
                RECT 368.360 182.720 401.320 183.040 ; 
                RECT 1196.600 182.720 1206.080 183.040 ; 
                RECT 0.160 184.080 134.080 184.400 ; 
                RECT 152.800 184.080 263.960 184.400 ; 
                RECT 368.360 184.080 401.320 184.400 ; 
                RECT 1196.600 184.080 1206.080 184.400 ; 
                RECT 0.160 185.440 134.080 185.760 ; 
                RECT 152.800 185.440 180.320 185.760 ; 
                RECT 186.120 185.440 263.960 185.760 ; 
                RECT 368.360 185.440 401.320 185.760 ; 
                RECT 1196.600 185.440 1206.080 185.760 ; 
                RECT 0.160 186.800 134.080 187.120 ; 
                RECT 152.800 186.800 159.240 187.120 ; 
                RECT 166.400 186.800 263.960 187.120 ; 
                RECT 1196.600 186.800 1206.080 187.120 ; 
                RECT 0.160 188.160 134.080 188.480 ; 
                RECT 152.800 188.160 153.800 188.480 ; 
                RECT 171.160 188.160 263.960 188.480 ; 
                RECT 1196.600 188.160 1206.080 188.480 ; 
                RECT 0.160 189.520 134.080 189.840 ; 
                RECT 152.800 189.520 263.960 189.840 ; 
                RECT 1196.600 189.520 1206.080 189.840 ; 
                RECT 0.160 190.880 128.640 191.200 ; 
                RECT 166.400 190.880 173.520 191.200 ; 
                RECT 184.760 190.880 263.960 191.200 ; 
                RECT 368.360 190.880 401.320 191.200 ; 
                RECT 1196.600 190.880 1206.080 191.200 ; 
                RECT 0.160 192.240 159.240 192.560 ; 
                RECT 179.320 192.240 1206.080 192.560 ; 
                RECT 0.160 193.600 32.080 193.920 ; 
                RECT 177.960 193.600 1206.080 193.920 ; 
                RECT 0.160 194.960 398.600 195.280 ; 
                RECT 1199.320 194.960 1206.080 195.280 ; 
                RECT 0.160 196.320 398.600 196.640 ; 
                RECT 1199.320 196.320 1206.080 196.640 ; 
                RECT 0.160 197.680 27.320 198.000 ; 
                RECT 33.800 197.680 99.400 198.000 ; 
                RECT 1199.320 197.680 1206.080 198.000 ; 
                RECT 0.160 199.040 25.280 199.360 ; 
                RECT 35.840 199.040 36.840 199.360 ; 
                RECT 48.760 199.040 99.400 199.360 ; 
                RECT 1199.320 199.040 1206.080 199.360 ; 
                RECT 0.160 200.400 25.280 200.720 ; 
                RECT 35.840 200.400 38.200 200.720 ; 
                RECT 47.400 200.400 59.280 200.720 ; 
                RECT 61.000 200.400 75.600 200.720 ; 
                RECT 89.560 200.400 99.400 200.720 ; 
                RECT 1199.320 200.400 1206.080 200.720 ; 
                RECT 0.160 201.760 59.280 202.080 ; 
                RECT 61.000 201.760 75.600 202.080 ; 
                RECT 89.560 201.760 99.400 202.080 ; 
                RECT 1199.320 201.760 1206.080 202.080 ; 
                RECT 0.160 203.120 25.280 203.440 ; 
                RECT 35.840 203.120 59.280 203.440 ; 
                RECT 63.720 203.120 75.600 203.440 ; 
                RECT 89.560 203.120 99.400 203.440 ; 
                RECT 1199.320 203.120 1206.080 203.440 ; 
                RECT 0.160 204.480 25.280 204.800 ; 
                RECT 35.840 204.480 59.280 204.800 ; 
                RECT 64.400 204.480 75.600 204.800 ; 
                RECT 89.560 204.480 99.400 204.800 ; 
                RECT 1199.320 204.480 1206.080 204.800 ; 
                RECT 0.160 205.840 25.280 206.160 ; 
                RECT 35.840 205.840 59.280 206.160 ; 
                RECT 65.080 205.840 75.600 206.160 ; 
                RECT 89.560 205.840 99.400 206.160 ; 
                RECT 1199.320 205.840 1206.080 206.160 ; 
                RECT 0.160 207.200 25.280 207.520 ; 
                RECT 35.840 207.200 99.400 207.520 ; 
                RECT 1199.320 207.200 1206.080 207.520 ; 
                RECT 0.160 208.560 75.600 208.880 ; 
                RECT 89.560 208.560 99.400 208.880 ; 
                RECT 1199.320 208.560 1206.080 208.880 ; 
                RECT 0.160 209.920 75.600 210.240 ; 
                RECT 89.560 209.920 99.400 210.240 ; 
                RECT 1199.320 209.920 1206.080 210.240 ; 
                RECT 0.160 211.280 18.480 211.600 ; 
                RECT 20.880 211.280 75.600 211.600 ; 
                RECT 89.560 211.280 99.400 211.600 ; 
                RECT 1199.320 211.280 1206.080 211.600 ; 
                RECT 0.160 212.640 17.800 212.960 ; 
                RECT 20.880 212.640 75.600 212.960 ; 
                RECT 89.560 212.640 99.400 212.960 ; 
                RECT 1199.320 212.640 1206.080 212.960 ; 
                RECT 0.160 214.000 38.880 214.320 ; 
                RECT 48.760 214.000 75.600 214.320 ; 
                RECT 83.440 214.000 99.400 214.320 ; 
                RECT 1199.320 214.000 1206.080 214.320 ; 
                RECT 0.160 215.360 17.120 215.680 ; 
                RECT 20.880 215.360 34.120 215.680 ; 
                RECT 48.080 215.360 83.760 215.680 ; 
                RECT 89.560 215.360 99.400 215.680 ; 
                RECT 1199.320 215.360 1206.080 215.680 ; 
                RECT 0.160 216.720 16.440 217.040 ; 
                RECT 20.880 216.720 34.120 217.040 ; 
                RECT 39.240 216.720 59.280 217.040 ; 
                RECT 61.680 216.720 75.600 217.040 ; 
                RECT 89.560 216.720 99.400 217.040 ; 
                RECT 1199.320 216.720 1206.080 217.040 ; 
                RECT 0.160 218.080 59.280 218.400 ; 
                RECT 61.680 218.080 75.600 218.400 ; 
                RECT 89.560 218.080 99.400 218.400 ; 
                RECT 1199.320 218.080 1206.080 218.400 ; 
                RECT 0.160 219.440 15.760 219.760 ; 
                RECT 20.880 219.440 34.120 219.760 ; 
                RECT 39.920 219.440 59.280 219.760 ; 
                RECT 62.360 219.440 75.600 219.760 ; 
                RECT 89.560 219.440 99.400 219.760 ; 
                RECT 1199.320 219.440 1206.080 219.760 ; 
                RECT 0.160 220.800 15.080 221.120 ; 
                RECT 20.880 220.800 34.120 221.120 ; 
                RECT 40.600 220.800 59.280 221.120 ; 
                RECT 61.000 220.800 75.600 221.120 ; 
                RECT 89.560 220.800 99.400 221.120 ; 
                RECT 1199.320 220.800 1206.080 221.120 ; 
                RECT 0.160 222.160 14.400 222.480 ; 
                RECT 20.880 222.160 34.120 222.480 ; 
                RECT 41.280 222.160 59.280 222.480 ; 
                RECT 63.040 222.160 75.600 222.480 ; 
                RECT 84.120 222.160 99.400 222.480 ; 
                RECT 1199.320 222.160 1206.080 222.480 ; 
                RECT 0.160 223.520 13.720 223.840 ; 
                RECT 20.880 223.520 75.600 223.840 ; 
                RECT 89.560 223.520 99.400 223.840 ; 
                RECT 1199.320 223.520 1206.080 223.840 ; 
                RECT 0.160 224.880 75.600 225.200 ; 
                RECT 89.560 224.880 99.400 225.200 ; 
                RECT 1199.320 224.880 1206.080 225.200 ; 
                RECT 0.160 226.240 13.040 226.560 ; 
                RECT 20.880 226.240 75.600 226.560 ; 
                RECT 89.560 226.240 99.400 226.560 ; 
                RECT 1199.320 226.240 1206.080 226.560 ; 
                RECT 0.160 227.600 12.360 227.920 ; 
                RECT 20.880 227.600 75.600 227.920 ; 
                RECT 89.560 227.600 99.400 227.920 ; 
                RECT 1199.320 227.600 1206.080 227.920 ; 
                RECT 0.160 228.960 11.680 229.280 ; 
                RECT 20.880 228.960 75.600 229.280 ; 
                RECT 89.560 228.960 99.400 229.280 ; 
                RECT 1199.320 228.960 1206.080 229.280 ; 
                RECT 0.160 230.320 99.400 230.640 ; 
                RECT 1199.320 230.320 1206.080 230.640 ; 
                RECT 0.160 231.680 11.000 232.000 ; 
                RECT 20.880 231.680 34.120 232.000 ; 
                RECT 38.560 231.680 75.600 232.000 ; 
                RECT 89.560 231.680 99.400 232.000 ; 
                RECT 1199.320 231.680 1206.080 232.000 ; 
                RECT 0.160 233.040 10.320 233.360 ; 
                RECT 20.880 233.040 75.600 233.360 ; 
                RECT 89.560 233.040 99.400 233.360 ; 
                RECT 1199.320 233.040 1206.080 233.360 ; 
                RECT 0.160 234.400 75.600 234.720 ; 
                RECT 89.560 234.400 99.400 234.720 ; 
                RECT 1199.320 234.400 1206.080 234.720 ; 
                RECT 0.160 235.760 9.640 236.080 ; 
                RECT 20.880 235.760 34.120 236.080 ; 
                RECT 37.200 235.760 75.600 236.080 ; 
                RECT 89.560 235.760 99.400 236.080 ; 
                RECT 1199.320 235.760 1206.080 236.080 ; 
                RECT 0.160 237.120 75.600 237.440 ; 
                RECT 89.560 237.120 99.400 237.440 ; 
                RECT 1199.320 237.120 1206.080 237.440 ; 
                RECT 0.160 238.480 99.400 238.800 ; 
                RECT 1199.320 238.480 1206.080 238.800 ; 
                RECT 0.160 239.840 75.600 240.160 ; 
                RECT 89.560 239.840 99.400 240.160 ; 
                RECT 1199.320 239.840 1206.080 240.160 ; 
                RECT 0.160 241.200 75.600 241.520 ; 
                RECT 89.560 241.200 99.400 241.520 ; 
                RECT 1199.320 241.200 1206.080 241.520 ; 
                RECT 0.160 242.560 75.600 242.880 ; 
                RECT 89.560 242.560 99.400 242.880 ; 
                RECT 1199.320 242.560 1206.080 242.880 ; 
                RECT 0.160 243.920 75.600 244.240 ; 
                RECT 89.560 243.920 99.400 244.240 ; 
                RECT 1199.320 243.920 1206.080 244.240 ; 
                RECT 0.160 245.280 75.600 245.600 ; 
                RECT 89.560 245.280 99.400 245.600 ; 
                RECT 1199.320 245.280 1206.080 245.600 ; 
                RECT 0.160 246.640 99.400 246.960 ; 
                RECT 1199.320 246.640 1206.080 246.960 ; 
                RECT 0.160 248.000 75.600 248.320 ; 
                RECT 89.560 248.000 99.400 248.320 ; 
                RECT 1199.320 248.000 1206.080 248.320 ; 
                RECT 0.160 249.360 75.600 249.680 ; 
                RECT 89.560 249.360 99.400 249.680 ; 
                RECT 1199.320 249.360 1206.080 249.680 ; 
                RECT 0.160 250.720 75.600 251.040 ; 
                RECT 89.560 250.720 99.400 251.040 ; 
                RECT 1199.320 250.720 1206.080 251.040 ; 
                RECT 0.160 252.080 75.600 252.400 ; 
                RECT 89.560 252.080 99.400 252.400 ; 
                RECT 1199.320 252.080 1206.080 252.400 ; 
                RECT 0.160 253.440 75.600 253.760 ; 
                RECT 88.200 253.440 99.400 253.760 ; 
                RECT 1199.320 253.440 1206.080 253.760 ; 
                RECT 0.160 254.800 85.800 255.120 ; 
                RECT 89.560 254.800 99.400 255.120 ; 
                RECT 1199.320 254.800 1206.080 255.120 ; 
                RECT 0.160 256.160 75.600 256.480 ; 
                RECT 89.560 256.160 99.400 256.480 ; 
                RECT 1199.320 256.160 1206.080 256.480 ; 
                RECT 0.160 257.520 75.600 257.840 ; 
                RECT 89.560 257.520 99.400 257.840 ; 
                RECT 1199.320 257.520 1206.080 257.840 ; 
                RECT 0.160 258.880 75.600 259.200 ; 
                RECT 89.560 258.880 99.400 259.200 ; 
                RECT 1199.320 258.880 1206.080 259.200 ; 
                RECT 0.160 260.240 75.600 260.560 ; 
                RECT 89.560 260.240 99.400 260.560 ; 
                RECT 1199.320 260.240 1206.080 260.560 ; 
                RECT 0.160 261.600 75.600 261.920 ; 
                RECT 88.880 261.600 99.400 261.920 ; 
                RECT 1199.320 261.600 1206.080 261.920 ; 
                RECT 0.160 262.960 80.360 263.280 ; 
                RECT 89.560 262.960 99.400 263.280 ; 
                RECT 1199.320 262.960 1206.080 263.280 ; 
                RECT 0.160 264.320 76.960 264.640 ; 
                RECT 89.560 264.320 99.400 264.640 ; 
                RECT 1199.320 264.320 1206.080 264.640 ; 
                RECT 0.160 265.680 76.960 266.000 ; 
                RECT 89.560 265.680 99.400 266.000 ; 
                RECT 1199.320 265.680 1206.080 266.000 ; 
                RECT 0.160 267.040 76.960 267.360 ; 
                RECT 89.560 267.040 99.400 267.360 ; 
                RECT 1199.320 267.040 1206.080 267.360 ; 
                RECT 0.160 268.400 76.960 268.720 ; 
                RECT 89.560 268.400 99.400 268.720 ; 
                RECT 1199.320 268.400 1206.080 268.720 ; 
                RECT 0.160 269.760 39.560 270.080 ; 
                RECT 65.080 269.760 99.400 270.080 ; 
                RECT 1199.320 269.760 1206.080 270.080 ; 
                RECT 0.160 271.120 38.200 271.440 ; 
                RECT 64.400 271.120 76.960 271.440 ; 
                RECT 89.560 271.120 99.400 271.440 ; 
                RECT 1199.320 271.120 1206.080 271.440 ; 
                RECT 0.160 272.480 36.840 272.800 ; 
                RECT 63.040 272.480 75.600 272.800 ; 
                RECT 89.560 272.480 99.400 272.800 ; 
                RECT 1199.320 272.480 1206.080 272.800 ; 
                RECT 0.160 273.840 75.600 274.160 ; 
                RECT 89.560 273.840 99.400 274.160 ; 
                RECT 1199.320 273.840 1206.080 274.160 ; 
                RECT 0.160 275.200 75.600 275.520 ; 
                RECT 89.560 275.200 99.400 275.520 ; 
                RECT 1199.320 275.200 1206.080 275.520 ; 
                RECT 0.160 276.560 75.600 276.880 ; 
                RECT 89.560 276.560 99.400 276.880 ; 
                RECT 1199.320 276.560 1206.080 276.880 ; 
                RECT 0.160 277.920 99.400 278.240 ; 
                RECT 1199.320 277.920 1206.080 278.240 ; 
                RECT 0.160 279.280 76.960 279.600 ; 
                RECT 89.560 279.280 99.400 279.600 ; 
                RECT 1199.320 279.280 1206.080 279.600 ; 
                RECT 0.160 280.640 75.600 280.960 ; 
                RECT 89.560 280.640 99.400 280.960 ; 
                RECT 1199.320 280.640 1206.080 280.960 ; 
                RECT 0.160 282.000 75.600 282.320 ; 
                RECT 89.560 282.000 99.400 282.320 ; 
                RECT 1199.320 282.000 1206.080 282.320 ; 
                RECT 0.160 283.360 75.600 283.680 ; 
                RECT 89.560 283.360 99.400 283.680 ; 
                RECT 1199.320 283.360 1206.080 283.680 ; 
                RECT 0.160 284.720 75.600 285.040 ; 
                RECT 89.560 284.720 99.400 285.040 ; 
                RECT 1199.320 284.720 1206.080 285.040 ; 
                RECT 0.160 286.080 99.400 286.400 ; 
                RECT 1199.320 286.080 1206.080 286.400 ; 
                RECT 0.160 287.440 75.600 287.760 ; 
                RECT 89.560 287.440 99.400 287.760 ; 
                RECT 1199.320 287.440 1206.080 287.760 ; 
                RECT 0.160 288.800 75.600 289.120 ; 
                RECT 89.560 288.800 99.400 289.120 ; 
                RECT 1199.320 288.800 1206.080 289.120 ; 
                RECT 0.160 290.160 75.600 290.480 ; 
                RECT 89.560 290.160 99.400 290.480 ; 
                RECT 1199.320 290.160 1206.080 290.480 ; 
                RECT 0.160 291.520 75.600 291.840 ; 
                RECT 89.560 291.520 99.400 291.840 ; 
                RECT 1199.320 291.520 1206.080 291.840 ; 
                RECT 0.160 292.880 75.600 293.200 ; 
                RECT 78.680 292.880 99.400 293.200 ; 
                RECT 1199.320 292.880 1206.080 293.200 ; 
                RECT 0.160 294.240 80.360 294.560 ; 
                RECT 89.560 294.240 99.400 294.560 ; 
                RECT 1199.320 294.240 1206.080 294.560 ; 
                RECT 0.160 295.600 75.600 295.920 ; 
                RECT 89.560 295.600 99.400 295.920 ; 
                RECT 1199.320 295.600 1206.080 295.920 ; 
                RECT 0.160 296.960 75.600 297.280 ; 
                RECT 89.560 296.960 99.400 297.280 ; 
                RECT 1199.320 296.960 1206.080 297.280 ; 
                RECT 0.160 298.320 77.640 298.640 ; 
                RECT 89.560 298.320 99.400 298.640 ; 
                RECT 1199.320 298.320 1206.080 298.640 ; 
                RECT 0.160 299.680 75.600 300.000 ; 
                RECT 89.560 299.680 99.400 300.000 ; 
                RECT 1199.320 299.680 1206.080 300.000 ; 
                RECT 0.160 301.040 75.600 301.360 ; 
                RECT 79.360 301.040 99.400 301.360 ; 
                RECT 1199.320 301.040 1206.080 301.360 ; 
                RECT 0.160 302.400 81.720 302.720 ; 
                RECT 89.560 302.400 99.400 302.720 ; 
                RECT 1199.320 302.400 1206.080 302.720 ; 
                RECT 0.160 303.760 75.600 304.080 ; 
                RECT 89.560 303.760 99.400 304.080 ; 
                RECT 1199.320 303.760 1206.080 304.080 ; 
                RECT 0.160 305.120 75.600 305.440 ; 
                RECT 89.560 305.120 99.400 305.440 ; 
                RECT 1199.320 305.120 1206.080 305.440 ; 
                RECT 0.160 306.480 75.600 306.800 ; 
                RECT 89.560 306.480 99.400 306.800 ; 
                RECT 1199.320 306.480 1206.080 306.800 ; 
                RECT 0.160 307.840 75.600 308.160 ; 
                RECT 89.560 307.840 99.400 308.160 ; 
                RECT 1199.320 307.840 1206.080 308.160 ; 
                RECT 0.160 309.200 99.400 309.520 ; 
                RECT 1199.320 309.200 1206.080 309.520 ; 
                RECT 0.160 310.560 77.640 310.880 ; 
                RECT 89.560 310.560 99.400 310.880 ; 
                RECT 1199.320 310.560 1206.080 310.880 ; 
                RECT 0.160 311.920 75.600 312.240 ; 
                RECT 89.560 311.920 99.400 312.240 ; 
                RECT 1199.320 311.920 1206.080 312.240 ; 
                RECT 0.160 313.280 75.600 313.600 ; 
                RECT 89.560 313.280 99.400 313.600 ; 
                RECT 1199.320 313.280 1206.080 313.600 ; 
                RECT 0.160 314.640 75.600 314.960 ; 
                RECT 89.560 314.640 99.400 314.960 ; 
                RECT 1199.320 314.640 1206.080 314.960 ; 
                RECT 0.160 316.000 75.600 316.320 ; 
                RECT 89.560 316.000 99.400 316.320 ; 
                RECT 1199.320 316.000 1206.080 316.320 ; 
                RECT 0.160 317.360 99.400 317.680 ; 
                RECT 1199.320 317.360 1206.080 317.680 ; 
                RECT 0.160 318.720 77.640 319.040 ; 
                RECT 89.560 318.720 99.400 319.040 ; 
                RECT 1199.320 318.720 1206.080 319.040 ; 
                RECT 0.160 320.080 75.600 320.400 ; 
                RECT 89.560 320.080 99.400 320.400 ; 
                RECT 1199.320 320.080 1206.080 320.400 ; 
                RECT 0.160 321.440 75.600 321.760 ; 
                RECT 89.560 321.440 99.400 321.760 ; 
                RECT 1199.320 321.440 1206.080 321.760 ; 
                RECT 0.160 322.800 75.600 323.120 ; 
                RECT 89.560 322.800 99.400 323.120 ; 
                RECT 1199.320 322.800 1206.080 323.120 ; 
                RECT 0.160 324.160 75.600 324.480 ; 
                RECT 89.560 324.160 99.400 324.480 ; 
                RECT 1199.320 324.160 1206.080 324.480 ; 
                RECT 0.160 325.520 99.400 325.840 ; 
                RECT 1199.320 325.520 1206.080 325.840 ; 
                RECT 0.160 326.880 75.600 327.200 ; 
                RECT 89.560 326.880 99.400 327.200 ; 
                RECT 1199.320 326.880 1206.080 327.200 ; 
                RECT 0.160 328.240 75.600 328.560 ; 
                RECT 89.560 328.240 99.400 328.560 ; 
                RECT 1199.320 328.240 1206.080 328.560 ; 
                RECT 0.160 329.600 75.600 329.920 ; 
                RECT 89.560 329.600 99.400 329.920 ; 
                RECT 1199.320 329.600 1206.080 329.920 ; 
                RECT 0.160 330.960 75.600 331.280 ; 
                RECT 89.560 330.960 99.400 331.280 ; 
                RECT 1199.320 330.960 1206.080 331.280 ; 
                RECT 0.160 332.320 75.600 332.640 ; 
                RECT 81.400 332.320 99.400 332.640 ; 
                RECT 1199.320 332.320 1206.080 332.640 ; 
                RECT 0.160 333.680 99.400 334.000 ; 
                RECT 1199.320 333.680 1206.080 334.000 ; 
                RECT 0.160 335.040 78.320 335.360 ; 
                RECT 89.560 335.040 99.400 335.360 ; 
                RECT 1199.320 335.040 1206.080 335.360 ; 
                RECT 0.160 336.400 78.320 336.720 ; 
                RECT 89.560 336.400 99.400 336.720 ; 
                RECT 1199.320 336.400 1206.080 336.720 ; 
                RECT 0.160 337.760 78.320 338.080 ; 
                RECT 89.560 337.760 99.400 338.080 ; 
                RECT 1199.320 337.760 1206.080 338.080 ; 
                RECT 0.160 339.120 78.320 339.440 ; 
                RECT 89.560 339.120 99.400 339.440 ; 
                RECT 1199.320 339.120 1206.080 339.440 ; 
                RECT 0.160 340.480 99.400 340.800 ; 
                RECT 1199.320 340.480 1206.080 340.800 ; 
                RECT 0.160 341.840 83.760 342.160 ; 
                RECT 89.560 341.840 99.400 342.160 ; 
                RECT 1199.320 341.840 1206.080 342.160 ; 
                RECT 0.160 343.200 78.320 343.520 ; 
                RECT 89.560 343.200 99.400 343.520 ; 
                RECT 1199.320 343.200 1206.080 343.520 ; 
                RECT 0.160 344.560 78.320 344.880 ; 
                RECT 89.560 344.560 99.400 344.880 ; 
                RECT 1199.320 344.560 1206.080 344.880 ; 
                RECT 0.160 345.920 78.320 346.240 ; 
                RECT 89.560 345.920 99.400 346.240 ; 
                RECT 1199.320 345.920 1206.080 346.240 ; 
                RECT 0.160 347.280 78.320 347.600 ; 
                RECT 89.560 347.280 99.400 347.600 ; 
                RECT 1199.320 347.280 1206.080 347.600 ; 
                RECT 0.160 348.640 99.400 348.960 ; 
                RECT 1199.320 348.640 1206.080 348.960 ; 
                RECT 0.160 350.000 78.320 350.320 ; 
                RECT 89.560 350.000 99.400 350.320 ; 
                RECT 1199.320 350.000 1206.080 350.320 ; 
                RECT 0.160 351.360 86.480 351.680 ; 
                RECT 89.560 351.360 99.400 351.680 ; 
                RECT 1199.320 351.360 1206.080 351.680 ; 
                RECT 0.160 352.720 78.320 353.040 ; 
                RECT 89.560 352.720 99.400 353.040 ; 
                RECT 1199.320 352.720 1206.080 353.040 ; 
                RECT 0.160 354.080 78.320 354.400 ; 
                RECT 89.560 354.080 99.400 354.400 ; 
                RECT 1199.320 354.080 1206.080 354.400 ; 
                RECT 0.160 355.440 78.320 355.760 ; 
                RECT 89.560 355.440 99.400 355.760 ; 
                RECT 1199.320 355.440 1206.080 355.760 ; 
                RECT 0.160 356.800 99.400 357.120 ; 
                RECT 1199.320 356.800 1206.080 357.120 ; 
                RECT 0.160 358.160 79.000 358.480 ; 
                RECT 89.560 358.160 99.400 358.480 ; 
                RECT 1199.320 358.160 1206.080 358.480 ; 
                RECT 0.160 359.520 79.000 359.840 ; 
                RECT 89.560 359.520 99.400 359.840 ; 
                RECT 1199.320 359.520 1206.080 359.840 ; 
                RECT 0.160 360.880 81.040 361.200 ; 
                RECT 89.560 360.880 99.400 361.200 ; 
                RECT 1199.320 360.880 1206.080 361.200 ; 
                RECT 0.160 362.240 79.000 362.560 ; 
                RECT 89.560 362.240 99.400 362.560 ; 
                RECT 1199.320 362.240 1206.080 362.560 ; 
                RECT 0.160 363.600 79.000 363.920 ; 
                RECT 89.560 363.600 99.400 363.920 ; 
                RECT 1199.320 363.600 1206.080 363.920 ; 
                RECT 0.160 364.960 99.400 365.280 ; 
                RECT 1199.320 364.960 1206.080 365.280 ; 
                RECT 0.160 366.320 79.000 366.640 ; 
                RECT 89.560 366.320 99.400 366.640 ; 
                RECT 1199.320 366.320 1206.080 366.640 ; 
                RECT 0.160 367.680 79.000 368.000 ; 
                RECT 89.560 367.680 99.400 368.000 ; 
                RECT 1199.320 367.680 1206.080 368.000 ; 
                RECT 0.160 369.040 79.000 369.360 ; 
                RECT 89.560 369.040 99.400 369.360 ; 
                RECT 1199.320 369.040 1206.080 369.360 ; 
                RECT 0.160 370.400 83.760 370.720 ; 
                RECT 89.560 370.400 99.400 370.720 ; 
                RECT 1199.320 370.400 1206.080 370.720 ; 
                RECT 0.160 371.760 79.000 372.080 ; 
                RECT 89.560 371.760 99.400 372.080 ; 
                RECT 1199.320 371.760 1206.080 372.080 ; 
                RECT 0.160 373.120 99.400 373.440 ; 
                RECT 1199.320 373.120 1206.080 373.440 ; 
                RECT 0.160 374.480 79.000 374.800 ; 
                RECT 89.560 374.480 99.400 374.800 ; 
                RECT 1199.320 374.480 1206.080 374.800 ; 
                RECT 0.160 375.840 79.000 376.160 ; 
                RECT 89.560 375.840 99.400 376.160 ; 
                RECT 1199.320 375.840 1206.080 376.160 ; 
                RECT 0.160 377.200 79.000 377.520 ; 
                RECT 89.560 377.200 99.400 377.520 ; 
                RECT 1199.320 377.200 1206.080 377.520 ; 
                RECT 0.160 378.560 79.000 378.880 ; 
                RECT 89.560 378.560 99.400 378.880 ; 
                RECT 1199.320 378.560 1206.080 378.880 ; 
                RECT 0.160 379.920 99.400 380.240 ; 
                RECT 1199.320 379.920 1206.080 380.240 ; 
                RECT 0.160 381.280 85.800 381.600 ; 
                RECT 89.560 381.280 99.400 381.600 ; 
                RECT 1199.320 381.280 1206.080 381.600 ; 
                RECT 0.160 382.640 79.000 382.960 ; 
                RECT 89.560 382.640 99.400 382.960 ; 
                RECT 1199.320 382.640 1206.080 382.960 ; 
                RECT 0.160 384.000 79.000 384.320 ; 
                RECT 89.560 384.000 99.400 384.320 ; 
                RECT 1199.320 384.000 1206.080 384.320 ; 
                RECT 0.160 385.360 79.000 385.680 ; 
                RECT 89.560 385.360 99.400 385.680 ; 
                RECT 1199.320 385.360 1206.080 385.680 ; 
                RECT 0.160 386.720 79.000 387.040 ; 
                RECT 89.560 386.720 99.400 387.040 ; 
                RECT 1199.320 386.720 1206.080 387.040 ; 
                RECT 0.160 388.080 99.400 388.400 ; 
                RECT 1199.320 388.080 1206.080 388.400 ; 
                RECT 0.160 389.440 80.360 389.760 ; 
                RECT 89.560 389.440 99.400 389.760 ; 
                RECT 1199.320 389.440 1206.080 389.760 ; 
                RECT 0.160 390.800 80.360 391.120 ; 
                RECT 89.560 390.800 99.400 391.120 ; 
                RECT 1199.320 390.800 1206.080 391.120 ; 
                RECT 0.160 392.160 79.000 392.480 ; 
                RECT 89.560 392.160 99.400 392.480 ; 
                RECT 1199.320 392.160 1206.080 392.480 ; 
                RECT 0.160 393.520 79.000 393.840 ; 
                RECT 89.560 393.520 99.400 393.840 ; 
                RECT 1199.320 393.520 1206.080 393.840 ; 
                RECT 0.160 394.880 79.000 395.200 ; 
                RECT 89.560 394.880 99.400 395.200 ; 
                RECT 1199.320 394.880 1206.080 395.200 ; 
                RECT 0.160 396.240 99.400 396.560 ; 
                RECT 1199.320 396.240 1206.080 396.560 ; 
                RECT 0.160 397.600 79.000 397.920 ; 
                RECT 89.560 397.600 99.400 397.920 ; 
                RECT 1199.320 397.600 1206.080 397.920 ; 
                RECT 0.160 398.960 79.000 399.280 ; 
                RECT 89.560 398.960 99.400 399.280 ; 
                RECT 1199.320 398.960 1206.080 399.280 ; 
                RECT 0.160 400.320 83.080 400.640 ; 
                RECT 89.560 400.320 99.400 400.640 ; 
                RECT 1199.320 400.320 1206.080 400.640 ; 
                RECT 0.160 401.680 79.000 402.000 ; 
                RECT 89.560 401.680 99.400 402.000 ; 
                RECT 1199.320 401.680 1206.080 402.000 ; 
                RECT 0.160 403.040 79.000 403.360 ; 
                RECT 89.560 403.040 99.400 403.360 ; 
                RECT 1199.320 403.040 1206.080 403.360 ; 
                RECT 0.160 404.400 99.400 404.720 ; 
                RECT 1199.320 404.400 1206.080 404.720 ; 
                RECT 0.160 405.760 79.000 406.080 ; 
                RECT 89.560 405.760 99.400 406.080 ; 
                RECT 1199.320 405.760 1206.080 406.080 ; 
                RECT 0.160 407.120 79.000 407.440 ; 
                RECT 89.560 407.120 99.400 407.440 ; 
                RECT 1199.320 407.120 1206.080 407.440 ; 
                RECT 0.160 408.480 79.000 408.800 ; 
                RECT 89.560 408.480 99.400 408.800 ; 
                RECT 1199.320 408.480 1206.080 408.800 ; 
                RECT 0.160 409.840 85.120 410.160 ; 
                RECT 89.560 409.840 99.400 410.160 ; 
                RECT 1199.320 409.840 1206.080 410.160 ; 
                RECT 0.160 411.200 79.000 411.520 ; 
                RECT 89.560 411.200 99.400 411.520 ; 
                RECT 1199.320 411.200 1206.080 411.520 ; 
                RECT 0.160 412.560 99.400 412.880 ; 
                RECT 1199.320 412.560 1206.080 412.880 ; 
                RECT 0.160 413.920 79.000 414.240 ; 
                RECT 89.560 413.920 99.400 414.240 ; 
                RECT 1199.320 413.920 1206.080 414.240 ; 
                RECT 0.160 415.280 79.000 415.600 ; 
                RECT 89.560 415.280 99.400 415.600 ; 
                RECT 1199.320 415.280 1206.080 415.600 ; 
                RECT 0.160 416.640 79.000 416.960 ; 
                RECT 89.560 416.640 99.400 416.960 ; 
                RECT 1199.320 416.640 1206.080 416.960 ; 
                RECT 0.160 418.000 79.000 418.320 ; 
                RECT 89.560 418.000 99.400 418.320 ; 
                RECT 1199.320 418.000 1206.080 418.320 ; 
                RECT 0.160 419.360 99.400 419.680 ; 
                RECT 1199.320 419.360 1206.080 419.680 ; 
                RECT 0.160 420.720 80.360 421.040 ; 
                RECT 89.560 420.720 99.400 421.040 ; 
                RECT 1199.320 420.720 1206.080 421.040 ; 
                RECT 0.160 422.080 79.680 422.400 ; 
                RECT 89.560 422.080 99.400 422.400 ; 
                RECT 1199.320 422.080 1206.080 422.400 ; 
                RECT 0.160 423.440 79.680 423.760 ; 
                RECT 89.560 423.440 99.400 423.760 ; 
                RECT 1199.320 423.440 1206.080 423.760 ; 
                RECT 0.160 424.800 79.680 425.120 ; 
                RECT 89.560 424.800 99.400 425.120 ; 
                RECT 1199.320 424.800 1206.080 425.120 ; 
                RECT 0.160 426.160 79.680 426.480 ; 
                RECT 89.560 426.160 99.400 426.480 ; 
                RECT 1199.320 426.160 1206.080 426.480 ; 
                RECT 0.160 427.520 99.400 427.840 ; 
                RECT 1199.320 427.520 1206.080 427.840 ; 
                RECT 0.160 428.880 81.720 429.200 ; 
                RECT 89.560 428.880 99.400 429.200 ; 
                RECT 1199.320 428.880 1206.080 429.200 ; 
                RECT 0.160 430.240 79.680 430.560 ; 
                RECT 89.560 430.240 99.400 430.560 ; 
                RECT 1199.320 430.240 1206.080 430.560 ; 
                RECT 0.160 431.600 79.680 431.920 ; 
                RECT 89.560 431.600 99.400 431.920 ; 
                RECT 1199.320 431.600 1206.080 431.920 ; 
                RECT 0.160 432.960 79.680 433.280 ; 
                RECT 89.560 432.960 99.400 433.280 ; 
                RECT 1199.320 432.960 1206.080 433.280 ; 
                RECT 0.160 434.320 79.680 434.640 ; 
                RECT 89.560 434.320 99.400 434.640 ; 
                RECT 1199.320 434.320 1206.080 434.640 ; 
                RECT 0.160 435.680 99.400 436.000 ; 
                RECT 1199.320 435.680 1206.080 436.000 ; 
                RECT 0.160 437.040 79.680 437.360 ; 
                RECT 89.560 437.040 99.400 437.360 ; 
                RECT 1199.320 437.040 1206.080 437.360 ; 
                RECT 0.160 438.400 84.440 438.720 ; 
                RECT 89.560 438.400 99.400 438.720 ; 
                RECT 1199.320 438.400 1206.080 438.720 ; 
                RECT 0.160 439.760 85.120 440.080 ; 
                RECT 89.560 439.760 99.400 440.080 ; 
                RECT 1199.320 439.760 1206.080 440.080 ; 
                RECT 0.160 441.120 79.680 441.440 ; 
                RECT 89.560 441.120 99.400 441.440 ; 
                RECT 1199.320 441.120 1206.080 441.440 ; 
                RECT 0.160 442.480 79.680 442.800 ; 
                RECT 89.560 442.480 99.400 442.800 ; 
                RECT 1199.320 442.480 1206.080 442.800 ; 
                RECT 0.160 443.840 99.400 444.160 ; 
                RECT 1199.320 443.840 1206.080 444.160 ; 
                RECT 0.160 445.200 79.680 445.520 ; 
                RECT 89.560 445.200 99.400 445.520 ; 
                RECT 1199.320 445.200 1206.080 445.520 ; 
                RECT 0.160 446.560 79.680 446.880 ; 
                RECT 89.560 446.560 99.400 446.880 ; 
                RECT 1199.320 446.560 1206.080 446.880 ; 
                RECT 0.160 447.920 87.160 448.240 ; 
                RECT 89.560 447.920 99.400 448.240 ; 
                RECT 1199.320 447.920 1206.080 448.240 ; 
                RECT 0.160 449.280 87.160 449.600 ; 
                RECT 89.560 449.280 99.400 449.600 ; 
                RECT 1199.320 449.280 1206.080 449.600 ; 
                RECT 0.160 450.640 79.680 450.960 ; 
                RECT 89.560 450.640 99.400 450.960 ; 
                RECT 1199.320 450.640 1206.080 450.960 ; 
                RECT 0.160 452.000 99.400 452.320 ; 
                RECT 1199.320 452.000 1206.080 452.320 ; 
                RECT 0.160 453.360 398.600 453.680 ; 
                RECT 1199.320 453.360 1206.080 453.680 ; 
                RECT 0.160 454.720 398.600 455.040 ; 
                RECT 1199.320 454.720 1206.080 455.040 ; 
                RECT 0.160 456.080 398.600 456.400 ; 
                RECT 1199.320 456.080 1206.080 456.400 ; 
                RECT 0.160 457.440 1206.080 457.760 ; 
                RECT 0.160 458.800 1206.080 459.120 ; 
                RECT 0.160 460.160 1206.080 460.480 ; 
                RECT 0.160 461.520 1206.080 461.840 ; 
                RECT 0.160 0.160 1206.080 1.520 ; 
                RECT 0.160 466.240 1206.080 467.600 ; 
                RECT 402.740 32.110 408.540 33.480 ; 
                RECT 1189.040 32.110 1194.840 33.480 ; 
                RECT 402.740 37.145 408.540 38.505 ; 
                RECT 1189.040 37.145 1194.840 38.505 ; 
                RECT 402.740 42.210 408.540 43.610 ; 
                RECT 1189.040 42.210 1194.840 43.610 ; 
                RECT 402.740 47.385 408.540 48.825 ; 
                RECT 1189.040 47.385 1194.840 48.825 ; 
                RECT 402.740 52.480 408.540 53.810 ; 
                RECT 1189.040 52.480 1194.840 53.810 ; 
                RECT 402.740 57.410 408.540 58.740 ; 
                RECT 1189.040 57.410 1194.840 58.740 ; 
                RECT 402.740 84.920 1194.840 85.720 ; 
                RECT 402.740 178.865 1194.840 182.465 ; 
                RECT 402.740 95.445 1194.840 99.045 ; 
                RECT 402.740 102.825 1194.840 103.115 ; 
                RECT 402.740 136.325 1194.840 138.125 ; 
                RECT 402.740 80.030 1194.840 80.830 ; 
                RECT 402.740 77.020 1194.840 77.820 ; 
                RECT 402.740 65.550 1194.840 67.350 ; 
                RECT 402.740 16.355 1194.840 18.155 ; 
                RECT 103.900 198.075 105.820 452.455 ; 
                RECT 114.115 198.075 116.035 452.455 ; 
                RECT 117.955 198.075 119.875 452.455 ; 
                RECT 131.010 198.075 132.930 452.455 ; 
                RECT 134.850 198.075 136.770 452.455 ; 
                RECT 138.690 198.075 140.610 452.455 ; 
                RECT 142.530 198.075 144.450 452.455 ; 
                RECT 161.250 198.075 163.170 452.455 ; 
                RECT 165.090 198.075 167.010 452.455 ; 
                RECT 168.930 198.075 170.850 452.455 ; 
                RECT 172.770 198.075 174.690 452.455 ; 
                RECT 176.610 198.075 178.530 452.455 ; 
                RECT 180.450 198.075 182.370 452.455 ; 
                RECT 184.290 198.075 186.210 452.455 ; 
                RECT 213.250 198.075 215.170 452.455 ; 
                RECT 217.090 198.075 219.010 452.455 ; 
                RECT 220.930 198.075 222.850 452.455 ; 
                RECT 224.770 198.075 226.690 452.455 ; 
                RECT 228.610 198.075 230.530 452.455 ; 
                RECT 232.450 198.075 234.370 452.455 ; 
                RECT 236.290 198.075 238.210 452.455 ; 
                RECT 240.130 198.075 242.050 452.455 ; 
                RECT 243.970 198.075 245.890 452.455 ; 
                RECT 247.810 198.075 249.730 452.455 ; 
                RECT 251.650 198.075 253.570 452.455 ; 
                RECT 255.490 198.075 257.410 452.455 ; 
                RECT 259.330 198.075 261.250 452.455 ; 
                RECT 305.315 198.075 307.235 452.455 ; 
                RECT 309.155 198.075 311.075 452.455 ; 
                RECT 312.995 198.075 314.915 452.455 ; 
                RECT 316.835 198.075 318.755 452.455 ; 
                RECT 320.675 198.075 322.595 452.455 ; 
                RECT 324.515 198.075 326.435 452.455 ; 
                RECT 328.355 198.075 330.275 452.455 ; 
                RECT 332.195 198.075 334.115 452.455 ; 
                RECT 336.035 198.075 337.955 452.455 ; 
                RECT 339.875 198.075 341.795 452.455 ; 
                RECT 343.715 198.075 345.635 452.455 ; 
                RECT 347.555 198.075 349.475 452.455 ; 
                RECT 351.395 198.075 353.315 452.455 ; 
                RECT 355.235 198.075 357.155 452.455 ; 
                RECT 359.075 198.075 360.995 452.455 ; 
                RECT 362.915 198.075 364.835 452.455 ; 
                RECT 366.755 198.075 368.675 452.455 ; 
                RECT 370.595 198.075 372.515 452.455 ; 
                RECT 374.435 198.075 376.355 452.455 ; 
                RECT 378.275 198.075 380.195 452.455 ; 
                RECT 382.115 198.075 384.035 452.455 ; 
                RECT 385.955 198.075 387.875 452.455 ; 
                RECT 389.795 198.075 391.715 452.455 ; 
                RECT 393.635 198.075 395.555 452.455 ; 
                RECT 213.305 61.225 215.055 113.825 ; 
                RECT 219.765 61.225 221.685 113.825 ; 
                RECT 226.395 61.225 228.145 113.825 ; 
                RECT 234.575 61.225 236.495 113.825 ; 
                RECT 246.940 61.225 248.860 113.825 ; 
                RECT 250.780 61.225 252.700 113.825 ; 
                RECT 267.950 61.225 269.870 113.825 ; 
                RECT 271.790 61.225 273.710 113.825 ; 
                RECT 275.630 61.225 277.550 113.825 ; 
                RECT 279.470 61.225 281.390 113.825 ; 
                RECT 283.310 61.225 285.230 113.825 ; 
                RECT 287.150 61.225 289.070 113.825 ; 
                RECT 315.895 61.225 317.815 113.825 ; 
                RECT 319.735 61.225 321.655 113.825 ; 
                RECT 323.575 61.225 325.495 113.825 ; 
                RECT 327.415 61.225 329.335 113.825 ; 
                RECT 331.255 61.225 333.175 113.825 ; 
                RECT 335.095 61.225 337.015 113.825 ; 
                RECT 338.935 61.225 340.855 113.825 ; 
                RECT 342.775 61.225 344.695 113.825 ; 
                RECT 346.615 61.225 348.535 113.825 ; 
                RECT 350.455 61.225 352.375 113.825 ; 
                RECT 354.295 61.225 356.215 113.825 ; 
                RECT 358.135 61.225 360.055 113.825 ; 
                RECT 361.975 61.225 363.895 113.825 ; 
                RECT 365.815 61.225 367.735 113.825 ; 
                RECT 268.645 164.320 270.565 191.440 ; 
                RECT 276.135 164.320 277.885 191.440 ; 
                RECT 283.240 164.320 285.160 191.440 ; 
                RECT 295.190 164.320 297.110 191.440 ; 
                RECT 299.030 164.320 300.950 191.440 ; 
                RECT 302.870 164.320 304.790 191.440 ; 
                RECT 327.440 164.320 329.360 191.440 ; 
                RECT 331.280 164.320 333.200 191.440 ; 
                RECT 335.120 164.320 337.040 191.440 ; 
                RECT 338.960 164.320 340.880 191.440 ; 
                RECT 342.800 164.320 344.720 191.440 ; 
                RECT 346.640 164.320 348.560 191.440 ; 
                RECT 350.480 164.320 352.400 191.440 ; 
                RECT 354.320 164.320 356.240 191.440 ; 
                RECT 358.160 164.320 360.080 191.440 ; 
                RECT 362.000 164.320 363.920 191.440 ; 
                RECT 365.840 164.320 367.760 191.440 ; 
                RECT 267.355 147.420 269.275 158.320 ; 
                RECT 274.545 147.420 276.465 158.320 ; 
                RECT 283.240 147.420 285.160 158.320 ; 
                RECT 296.065 147.420 297.985 158.320 ; 
                RECT 299.905 147.420 301.825 158.320 ; 
                RECT 303.745 147.420 305.665 158.320 ; 
                RECT 307.585 147.420 309.505 158.320 ; 
                RECT 330.865 147.420 332.785 158.320 ; 
                RECT 334.705 147.420 336.625 158.320 ; 
                RECT 338.545 147.420 340.465 158.320 ; 
                RECT 342.385 147.420 344.305 158.320 ; 
                RECT 346.225 147.420 348.145 158.320 ; 
                RECT 350.065 147.420 351.985 158.320 ; 
                RECT 353.905 147.420 355.825 158.320 ; 
                RECT 357.745 147.420 359.665 158.320 ; 
                RECT 361.585 147.420 363.505 158.320 ; 
                RECT 365.425 147.420 367.345 158.320 ; 
                RECT 341.720 50.065 343.640 55.225 ; 
                RECT 349.555 50.065 351.475 55.225 ; 
                RECT 361.275 50.065 363.195 55.225 ; 
                RECT 365.115 50.065 367.035 55.225 ; 
                RECT 26.110 200.345 35.270 201.095 ; 
                RECT 26.110 205.100 35.270 207.020 ; 
                RECT 154.180 188.055 170.220 188.905 ; 
                RECT 134.980 188.395 152.220 190.425 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 411.520 5.560 ; 
                RECT 1187.760 5.240 1203.360 5.560 ; 
                RECT 2.880 6.600 1203.360 6.920 ; 
                RECT 2.880 7.960 1203.360 8.280 ; 
                RECT 2.880 9.320 370.720 9.640 ; 
                RECT 407.120 9.320 1203.360 9.640 ; 
                RECT 2.880 10.680 401.320 11.000 ; 
                RECT 1196.600 10.680 1203.360 11.000 ; 
                RECT 2.880 12.040 401.320 12.360 ; 
                RECT 1196.600 12.040 1203.360 12.360 ; 
                RECT 2.880 13.400 401.320 13.720 ; 
                RECT 1196.600 13.400 1203.360 13.720 ; 
                RECT 2.880 14.760 401.320 15.080 ; 
                RECT 1196.600 14.760 1203.360 15.080 ; 
                RECT 2.880 16.120 401.320 16.440 ; 
                RECT 1196.600 16.120 1203.360 16.440 ; 
                RECT 2.880 17.480 401.320 17.800 ; 
                RECT 1196.600 17.480 1203.360 17.800 ; 
                RECT 2.880 18.840 401.320 19.160 ; 
                RECT 1196.600 18.840 1203.360 19.160 ; 
                RECT 2.880 20.200 302.040 20.520 ; 
                RECT 371.760 20.200 401.320 20.520 ; 
                RECT 1196.600 20.200 1203.360 20.520 ; 
                RECT 2.880 21.560 401.320 21.880 ; 
                RECT 1196.600 21.560 1203.360 21.880 ; 
                RECT 2.880 22.920 401.320 23.240 ; 
                RECT 1196.600 22.920 1203.360 23.240 ; 
                RECT 2.880 24.280 302.040 24.600 ; 
                RECT 371.080 24.280 401.320 24.600 ; 
                RECT 1196.600 24.280 1203.360 24.600 ; 
                RECT 2.880 25.640 401.320 25.960 ; 
                RECT 1196.600 25.640 1203.360 25.960 ; 
                RECT 2.880 27.000 401.320 27.320 ; 
                RECT 1196.600 27.000 1203.360 27.320 ; 
                RECT 2.880 28.360 400.640 28.680 ; 
                RECT 1196.600 28.360 1203.360 28.680 ; 
                RECT 2.880 29.720 401.320 30.040 ; 
                RECT 1196.600 29.720 1203.360 30.040 ; 
                RECT 2.880 31.080 401.320 31.400 ; 
                RECT 1196.600 31.080 1203.360 31.400 ; 
                RECT 2.880 32.440 401.320 32.760 ; 
                RECT 1196.600 32.440 1203.360 32.760 ; 
                RECT 2.880 33.800 401.320 34.120 ; 
                RECT 1196.600 33.800 1203.360 34.120 ; 
                RECT 2.880 35.160 401.320 35.480 ; 
                RECT 1196.600 35.160 1203.360 35.480 ; 
                RECT 2.880 36.520 401.320 36.840 ; 
                RECT 1196.600 36.520 1203.360 36.840 ; 
                RECT 2.880 37.880 401.320 38.200 ; 
                RECT 1196.600 37.880 1203.360 38.200 ; 
                RECT 2.880 39.240 401.320 39.560 ; 
                RECT 1196.600 39.240 1203.360 39.560 ; 
                RECT 2.880 40.600 401.320 40.920 ; 
                RECT 1196.600 40.600 1203.360 40.920 ; 
                RECT 2.880 41.960 200.720 42.280 ; 
                RECT 350.000 41.960 401.320 42.280 ; 
                RECT 1196.600 41.960 1203.360 42.280 ; 
                RECT 2.880 43.320 199.360 43.640 ; 
                RECT 356.120 43.320 401.320 43.640 ; 
                RECT 1196.600 43.320 1203.360 43.640 ; 
                RECT 2.880 44.680 176.240 45.000 ; 
                RECT 371.080 44.680 401.320 45.000 ; 
                RECT 1196.600 44.680 1203.360 45.000 ; 
                RECT 2.880 46.040 177.600 46.360 ; 
                RECT 360.880 46.040 401.320 46.360 ; 
                RECT 1196.600 46.040 1203.360 46.360 ; 
                RECT 2.880 47.400 401.320 47.720 ; 
                RECT 1196.600 47.400 1203.360 47.720 ; 
                RECT 2.880 48.760 401.320 49.080 ; 
                RECT 1196.600 48.760 1203.360 49.080 ; 
                RECT 2.880 50.120 338.080 50.440 ; 
                RECT 367.680 50.120 401.320 50.440 ; 
                RECT 1196.600 50.120 1203.360 50.440 ; 
                RECT 2.880 51.480 338.080 51.800 ; 
                RECT 1196.600 51.480 1203.360 51.800 ; 
                RECT 2.880 52.840 338.080 53.160 ; 
                RECT 1196.600 52.840 1203.360 53.160 ; 
                RECT 2.880 54.200 338.080 54.520 ; 
                RECT 367.680 54.200 401.320 54.520 ; 
                RECT 1196.600 54.200 1203.360 54.520 ; 
                RECT 2.880 55.560 338.080 55.880 ; 
                RECT 367.680 55.560 401.320 55.880 ; 
                RECT 1196.600 55.560 1203.360 55.880 ; 
                RECT 2.880 56.920 401.320 57.240 ; 
                RECT 1196.600 56.920 1203.360 57.240 ; 
                RECT 2.880 58.280 401.320 58.600 ; 
                RECT 1196.600 58.280 1203.360 58.600 ; 
                RECT 2.880 59.640 401.320 59.960 ; 
                RECT 1196.600 59.640 1203.360 59.960 ; 
                RECT 2.880 61.000 210.240 61.320 ; 
                RECT 368.360 61.000 401.320 61.320 ; 
                RECT 1196.600 61.000 1203.360 61.320 ; 
                RECT 2.880 62.360 199.360 62.680 ; 
                RECT 204.480 62.360 210.240 62.680 ; 
                RECT 368.360 62.360 401.320 62.680 ; 
                RECT 1196.600 62.360 1203.360 62.680 ; 
                RECT 2.880 63.720 200.720 64.040 ; 
                RECT 203.120 63.720 210.240 64.040 ; 
                RECT 382.640 63.720 401.320 64.040 ; 
                RECT 1196.600 63.720 1203.360 64.040 ; 
                RECT 2.880 65.080 210.240 65.400 ; 
                RECT 385.360 65.080 401.320 65.400 ; 
                RECT 1196.600 65.080 1203.360 65.400 ; 
                RECT 2.880 66.440 210.240 66.760 ; 
                RECT 385.360 66.440 401.320 66.760 ; 
                RECT 1196.600 66.440 1203.360 66.760 ; 
                RECT 2.880 67.800 210.240 68.120 ; 
                RECT 382.640 67.800 401.320 68.120 ; 
                RECT 1196.600 67.800 1203.360 68.120 ; 
                RECT 2.880 69.160 210.240 69.480 ; 
                RECT 385.360 69.160 401.320 69.480 ; 
                RECT 1196.600 69.160 1203.360 69.480 ; 
                RECT 2.880 70.520 210.240 70.840 ; 
                RECT 368.360 70.520 401.320 70.840 ; 
                RECT 1196.600 70.520 1203.360 70.840 ; 
                RECT 2.880 71.880 210.240 72.200 ; 
                RECT 385.360 71.880 401.320 72.200 ; 
                RECT 1196.600 71.880 1203.360 72.200 ; 
                RECT 2.880 73.240 210.240 73.560 ; 
                RECT 385.360 73.240 401.320 73.560 ; 
                RECT 1196.600 73.240 1203.360 73.560 ; 
                RECT 2.880 74.600 210.240 74.920 ; 
                RECT 382.640 74.600 401.320 74.920 ; 
                RECT 1196.600 74.600 1203.360 74.920 ; 
                RECT 2.880 75.960 174.880 76.280 ; 
                RECT 185.440 75.960 210.240 76.280 ; 
                RECT 390.800 75.960 401.320 76.280 ; 
                RECT 1196.600 75.960 1203.360 76.280 ; 
                RECT 2.880 77.320 176.240 77.640 ; 
                RECT 182.040 77.320 189.160 77.640 ; 
                RECT 192.240 77.320 210.240 77.640 ; 
                RECT 390.800 77.320 401.320 77.640 ; 
                RECT 1196.600 77.320 1203.360 77.640 ; 
                RECT 2.880 78.680 177.600 79.000 ; 
                RECT 180.680 78.680 210.240 79.000 ; 
                RECT 368.360 78.680 401.320 79.000 ; 
                RECT 1196.600 78.680 1203.360 79.000 ; 
                RECT 2.880 80.040 183.720 80.360 ; 
                RECT 190.880 80.040 210.240 80.360 ; 
                RECT 390.800 80.040 401.320 80.360 ; 
                RECT 1196.600 80.040 1203.360 80.360 ; 
                RECT 2.880 81.400 178.960 81.720 ; 
                RECT 185.440 81.400 186.440 81.720 ; 
                RECT 192.240 81.400 210.240 81.720 ; 
                RECT 388.080 81.400 401.320 81.720 ; 
                RECT 1196.600 81.400 1203.360 81.720 ; 
                RECT 2.880 82.760 176.240 83.080 ; 
                RECT 185.440 82.760 210.240 83.080 ; 
                RECT 390.800 82.760 401.320 83.080 ; 
                RECT 1196.600 82.760 1203.360 83.080 ; 
                RECT 2.880 84.120 210.240 84.440 ; 
                RECT 390.800 84.120 401.320 84.440 ; 
                RECT 1196.600 84.120 1203.360 84.440 ; 
                RECT 2.880 85.480 176.240 85.800 ; 
                RECT 178.640 85.480 183.720 85.800 ; 
                RECT 192.920 85.480 210.240 85.800 ; 
                RECT 390.800 85.480 401.320 85.800 ; 
                RECT 1196.600 85.480 1203.360 85.800 ; 
                RECT 2.880 86.840 183.720 87.160 ; 
                RECT 191.560 86.840 210.240 87.160 ; 
                RECT 388.080 86.840 401.320 87.160 ; 
                RECT 1196.600 86.840 1203.360 87.160 ; 
                RECT 2.880 88.200 183.040 88.520 ; 
                RECT 185.440 88.200 210.240 88.520 ; 
                RECT 368.360 88.200 401.320 88.520 ; 
                RECT 1196.600 88.200 1203.360 88.520 ; 
                RECT 2.880 89.560 210.240 89.880 ; 
                RECT 393.520 89.560 401.320 89.880 ; 
                RECT 1196.600 89.560 1203.360 89.880 ; 
                RECT 2.880 90.920 183.720 91.240 ; 
                RECT 192.240 90.920 210.240 91.240 ; 
                RECT 396.240 90.920 401.320 91.240 ; 
                RECT 1196.600 90.920 1203.360 91.240 ; 
                RECT 2.880 92.280 181.000 92.600 ; 
                RECT 185.440 92.280 210.240 92.600 ; 
                RECT 396.240 92.280 401.320 92.600 ; 
                RECT 1196.600 92.280 1203.360 92.600 ; 
                RECT 2.880 93.640 183.040 93.960 ; 
                RECT 185.440 93.640 210.240 93.960 ; 
                RECT 393.520 93.640 401.320 93.960 ; 
                RECT 1196.600 93.640 1203.360 93.960 ; 
                RECT 2.880 95.000 210.240 95.320 ; 
                RECT 396.240 95.000 401.320 95.320 ; 
                RECT 1196.600 95.000 1203.360 95.320 ; 
                RECT 2.880 96.360 174.200 96.680 ; 
                RECT 197.000 96.360 210.240 96.680 ; 
                RECT 368.360 96.360 401.320 96.680 ; 
                RECT 1196.600 96.360 1203.360 96.680 ; 
                RECT 2.880 97.720 192.560 98.040 ; 
                RECT 198.360 97.720 210.240 98.040 ; 
                RECT 396.240 97.720 401.320 98.040 ; 
                RECT 1196.600 97.720 1203.360 98.040 ; 
                RECT 2.880 99.080 183.040 99.400 ; 
                RECT 185.440 99.080 195.280 99.400 ; 
                RECT 199.040 99.080 210.240 99.400 ; 
                RECT 396.240 99.080 401.320 99.400 ; 
                RECT 1196.600 99.080 1203.360 99.400 ; 
                RECT 2.880 100.440 174.880 100.760 ; 
                RECT 188.160 100.440 210.240 100.760 ; 
                RECT 393.520 100.440 401.320 100.760 ; 
                RECT 1196.600 100.440 1203.360 100.760 ; 
                RECT 2.880 101.800 183.720 102.120 ; 
                RECT 192.240 101.800 210.240 102.120 ; 
                RECT 1196.600 101.800 1203.360 102.120 ; 
                RECT 2.880 103.160 181.000 103.480 ; 
                RECT 185.440 103.160 187.800 103.480 ; 
                RECT 192.920 103.160 210.240 103.480 ; 
                RECT 1196.600 103.160 1203.360 103.480 ; 
                RECT 2.880 104.520 183.720 104.840 ; 
                RECT 192.240 104.520 210.240 104.840 ; 
                RECT 368.360 104.520 401.320 104.840 ; 
                RECT 1196.600 104.520 1203.360 104.840 ; 
                RECT 2.880 105.880 210.240 106.200 ; 
                RECT 1196.600 105.880 1203.360 106.200 ; 
                RECT 2.880 107.240 176.920 107.560 ; 
                RECT 179.320 107.240 210.240 107.560 ; 
                RECT 368.360 107.240 401.320 107.560 ; 
                RECT 1196.600 107.240 1203.360 107.560 ; 
                RECT 2.880 108.600 176.240 108.920 ; 
                RECT 185.440 108.600 210.240 108.920 ; 
                RECT 1196.600 108.600 1203.360 108.920 ; 
                RECT 2.880 109.960 210.240 110.280 ; 
                RECT 1196.600 109.960 1203.360 110.280 ; 
                RECT 2.880 111.320 183.040 111.640 ; 
                RECT 185.440 111.320 210.240 111.640 ; 
                RECT 1196.600 111.320 1203.360 111.640 ; 
                RECT 2.880 112.680 183.720 113.000 ; 
                RECT 186.120 112.680 210.240 113.000 ; 
                RECT 1196.600 112.680 1203.360 113.000 ; 
                RECT 2.880 114.040 210.240 114.360 ; 
                RECT 368.360 114.040 401.320 114.360 ; 
                RECT 1196.600 114.040 1203.360 114.360 ; 
                RECT 2.880 115.400 183.040 115.720 ; 
                RECT 185.440 115.400 401.320 115.720 ; 
                RECT 1196.600 115.400 1203.360 115.720 ; 
                RECT 2.880 116.760 173.520 117.080 ; 
                RECT 185.440 116.760 375.480 117.080 ; 
                RECT 1196.600 116.760 1203.360 117.080 ; 
                RECT 2.880 118.120 183.720 118.440 ; 
                RECT 186.120 118.120 395.880 118.440 ; 
                RECT 1196.600 118.120 1203.360 118.440 ; 
                RECT 2.880 119.480 395.880 119.800 ; 
                RECT 1196.600 119.480 1203.360 119.800 ; 
                RECT 2.880 120.840 390.440 121.160 ; 
                RECT 1196.600 120.840 1203.360 121.160 ; 
                RECT 2.880 122.200 170.800 122.520 ; 
                RECT 184.760 122.200 390.440 122.520 ; 
                RECT 1196.600 122.200 1203.360 122.520 ; 
                RECT 2.880 123.560 176.240 123.880 ; 
                RECT 188.160 123.560 385.000 123.880 ; 
                RECT 1196.600 123.560 1203.360 123.880 ; 
                RECT 2.880 124.920 178.960 125.240 ; 
                RECT 192.240 124.920 385.000 125.240 ; 
                RECT 1196.600 124.920 1203.360 125.240 ; 
                RECT 2.880 126.280 385.000 126.600 ; 
                RECT 1196.600 126.280 1203.360 126.600 ; 
                RECT 2.880 127.640 176.240 127.960 ; 
                RECT 194.280 127.640 379.560 127.960 ; 
                RECT 1196.600 127.640 1203.360 127.960 ; 
                RECT 2.880 129.000 180.320 129.320 ; 
                RECT 190.880 129.000 379.560 129.320 ; 
                RECT 1196.600 129.000 1203.360 129.320 ; 
                RECT 2.880 130.360 401.320 130.680 ; 
                RECT 1196.600 130.360 1203.360 130.680 ; 
                RECT 2.880 131.720 401.320 132.040 ; 
                RECT 1196.600 131.720 1203.360 132.040 ; 
                RECT 2.880 133.080 174.200 133.400 ; 
                RECT 177.960 133.080 401.320 133.400 ; 
                RECT 1196.600 133.080 1203.360 133.400 ; 
                RECT 2.880 134.440 174.880 134.760 ; 
                RECT 182.040 134.440 401.320 134.760 ; 
                RECT 1196.600 134.440 1203.360 134.760 ; 
                RECT 2.880 135.800 180.320 136.120 ; 
                RECT 182.720 135.800 401.320 136.120 ; 
                RECT 1196.600 135.800 1203.360 136.120 ; 
                RECT 2.880 137.160 179.640 137.480 ; 
                RECT 192.240 137.160 401.320 137.480 ; 
                RECT 1196.600 137.160 1203.360 137.480 ; 
                RECT 2.880 138.520 401.320 138.840 ; 
                RECT 1196.600 138.520 1203.360 138.840 ; 
                RECT 2.880 139.880 401.320 140.200 ; 
                RECT 1196.600 139.880 1203.360 140.200 ; 
                RECT 2.880 141.240 153.120 141.560 ; 
                RECT 171.160 141.240 401.320 141.560 ; 
                RECT 1196.600 141.240 1203.360 141.560 ; 
                RECT 2.880 142.600 153.120 142.920 ; 
                RECT 171.160 142.600 176.240 142.920 ; 
                RECT 181.360 142.600 401.320 142.920 ; 
                RECT 1196.600 142.600 1203.360 142.920 ; 
                RECT 2.880 143.960 153.120 144.280 ; 
                RECT 171.160 143.960 401.320 144.280 ; 
                RECT 1196.600 143.960 1203.360 144.280 ; 
                RECT 2.880 145.320 153.120 145.640 ; 
                RECT 171.160 145.320 189.840 145.640 ; 
                RECT 192.240 145.320 401.320 145.640 ; 
                RECT 1196.600 145.320 1203.360 145.640 ; 
                RECT 2.880 146.680 153.120 147.000 ; 
                RECT 171.160 146.680 401.320 147.000 ; 
                RECT 1196.600 146.680 1203.360 147.000 ; 
                RECT 2.880 148.040 153.120 148.360 ; 
                RECT 171.160 148.040 198.000 148.360 ; 
                RECT 260.240 148.040 263.280 148.360 ; 
                RECT 368.360 148.040 401.320 148.360 ; 
                RECT 1196.600 148.040 1203.360 148.360 ; 
                RECT 2.880 149.400 153.120 149.720 ; 
                RECT 171.160 149.400 177.600 149.720 ; 
                RECT 179.320 149.400 263.280 149.720 ; 
                RECT 368.360 149.400 401.320 149.720 ; 
                RECT 1196.600 149.400 1203.360 149.720 ; 
                RECT 2.880 150.760 153.120 151.080 ; 
                RECT 171.160 150.760 263.280 151.080 ; 
                RECT 368.360 150.760 401.320 151.080 ; 
                RECT 1196.600 150.760 1203.360 151.080 ; 
                RECT 2.880 152.120 153.120 152.440 ; 
                RECT 171.160 152.120 263.280 152.440 ; 
                RECT 368.360 152.120 401.320 152.440 ; 
                RECT 1196.600 152.120 1203.360 152.440 ; 
                RECT 2.880 153.480 153.120 153.800 ; 
                RECT 171.160 153.480 183.040 153.800 ; 
                RECT 191.560 153.480 263.280 153.800 ; 
                RECT 368.360 153.480 401.320 153.800 ; 
                RECT 1196.600 153.480 1203.360 153.800 ; 
                RECT 2.880 154.840 153.120 155.160 ; 
                RECT 171.160 154.840 263.280 155.160 ; 
                RECT 368.360 154.840 382.280 155.160 ; 
                RECT 1196.600 154.840 1203.360 155.160 ; 
                RECT 2.880 156.200 153.120 156.520 ; 
                RECT 171.160 156.200 263.280 156.520 ; 
                RECT 368.360 156.200 382.280 156.520 ; 
                RECT 1196.600 156.200 1203.360 156.520 ; 
                RECT 2.880 157.560 153.120 157.880 ; 
                RECT 171.160 157.560 263.280 157.880 ; 
                RECT 368.360 157.560 382.280 157.880 ; 
                RECT 1196.600 157.560 1203.360 157.880 ; 
                RECT 2.880 158.920 153.120 159.240 ; 
                RECT 171.840 158.920 387.720 159.240 ; 
                RECT 1196.600 158.920 1203.360 159.240 ; 
                RECT 2.880 160.280 153.120 160.600 ; 
                RECT 171.160 160.280 387.720 160.600 ; 
                RECT 1196.600 160.280 1203.360 160.600 ; 
                RECT 2.880 161.640 153.120 161.960 ; 
                RECT 171.160 161.640 393.160 161.960 ; 
                RECT 1196.600 161.640 1203.360 161.960 ; 
                RECT 2.880 163.000 153.120 163.320 ; 
                RECT 171.160 163.000 393.160 163.320 ; 
                RECT 1196.600 163.000 1203.360 163.320 ; 
                RECT 2.880 164.360 153.120 164.680 ; 
                RECT 171.160 164.360 263.960 164.680 ; 
                RECT 368.360 164.360 398.600 164.680 ; 
                RECT 1196.600 164.360 1203.360 164.680 ; 
                RECT 2.880 165.720 153.120 166.040 ; 
                RECT 171.160 165.720 263.960 166.040 ; 
                RECT 368.360 165.720 398.600 166.040 ; 
                RECT 1196.600 165.720 1203.360 166.040 ; 
                RECT 2.880 167.080 153.120 167.400 ; 
                RECT 171.160 167.080 263.960 167.400 ; 
                RECT 368.360 167.080 401.320 167.400 ; 
                RECT 1196.600 167.080 1203.360 167.400 ; 
                RECT 2.880 168.440 153.120 168.760 ; 
                RECT 171.160 168.440 263.960 168.760 ; 
                RECT 1196.600 168.440 1203.360 168.760 ; 
                RECT 2.880 169.800 153.120 170.120 ; 
                RECT 171.160 169.800 178.960 170.120 ; 
                RECT 182.040 169.800 263.960 170.120 ; 
                RECT 1196.600 169.800 1203.360 170.120 ; 
                RECT 2.880 171.160 153.120 171.480 ; 
                RECT 171.160 171.160 263.960 171.480 ; 
                RECT 1196.600 171.160 1203.360 171.480 ; 
                RECT 2.880 172.520 153.120 172.840 ; 
                RECT 171.160 172.520 263.960 172.840 ; 
                RECT 368.360 172.520 401.320 172.840 ; 
                RECT 1196.600 172.520 1203.360 172.840 ; 
                RECT 2.880 173.880 153.120 174.200 ; 
                RECT 171.160 173.880 263.960 174.200 ; 
                RECT 368.360 173.880 401.320 174.200 ; 
                RECT 1196.600 173.880 1203.360 174.200 ; 
                RECT 2.880 175.240 153.120 175.560 ; 
                RECT 171.160 175.240 263.960 175.560 ; 
                RECT 368.360 175.240 401.320 175.560 ; 
                RECT 1196.600 175.240 1203.360 175.560 ; 
                RECT 2.880 176.600 153.120 176.920 ; 
                RECT 171.160 176.600 263.960 176.920 ; 
                RECT 368.360 176.600 401.320 176.920 ; 
                RECT 1196.600 176.600 1203.360 176.920 ; 
                RECT 2.880 177.960 153.120 178.280 ; 
                RECT 171.160 177.960 263.960 178.280 ; 
                RECT 368.360 177.960 401.320 178.280 ; 
                RECT 1196.600 177.960 1203.360 178.280 ; 
                RECT 2.880 179.320 153.120 179.640 ; 
                RECT 171.160 179.320 263.960 179.640 ; 
                RECT 368.360 179.320 401.320 179.640 ; 
                RECT 1196.600 179.320 1203.360 179.640 ; 
                RECT 2.880 180.680 176.240 181.000 ; 
                RECT 182.040 180.680 263.960 181.000 ; 
                RECT 368.360 180.680 401.320 181.000 ; 
                RECT 1196.600 180.680 1203.360 181.000 ; 
                RECT 2.880 182.040 263.960 182.360 ; 
                RECT 368.360 182.040 401.320 182.360 ; 
                RECT 1196.600 182.040 1203.360 182.360 ; 
                RECT 2.880 183.400 263.960 183.720 ; 
                RECT 368.360 183.400 401.320 183.720 ; 
                RECT 1196.600 183.400 1203.360 183.720 ; 
                RECT 2.880 184.760 134.080 185.080 ; 
                RECT 152.800 184.760 180.320 185.080 ; 
                RECT 186.120 184.760 263.960 185.080 ; 
                RECT 368.360 184.760 401.320 185.080 ; 
                RECT 1196.600 184.760 1203.360 185.080 ; 
                RECT 2.880 186.120 134.080 186.440 ; 
                RECT 152.800 186.120 159.240 186.440 ; 
                RECT 166.400 186.120 263.960 186.440 ; 
                RECT 1196.600 186.120 1203.360 186.440 ; 
                RECT 2.880 187.480 134.080 187.800 ; 
                RECT 152.800 187.480 153.800 187.800 ; 
                RECT 171.160 187.480 263.960 187.800 ; 
                RECT 1196.600 187.480 1203.360 187.800 ; 
                RECT 2.880 188.840 134.080 189.160 ; 
                RECT 152.800 188.840 153.800 189.160 ; 
                RECT 171.160 188.840 263.960 189.160 ; 
                RECT 1196.600 188.840 1203.360 189.160 ; 
                RECT 2.880 190.200 134.080 190.520 ; 
                RECT 152.800 190.200 159.240 190.520 ; 
                RECT 166.400 190.200 173.520 190.520 ; 
                RECT 184.760 190.200 263.960 190.520 ; 
                RECT 1196.600 190.200 1203.360 190.520 ; 
                RECT 2.880 191.560 128.640 191.880 ; 
                RECT 165.720 191.560 263.960 191.880 ; 
                RECT 368.360 191.560 1203.360 191.880 ; 
                RECT 2.880 192.920 165.360 193.240 ; 
                RECT 260.920 192.920 1203.360 193.240 ; 
                RECT 2.880 194.280 398.600 194.600 ; 
                RECT 1199.320 194.280 1203.360 194.600 ; 
                RECT 2.880 195.640 398.600 195.960 ; 
                RECT 1199.320 195.640 1203.360 195.960 ; 
                RECT 2.880 197.000 398.600 197.320 ; 
                RECT 1199.320 197.000 1203.360 197.320 ; 
                RECT 2.880 198.360 27.320 198.680 ; 
                RECT 33.800 198.360 36.160 198.680 ; 
                RECT 48.760 198.360 99.400 198.680 ; 
                RECT 1199.320 198.360 1203.360 198.680 ; 
                RECT 2.880 199.720 25.280 200.040 ; 
                RECT 48.080 199.720 59.280 200.040 ; 
                RECT 61.000 199.720 75.600 200.040 ; 
                RECT 89.560 199.720 99.400 200.040 ; 
                RECT 1199.320 199.720 1203.360 200.040 ; 
                RECT 2.880 201.080 25.280 201.400 ; 
                RECT 35.840 201.080 59.280 201.400 ; 
                RECT 63.720 201.080 75.600 201.400 ; 
                RECT 89.560 201.080 99.400 201.400 ; 
                RECT 1199.320 201.080 1203.360 201.400 ; 
                RECT 2.880 202.440 25.280 202.760 ; 
                RECT 35.840 202.440 59.280 202.760 ; 
                RECT 63.720 202.440 75.600 202.760 ; 
                RECT 89.560 202.440 99.400 202.760 ; 
                RECT 1199.320 202.440 1203.360 202.760 ; 
                RECT 2.880 203.800 59.280 204.120 ; 
                RECT 64.400 203.800 75.600 204.120 ; 
                RECT 89.560 203.800 99.400 204.120 ; 
                RECT 1199.320 203.800 1203.360 204.120 ; 
                RECT 2.880 205.160 25.280 205.480 ; 
                RECT 35.840 205.160 59.280 205.480 ; 
                RECT 61.000 205.160 75.600 205.480 ; 
                RECT 89.560 205.160 99.400 205.480 ; 
                RECT 1199.320 205.160 1203.360 205.480 ; 
                RECT 2.880 206.520 25.280 206.840 ; 
                RECT 35.840 206.520 99.400 206.840 ; 
                RECT 1199.320 206.520 1203.360 206.840 ; 
                RECT 2.880 207.880 75.600 208.200 ; 
                RECT 89.560 207.880 99.400 208.200 ; 
                RECT 1199.320 207.880 1203.360 208.200 ; 
                RECT 2.880 209.240 75.600 209.560 ; 
                RECT 89.560 209.240 99.400 209.560 ; 
                RECT 1199.320 209.240 1203.360 209.560 ; 
                RECT 2.880 210.600 75.600 210.920 ; 
                RECT 89.560 210.600 99.400 210.920 ; 
                RECT 1199.320 210.600 1203.360 210.920 ; 
                RECT 2.880 211.960 18.480 212.280 ; 
                RECT 20.880 211.960 34.120 212.280 ; 
                RECT 37.200 211.960 75.600 212.280 ; 
                RECT 89.560 211.960 99.400 212.280 ; 
                RECT 1199.320 211.960 1203.360 212.280 ; 
                RECT 2.880 213.320 17.800 213.640 ; 
                RECT 20.880 213.320 34.120 213.640 ; 
                RECT 37.880 213.320 75.600 213.640 ; 
                RECT 89.560 213.320 99.400 213.640 ; 
                RECT 1199.320 213.320 1203.360 213.640 ; 
                RECT 2.880 214.680 17.120 215.000 ; 
                RECT 20.880 214.680 39.560 215.000 ; 
                RECT 48.760 214.680 99.400 215.000 ; 
                RECT 1199.320 214.680 1203.360 215.000 ; 
                RECT 2.880 216.040 16.440 216.360 ; 
                RECT 20.880 216.040 40.920 216.360 ; 
                RECT 47.400 216.040 59.280 216.360 ; 
                RECT 61.000 216.040 75.600 216.360 ; 
                RECT 89.560 216.040 99.400 216.360 ; 
                RECT 1199.320 216.040 1203.360 216.360 ; 
                RECT 2.880 217.400 59.280 217.720 ; 
                RECT 61.680 217.400 75.600 217.720 ; 
                RECT 89.560 217.400 99.400 217.720 ; 
                RECT 1199.320 217.400 1203.360 217.720 ; 
                RECT 2.880 218.760 15.760 219.080 ; 
                RECT 20.880 218.760 59.280 219.080 ; 
                RECT 61.680 218.760 75.600 219.080 ; 
                RECT 89.560 218.760 99.400 219.080 ; 
                RECT 1199.320 218.760 1203.360 219.080 ; 
                RECT 2.880 220.120 15.080 220.440 ; 
                RECT 20.880 220.120 59.280 220.440 ; 
                RECT 62.360 220.120 75.600 220.440 ; 
                RECT 89.560 220.120 99.400 220.440 ; 
                RECT 1199.320 220.120 1203.360 220.440 ; 
                RECT 2.880 221.480 59.280 221.800 ; 
                RECT 63.040 221.480 75.600 221.800 ; 
                RECT 89.560 221.480 99.400 221.800 ; 
                RECT 1199.320 221.480 1203.360 221.800 ; 
                RECT 2.880 222.840 14.400 223.160 ; 
                RECT 20.880 222.840 99.400 223.160 ; 
                RECT 1199.320 222.840 1203.360 223.160 ; 
                RECT 2.880 224.200 13.720 224.520 ; 
                RECT 20.880 224.200 34.120 224.520 ; 
                RECT 41.960 224.200 75.600 224.520 ; 
                RECT 89.560 224.200 99.400 224.520 ; 
                RECT 1199.320 224.200 1203.360 224.520 ; 
                RECT 2.880 225.560 75.600 225.880 ; 
                RECT 89.560 225.560 99.400 225.880 ; 
                RECT 1199.320 225.560 1203.360 225.880 ; 
                RECT 2.880 226.920 13.040 227.240 ; 
                RECT 20.880 226.920 34.120 227.240 ; 
                RECT 40.600 226.920 75.600 227.240 ; 
                RECT 89.560 226.920 99.400 227.240 ; 
                RECT 1199.320 226.920 1203.360 227.240 ; 
                RECT 2.880 228.280 12.360 228.600 ; 
                RECT 20.880 228.280 34.120 228.600 ; 
                RECT 39.920 228.280 75.600 228.600 ; 
                RECT 89.560 228.280 99.400 228.600 ; 
                RECT 1199.320 228.280 1203.360 228.600 ; 
                RECT 2.880 229.640 11.680 229.960 ; 
                RECT 20.880 229.640 34.120 229.960 ; 
                RECT 39.240 229.640 75.600 229.960 ; 
                RECT 85.480 229.640 99.400 229.960 ; 
                RECT 1199.320 229.640 1203.360 229.960 ; 
                RECT 2.880 231.000 11.000 231.320 ; 
                RECT 20.880 231.000 80.360 231.320 ; 
                RECT 89.560 231.000 99.400 231.320 ; 
                RECT 1199.320 231.000 1203.360 231.320 ; 
                RECT 2.880 232.360 75.600 232.680 ; 
                RECT 89.560 232.360 99.400 232.680 ; 
                RECT 1199.320 232.360 1203.360 232.680 ; 
                RECT 2.880 233.720 10.320 234.040 ; 
                RECT 20.880 233.720 34.120 234.040 ; 
                RECT 37.880 233.720 75.600 234.040 ; 
                RECT 89.560 233.720 99.400 234.040 ; 
                RECT 1199.320 233.720 1203.360 234.040 ; 
                RECT 2.880 235.080 9.640 235.400 ; 
                RECT 20.880 235.080 75.600 235.400 ; 
                RECT 89.560 235.080 99.400 235.400 ; 
                RECT 1199.320 235.080 1203.360 235.400 ; 
                RECT 2.880 236.440 75.600 236.760 ; 
                RECT 89.560 236.440 99.400 236.760 ; 
                RECT 1199.320 236.440 1203.360 236.760 ; 
                RECT 2.880 237.800 75.600 238.120 ; 
                RECT 86.160 237.800 99.400 238.120 ; 
                RECT 1199.320 237.800 1203.360 238.120 ; 
                RECT 2.880 239.160 75.600 239.480 ; 
                RECT 89.560 239.160 99.400 239.480 ; 
                RECT 1199.320 239.160 1203.360 239.480 ; 
                RECT 2.880 240.520 75.600 240.840 ; 
                RECT 89.560 240.520 99.400 240.840 ; 
                RECT 1199.320 240.520 1203.360 240.840 ; 
                RECT 2.880 241.880 75.600 242.200 ; 
                RECT 89.560 241.880 99.400 242.200 ; 
                RECT 1199.320 241.880 1203.360 242.200 ; 
                RECT 2.880 243.240 75.600 243.560 ; 
                RECT 89.560 243.240 99.400 243.560 ; 
                RECT 1199.320 243.240 1203.360 243.560 ; 
                RECT 2.880 244.600 75.600 244.920 ; 
                RECT 89.560 244.600 99.400 244.920 ; 
                RECT 1199.320 244.600 1203.360 244.920 ; 
                RECT 2.880 245.960 75.600 246.280 ; 
                RECT 86.840 245.960 99.400 246.280 ; 
                RECT 1199.320 245.960 1203.360 246.280 ; 
                RECT 2.880 247.320 75.600 247.640 ; 
                RECT 89.560 247.320 99.400 247.640 ; 
                RECT 1199.320 247.320 1203.360 247.640 ; 
                RECT 2.880 248.680 75.600 249.000 ; 
                RECT 89.560 248.680 99.400 249.000 ; 
                RECT 1199.320 248.680 1203.360 249.000 ; 
                RECT 2.880 250.040 75.600 250.360 ; 
                RECT 89.560 250.040 99.400 250.360 ; 
                RECT 1199.320 250.040 1203.360 250.360 ; 
                RECT 2.880 251.400 75.600 251.720 ; 
                RECT 89.560 251.400 99.400 251.720 ; 
                RECT 1199.320 251.400 1203.360 251.720 ; 
                RECT 2.880 252.760 75.600 253.080 ; 
                RECT 89.560 252.760 99.400 253.080 ; 
                RECT 1199.320 252.760 1203.360 253.080 ; 
                RECT 2.880 254.120 99.400 254.440 ; 
                RECT 1199.320 254.120 1203.360 254.440 ; 
                RECT 2.880 255.480 75.600 255.800 ; 
                RECT 89.560 255.480 99.400 255.800 ; 
                RECT 1199.320 255.480 1203.360 255.800 ; 
                RECT 2.880 256.840 75.600 257.160 ; 
                RECT 89.560 256.840 99.400 257.160 ; 
                RECT 1199.320 256.840 1203.360 257.160 ; 
                RECT 2.880 258.200 75.600 258.520 ; 
                RECT 89.560 258.200 99.400 258.520 ; 
                RECT 1199.320 258.200 1203.360 258.520 ; 
                RECT 2.880 259.560 75.600 259.880 ; 
                RECT 89.560 259.560 99.400 259.880 ; 
                RECT 1199.320 259.560 1203.360 259.880 ; 
                RECT 2.880 260.920 75.600 261.240 ; 
                RECT 89.560 260.920 99.400 261.240 ; 
                RECT 1199.320 260.920 1203.360 261.240 ; 
                RECT 2.880 262.280 99.400 262.600 ; 
                RECT 1199.320 262.280 1203.360 262.600 ; 
                RECT 2.880 263.640 76.960 263.960 ; 
                RECT 89.560 263.640 99.400 263.960 ; 
                RECT 1199.320 263.640 1203.360 263.960 ; 
                RECT 2.880 265.000 76.960 265.320 ; 
                RECT 89.560 265.000 99.400 265.320 ; 
                RECT 1199.320 265.000 1203.360 265.320 ; 
                RECT 2.880 266.360 76.960 266.680 ; 
                RECT 89.560 266.360 99.400 266.680 ; 
                RECT 1199.320 266.360 1203.360 266.680 ; 
                RECT 2.880 267.720 81.720 268.040 ; 
                RECT 89.560 267.720 99.400 268.040 ; 
                RECT 1199.320 267.720 1203.360 268.040 ; 
                RECT 2.880 269.080 76.960 269.400 ; 
                RECT 89.560 269.080 99.400 269.400 ; 
                RECT 1199.320 269.080 1203.360 269.400 ; 
                RECT 2.880 270.440 38.880 270.760 ; 
                RECT 64.400 270.440 99.400 270.760 ; 
                RECT 1199.320 270.440 1203.360 270.760 ; 
                RECT 2.880 271.800 37.520 272.120 ; 
                RECT 63.720 271.800 75.600 272.120 ; 
                RECT 89.560 271.800 99.400 272.120 ; 
                RECT 1199.320 271.800 1203.360 272.120 ; 
                RECT 2.880 273.160 36.160 273.480 ; 
                RECT 63.040 273.160 75.600 273.480 ; 
                RECT 89.560 273.160 99.400 273.480 ; 
                RECT 1199.320 273.160 1203.360 273.480 ; 
                RECT 2.880 274.520 76.960 274.840 ; 
                RECT 89.560 274.520 99.400 274.840 ; 
                RECT 1199.320 274.520 1203.360 274.840 ; 
                RECT 2.880 275.880 75.600 276.200 ; 
                RECT 89.560 275.880 99.400 276.200 ; 
                RECT 1199.320 275.880 1203.360 276.200 ; 
                RECT 2.880 277.240 75.600 277.560 ; 
                RECT 78.000 277.240 99.400 277.560 ; 
                RECT 1199.320 277.240 1203.360 277.560 ; 
                RECT 2.880 278.600 83.760 278.920 ; 
                RECT 89.560 278.600 99.400 278.920 ; 
                RECT 1199.320 278.600 1203.360 278.920 ; 
                RECT 2.880 279.960 75.600 280.280 ; 
                RECT 89.560 279.960 99.400 280.280 ; 
                RECT 1199.320 279.960 1203.360 280.280 ; 
                RECT 2.880 281.320 75.600 281.640 ; 
                RECT 89.560 281.320 99.400 281.640 ; 
                RECT 1199.320 281.320 1203.360 281.640 ; 
                RECT 2.880 282.680 75.600 283.000 ; 
                RECT 89.560 282.680 99.400 283.000 ; 
                RECT 1199.320 282.680 1203.360 283.000 ; 
                RECT 2.880 284.040 75.600 284.360 ; 
                RECT 89.560 284.040 99.400 284.360 ; 
                RECT 1199.320 284.040 1203.360 284.360 ; 
                RECT 2.880 285.400 75.600 285.720 ; 
                RECT 78.680 285.400 99.400 285.720 ; 
                RECT 1199.320 285.400 1203.360 285.720 ; 
                RECT 2.880 286.760 85.800 287.080 ; 
                RECT 89.560 286.760 99.400 287.080 ; 
                RECT 1199.320 286.760 1203.360 287.080 ; 
                RECT 2.880 288.120 75.600 288.440 ; 
                RECT 89.560 288.120 99.400 288.440 ; 
                RECT 1199.320 288.120 1203.360 288.440 ; 
                RECT 2.880 289.480 75.600 289.800 ; 
                RECT 89.560 289.480 99.400 289.800 ; 
                RECT 1199.320 289.480 1203.360 289.800 ; 
                RECT 2.880 290.840 75.600 291.160 ; 
                RECT 89.560 290.840 99.400 291.160 ; 
                RECT 1199.320 290.840 1203.360 291.160 ; 
                RECT 2.880 292.200 75.600 292.520 ; 
                RECT 89.560 292.200 99.400 292.520 ; 
                RECT 1199.320 292.200 1203.360 292.520 ; 
                RECT 2.880 293.560 99.400 293.880 ; 
                RECT 1199.320 293.560 1203.360 293.880 ; 
                RECT 2.880 294.920 77.640 295.240 ; 
                RECT 89.560 294.920 99.400 295.240 ; 
                RECT 1199.320 294.920 1203.360 295.240 ; 
                RECT 2.880 296.280 75.600 296.600 ; 
                RECT 89.560 296.280 99.400 296.600 ; 
                RECT 1199.320 296.280 1203.360 296.600 ; 
                RECT 2.880 297.640 75.600 297.960 ; 
                RECT 89.560 297.640 99.400 297.960 ; 
                RECT 1199.320 297.640 1203.360 297.960 ; 
                RECT 2.880 299.000 75.600 299.320 ; 
                RECT 89.560 299.000 99.400 299.320 ; 
                RECT 1199.320 299.000 1203.360 299.320 ; 
                RECT 2.880 300.360 75.600 300.680 ; 
                RECT 89.560 300.360 99.400 300.680 ; 
                RECT 1199.320 300.360 1203.360 300.680 ; 
                RECT 2.880 301.720 99.400 302.040 ; 
                RECT 1199.320 301.720 1203.360 302.040 ; 
                RECT 2.880 303.080 77.640 303.400 ; 
                RECT 89.560 303.080 99.400 303.400 ; 
                RECT 1199.320 303.080 1203.360 303.400 ; 
                RECT 2.880 304.440 75.600 304.760 ; 
                RECT 89.560 304.440 99.400 304.760 ; 
                RECT 1199.320 304.440 1203.360 304.760 ; 
                RECT 2.880 305.800 75.600 306.120 ; 
                RECT 89.560 305.800 99.400 306.120 ; 
                RECT 1199.320 305.800 1203.360 306.120 ; 
                RECT 2.880 307.160 75.600 307.480 ; 
                RECT 89.560 307.160 99.400 307.480 ; 
                RECT 1199.320 307.160 1203.360 307.480 ; 
                RECT 2.880 308.520 75.600 308.840 ; 
                RECT 89.560 308.520 99.400 308.840 ; 
                RECT 1199.320 308.520 1203.360 308.840 ; 
                RECT 2.880 309.880 99.400 310.200 ; 
                RECT 1199.320 309.880 1203.360 310.200 ; 
                RECT 2.880 311.240 75.600 311.560 ; 
                RECT 89.560 311.240 99.400 311.560 ; 
                RECT 1199.320 311.240 1203.360 311.560 ; 
                RECT 2.880 312.600 75.600 312.920 ; 
                RECT 89.560 312.600 99.400 312.920 ; 
                RECT 1199.320 312.600 1203.360 312.920 ; 
                RECT 2.880 313.960 77.640 314.280 ; 
                RECT 89.560 313.960 99.400 314.280 ; 
                RECT 1199.320 313.960 1203.360 314.280 ; 
                RECT 2.880 315.320 75.600 315.640 ; 
                RECT 89.560 315.320 99.400 315.640 ; 
                RECT 1199.320 315.320 1203.360 315.640 ; 
                RECT 2.880 316.680 75.600 317.000 ; 
                RECT 80.720 316.680 99.400 317.000 ; 
                RECT 1199.320 316.680 1203.360 317.000 ; 
                RECT 2.880 318.040 85.800 318.360 ; 
                RECT 89.560 318.040 99.400 318.360 ; 
                RECT 1199.320 318.040 1203.360 318.360 ; 
                RECT 2.880 319.400 75.600 319.720 ; 
                RECT 89.560 319.400 99.400 319.720 ; 
                RECT 1199.320 319.400 1203.360 319.720 ; 
                RECT 2.880 320.760 75.600 321.080 ; 
                RECT 89.560 320.760 99.400 321.080 ; 
                RECT 1199.320 320.760 1203.360 321.080 ; 
                RECT 2.880 322.120 75.600 322.440 ; 
                RECT 89.560 322.120 99.400 322.440 ; 
                RECT 1199.320 322.120 1203.360 322.440 ; 
                RECT 2.880 323.480 75.600 323.800 ; 
                RECT 89.560 323.480 99.400 323.800 ; 
                RECT 1199.320 323.480 1203.360 323.800 ; 
                RECT 2.880 324.840 75.600 325.160 ; 
                RECT 80.720 324.840 99.400 325.160 ; 
                RECT 1199.320 324.840 1203.360 325.160 ; 
                RECT 2.880 326.200 80.360 326.520 ; 
                RECT 89.560 326.200 99.400 326.520 ; 
                RECT 1199.320 326.200 1203.360 326.520 ; 
                RECT 2.880 327.560 75.600 327.880 ; 
                RECT 89.560 327.560 99.400 327.880 ; 
                RECT 1199.320 327.560 1203.360 327.880 ; 
                RECT 2.880 328.920 75.600 329.240 ; 
                RECT 89.560 328.920 99.400 329.240 ; 
                RECT 1199.320 328.920 1203.360 329.240 ; 
                RECT 2.880 330.280 75.600 330.600 ; 
                RECT 89.560 330.280 99.400 330.600 ; 
                RECT 1199.320 330.280 1203.360 330.600 ; 
                RECT 2.880 331.640 75.600 331.960 ; 
                RECT 89.560 331.640 99.400 331.960 ; 
                RECT 1199.320 331.640 1203.360 331.960 ; 
                RECT 2.880 333.000 99.400 333.320 ; 
                RECT 1199.320 333.000 1203.360 333.320 ; 
                RECT 2.880 334.360 78.320 334.680 ; 
                RECT 89.560 334.360 99.400 334.680 ; 
                RECT 1199.320 334.360 1203.360 334.680 ; 
                RECT 2.880 335.720 82.400 336.040 ; 
                RECT 89.560 335.720 99.400 336.040 ; 
                RECT 1199.320 335.720 1203.360 336.040 ; 
                RECT 2.880 337.080 83.080 337.400 ; 
                RECT 89.560 337.080 99.400 337.400 ; 
                RECT 1199.320 337.080 1203.360 337.400 ; 
                RECT 2.880 338.440 78.320 338.760 ; 
                RECT 89.560 338.440 99.400 338.760 ; 
                RECT 1199.320 338.440 1203.360 338.760 ; 
                RECT 2.880 339.800 78.320 340.120 ; 
                RECT 89.560 339.800 99.400 340.120 ; 
                RECT 1199.320 339.800 1203.360 340.120 ; 
                RECT 2.880 341.160 99.400 341.480 ; 
                RECT 1199.320 341.160 1203.360 341.480 ; 
                RECT 2.880 342.520 78.320 342.840 ; 
                RECT 89.560 342.520 99.400 342.840 ; 
                RECT 1199.320 342.520 1203.360 342.840 ; 
                RECT 2.880 343.880 78.320 344.200 ; 
                RECT 89.560 343.880 99.400 344.200 ; 
                RECT 1199.320 343.880 1203.360 344.200 ; 
                RECT 2.880 345.240 78.320 345.560 ; 
                RECT 89.560 345.240 99.400 345.560 ; 
                RECT 1199.320 345.240 1203.360 345.560 ; 
                RECT 2.880 346.600 85.120 346.920 ; 
                RECT 89.560 346.600 99.400 346.920 ; 
                RECT 1199.320 346.600 1203.360 346.920 ; 
                RECT 2.880 347.960 78.320 348.280 ; 
                RECT 89.560 347.960 99.400 348.280 ; 
                RECT 1199.320 347.960 1203.360 348.280 ; 
                RECT 2.880 349.320 99.400 349.640 ; 
                RECT 1199.320 349.320 1203.360 349.640 ; 
                RECT 2.880 350.680 78.320 351.000 ; 
                RECT 89.560 350.680 99.400 351.000 ; 
                RECT 1199.320 350.680 1203.360 351.000 ; 
                RECT 2.880 352.040 78.320 352.360 ; 
                RECT 89.560 352.040 99.400 352.360 ; 
                RECT 1199.320 352.040 1203.360 352.360 ; 
                RECT 2.880 353.400 78.320 353.720 ; 
                RECT 89.560 353.400 99.400 353.720 ; 
                RECT 1199.320 353.400 1203.360 353.720 ; 
                RECT 2.880 354.760 78.320 355.080 ; 
                RECT 89.560 354.760 99.400 355.080 ; 
                RECT 1199.320 354.760 1203.360 355.080 ; 
                RECT 2.880 356.120 99.400 356.440 ; 
                RECT 1199.320 356.120 1203.360 356.440 ; 
                RECT 2.880 357.480 80.360 357.800 ; 
                RECT 89.560 357.480 99.400 357.800 ; 
                RECT 1199.320 357.480 1203.360 357.800 ; 
                RECT 2.880 358.840 79.000 359.160 ; 
                RECT 89.560 358.840 99.400 359.160 ; 
                RECT 1199.320 358.840 1203.360 359.160 ; 
                RECT 2.880 360.200 79.000 360.520 ; 
                RECT 89.560 360.200 99.400 360.520 ; 
                RECT 1199.320 360.200 1203.360 360.520 ; 
                RECT 2.880 361.560 79.000 361.880 ; 
                RECT 89.560 361.560 99.400 361.880 ; 
                RECT 1199.320 361.560 1203.360 361.880 ; 
                RECT 2.880 362.920 79.000 363.240 ; 
                RECT 89.560 362.920 99.400 363.240 ; 
                RECT 1199.320 362.920 1203.360 363.240 ; 
                RECT 2.880 364.280 99.400 364.600 ; 
                RECT 1199.320 364.280 1203.360 364.600 ; 
                RECT 2.880 365.640 81.720 365.960 ; 
                RECT 89.560 365.640 99.400 365.960 ; 
                RECT 1199.320 365.640 1203.360 365.960 ; 
                RECT 2.880 367.000 79.000 367.320 ; 
                RECT 89.560 367.000 99.400 367.320 ; 
                RECT 1199.320 367.000 1203.360 367.320 ; 
                RECT 2.880 368.360 79.000 368.680 ; 
                RECT 89.560 368.360 99.400 368.680 ; 
                RECT 1199.320 368.360 1203.360 368.680 ; 
                RECT 2.880 369.720 79.000 370.040 ; 
                RECT 89.560 369.720 99.400 370.040 ; 
                RECT 1199.320 369.720 1203.360 370.040 ; 
                RECT 2.880 371.080 79.000 371.400 ; 
                RECT 89.560 371.080 99.400 371.400 ; 
                RECT 1199.320 371.080 1203.360 371.400 ; 
                RECT 2.880 372.440 99.400 372.760 ; 
                RECT 1199.320 372.440 1203.360 372.760 ; 
                RECT 2.880 373.800 79.000 374.120 ; 
                RECT 89.560 373.800 99.400 374.120 ; 
                RECT 1199.320 373.800 1203.360 374.120 ; 
                RECT 2.880 375.160 84.440 375.480 ; 
                RECT 89.560 375.160 99.400 375.480 ; 
                RECT 1199.320 375.160 1203.360 375.480 ; 
                RECT 2.880 376.520 79.000 376.840 ; 
                RECT 89.560 376.520 99.400 376.840 ; 
                RECT 1199.320 376.520 1203.360 376.840 ; 
                RECT 2.880 377.880 79.000 378.200 ; 
                RECT 89.560 377.880 99.400 378.200 ; 
                RECT 1199.320 377.880 1203.360 378.200 ; 
                RECT 2.880 379.240 79.000 379.560 ; 
                RECT 89.560 379.240 99.400 379.560 ; 
                RECT 1199.320 379.240 1203.360 379.560 ; 
                RECT 2.880 380.600 99.400 380.920 ; 
                RECT 1199.320 380.600 1203.360 380.920 ; 
                RECT 2.880 381.960 79.000 382.280 ; 
                RECT 89.560 381.960 99.400 382.280 ; 
                RECT 1199.320 381.960 1203.360 382.280 ; 
                RECT 2.880 383.320 79.000 383.640 ; 
                RECT 89.560 383.320 99.400 383.640 ; 
                RECT 1199.320 383.320 1203.360 383.640 ; 
                RECT 2.880 384.680 87.160 385.000 ; 
                RECT 89.560 384.680 99.400 385.000 ; 
                RECT 1199.320 384.680 1203.360 385.000 ; 
                RECT 2.880 386.040 87.160 386.360 ; 
                RECT 89.560 386.040 99.400 386.360 ; 
                RECT 1199.320 386.040 1203.360 386.360 ; 
                RECT 2.880 387.400 79.000 387.720 ; 
                RECT 89.560 387.400 99.400 387.720 ; 
                RECT 1199.320 387.400 1203.360 387.720 ; 
                RECT 2.880 388.760 99.400 389.080 ; 
                RECT 1199.320 388.760 1203.360 389.080 ; 
                RECT 2.880 390.120 79.000 390.440 ; 
                RECT 89.560 390.120 99.400 390.440 ; 
                RECT 1199.320 390.120 1203.360 390.440 ; 
                RECT 2.880 391.480 79.000 391.800 ; 
                RECT 89.560 391.480 99.400 391.800 ; 
                RECT 1199.320 391.480 1203.360 391.800 ; 
                RECT 2.880 392.840 79.000 393.160 ; 
                RECT 89.560 392.840 99.400 393.160 ; 
                RECT 1199.320 392.840 1203.360 393.160 ; 
                RECT 2.880 394.200 81.720 394.520 ; 
                RECT 89.560 394.200 99.400 394.520 ; 
                RECT 1199.320 394.200 1203.360 394.520 ; 
                RECT 2.880 395.560 99.400 395.880 ; 
                RECT 1199.320 395.560 1203.360 395.880 ; 
                RECT 2.880 396.920 81.720 397.240 ; 
                RECT 89.560 396.920 99.400 397.240 ; 
                RECT 1199.320 396.920 1203.360 397.240 ; 
                RECT 2.880 398.280 79.000 398.600 ; 
                RECT 89.560 398.280 99.400 398.600 ; 
                RECT 1199.320 398.280 1203.360 398.600 ; 
                RECT 2.880 399.640 79.000 399.960 ; 
                RECT 89.560 399.640 99.400 399.960 ; 
                RECT 1199.320 399.640 1203.360 399.960 ; 
                RECT 2.880 401.000 79.000 401.320 ; 
                RECT 89.560 401.000 99.400 401.320 ; 
                RECT 1199.320 401.000 1203.360 401.320 ; 
                RECT 2.880 402.360 79.000 402.680 ; 
                RECT 89.560 402.360 99.400 402.680 ; 
                RECT 1199.320 402.360 1203.360 402.680 ; 
                RECT 2.880 403.720 99.400 404.040 ; 
                RECT 1199.320 403.720 1203.360 404.040 ; 
                RECT 2.880 405.080 83.760 405.400 ; 
                RECT 89.560 405.080 99.400 405.400 ; 
                RECT 1199.320 405.080 1203.360 405.400 ; 
                RECT 2.880 406.440 79.000 406.760 ; 
                RECT 89.560 406.440 99.400 406.760 ; 
                RECT 1199.320 406.440 1203.360 406.760 ; 
                RECT 2.880 407.800 79.000 408.120 ; 
                RECT 89.560 407.800 99.400 408.120 ; 
                RECT 1199.320 407.800 1203.360 408.120 ; 
                RECT 2.880 409.160 79.000 409.480 ; 
                RECT 89.560 409.160 99.400 409.480 ; 
                RECT 1199.320 409.160 1203.360 409.480 ; 
                RECT 2.880 410.520 79.000 410.840 ; 
                RECT 89.560 410.520 99.400 410.840 ; 
                RECT 1199.320 410.520 1203.360 410.840 ; 
                RECT 2.880 411.880 99.400 412.200 ; 
                RECT 1199.320 411.880 1203.360 412.200 ; 
                RECT 2.880 413.240 79.000 413.560 ; 
                RECT 89.560 413.240 99.400 413.560 ; 
                RECT 1199.320 413.240 1203.360 413.560 ; 
                RECT 2.880 414.600 86.480 414.920 ; 
                RECT 89.560 414.600 99.400 414.920 ; 
                RECT 1199.320 414.600 1203.360 414.920 ; 
                RECT 2.880 415.960 79.000 416.280 ; 
                RECT 89.560 415.960 99.400 416.280 ; 
                RECT 1199.320 415.960 1203.360 416.280 ; 
                RECT 2.880 417.320 79.000 417.640 ; 
                RECT 89.560 417.320 99.400 417.640 ; 
                RECT 1199.320 417.320 1203.360 417.640 ; 
                RECT 2.880 418.680 79.000 419.000 ; 
                RECT 89.560 418.680 99.400 419.000 ; 
                RECT 1199.320 418.680 1203.360 419.000 ; 
                RECT 2.880 420.040 99.400 420.360 ; 
                RECT 1199.320 420.040 1203.360 420.360 ; 
                RECT 2.880 421.400 79.680 421.720 ; 
                RECT 89.560 421.400 99.400 421.720 ; 
                RECT 1199.320 421.400 1203.360 421.720 ; 
                RECT 2.880 422.760 79.680 423.080 ; 
                RECT 89.560 422.760 99.400 423.080 ; 
                RECT 1199.320 422.760 1203.360 423.080 ; 
                RECT 2.880 424.120 81.040 424.440 ; 
                RECT 89.560 424.120 99.400 424.440 ; 
                RECT 1199.320 424.120 1203.360 424.440 ; 
                RECT 2.880 425.480 79.680 425.800 ; 
                RECT 89.560 425.480 99.400 425.800 ; 
                RECT 1199.320 425.480 1203.360 425.800 ; 
                RECT 2.880 426.840 79.680 427.160 ; 
                RECT 89.560 426.840 99.400 427.160 ; 
                RECT 1199.320 426.840 1203.360 427.160 ; 
                RECT 2.880 428.200 99.400 428.520 ; 
                RECT 1199.320 428.200 1203.360 428.520 ; 
                RECT 2.880 429.560 79.680 429.880 ; 
                RECT 89.560 429.560 99.400 429.880 ; 
                RECT 1199.320 429.560 1203.360 429.880 ; 
                RECT 2.880 430.920 79.680 431.240 ; 
                RECT 89.560 430.920 99.400 431.240 ; 
                RECT 1199.320 430.920 1203.360 431.240 ; 
                RECT 2.880 432.280 79.680 432.600 ; 
                RECT 89.560 432.280 99.400 432.600 ; 
                RECT 1199.320 432.280 1203.360 432.600 ; 
                RECT 2.880 433.640 83.760 433.960 ; 
                RECT 89.560 433.640 99.400 433.960 ; 
                RECT 1199.320 433.640 1203.360 433.960 ; 
                RECT 2.880 435.000 79.680 435.320 ; 
                RECT 89.560 435.000 99.400 435.320 ; 
                RECT 1199.320 435.000 1203.360 435.320 ; 
                RECT 2.880 436.360 99.400 436.680 ; 
                RECT 1199.320 436.360 1203.360 436.680 ; 
                RECT 2.880 437.720 79.680 438.040 ; 
                RECT 89.560 437.720 99.400 438.040 ; 
                RECT 1199.320 437.720 1203.360 438.040 ; 
                RECT 2.880 439.080 79.680 439.400 ; 
                RECT 89.560 439.080 99.400 439.400 ; 
                RECT 1199.320 439.080 1203.360 439.400 ; 
                RECT 2.880 440.440 79.680 440.760 ; 
                RECT 89.560 440.440 99.400 440.760 ; 
                RECT 1199.320 440.440 1203.360 440.760 ; 
                RECT 2.880 441.800 79.680 442.120 ; 
                RECT 89.560 441.800 99.400 442.120 ; 
                RECT 1199.320 441.800 1203.360 442.120 ; 
                RECT 2.880 443.160 99.400 443.480 ; 
                RECT 1199.320 443.160 1203.360 443.480 ; 
                RECT 2.880 444.520 85.800 444.840 ; 
                RECT 89.560 444.520 99.400 444.840 ; 
                RECT 1199.320 444.520 1203.360 444.840 ; 
                RECT 2.880 445.880 79.680 446.200 ; 
                RECT 89.560 445.880 99.400 446.200 ; 
                RECT 1199.320 445.880 1203.360 446.200 ; 
                RECT 2.880 447.240 79.680 447.560 ; 
                RECT 89.560 447.240 99.400 447.560 ; 
                RECT 1199.320 447.240 1203.360 447.560 ; 
                RECT 2.880 448.600 79.680 448.920 ; 
                RECT 89.560 448.600 99.400 448.920 ; 
                RECT 1199.320 448.600 1203.360 448.920 ; 
                RECT 2.880 449.960 79.680 450.280 ; 
                RECT 89.560 449.960 99.400 450.280 ; 
                RECT 1199.320 449.960 1203.360 450.280 ; 
                RECT 2.880 451.320 99.400 451.640 ; 
                RECT 1199.320 451.320 1203.360 451.640 ; 
                RECT 2.880 452.680 99.400 453.000 ; 
                RECT 1199.320 452.680 1203.360 453.000 ; 
                RECT 2.880 454.040 398.600 454.360 ; 
                RECT 1199.320 454.040 1203.360 454.360 ; 
                RECT 2.880 455.400 398.600 455.720 ; 
                RECT 1199.320 455.400 1203.360 455.720 ; 
                RECT 2.880 456.760 1203.360 457.080 ; 
                RECT 2.880 458.120 1203.360 458.440 ; 
                RECT 2.880 459.480 1203.360 459.800 ; 
                RECT 2.880 460.840 1203.360 461.160 ; 
                RECT 2.880 462.200 1203.360 462.520 ; 
                RECT 2.880 2.880 1203.360 4.240 ; 
                RECT 2.880 463.520 1203.360 464.880 ; 
                RECT 402.740 29.465 408.540 30.585 ; 
                RECT 1189.040 29.465 1194.840 30.585 ; 
                RECT 402.740 35.255 408.540 35.875 ; 
                RECT 1189.040 35.255 1194.840 35.875 ; 
                RECT 402.740 40.280 408.540 40.920 ; 
                RECT 1189.040 40.280 1194.840 40.920 ; 
                RECT 402.740 45.410 408.540 46.060 ; 
                RECT 1189.040 45.410 1194.840 46.060 ; 
                RECT 402.740 50.625 408.540 51.235 ; 
                RECT 1189.040 50.625 1194.840 51.235 ; 
                RECT 402.740 55.555 408.540 56.165 ; 
                RECT 1189.040 55.555 1194.840 56.165 ; 
                RECT 402.740 149.055 1194.840 150.855 ; 
                RECT 402.740 89.925 1194.840 93.525 ; 
                RECT 402.740 115.385 1194.840 115.675 ; 
                RECT 402.740 81.350 1194.840 82.150 ; 
                RECT 402.740 69.290 1194.840 71.090 ; 
                RECT 402.740 86.240 1194.840 87.040 ; 
                RECT 402.740 83.030 1194.840 83.830 ; 
                RECT 402.740 78.340 1194.840 79.140 ; 
                RECT 402.740 20.095 1194.840 21.895 ; 
                RECT 99.985 198.075 101.305 452.455 ; 
                RECT 109.240 198.075 111.160 452.455 ; 
                RECT 124.815 198.075 126.735 452.455 ; 
                RECT 147.945 198.075 149.865 452.455 ; 
                RECT 151.785 198.075 153.705 452.455 ; 
                RECT 155.625 198.075 157.545 452.455 ; 
                RECT 191.285 198.075 193.205 452.455 ; 
                RECT 195.125 198.075 197.045 452.455 ; 
                RECT 198.965 198.075 200.885 452.455 ; 
                RECT 202.805 198.075 204.725 452.455 ; 
                RECT 206.645 198.075 208.565 452.455 ; 
                RECT 267.120 198.075 269.040 452.455 ; 
                RECT 270.960 198.075 272.880 452.455 ; 
                RECT 274.800 198.075 276.720 452.455 ; 
                RECT 278.640 198.075 280.560 452.455 ; 
                RECT 282.480 198.075 284.400 452.455 ; 
                RECT 286.320 198.075 288.240 452.455 ; 
                RECT 290.160 198.075 292.080 452.455 ; 
                RECT 294.000 198.075 295.920 452.455 ; 
                RECT 297.840 198.075 299.760 452.455 ; 
                RECT 210.810 61.225 211.700 113.825 ; 
                RECT 217.140 61.225 218.030 113.825 ; 
                RECT 223.900 61.225 224.790 113.825 ; 
                RECT 230.445 61.225 231.765 113.825 ; 
                RECT 240.560 61.225 242.480 113.825 ; 
                RECT 258.300 61.225 260.220 113.825 ; 
                RECT 262.140 61.225 264.060 113.825 ; 
                RECT 293.915 61.225 295.835 113.825 ; 
                RECT 297.755 61.225 299.675 113.825 ; 
                RECT 301.595 61.225 303.515 113.825 ; 
                RECT 305.435 61.225 307.355 113.825 ; 
                RECT 309.275 61.225 311.195 113.825 ; 
                RECT 264.515 164.320 265.835 191.440 ; 
                RECT 273.640 164.320 274.530 191.440 ; 
                RECT 280.075 164.320 281.185 191.440 ; 
                RECT 289.010 164.320 290.930 191.440 ; 
                RECT 309.790 164.320 311.710 191.440 ; 
                RECT 313.630 164.320 315.550 191.440 ; 
                RECT 317.470 164.320 319.390 191.440 ; 
                RECT 321.310 164.320 323.230 191.440 ; 
                RECT 263.975 147.420 265.085 158.320 ; 
                RECT 271.920 147.420 272.810 158.320 ; 
                RECT 278.895 147.420 280.215 158.320 ; 
                RECT 290.300 147.420 292.220 158.320 ; 
                RECT 313.230 147.420 315.150 158.320 ; 
                RECT 317.070 147.420 318.990 158.320 ; 
                RECT 320.910 147.420 322.830 158.320 ; 
                RECT 324.750 147.420 326.670 158.320 ; 
                RECT 338.880 50.065 339.770 55.225 ; 
                RECT 346.175 50.065 347.285 55.225 ; 
                RECT 355.110 50.065 357.030 55.225 ; 
                RECT 26.110 199.140 35.270 199.510 ; 
                RECT 26.110 202.475 35.270 203.365 ; 
                RECT 134.980 184.550 152.220 185.220 ; 
                RECT 134.980 185.880 152.220 187.230 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 1206.240 467.760 ; 
        LAYER met2 ;
            RECT 0.000 0.000 1206.240 467.760 ; 
    END 
END sram22_512x128m4w8 
END LIBRARY 

