VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_256x16m8w8
    CLASS BLOCK  ;
    FOREIGN sram22_256x16m8w8   ;
    SIZE 396.360 BY 225.680 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 210.910 0.000 211.050 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 221.810 0.000 221.950 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 232.710 0.000 232.850 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 243.610 0.000 243.750 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 254.510 0.000 254.650 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 265.410 0.000 265.550 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 276.310 0.000 276.450 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 287.210 0.000 287.350 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 298.110 0.000 298.250 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 309.010 0.000 309.150 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 319.910 0.000 320.050 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.810 0.000 330.950 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 341.710 0.000 341.850 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 352.610 0.000 352.750 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 363.510 0.000 363.650 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 374.410 0.000 374.550 0.140 ; 
        END 
    END dout[15] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 210.490 0.000 210.630 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 221.390 0.000 221.530 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 232.290 0.000 232.430 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 243.190 0.000 243.330 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 254.090 0.000 254.230 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 264.990 0.000 265.130 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 275.890 0.000 276.030 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 286.790 0.000 286.930 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 297.690 0.000 297.830 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 308.590 0.000 308.730 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 319.490 0.000 319.630 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.390 0.000 330.530 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 341.290 0.000 341.430 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 352.190 0.000 352.330 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 363.090 0.000 363.230 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.811200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 373.990 0.000 374.130 0.140 ; 
        END 
    END din[15] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.621600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 210.140 0.000 210.280 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.621600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 297.340 0.000 297.480 0.140 ; 
        END 
    END wmask[1] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 154.840 0.000 155.160 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 148.720 0.000 149.040 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 142.600 0.000 142.920 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 136.480 0.000 136.800 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 131.040 0.000 131.360 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 124.920 0.000 125.240 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 118.800 0.000 119.120 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 112.680 0.000 113.000 0.320 ; 
        END 
    END addr[7] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 167.080 0.000 167.400 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 160.960 0.000 161.280 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 12.834000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 170.480 0.000 170.800 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 16.740000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 171.160 0.000 171.480 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 210.240 6.240 ; 
                RECT 375.160 5.920 396.200 6.240 ; 
                RECT 0.160 7.280 396.200 7.600 ; 
                RECT 0.160 8.640 396.200 8.960 ; 
                RECT 0.160 10.000 170.120 10.320 ; 
                RECT 386.040 10.000 396.200 10.320 ; 
                RECT 0.160 11.360 197.320 11.680 ; 
                RECT 386.040 11.360 396.200 11.680 ; 
                RECT 0.160 12.720 197.320 13.040 ; 
                RECT 386.040 12.720 396.200 13.040 ; 
                RECT 0.160 14.080 197.320 14.400 ; 
                RECT 386.040 14.080 396.200 14.400 ; 
                RECT 0.160 15.440 197.320 15.760 ; 
                RECT 386.040 15.440 396.200 15.760 ; 
                RECT 0.160 16.800 197.320 17.120 ; 
                RECT 386.040 16.800 396.200 17.120 ; 
                RECT 0.160 18.160 197.320 18.480 ; 
                RECT 386.040 18.160 396.200 18.480 ; 
                RECT 0.160 19.520 197.320 19.840 ; 
                RECT 386.040 19.520 396.200 19.840 ; 
                RECT 0.160 20.880 108.240 21.200 ; 
                RECT 171.840 20.880 197.320 21.200 ; 
                RECT 386.040 20.880 396.200 21.200 ; 
                RECT 0.160 22.240 197.320 22.560 ; 
                RECT 386.040 22.240 396.200 22.560 ; 
                RECT 0.160 23.600 197.320 23.920 ; 
                RECT 386.040 23.600 396.200 23.920 ; 
                RECT 0.160 24.960 108.240 25.280 ; 
                RECT 171.160 24.960 197.320 25.280 ; 
                RECT 386.040 24.960 396.200 25.280 ; 
                RECT 0.160 26.320 197.320 26.640 ; 
                RECT 386.040 26.320 396.200 26.640 ; 
                RECT 0.160 27.680 196.640 28.000 ; 
                RECT 386.040 27.680 396.200 28.000 ; 
                RECT 0.160 29.040 197.320 29.360 ; 
                RECT 386.040 29.040 396.200 29.360 ; 
                RECT 0.160 30.400 197.320 30.720 ; 
                RECT 386.040 30.400 396.200 30.720 ; 
                RECT 0.160 31.760 197.320 32.080 ; 
                RECT 386.040 31.760 396.200 32.080 ; 
                RECT 0.160 33.120 197.320 33.440 ; 
                RECT 386.040 33.120 396.200 33.440 ; 
                RECT 0.160 34.480 197.320 34.800 ; 
                RECT 386.040 34.480 396.200 34.800 ; 
                RECT 0.160 35.840 197.320 36.160 ; 
                RECT 386.040 35.840 396.200 36.160 ; 
                RECT 0.160 37.200 197.320 37.520 ; 
                RECT 386.040 37.200 396.200 37.520 ; 
                RECT 0.160 38.560 197.320 38.880 ; 
                RECT 386.040 38.560 396.200 38.880 ; 
                RECT 0.160 39.920 132.040 40.240 ; 
                RECT 142.600 39.920 197.320 40.240 ; 
                RECT 386.040 39.920 396.200 40.240 ; 
                RECT 0.160 41.280 130.680 41.600 ; 
                RECT 148.720 41.280 197.320 41.600 ; 
                RECT 386.040 41.280 396.200 41.600 ; 
                RECT 0.160 42.640 129.320 42.960 ; 
                RECT 154.840 42.640 197.320 42.960 ; 
                RECT 386.040 42.640 396.200 42.960 ; 
                RECT 0.160 44.000 109.600 44.320 ; 
                RECT 171.840 44.000 197.320 44.320 ; 
                RECT 386.040 44.000 396.200 44.320 ; 
                RECT 0.160 45.360 108.920 45.680 ; 
                RECT 167.760 45.360 197.320 45.680 ; 
                RECT 386.040 45.360 396.200 45.680 ; 
                RECT 0.160 46.720 197.320 47.040 ; 
                RECT 386.040 46.720 396.200 47.040 ; 
                RECT 0.160 48.080 197.320 48.400 ; 
                RECT 386.040 48.080 396.200 48.400 ; 
                RECT 0.160 49.440 197.320 49.760 ; 
                RECT 386.040 49.440 396.200 49.760 ; 
                RECT 0.160 50.800 197.320 51.120 ; 
                RECT 386.040 50.800 396.200 51.120 ; 
                RECT 0.160 52.160 105.520 52.480 ; 
                RECT 116.080 52.160 164.000 52.480 ; 
                RECT 169.800 52.160 197.320 52.480 ; 
                RECT 386.040 52.160 396.200 52.480 ; 
                RECT 0.160 53.520 106.880 53.840 ; 
                RECT 109.960 53.520 164.000 53.840 ; 
                RECT 386.040 53.520 396.200 53.840 ; 
                RECT 0.160 54.880 108.240 55.200 ; 
                RECT 112.680 54.880 119.800 55.200 ; 
                RECT 122.880 54.880 164.000 55.200 ; 
                RECT 169.800 54.880 197.320 55.200 ; 
                RECT 386.040 54.880 396.200 55.200 ; 
                RECT 0.160 56.240 164.000 56.560 ; 
                RECT 169.800 56.240 197.320 56.560 ; 
                RECT 386.040 56.240 396.200 56.560 ; 
                RECT 0.160 57.600 114.360 57.920 ; 
                RECT 122.880 57.600 197.320 57.920 ; 
                RECT 386.040 57.600 396.200 57.920 ; 
                RECT 0.160 58.960 104.840 59.280 ; 
                RECT 116.080 58.960 197.320 59.280 ; 
                RECT 386.040 58.960 396.200 59.280 ; 
                RECT 0.160 60.320 110.960 60.640 ; 
                RECT 115.400 60.320 197.320 60.640 ; 
                RECT 386.040 60.320 396.200 60.640 ; 
                RECT 0.160 61.680 144.280 62.000 ; 
                RECT 169.120 61.680 197.320 62.000 ; 
                RECT 386.040 61.680 396.200 62.000 ; 
                RECT 0.160 63.040 106.880 63.360 ; 
                RECT 116.080 63.040 130.000 63.360 ; 
                RECT 137.160 63.040 144.280 63.360 ; 
                RECT 169.120 63.040 197.320 63.360 ; 
                RECT 386.040 63.040 396.200 63.360 ; 
                RECT 0.160 64.400 113.680 64.720 ; 
                RECT 122.200 64.400 131.360 64.720 ; 
                RECT 135.800 64.400 144.280 64.720 ; 
                RECT 178.640 64.400 197.320 64.720 ; 
                RECT 386.040 64.400 396.200 64.720 ; 
                RECT 0.160 65.760 132.720 66.080 ; 
                RECT 135.120 65.760 144.280 66.080 ; 
                RECT 178.640 65.760 197.320 66.080 ; 
                RECT 386.040 65.760 396.200 66.080 ; 
                RECT 0.160 67.120 114.360 67.440 ; 
                RECT 120.160 67.120 144.280 67.440 ; 
                RECT 181.360 67.120 197.320 67.440 ; 
                RECT 386.040 67.120 396.200 67.440 ; 
                RECT 0.160 68.480 117.080 68.800 ; 
                RECT 122.880 68.480 144.280 68.800 ; 
                RECT 180.000 68.480 197.320 68.800 ; 
                RECT 386.040 68.480 396.200 68.800 ; 
                RECT 0.160 69.840 110.960 70.160 ; 
                RECT 116.080 69.840 144.280 70.160 ; 
                RECT 181.360 69.840 197.320 70.160 ; 
                RECT 386.040 69.840 396.200 70.160 ; 
                RECT 0.160 71.200 144.280 71.520 ; 
                RECT 169.120 71.200 197.320 71.520 ; 
                RECT 386.040 71.200 396.200 71.520 ; 
                RECT 0.160 72.560 106.880 72.880 ; 
                RECT 127.640 72.560 144.280 72.880 ; 
                RECT 184.080 72.560 197.320 72.880 ; 
                RECT 386.040 72.560 396.200 72.880 ; 
                RECT 0.160 73.920 114.360 74.240 ; 
                RECT 122.880 73.920 144.280 74.240 ; 
                RECT 184.080 73.920 197.320 74.240 ; 
                RECT 386.040 73.920 396.200 74.240 ; 
                RECT 0.160 75.280 113.680 75.600 ; 
                RECT 116.080 75.280 123.200 75.600 ; 
                RECT 129.680 75.280 144.280 75.600 ; 
                RECT 182.720 75.280 197.320 75.600 ; 
                RECT 386.040 75.280 396.200 75.600 ; 
                RECT 0.160 76.640 105.520 76.960 ; 
                RECT 118.800 76.640 144.280 76.960 ; 
                RECT 186.800 76.640 197.320 76.960 ; 
                RECT 386.040 76.640 396.200 76.960 ; 
                RECT 0.160 78.000 113.680 78.320 ; 
                RECT 122.880 78.000 144.280 78.320 ; 
                RECT 186.800 78.000 197.320 78.320 ; 
                RECT 386.040 78.000 396.200 78.320 ; 
                RECT 0.160 79.360 144.280 79.680 ; 
                RECT 169.120 79.360 197.320 79.680 ; 
                RECT 386.040 79.360 396.200 79.680 ; 
                RECT 0.160 80.720 111.640 81.040 ; 
                RECT 122.880 80.720 144.280 81.040 ; 
                RECT 189.520 80.720 197.320 81.040 ; 
                RECT 386.040 80.720 396.200 81.040 ; 
                RECT 0.160 82.080 109.600 82.400 ; 
                RECT 113.360 82.080 144.280 82.400 ; 
                RECT 188.160 82.080 197.320 82.400 ; 
                RECT 386.040 82.080 396.200 82.400 ; 
                RECT 0.160 83.440 107.560 83.760 ; 
                RECT 109.960 83.440 144.280 83.760 ; 
                RECT 189.520 83.440 197.320 83.760 ; 
                RECT 386.040 83.440 396.200 83.760 ; 
                RECT 0.160 84.800 106.880 85.120 ; 
                RECT 116.080 84.800 144.280 85.120 ; 
                RECT 192.240 84.800 197.320 85.120 ; 
                RECT 386.040 84.800 396.200 85.120 ; 
                RECT 0.160 86.160 106.880 86.480 ; 
                RECT 121.520 86.160 144.280 86.480 ; 
                RECT 192.240 86.160 197.320 86.480 ; 
                RECT 386.040 86.160 396.200 86.480 ; 
                RECT 0.160 87.520 144.280 87.840 ; 
                RECT 190.880 87.520 197.320 87.840 ; 
                RECT 386.040 87.520 396.200 87.840 ; 
                RECT 0.160 88.880 113.680 89.200 ; 
                RECT 115.400 88.880 144.280 89.200 ; 
                RECT 169.120 88.880 197.320 89.200 ; 
                RECT 386.040 88.880 396.200 89.200 ; 
                RECT 0.160 90.240 114.360 90.560 ; 
                RECT 116.760 90.240 144.280 90.560 ; 
                RECT 193.600 90.240 197.320 90.560 ; 
                RECT 386.040 90.240 396.200 90.560 ; 
                RECT 0.160 91.600 105.520 91.920 ; 
                RECT 112.680 91.600 113.680 91.920 ; 
                RECT 115.400 91.600 144.280 91.920 ; 
                RECT 194.960 91.600 197.320 91.920 ; 
                RECT 386.040 91.600 396.200 91.920 ; 
                RECT 0.160 92.960 105.520 93.280 ; 
                RECT 116.080 92.960 144.280 93.280 ; 
                RECT 386.040 92.960 396.200 93.280 ; 
                RECT 0.160 94.320 108.240 94.640 ; 
                RECT 122.880 94.320 144.280 94.640 ; 
                RECT 386.040 94.320 396.200 94.640 ; 
                RECT 0.160 95.680 113.680 96.000 ; 
                RECT 116.760 95.680 120.480 96.000 ; 
                RECT 122.880 95.680 144.280 96.000 ; 
                RECT 386.040 95.680 396.200 96.000 ; 
                RECT 0.160 97.040 144.280 97.360 ; 
                RECT 169.120 97.040 197.320 97.360 ; 
                RECT 386.040 97.040 396.200 97.360 ; 
                RECT 0.160 98.400 197.320 98.720 ; 
                RECT 386.040 98.400 396.200 98.720 ; 
                RECT 0.160 99.760 101.440 100.080 ; 
                RECT 118.800 99.760 172.840 100.080 ; 
                RECT 386.040 99.760 396.200 100.080 ; 
                RECT 0.160 101.120 197.320 101.440 ; 
                RECT 386.040 101.120 396.200 101.440 ; 
                RECT 0.160 102.480 191.880 102.800 ; 
                RECT 386.040 102.480 396.200 102.800 ; 
                RECT 0.160 103.840 108.240 104.160 ; 
                RECT 112.000 103.840 189.160 104.160 ; 
                RECT 386.040 103.840 396.200 104.160 ; 
                RECT 0.160 105.200 117.080 105.520 ; 
                RECT 124.920 105.200 186.440 105.520 ; 
                RECT 386.040 105.200 396.200 105.520 ; 
                RECT 0.160 106.560 108.240 106.880 ; 
                RECT 122.880 106.560 183.720 106.880 ; 
                RECT 386.040 106.560 396.200 106.880 ; 
                RECT 0.160 107.920 181.000 108.240 ; 
                RECT 386.040 107.920 396.200 108.240 ; 
                RECT 0.160 109.280 105.520 109.600 ; 
                RECT 108.600 109.280 178.280 109.600 ; 
                RECT 386.040 109.280 396.200 109.600 ; 
                RECT 0.160 110.640 144.960 110.960 ; 
                RECT 167.760 110.640 175.560 110.960 ; 
                RECT 386.040 110.640 396.200 110.960 ; 
                RECT 0.160 112.000 83.760 112.320 ; 
                RECT 101.800 112.000 110.960 112.320 ; 
                RECT 113.360 112.000 144.960 112.320 ; 
                RECT 167.760 112.000 197.320 112.320 ; 
                RECT 386.040 112.000 396.200 112.320 ; 
                RECT 0.160 113.360 83.760 113.680 ; 
                RECT 101.800 113.360 144.960 113.680 ; 
                RECT 167.760 113.360 197.320 113.680 ; 
                RECT 386.040 113.360 396.200 113.680 ; 
                RECT 0.160 114.720 83.760 115.040 ; 
                RECT 101.800 114.720 144.960 115.040 ; 
                RECT 167.760 114.720 197.320 115.040 ; 
                RECT 386.040 114.720 396.200 115.040 ; 
                RECT 0.160 116.080 83.760 116.400 ; 
                RECT 101.800 116.080 120.480 116.400 ; 
                RECT 122.880 116.080 144.960 116.400 ; 
                RECT 167.760 116.080 197.320 116.400 ; 
                RECT 386.040 116.080 396.200 116.400 ; 
                RECT 0.160 117.440 83.760 117.760 ; 
                RECT 101.800 117.440 109.600 117.760 ; 
                RECT 112.680 117.440 144.960 117.760 ; 
                RECT 167.760 117.440 197.320 117.760 ; 
                RECT 386.040 117.440 396.200 117.760 ; 
                RECT 0.160 118.800 83.760 119.120 ; 
                RECT 101.800 118.800 106.880 119.120 ; 
                RECT 113.360 118.800 144.960 119.120 ; 
                RECT 167.760 118.800 197.320 119.120 ; 
                RECT 386.040 118.800 396.200 119.120 ; 
                RECT 0.160 120.160 83.760 120.480 ; 
                RECT 101.800 120.160 176.920 120.480 ; 
                RECT 386.040 120.160 396.200 120.480 ; 
                RECT 0.160 121.520 83.760 121.840 ; 
                RECT 101.800 121.520 176.920 121.840 ; 
                RECT 386.040 121.520 396.200 121.840 ; 
                RECT 0.160 122.880 83.760 123.200 ; 
                RECT 101.800 122.880 179.640 123.200 ; 
                RECT 386.040 122.880 396.200 123.200 ; 
                RECT 0.160 124.240 83.760 124.560 ; 
                RECT 101.800 124.240 113.680 124.560 ; 
                RECT 122.200 124.240 185.080 124.560 ; 
                RECT 386.040 124.240 396.200 124.560 ; 
                RECT 0.160 125.600 83.760 125.920 ; 
                RECT 101.800 125.600 106.880 125.920 ; 
                RECT 109.960 125.600 144.280 125.920 ; 
                RECT 167.760 125.600 187.800 125.920 ; 
                RECT 386.040 125.600 396.200 125.920 ; 
                RECT 0.160 126.960 144.280 127.280 ; 
                RECT 167.760 126.960 190.520 127.280 ; 
                RECT 386.040 126.960 396.200 127.280 ; 
                RECT 0.160 128.320 104.840 128.640 ; 
                RECT 112.680 128.320 144.280 128.640 ; 
                RECT 167.760 128.320 193.240 128.640 ; 
                RECT 386.040 128.320 396.200 128.640 ; 
                RECT 0.160 129.680 144.280 130.000 ; 
                RECT 167.760 129.680 195.960 130.000 ; 
                RECT 386.040 129.680 396.200 130.000 ; 
                RECT 0.160 131.040 67.440 131.360 ; 
                RECT 83.440 131.040 144.280 131.360 ; 
                RECT 386.040 131.040 396.200 131.360 ; 
                RECT 0.160 132.400 67.440 132.720 ; 
                RECT 83.440 132.400 110.960 132.720 ; 
                RECT 116.760 132.400 144.280 132.720 ; 
                RECT 167.760 132.400 197.320 132.720 ; 
                RECT 386.040 132.400 396.200 132.720 ; 
                RECT 0.160 133.760 67.440 134.080 ; 
                RECT 83.440 133.760 89.200 134.080 ; 
                RECT 97.040 133.760 144.280 134.080 ; 
                RECT 167.760 133.760 197.320 134.080 ; 
                RECT 386.040 133.760 396.200 134.080 ; 
                RECT 0.160 135.120 67.440 135.440 ; 
                RECT 101.120 135.120 144.280 135.440 ; 
                RECT 167.760 135.120 197.320 135.440 ; 
                RECT 386.040 135.120 396.200 135.440 ; 
                RECT 0.160 136.480 67.440 136.800 ; 
                RECT 101.120 136.480 144.280 136.800 ; 
                RECT 386.040 136.480 396.200 136.800 ; 
                RECT 0.160 137.840 67.440 138.160 ; 
                RECT 83.440 137.840 89.200 138.160 ; 
                RECT 97.040 137.840 106.880 138.160 ; 
                RECT 115.400 137.840 144.280 138.160 ; 
                RECT 386.040 137.840 396.200 138.160 ; 
                RECT 0.160 139.200 62.000 139.520 ; 
                RECT 96.360 139.200 144.280 139.520 ; 
                RECT 167.760 139.200 396.200 139.520 ; 
                RECT 0.160 140.560 96.000 140.880 ; 
                RECT 141.920 140.560 396.200 140.880 ; 
                RECT 0.160 141.920 194.600 142.240 ; 
                RECT 388.760 141.920 396.200 142.240 ; 
                RECT 0.160 143.280 194.600 143.600 ; 
                RECT 388.760 143.280 396.200 143.600 ; 
                RECT 0.160 144.640 194.600 144.960 ; 
                RECT 388.760 144.640 396.200 144.960 ; 
                RECT 0.160 146.000 24.600 146.320 ; 
                RECT 31.080 146.000 33.440 146.320 ; 
                RECT 44.680 146.000 72.880 146.320 ; 
                RECT 388.760 146.000 396.200 146.320 ; 
                RECT 0.160 147.360 22.560 147.680 ; 
                RECT 33.120 147.360 34.800 147.680 ; 
                RECT 43.320 147.360 57.240 147.680 ; 
                RECT 63.040 147.360 72.880 147.680 ; 
                RECT 388.760 147.360 396.200 147.680 ; 
                RECT 0.160 148.720 22.560 149.040 ; 
                RECT 33.120 148.720 36.160 149.040 ; 
                RECT 42.640 148.720 55.200 149.040 ; 
                RECT 63.040 148.720 72.880 149.040 ; 
                RECT 388.760 148.720 396.200 149.040 ; 
                RECT 0.160 150.080 22.560 150.400 ; 
                RECT 33.120 150.080 55.200 150.400 ; 
                RECT 58.960 150.080 72.880 150.400 ; 
                RECT 388.760 150.080 396.200 150.400 ; 
                RECT 0.160 151.440 55.200 151.760 ; 
                RECT 63.040 151.440 72.880 151.760 ; 
                RECT 388.760 151.440 396.200 151.760 ; 
                RECT 0.160 152.800 22.560 153.120 ; 
                RECT 33.120 152.800 55.200 153.120 ; 
                RECT 63.040 152.800 72.880 153.120 ; 
                RECT 388.760 152.800 396.200 153.120 ; 
                RECT 0.160 154.160 22.560 154.480 ; 
                RECT 33.120 154.160 72.880 154.480 ; 
                RECT 388.760 154.160 396.200 154.480 ; 
                RECT 0.160 155.520 59.280 155.840 ; 
                RECT 63.040 155.520 72.880 155.840 ; 
                RECT 388.760 155.520 396.200 155.840 ; 
                RECT 0.160 156.880 55.200 157.200 ; 
                RECT 63.040 156.880 72.880 157.200 ; 
                RECT 388.760 156.880 396.200 157.200 ; 
                RECT 0.160 158.240 55.200 158.560 ; 
                RECT 63.040 158.240 72.880 158.560 ; 
                RECT 388.760 158.240 396.200 158.560 ; 
                RECT 0.160 159.600 15.760 159.920 ; 
                RECT 18.160 159.600 31.400 159.920 ; 
                RECT 34.480 159.600 55.200 159.920 ; 
                RECT 56.920 159.600 72.880 159.920 ; 
                RECT 388.760 159.600 396.200 159.920 ; 
                RECT 0.160 160.960 15.080 161.280 ; 
                RECT 18.160 160.960 31.400 161.280 ; 
                RECT 35.160 160.960 55.200 161.280 ; 
                RECT 63.040 160.960 72.880 161.280 ; 
                RECT 388.760 160.960 396.200 161.280 ; 
                RECT 0.160 162.320 14.400 162.640 ; 
                RECT 18.160 162.320 72.880 162.640 ; 
                RECT 388.760 162.320 396.200 162.640 ; 
                RECT 0.160 163.680 13.720 164.000 ; 
                RECT 18.160 163.680 57.240 164.000 ; 
                RECT 63.040 163.680 72.880 164.000 ; 
                RECT 388.760 163.680 396.200 164.000 ; 
                RECT 0.160 165.040 55.200 165.360 ; 
                RECT 63.040 165.040 72.880 165.360 ; 
                RECT 388.760 165.040 396.200 165.360 ; 
                RECT 0.160 166.400 13.040 166.720 ; 
                RECT 18.160 166.400 55.200 166.720 ; 
                RECT 63.040 166.400 72.880 166.720 ; 
                RECT 388.760 166.400 396.200 166.720 ; 
                RECT 0.160 167.760 12.360 168.080 ; 
                RECT 18.160 167.760 55.200 168.080 ; 
                RECT 63.040 167.760 72.880 168.080 ; 
                RECT 388.760 167.760 396.200 168.080 ; 
                RECT 0.160 169.120 55.200 169.440 ; 
                RECT 61.680 169.120 72.880 169.440 ; 
                RECT 388.760 169.120 396.200 169.440 ; 
                RECT 0.160 170.480 11.680 170.800 ; 
                RECT 18.160 170.480 72.880 170.800 ; 
                RECT 388.760 170.480 396.200 170.800 ; 
                RECT 0.160 171.840 11.000 172.160 ; 
                RECT 18.160 171.840 31.400 172.160 ; 
                RECT 35.840 171.840 55.200 172.160 ; 
                RECT 63.040 171.840 72.880 172.160 ; 
                RECT 388.760 171.840 396.200 172.160 ; 
                RECT 0.160 173.200 55.200 173.520 ; 
                RECT 63.040 173.200 72.880 173.520 ; 
                RECT 388.760 173.200 396.200 173.520 ; 
                RECT 0.160 174.560 10.320 174.880 ; 
                RECT 18.160 174.560 31.400 174.880 ; 
                RECT 35.160 174.560 55.200 174.880 ; 
                RECT 63.040 174.560 72.880 174.880 ; 
                RECT 388.760 174.560 396.200 174.880 ; 
                RECT 0.160 175.920 9.640 176.240 ; 
                RECT 18.160 175.920 31.400 176.240 ; 
                RECT 34.480 175.920 55.200 176.240 ; 
                RECT 63.040 175.920 72.880 176.240 ; 
                RECT 388.760 175.920 396.200 176.240 ; 
                RECT 0.160 177.280 55.200 177.600 ; 
                RECT 62.360 177.280 72.880 177.600 ; 
                RECT 388.760 177.280 396.200 177.600 ; 
                RECT 0.160 178.640 57.240 178.960 ; 
                RECT 63.040 178.640 72.880 178.960 ; 
                RECT 388.760 178.640 396.200 178.960 ; 
                RECT 0.160 180.000 72.880 180.320 ; 
                RECT 388.760 180.000 396.200 180.320 ; 
                RECT 0.160 181.360 57.920 181.680 ; 
                RECT 63.040 181.360 72.880 181.680 ; 
                RECT 388.760 181.360 396.200 181.680 ; 
                RECT 0.160 182.720 58.600 183.040 ; 
                RECT 63.040 182.720 72.880 183.040 ; 
                RECT 388.760 182.720 396.200 183.040 ; 
                RECT 0.160 184.080 59.280 184.400 ; 
                RECT 63.040 184.080 72.880 184.400 ; 
                RECT 388.760 184.080 396.200 184.400 ; 
                RECT 0.160 185.440 35.480 185.760 ; 
                RECT 44.000 185.440 72.880 185.760 ; 
                RECT 388.760 185.440 396.200 185.760 ; 
                RECT 0.160 186.800 34.120 187.120 ; 
                RECT 42.640 186.800 55.200 187.120 ; 
                RECT 63.040 186.800 72.880 187.120 ; 
                RECT 388.760 186.800 396.200 187.120 ; 
                RECT 0.160 188.160 55.200 188.480 ; 
                RECT 63.040 188.160 72.880 188.480 ; 
                RECT 388.760 188.160 396.200 188.480 ; 
                RECT 0.160 189.520 55.200 189.840 ; 
                RECT 57.600 189.520 72.880 189.840 ; 
                RECT 388.760 189.520 396.200 189.840 ; 
                RECT 0.160 190.880 55.200 191.200 ; 
                RECT 63.040 190.880 72.880 191.200 ; 
                RECT 388.760 190.880 396.200 191.200 ; 
                RECT 0.160 192.240 55.200 192.560 ; 
                RECT 63.040 192.240 72.880 192.560 ; 
                RECT 388.760 192.240 396.200 192.560 ; 
                RECT 0.160 193.600 55.200 193.920 ; 
                RECT 58.960 193.600 72.880 193.920 ; 
                RECT 388.760 193.600 396.200 193.920 ; 
                RECT 0.160 194.960 57.240 195.280 ; 
                RECT 63.040 194.960 72.880 195.280 ; 
                RECT 388.760 194.960 396.200 195.280 ; 
                RECT 0.160 196.320 57.920 196.640 ; 
                RECT 63.040 196.320 72.880 196.640 ; 
                RECT 388.760 196.320 396.200 196.640 ; 
                RECT 0.160 197.680 58.600 198.000 ; 
                RECT 63.040 197.680 72.880 198.000 ; 
                RECT 388.760 197.680 396.200 198.000 ; 
                RECT 0.160 199.040 72.880 199.360 ; 
                RECT 388.760 199.040 396.200 199.360 ; 
                RECT 0.160 200.400 59.280 200.720 ; 
                RECT 63.040 200.400 72.880 200.720 ; 
                RECT 388.760 200.400 396.200 200.720 ; 
                RECT 0.160 201.760 72.880 202.080 ; 
                RECT 388.760 201.760 396.200 202.080 ; 
                RECT 0.160 203.120 59.280 203.440 ; 
                RECT 63.040 203.120 72.880 203.440 ; 
                RECT 388.760 203.120 396.200 203.440 ; 
                RECT 0.160 204.480 59.960 204.800 ; 
                RECT 63.040 204.480 72.880 204.800 ; 
                RECT 388.760 204.480 396.200 204.800 ; 
                RECT 0.160 205.840 60.640 206.160 ; 
                RECT 63.040 205.840 72.880 206.160 ; 
                RECT 388.760 205.840 396.200 206.160 ; 
                RECT 0.160 207.200 60.640 207.520 ; 
                RECT 63.040 207.200 72.880 207.520 ; 
                RECT 388.760 207.200 396.200 207.520 ; 
                RECT 0.160 208.560 72.880 208.880 ; 
                RECT 388.760 208.560 396.200 208.880 ; 
                RECT 0.160 209.920 72.880 210.240 ; 
                RECT 388.760 209.920 396.200 210.240 ; 
                RECT 0.160 211.280 194.600 211.600 ; 
                RECT 388.760 211.280 396.200 211.600 ; 
                RECT 0.160 212.640 194.600 212.960 ; 
                RECT 388.760 212.640 396.200 212.960 ; 
                RECT 0.160 214.000 194.600 214.320 ; 
                RECT 388.760 214.000 396.200 214.320 ; 
                RECT 0.160 215.360 396.200 215.680 ; 
                RECT 0.160 216.720 396.200 217.040 ; 
                RECT 0.160 218.080 396.200 218.400 ; 
                RECT 0.160 219.440 396.200 219.760 ; 
                RECT 0.160 0.160 396.200 1.520 ; 
                RECT 0.160 224.160 396.200 225.520 ; 
                RECT 198.740 32.080 204.540 33.450 ; 
                RECT 378.640 32.080 384.440 33.450 ; 
                RECT 198.740 37.195 204.540 38.615 ; 
                RECT 378.640 37.195 384.440 38.615 ; 
                RECT 198.740 42.515 204.540 44.035 ; 
                RECT 378.640 42.515 384.440 44.035 ; 
                RECT 198.740 47.985 204.540 49.505 ; 
                RECT 378.640 47.985 384.440 49.505 ; 
                RECT 198.740 75.760 384.440 76.560 ; 
                RECT 198.740 67.860 384.440 68.660 ; 
                RECT 198.740 82.075 384.440 83.145 ; 
                RECT 198.740 70.870 384.440 71.670 ; 
                RECT 198.740 133.920 384.440 135.270 ; 
                RECT 198.740 113.670 384.440 114.640 ; 
                RECT 198.740 86.365 384.440 86.655 ; 
                RECT 198.740 56.390 384.440 58.190 ; 
                RECT 198.740 16.325 384.440 18.125 ; 
                RECT 78.110 145.715 80.030 210.495 ; 
                RECT 88.985 145.715 90.905 210.495 ; 
                RECT 92.825 145.715 94.745 210.495 ; 
                RECT 96.665 145.715 98.585 210.495 ; 
                RECT 112.330 145.715 114.250 210.495 ; 
                RECT 116.170 145.715 118.090 210.495 ; 
                RECT 120.010 145.715 121.930 210.495 ; 
                RECT 123.850 145.715 125.770 210.495 ; 
                RECT 127.690 145.715 129.610 210.495 ; 
                RECT 152.290 145.715 154.210 210.495 ; 
                RECT 156.130 145.715 158.050 210.495 ; 
                RECT 159.970 145.715 161.890 210.495 ; 
                RECT 163.810 145.715 165.730 210.495 ; 
                RECT 167.650 145.715 169.570 210.495 ; 
                RECT 171.490 145.715 173.410 210.495 ; 
                RECT 175.330 145.715 177.250 210.495 ; 
                RECT 179.170 145.715 181.090 210.495 ; 
                RECT 183.010 145.715 184.930 210.495 ; 
                RECT 186.850 145.715 188.770 210.495 ; 
                RECT 190.690 145.715 192.610 210.495 ; 
                RECT 147.315 61.965 149.235 97.365 ; 
                RECT 154.075 61.965 155.995 97.365 ; 
                RECT 162.785 61.965 164.705 97.365 ; 
                RECT 166.625 61.965 168.545 97.365 ; 
                RECT 148.800 125.020 150.720 139.080 ; 
                RECT 156.075 125.020 157.825 139.080 ; 
                RECT 165.330 125.020 167.250 139.080 ; 
                RECT 148.800 110.700 150.720 119.020 ; 
                RECT 155.775 110.700 157.695 119.020 ; 
                RECT 165.330 110.700 167.250 119.020 ; 
                RECT 167.155 52.385 168.905 55.965 ; 
                RECT 23.460 147.985 32.620 148.735 ; 
                RECT 23.460 152.740 32.620 154.660 ; 
                RECT 84.700 135.770 100.740 136.570 ; 
                RECT 67.900 135.125 82.740 138.175 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 210.240 5.560 ; 
                RECT 375.160 5.240 393.480 5.560 ; 
                RECT 2.880 6.600 393.480 6.920 ; 
                RECT 2.880 7.960 393.480 8.280 ; 
                RECT 2.880 9.320 170.800 9.640 ; 
                RECT 203.120 9.320 393.480 9.640 ; 
                RECT 2.880 10.680 197.320 11.000 ; 
                RECT 386.040 10.680 393.480 11.000 ; 
                RECT 2.880 12.040 197.320 12.360 ; 
                RECT 386.040 12.040 393.480 12.360 ; 
                RECT 2.880 13.400 197.320 13.720 ; 
                RECT 386.040 13.400 393.480 13.720 ; 
                RECT 2.880 14.760 197.320 15.080 ; 
                RECT 386.040 14.760 393.480 15.080 ; 
                RECT 2.880 16.120 197.320 16.440 ; 
                RECT 386.040 16.120 393.480 16.440 ; 
                RECT 2.880 17.480 197.320 17.800 ; 
                RECT 386.040 17.480 393.480 17.800 ; 
                RECT 2.880 18.840 197.320 19.160 ; 
                RECT 386.040 18.840 393.480 19.160 ; 
                RECT 2.880 20.200 108.240 20.520 ; 
                RECT 171.840 20.200 197.320 20.520 ; 
                RECT 386.040 20.200 393.480 20.520 ; 
                RECT 2.880 21.560 197.320 21.880 ; 
                RECT 386.040 21.560 393.480 21.880 ; 
                RECT 2.880 22.920 197.320 23.240 ; 
                RECT 386.040 22.920 393.480 23.240 ; 
                RECT 2.880 24.280 108.240 24.600 ; 
                RECT 171.160 24.280 197.320 24.600 ; 
                RECT 386.040 24.280 393.480 24.600 ; 
                RECT 2.880 25.640 197.320 25.960 ; 
                RECT 386.040 25.640 393.480 25.960 ; 
                RECT 2.880 27.000 197.320 27.320 ; 
                RECT 386.040 27.000 393.480 27.320 ; 
                RECT 2.880 28.360 196.640 28.680 ; 
                RECT 386.040 28.360 393.480 28.680 ; 
                RECT 2.880 29.720 197.320 30.040 ; 
                RECT 386.040 29.720 393.480 30.040 ; 
                RECT 2.880 31.080 197.320 31.400 ; 
                RECT 386.040 31.080 393.480 31.400 ; 
                RECT 2.880 32.440 197.320 32.760 ; 
                RECT 386.040 32.440 393.480 32.760 ; 
                RECT 2.880 33.800 197.320 34.120 ; 
                RECT 386.040 33.800 393.480 34.120 ; 
                RECT 2.880 35.160 197.320 35.480 ; 
                RECT 386.040 35.160 393.480 35.480 ; 
                RECT 2.880 36.520 197.320 36.840 ; 
                RECT 386.040 36.520 393.480 36.840 ; 
                RECT 2.880 37.880 197.320 38.200 ; 
                RECT 386.040 37.880 393.480 38.200 ; 
                RECT 2.880 39.240 132.720 39.560 ; 
                RECT 143.960 39.240 197.320 39.560 ; 
                RECT 386.040 39.240 393.480 39.560 ; 
                RECT 2.880 40.600 131.360 40.920 ; 
                RECT 150.080 40.600 197.320 40.920 ; 
                RECT 386.040 40.600 393.480 40.920 ; 
                RECT 2.880 41.960 130.000 42.280 ; 
                RECT 156.200 41.960 197.320 42.280 ; 
                RECT 386.040 41.960 393.480 42.280 ; 
                RECT 2.880 43.320 106.880 43.640 ; 
                RECT 171.160 43.320 197.320 43.640 ; 
                RECT 386.040 43.320 393.480 43.640 ; 
                RECT 2.880 44.680 108.240 45.000 ; 
                RECT 161.640 44.680 197.320 45.000 ; 
                RECT 386.040 44.680 393.480 45.000 ; 
                RECT 2.880 46.040 197.320 46.360 ; 
                RECT 386.040 46.040 393.480 46.360 ; 
                RECT 2.880 47.400 197.320 47.720 ; 
                RECT 386.040 47.400 393.480 47.720 ; 
                RECT 2.880 48.760 197.320 49.080 ; 
                RECT 386.040 48.760 393.480 49.080 ; 
                RECT 2.880 50.120 197.320 50.440 ; 
                RECT 386.040 50.120 393.480 50.440 ; 
                RECT 2.880 51.480 105.520 51.800 ; 
                RECT 116.080 51.480 197.320 51.800 ; 
                RECT 386.040 51.480 393.480 51.800 ; 
                RECT 2.880 52.840 106.880 53.160 ; 
                RECT 108.600 52.840 164.000 53.160 ; 
                RECT 169.800 52.840 197.320 53.160 ; 
                RECT 386.040 52.840 393.480 53.160 ; 
                RECT 2.880 54.200 108.240 54.520 ; 
                RECT 112.680 54.200 119.800 54.520 ; 
                RECT 122.880 54.200 164.000 54.520 ; 
                RECT 386.040 54.200 393.480 54.520 ; 
                RECT 2.880 55.560 108.240 55.880 ; 
                RECT 111.320 55.560 127.960 55.880 ; 
                RECT 160.960 55.560 164.000 55.880 ; 
                RECT 169.800 55.560 197.320 55.880 ; 
                RECT 386.040 55.560 393.480 55.880 ; 
                RECT 2.880 56.920 114.360 57.240 ; 
                RECT 122.880 56.920 197.320 57.240 ; 
                RECT 386.040 56.920 393.480 57.240 ; 
                RECT 2.880 58.280 104.840 58.600 ; 
                RECT 116.080 58.280 197.320 58.600 ; 
                RECT 386.040 58.280 393.480 58.600 ; 
                RECT 2.880 59.640 106.880 59.960 ; 
                RECT 116.080 59.640 197.320 59.960 ; 
                RECT 386.040 59.640 393.480 59.960 ; 
                RECT 2.880 61.000 197.320 61.320 ; 
                RECT 386.040 61.000 393.480 61.320 ; 
                RECT 2.880 62.360 106.880 62.680 ; 
                RECT 116.080 62.360 129.320 62.680 ; 
                RECT 137.840 62.360 144.280 62.680 ; 
                RECT 169.120 62.360 197.320 62.680 ; 
                RECT 386.040 62.360 393.480 62.680 ; 
                RECT 2.880 63.720 114.360 64.040 ; 
                RECT 122.200 63.720 130.680 64.040 ; 
                RECT 136.480 63.720 144.280 64.040 ; 
                RECT 178.640 63.720 197.320 64.040 ; 
                RECT 386.040 63.720 393.480 64.040 ; 
                RECT 2.880 65.080 113.680 65.400 ; 
                RECT 116.080 65.080 132.040 65.400 ; 
                RECT 135.800 65.080 144.280 65.400 ; 
                RECT 178.640 65.080 197.320 65.400 ; 
                RECT 386.040 65.080 393.480 65.400 ; 
                RECT 2.880 66.440 144.280 66.760 ; 
                RECT 177.280 66.440 197.320 66.760 ; 
                RECT 386.040 66.440 393.480 66.760 ; 
                RECT 2.880 67.800 114.360 68.120 ; 
                RECT 122.880 67.800 144.280 68.120 ; 
                RECT 181.360 67.800 197.320 68.120 ; 
                RECT 386.040 67.800 393.480 68.120 ; 
                RECT 2.880 69.160 110.960 69.480 ; 
                RECT 116.080 69.160 144.280 69.480 ; 
                RECT 181.360 69.160 197.320 69.480 ; 
                RECT 386.040 69.160 393.480 69.480 ; 
                RECT 2.880 70.520 113.680 70.840 ; 
                RECT 116.080 70.520 144.280 70.840 ; 
                RECT 180.000 70.520 197.320 70.840 ; 
                RECT 386.040 70.520 393.480 70.840 ; 
                RECT 2.880 71.880 144.280 72.200 ; 
                RECT 184.080 71.880 197.320 72.200 ; 
                RECT 386.040 71.880 393.480 72.200 ; 
                RECT 2.880 73.240 106.880 73.560 ; 
                RECT 127.640 73.240 144.280 73.560 ; 
                RECT 182.720 73.240 197.320 73.560 ; 
                RECT 386.040 73.240 393.480 73.560 ; 
                RECT 2.880 74.600 123.200 74.920 ; 
                RECT 129.000 74.600 144.280 74.920 ; 
                RECT 184.080 74.600 197.320 74.920 ; 
                RECT 386.040 74.600 393.480 74.920 ; 
                RECT 2.880 75.960 113.680 76.280 ; 
                RECT 116.080 75.960 125.920 76.280 ; 
                RECT 129.680 75.960 144.280 76.280 ; 
                RECT 186.800 75.960 197.320 76.280 ; 
                RECT 386.040 75.960 393.480 76.280 ; 
                RECT 2.880 77.320 105.520 77.640 ; 
                RECT 118.800 77.320 144.280 77.640 ; 
                RECT 185.440 77.320 197.320 77.640 ; 
                RECT 386.040 77.320 393.480 77.640 ; 
                RECT 2.880 78.680 113.680 79.000 ; 
                RECT 122.880 78.680 144.280 79.000 ; 
                RECT 186.800 78.680 197.320 79.000 ; 
                RECT 386.040 78.680 393.480 79.000 ; 
                RECT 2.880 80.040 111.640 80.360 ; 
                RECT 122.880 80.040 144.280 80.360 ; 
                RECT 169.120 80.040 197.320 80.360 ; 
                RECT 386.040 80.040 393.480 80.360 ; 
                RECT 2.880 81.400 109.600 81.720 ; 
                RECT 113.360 81.400 144.280 81.720 ; 
                RECT 189.520 81.400 197.320 81.720 ; 
                RECT 386.040 81.400 393.480 81.720 ; 
                RECT 2.880 82.760 144.280 83.080 ; 
                RECT 189.520 82.760 197.320 83.080 ; 
                RECT 386.040 82.760 393.480 83.080 ; 
                RECT 2.880 84.120 106.880 84.440 ; 
                RECT 109.960 84.120 144.280 84.440 ; 
                RECT 169.120 84.120 197.320 84.440 ; 
                RECT 386.040 84.120 393.480 84.440 ; 
                RECT 2.880 85.480 106.880 85.800 ; 
                RECT 116.080 85.480 144.280 85.800 ; 
                RECT 190.880 85.480 197.320 85.800 ; 
                RECT 386.040 85.480 393.480 85.800 ; 
                RECT 2.880 86.840 110.960 87.160 ; 
                RECT 121.520 86.840 144.280 87.160 ; 
                RECT 192.240 86.840 197.320 87.160 ; 
                RECT 386.040 86.840 393.480 87.160 ; 
                RECT 2.880 88.200 113.680 88.520 ; 
                RECT 115.400 88.200 144.280 88.520 ; 
                RECT 169.120 88.200 197.320 88.520 ; 
                RECT 386.040 88.200 393.480 88.520 ; 
                RECT 2.880 89.560 114.360 89.880 ; 
                RECT 116.760 89.560 144.280 89.880 ; 
                RECT 194.960 89.560 197.320 89.880 ; 
                RECT 386.040 89.560 393.480 89.880 ; 
                RECT 2.880 90.920 144.280 91.240 ; 
                RECT 194.960 90.920 197.320 91.240 ; 
                RECT 386.040 90.920 393.480 91.240 ; 
                RECT 2.880 92.280 105.520 92.600 ; 
                RECT 115.400 92.280 144.280 92.600 ; 
                RECT 193.600 92.280 197.320 92.600 ; 
                RECT 386.040 92.280 393.480 92.600 ; 
                RECT 2.880 93.640 108.240 93.960 ; 
                RECT 122.880 93.640 144.280 93.960 ; 
                RECT 386.040 93.640 393.480 93.960 ; 
                RECT 2.880 95.000 113.680 95.320 ; 
                RECT 116.760 95.000 144.280 95.320 ; 
                RECT 386.040 95.000 393.480 95.320 ; 
                RECT 2.880 96.360 120.480 96.680 ; 
                RECT 122.880 96.360 144.280 96.680 ; 
                RECT 386.040 96.360 393.480 96.680 ; 
                RECT 2.880 97.720 144.280 98.040 ; 
                RECT 169.120 97.720 197.320 98.040 ; 
                RECT 386.040 97.720 393.480 98.040 ; 
                RECT 2.880 99.080 101.440 99.400 ; 
                RECT 115.400 99.080 197.320 99.400 ; 
                RECT 386.040 99.080 393.480 99.400 ; 
                RECT 2.880 100.440 111.640 100.760 ; 
                RECT 118.800 100.440 172.840 100.760 ; 
                RECT 386.040 100.440 393.480 100.760 ; 
                RECT 2.880 101.800 194.600 102.120 ; 
                RECT 386.040 101.800 393.480 102.120 ; 
                RECT 2.880 103.160 108.240 103.480 ; 
                RECT 112.000 103.160 191.880 103.480 ; 
                RECT 386.040 103.160 393.480 103.480 ; 
                RECT 2.880 104.520 117.080 104.840 ; 
                RECT 124.920 104.520 189.160 104.840 ; 
                RECT 386.040 104.520 393.480 104.840 ; 
                RECT 2.880 105.880 186.440 106.200 ; 
                RECT 386.040 105.880 393.480 106.200 ; 
                RECT 2.880 107.240 108.240 107.560 ; 
                RECT 122.880 107.240 183.720 107.560 ; 
                RECT 386.040 107.240 393.480 107.560 ; 
                RECT 2.880 108.600 181.000 108.920 ; 
                RECT 386.040 108.600 393.480 108.920 ; 
                RECT 2.880 109.960 105.520 110.280 ; 
                RECT 108.600 109.960 175.560 110.280 ; 
                RECT 386.040 109.960 393.480 110.280 ; 
                RECT 2.880 111.320 110.960 111.640 ; 
                RECT 113.360 111.320 128.640 111.640 ; 
                RECT 141.920 111.320 144.960 111.640 ; 
                RECT 167.760 111.320 175.560 111.640 ; 
                RECT 386.040 111.320 393.480 111.640 ; 
                RECT 2.880 112.680 83.760 113.000 ; 
                RECT 101.800 112.680 144.960 113.000 ; 
                RECT 167.760 112.680 197.320 113.000 ; 
                RECT 386.040 112.680 393.480 113.000 ; 
                RECT 2.880 114.040 83.760 114.360 ; 
                RECT 101.800 114.040 144.960 114.360 ; 
                RECT 167.760 114.040 197.320 114.360 ; 
                RECT 386.040 114.040 393.480 114.360 ; 
                RECT 2.880 115.400 83.760 115.720 ; 
                RECT 101.800 115.400 120.480 115.720 ; 
                RECT 122.880 115.400 144.960 115.720 ; 
                RECT 167.760 115.400 197.320 115.720 ; 
                RECT 386.040 115.400 393.480 115.720 ; 
                RECT 2.880 116.760 83.760 117.080 ; 
                RECT 101.800 116.760 109.600 117.080 ; 
                RECT 112.680 116.760 144.960 117.080 ; 
                RECT 167.760 116.760 197.320 117.080 ; 
                RECT 386.040 116.760 393.480 117.080 ; 
                RECT 2.880 118.120 83.760 118.440 ; 
                RECT 102.480 118.120 106.880 118.440 ; 
                RECT 109.960 118.120 144.960 118.440 ; 
                RECT 167.760 118.120 197.320 118.440 ; 
                RECT 386.040 118.120 393.480 118.440 ; 
                RECT 2.880 119.480 83.760 119.800 ; 
                RECT 101.800 119.480 108.240 119.800 ; 
                RECT 113.360 119.480 197.320 119.800 ; 
                RECT 386.040 119.480 393.480 119.800 ; 
                RECT 2.880 120.840 83.760 121.160 ; 
                RECT 101.800 120.840 176.920 121.160 ; 
                RECT 386.040 120.840 393.480 121.160 ; 
                RECT 2.880 122.200 83.760 122.520 ; 
                RECT 101.800 122.200 179.640 122.520 ; 
                RECT 386.040 122.200 393.480 122.520 ; 
                RECT 2.880 123.560 83.760 123.880 ; 
                RECT 101.800 123.560 182.360 123.880 ; 
                RECT 386.040 123.560 393.480 123.880 ; 
                RECT 2.880 124.920 83.760 125.240 ; 
                RECT 101.800 124.920 106.880 125.240 ; 
                RECT 122.200 124.920 144.280 125.240 ; 
                RECT 167.760 124.920 185.080 125.240 ; 
                RECT 386.040 124.920 393.480 125.240 ; 
                RECT 2.880 126.280 83.760 126.600 ; 
                RECT 101.800 126.280 144.280 126.600 ; 
                RECT 167.760 126.280 187.800 126.600 ; 
                RECT 386.040 126.280 393.480 126.600 ; 
                RECT 2.880 127.640 104.840 127.960 ; 
                RECT 112.680 127.640 144.280 127.960 ; 
                RECT 167.760 127.640 190.520 127.960 ; 
                RECT 386.040 127.640 393.480 127.960 ; 
                RECT 2.880 129.000 144.280 129.320 ; 
                RECT 167.760 129.000 193.240 129.320 ; 
                RECT 386.040 129.000 393.480 129.320 ; 
                RECT 2.880 130.360 67.440 130.680 ; 
                RECT 83.440 130.360 144.280 130.680 ; 
                RECT 386.040 130.360 393.480 130.680 ; 
                RECT 2.880 131.720 67.440 132.040 ; 
                RECT 83.440 131.720 144.280 132.040 ; 
                RECT 386.040 131.720 393.480 132.040 ; 
                RECT 2.880 133.080 67.440 133.400 ; 
                RECT 83.440 133.080 110.960 133.400 ; 
                RECT 116.760 133.080 144.280 133.400 ; 
                RECT 167.760 133.080 197.320 133.400 ; 
                RECT 386.040 133.080 393.480 133.400 ; 
                RECT 2.880 134.440 67.440 134.760 ; 
                RECT 83.440 134.440 89.200 134.760 ; 
                RECT 97.040 134.440 144.280 134.760 ; 
                RECT 167.760 134.440 197.320 134.760 ; 
                RECT 386.040 134.440 393.480 134.760 ; 
                RECT 2.880 135.800 67.440 136.120 ; 
                RECT 101.120 135.800 144.280 136.120 ; 
                RECT 167.760 135.800 197.320 136.120 ; 
                RECT 386.040 135.800 393.480 136.120 ; 
                RECT 2.880 137.160 67.440 137.480 ; 
                RECT 83.440 137.160 144.280 137.480 ; 
                RECT 386.040 137.160 393.480 137.480 ; 
                RECT 2.880 138.520 62.000 138.840 ; 
                RECT 97.040 138.520 106.880 138.840 ; 
                RECT 115.400 138.520 144.280 138.840 ; 
                RECT 167.760 138.520 197.320 138.840 ; 
                RECT 386.040 138.520 393.480 138.840 ; 
                RECT 2.880 139.880 89.200 140.200 ; 
                RECT 109.960 139.880 393.480 140.200 ; 
                RECT 2.880 141.240 29.360 141.560 ; 
                RECT 108.600 141.240 393.480 141.560 ; 
                RECT 2.880 142.600 194.600 142.920 ; 
                RECT 388.760 142.600 393.480 142.920 ; 
                RECT 2.880 143.960 194.600 144.280 ; 
                RECT 388.760 143.960 393.480 144.280 ; 
                RECT 2.880 145.320 24.600 145.640 ; 
                RECT 31.080 145.320 72.880 145.640 ; 
                RECT 388.760 145.320 393.480 145.640 ; 
                RECT 2.880 146.680 22.560 147.000 ; 
                RECT 44.000 146.680 72.880 147.000 ; 
                RECT 388.760 146.680 393.480 147.000 ; 
                RECT 2.880 148.040 22.560 148.360 ; 
                RECT 43.320 148.040 55.200 148.360 ; 
                RECT 63.040 148.040 72.880 148.360 ; 
                RECT 388.760 148.040 393.480 148.360 ; 
                RECT 2.880 149.400 36.840 149.720 ; 
                RECT 41.960 149.400 55.200 149.720 ; 
                RECT 63.040 149.400 72.880 149.720 ; 
                RECT 388.760 149.400 393.480 149.720 ; 
                RECT 2.880 150.760 22.560 151.080 ; 
                RECT 33.120 150.760 55.200 151.080 ; 
                RECT 63.040 150.760 72.880 151.080 ; 
                RECT 388.760 150.760 393.480 151.080 ; 
                RECT 2.880 152.120 22.560 152.440 ; 
                RECT 33.120 152.120 55.200 152.440 ; 
                RECT 63.040 152.120 72.880 152.440 ; 
                RECT 388.760 152.120 393.480 152.440 ; 
                RECT 2.880 153.480 22.560 153.800 ; 
                RECT 33.120 153.480 55.200 153.800 ; 
                RECT 59.640 153.480 72.880 153.800 ; 
                RECT 388.760 153.480 393.480 153.800 ; 
                RECT 2.880 154.840 22.560 155.160 ; 
                RECT 33.120 154.840 72.880 155.160 ; 
                RECT 388.760 154.840 393.480 155.160 ; 
                RECT 2.880 156.200 55.200 156.520 ; 
                RECT 63.040 156.200 72.880 156.520 ; 
                RECT 388.760 156.200 393.480 156.520 ; 
                RECT 2.880 157.560 55.200 157.880 ; 
                RECT 63.040 157.560 72.880 157.880 ; 
                RECT 388.760 157.560 393.480 157.880 ; 
                RECT 2.880 158.920 15.760 159.240 ; 
                RECT 18.160 158.920 60.640 159.240 ; 
                RECT 63.040 158.920 72.880 159.240 ; 
                RECT 388.760 158.920 393.480 159.240 ; 
                RECT 2.880 160.280 15.080 160.600 ; 
                RECT 18.160 160.280 55.200 160.600 ; 
                RECT 63.040 160.280 72.880 160.600 ; 
                RECT 388.760 160.280 393.480 160.600 ; 
                RECT 2.880 161.640 55.200 161.960 ; 
                RECT 60.320 161.640 72.880 161.960 ; 
                RECT 388.760 161.640 393.480 161.960 ; 
                RECT 2.880 163.000 14.400 163.320 ; 
                RECT 18.160 163.000 31.400 163.320 ; 
                RECT 35.840 163.000 57.240 163.320 ; 
                RECT 63.040 163.000 72.880 163.320 ; 
                RECT 388.760 163.000 393.480 163.320 ; 
                RECT 2.880 164.360 13.720 164.680 ; 
                RECT 18.160 164.360 31.400 164.680 ; 
                RECT 36.520 164.360 55.200 164.680 ; 
                RECT 56.920 164.360 72.880 164.680 ; 
                RECT 388.760 164.360 393.480 164.680 ; 
                RECT 2.880 165.720 55.200 166.040 ; 
                RECT 61.000 165.720 72.880 166.040 ; 
                RECT 388.760 165.720 393.480 166.040 ; 
                RECT 2.880 167.080 13.040 167.400 ; 
                RECT 18.160 167.080 31.400 167.400 ; 
                RECT 37.200 167.080 55.200 167.400 ; 
                RECT 63.040 167.080 72.880 167.400 ; 
                RECT 388.760 167.080 393.480 167.400 ; 
                RECT 2.880 168.440 12.360 168.760 ; 
                RECT 18.160 168.440 31.400 168.760 ; 
                RECT 37.880 168.440 55.200 168.760 ; 
                RECT 63.040 168.440 72.880 168.760 ; 
                RECT 388.760 168.440 393.480 168.760 ; 
                RECT 2.880 169.800 11.680 170.120 ; 
                RECT 18.160 169.800 31.400 170.120 ; 
                RECT 36.520 169.800 55.200 170.120 ; 
                RECT 61.680 169.800 72.880 170.120 ; 
                RECT 388.760 169.800 393.480 170.120 ; 
                RECT 2.880 171.160 11.000 171.480 ; 
                RECT 18.160 171.160 59.280 171.480 ; 
                RECT 63.040 171.160 72.880 171.480 ; 
                RECT 388.760 171.160 393.480 171.480 ; 
                RECT 2.880 172.520 55.200 172.840 ; 
                RECT 63.040 172.520 72.880 172.840 ; 
                RECT 388.760 172.520 393.480 172.840 ; 
                RECT 2.880 173.880 10.320 174.200 ; 
                RECT 18.160 173.880 55.200 174.200 ; 
                RECT 62.360 173.880 72.880 174.200 ; 
                RECT 388.760 173.880 393.480 174.200 ; 
                RECT 2.880 175.240 9.640 175.560 ; 
                RECT 18.160 175.240 55.200 175.560 ; 
                RECT 56.920 175.240 72.880 175.560 ; 
                RECT 388.760 175.240 393.480 175.560 ; 
                RECT 2.880 176.600 55.200 176.920 ; 
                RECT 63.040 176.600 72.880 176.920 ; 
                RECT 388.760 176.600 393.480 176.920 ; 
                RECT 2.880 177.960 72.880 178.280 ; 
                RECT 388.760 177.960 393.480 178.280 ; 
                RECT 2.880 179.320 57.240 179.640 ; 
                RECT 63.040 179.320 72.880 179.640 ; 
                RECT 388.760 179.320 393.480 179.640 ; 
                RECT 2.880 180.680 57.920 181.000 ; 
                RECT 63.040 180.680 72.880 181.000 ; 
                RECT 388.760 180.680 393.480 181.000 ; 
                RECT 2.880 182.040 58.600 182.360 ; 
                RECT 63.040 182.040 72.880 182.360 ; 
                RECT 388.760 182.040 393.480 182.360 ; 
                RECT 2.880 183.400 59.280 183.720 ; 
                RECT 63.040 183.400 72.880 183.720 ; 
                RECT 388.760 183.400 393.480 183.720 ; 
                RECT 2.880 184.760 72.880 185.080 ; 
                RECT 388.760 184.760 393.480 185.080 ; 
                RECT 2.880 186.120 34.800 186.440 ; 
                RECT 43.320 186.120 72.880 186.440 ; 
                RECT 388.760 186.120 393.480 186.440 ; 
                RECT 2.880 187.480 33.440 187.800 ; 
                RECT 42.640 187.480 55.200 187.800 ; 
                RECT 63.040 187.480 72.880 187.800 ; 
                RECT 388.760 187.480 393.480 187.800 ; 
                RECT 2.880 188.840 55.200 189.160 ; 
                RECT 63.040 188.840 72.880 189.160 ; 
                RECT 388.760 188.840 393.480 189.160 ; 
                RECT 2.880 190.200 55.200 190.520 ; 
                RECT 63.040 190.200 72.880 190.520 ; 
                RECT 388.760 190.200 393.480 190.520 ; 
                RECT 2.880 191.560 55.200 191.880 ; 
                RECT 63.040 191.560 72.880 191.880 ; 
                RECT 388.760 191.560 393.480 191.880 ; 
                RECT 2.880 192.920 55.200 193.240 ; 
                RECT 58.960 192.920 72.880 193.240 ; 
                RECT 388.760 192.920 393.480 193.240 ; 
                RECT 2.880 194.280 72.880 194.600 ; 
                RECT 388.760 194.280 393.480 194.600 ; 
                RECT 2.880 195.640 57.240 195.960 ; 
                RECT 63.040 195.640 72.880 195.960 ; 
                RECT 388.760 195.640 393.480 195.960 ; 
                RECT 2.880 197.000 57.920 197.320 ; 
                RECT 63.040 197.000 72.880 197.320 ; 
                RECT 388.760 197.000 393.480 197.320 ; 
                RECT 2.880 198.360 58.600 198.680 ; 
                RECT 63.040 198.360 72.880 198.680 ; 
                RECT 388.760 198.360 393.480 198.680 ; 
                RECT 2.880 199.720 59.280 200.040 ; 
                RECT 63.040 199.720 72.880 200.040 ; 
                RECT 388.760 199.720 393.480 200.040 ; 
                RECT 2.880 201.080 72.880 201.400 ; 
                RECT 388.760 201.080 393.480 201.400 ; 
                RECT 2.880 202.440 59.280 202.760 ; 
                RECT 63.040 202.440 72.880 202.760 ; 
                RECT 388.760 202.440 393.480 202.760 ; 
                RECT 2.880 203.800 72.880 204.120 ; 
                RECT 388.760 203.800 393.480 204.120 ; 
                RECT 2.880 205.160 59.960 205.480 ; 
                RECT 63.040 205.160 72.880 205.480 ; 
                RECT 388.760 205.160 393.480 205.480 ; 
                RECT 2.880 206.520 60.640 206.840 ; 
                RECT 63.040 206.520 72.880 206.840 ; 
                RECT 388.760 206.520 393.480 206.840 ; 
                RECT 2.880 207.880 60.640 208.200 ; 
                RECT 63.040 207.880 72.880 208.200 ; 
                RECT 388.760 207.880 393.480 208.200 ; 
                RECT 2.880 209.240 72.880 209.560 ; 
                RECT 388.760 209.240 393.480 209.560 ; 
                RECT 2.880 210.600 72.880 210.920 ; 
                RECT 388.760 210.600 393.480 210.920 ; 
                RECT 2.880 211.960 194.600 212.280 ; 
                RECT 388.760 211.960 393.480 212.280 ; 
                RECT 2.880 213.320 194.600 213.640 ; 
                RECT 388.760 213.320 393.480 213.640 ; 
                RECT 2.880 214.680 393.480 215.000 ; 
                RECT 2.880 216.040 393.480 216.360 ; 
                RECT 2.880 217.400 393.480 217.720 ; 
                RECT 2.880 218.760 393.480 219.080 ; 
                RECT 2.880 220.120 393.480 220.440 ; 
                RECT 2.880 2.880 393.480 4.240 ; 
                RECT 2.880 221.440 393.480 222.800 ; 
                RECT 198.740 29.435 204.540 30.555 ; 
                RECT 378.640 29.435 384.440 30.555 ; 
                RECT 198.740 35.235 204.540 35.885 ; 
                RECT 378.640 35.235 384.440 35.885 ; 
                RECT 198.740 40.445 204.540 41.135 ; 
                RECT 378.640 40.445 384.440 41.135 ; 
                RECT 198.740 45.915 204.540 46.605 ; 
                RECT 378.640 45.915 384.440 46.605 ; 
                RECT 198.740 69.180 384.440 69.980 ; 
                RECT 198.740 98.925 384.440 99.215 ; 
                RECT 198.740 73.870 384.440 74.670 ; 
                RECT 198.740 60.130 384.440 61.930 ; 
                RECT 198.740 77.080 384.440 77.880 ; 
                RECT 198.740 80.205 384.440 81.275 ; 
                RECT 198.740 118.150 384.440 118.520 ; 
                RECT 198.740 72.190 384.440 72.990 ; 
                RECT 198.740 20.065 384.440 21.865 ; 
                RECT 73.765 145.715 75.085 210.495 ; 
                RECT 84.310 145.715 86.230 210.495 ; 
                RECT 102.050 145.715 103.970 210.495 ; 
                RECT 105.890 145.715 107.810 210.495 ; 
                RECT 135.070 145.715 136.990 210.495 ; 
                RECT 138.910 145.715 140.830 210.495 ; 
                RECT 142.750 145.715 144.670 210.495 ; 
                RECT 146.590 145.715 148.510 210.495 ; 
                RECT 144.690 61.965 145.580 97.365 ; 
                RECT 151.450 61.965 152.340 97.365 ; 
                RECT 158.640 61.965 160.390 97.365 ; 
                RECT 145.205 125.020 146.315 139.080 ; 
                RECT 153.580 125.020 154.470 139.080 ; 
                RECT 160.230 125.020 161.770 139.080 ; 
                RECT 145.635 110.700 146.745 119.020 ; 
                RECT 153.150 110.700 154.040 119.020 ; 
                RECT 160.230 110.700 161.770 119.020 ; 
                RECT 164.660 52.385 165.550 55.965 ; 
                RECT 23.460 146.780 32.620 147.150 ; 
                RECT 23.460 150.115 32.620 151.005 ; 
                RECT 67.900 130.840 82.740 131.510 ; 
                RECT 67.900 132.105 82.740 134.135 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 396.360 225.680 ; 
        LAYER met2 ;
            RECT 0.000 0.000 396.360 225.680 ; 
    END 
END sram22_256x16m8w8 
END LIBRARY 

