VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_1024x64m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_1024x64m4w8   ;
    SIZE 715.960 BY 776.480 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 312.550 0.000 312.690 0.140 ;
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 318.650 0.000 318.790 0.140 ;
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 324.750 0.000 324.890 0.140 ;
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.850 0.000 330.990 0.140 ;
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.950 0.000 337.090 0.140 ;
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 343.050 0.000 343.190 0.140 ;
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 349.150 0.000 349.290 0.140 ;
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 355.250 0.000 355.390 0.140 ;
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 361.350 0.000 361.490 0.140 ;
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 367.450 0.000 367.590 0.140 ;
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 373.550 0.000 373.690 0.140 ;
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 379.650 0.000 379.790 0.140 ;
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 385.750 0.000 385.890 0.140 ;
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 391.850 0.000 391.990 0.140 ;
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 397.950 0.000 398.090 0.140 ;
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 404.050 0.000 404.190 0.140 ;
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 410.150 0.000 410.290 0.140 ;
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 416.250 0.000 416.390 0.140 ;
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 422.350 0.000 422.490 0.140 ;
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 428.450 0.000 428.590 0.140 ;
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 434.550 0.000 434.690 0.140 ;
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 440.650 0.000 440.790 0.140 ;
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 446.750 0.000 446.890 0.140 ;
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 452.850 0.000 452.990 0.140 ;
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 458.950 0.000 459.090 0.140 ;
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 465.050 0.000 465.190 0.140 ;
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 471.150 0.000 471.290 0.140 ;
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 477.250 0.000 477.390 0.140 ;
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 483.350 0.000 483.490 0.140 ;
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 489.450 0.000 489.590 0.140 ;
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 495.550 0.000 495.690 0.140 ;
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 501.650 0.000 501.790 0.140 ;
        END 
    END dout[31] 
    PIN dout[32] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 507.750 0.000 507.890 0.140 ;
        END 
    END dout[32] 
    PIN dout[33] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 513.850 0.000 513.990 0.140 ;
        END 
    END dout[33] 
    PIN dout[34] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 519.950 0.000 520.090 0.140 ;
        END 
    END dout[34] 
    PIN dout[35] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 526.050 0.000 526.190 0.140 ;
        END 
    END dout[35] 
    PIN dout[36] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 532.150 0.000 532.290 0.140 ;
        END 
    END dout[36] 
    PIN dout[37] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 538.250 0.000 538.390 0.140 ;
        END 
    END dout[37] 
    PIN dout[38] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 544.350 0.000 544.490 0.140 ;
        END 
    END dout[38] 
    PIN dout[39] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 550.450 0.000 550.590 0.140 ;
        END 
    END dout[39] 
    PIN dout[40] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 556.550 0.000 556.690 0.140 ;
        END 
    END dout[40] 
    PIN dout[41] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 562.650 0.000 562.790 0.140 ;
        END 
    END dout[41] 
    PIN dout[42] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 568.750 0.000 568.890 0.140 ;
        END 
    END dout[42] 
    PIN dout[43] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 574.850 0.000 574.990 0.140 ;
        END 
    END dout[43] 
    PIN dout[44] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 580.950 0.000 581.090 0.140 ;
        END 
    END dout[44] 
    PIN dout[45] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 587.050 0.000 587.190 0.140 ;
        END 
    END dout[45] 
    PIN dout[46] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 593.150 0.000 593.290 0.140 ;
        END 
    END dout[46] 
    PIN dout[47] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 599.250 0.000 599.390 0.140 ;
        END 
    END dout[47] 
    PIN dout[48] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 605.350 0.000 605.490 0.140 ;
        END 
    END dout[48] 
    PIN dout[49] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 611.450 0.000 611.590 0.140 ;
        END 
    END dout[49] 
    PIN dout[50] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 617.550 0.000 617.690 0.140 ;
        END 
    END dout[50] 
    PIN dout[51] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 623.650 0.000 623.790 0.140 ;
        END 
    END dout[51] 
    PIN dout[52] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 629.750 0.000 629.890 0.140 ;
        END 
    END dout[52] 
    PIN dout[53] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 635.850 0.000 635.990 0.140 ;
        END 
    END dout[53] 
    PIN dout[54] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 641.950 0.000 642.090 0.140 ;
        END 
    END dout[54] 
    PIN dout[55] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 648.050 0.000 648.190 0.140 ;
        END 
    END dout[55] 
    PIN dout[56] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 654.150 0.000 654.290 0.140 ;
        END 
    END dout[56] 
    PIN dout[57] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 660.250 0.000 660.390 0.140 ;
        END 
    END dout[57] 
    PIN dout[58] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 666.350 0.000 666.490 0.140 ;
        END 
    END dout[58] 
    PIN dout[59] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 672.450 0.000 672.590 0.140 ;
        END 
    END dout[59] 
    PIN dout[60] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 678.550 0.000 678.690 0.140 ;
        END 
    END dout[60] 
    PIN dout[61] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 684.650 0.000 684.790 0.140 ;
        END 
    END dout[61] 
    PIN dout[62] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 690.750 0.000 690.890 0.140 ;
        END 
    END dout[62] 
    PIN dout[63] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 696.850 0.000 696.990 0.140 ;
        END 
    END dout[63] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 312.130 0.000 312.270 0.140 ;
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 318.230 0.000 318.370 0.140 ;
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 324.330 0.000 324.470 0.140 ;
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.430 0.000 330.570 0.140 ;
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.530 0.000 336.670 0.140 ;
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 342.630 0.000 342.770 0.140 ;
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 348.730 0.000 348.870 0.140 ;
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 354.830 0.000 354.970 0.140 ;
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 360.930 0.000 361.070 0.140 ;
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 367.030 0.000 367.170 0.140 ;
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 373.130 0.000 373.270 0.140 ;
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 379.230 0.000 379.370 0.140 ;
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 385.330 0.000 385.470 0.140 ;
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 391.430 0.000 391.570 0.140 ;
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 397.530 0.000 397.670 0.140 ;
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 403.630 0.000 403.770 0.140 ;
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 409.730 0.000 409.870 0.140 ;
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 415.830 0.000 415.970 0.140 ;
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 421.930 0.000 422.070 0.140 ;
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 428.030 0.000 428.170 0.140 ;
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 434.130 0.000 434.270 0.140 ;
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 440.230 0.000 440.370 0.140 ;
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 446.330 0.000 446.470 0.140 ;
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 452.430 0.000 452.570 0.140 ;
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 458.530 0.000 458.670 0.140 ;
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 464.630 0.000 464.770 0.140 ;
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 470.730 0.000 470.870 0.140 ;
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 476.830 0.000 476.970 0.140 ;
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 482.930 0.000 483.070 0.140 ;
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 489.030 0.000 489.170 0.140 ;
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 495.130 0.000 495.270 0.140 ;
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 501.230 0.000 501.370 0.140 ;
        END 
    END din[31] 
    PIN din[32] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 507.330 0.000 507.470 0.140 ;
        END 
    END din[32] 
    PIN din[33] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 513.430 0.000 513.570 0.140 ;
        END 
    END din[33] 
    PIN din[34] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 519.530 0.000 519.670 0.140 ;
        END 
    END din[34] 
    PIN din[35] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 525.630 0.000 525.770 0.140 ;
        END 
    END din[35] 
    PIN din[36] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 531.730 0.000 531.870 0.140 ;
        END 
    END din[36] 
    PIN din[37] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 537.830 0.000 537.970 0.140 ;
        END 
    END din[37] 
    PIN din[38] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 543.930 0.000 544.070 0.140 ;
        END 
    END din[38] 
    PIN din[39] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 550.030 0.000 550.170 0.140 ;
        END 
    END din[39] 
    PIN din[40] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 556.130 0.000 556.270 0.140 ;
        END 
    END din[40] 
    PIN din[41] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 562.230 0.000 562.370 0.140 ;
        END 
    END din[41] 
    PIN din[42] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 568.330 0.000 568.470 0.140 ;
        END 
    END din[42] 
    PIN din[43] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 574.430 0.000 574.570 0.140 ;
        END 
    END din[43] 
    PIN din[44] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 580.530 0.000 580.670 0.140 ;
        END 
    END din[44] 
    PIN din[45] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 586.630 0.000 586.770 0.140 ;
        END 
    END din[45] 
    PIN din[46] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 592.730 0.000 592.870 0.140 ;
        END 
    END din[46] 
    PIN din[47] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 598.830 0.000 598.970 0.140 ;
        END 
    END din[47] 
    PIN din[48] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 604.930 0.000 605.070 0.140 ;
        END 
    END din[48] 
    PIN din[49] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 611.030 0.000 611.170 0.140 ;
        END 
    END din[49] 
    PIN din[50] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 617.130 0.000 617.270 0.140 ;
        END 
    END din[50] 
    PIN din[51] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 623.230 0.000 623.370 0.140 ;
        END 
    END din[51] 
    PIN din[52] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 629.330 0.000 629.470 0.140 ;
        END 
    END din[52] 
    PIN din[53] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 635.430 0.000 635.570 0.140 ;
        END 
    END din[53] 
    PIN din[54] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 641.530 0.000 641.670 0.140 ;
        END 
    END din[54] 
    PIN din[55] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 647.630 0.000 647.770 0.140 ;
        END 
    END din[55] 
    PIN din[56] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 653.730 0.000 653.870 0.140 ;
        END 
    END din[56] 
    PIN din[57] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 659.830 0.000 659.970 0.140 ;
        END 
    END din[57] 
    PIN din[58] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 665.930 0.000 666.070 0.140 ;
        END 
    END din[58] 
    PIN din[59] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 672.030 0.000 672.170 0.140 ;
        END 
    END din[59] 
    PIN din[60] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 678.130 0.000 678.270 0.140 ;
        END 
    END din[60] 
    PIN din[61] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 684.230 0.000 684.370 0.140 ;
        END 
    END din[61] 
    PIN din[62] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 690.330 0.000 690.470 0.140 ;
        END 
    END din[62] 
    PIN din[63] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.184600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 696.430 0.000 696.570 0.140 ;
        END 
    END din[63] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.995000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 311.780 0.000 311.920 0.140 ;
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.995000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 360.580 0.000 360.720 0.140 ;
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.995000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 409.380 0.000 409.520 0.140 ;
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.995000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 458.180 0.000 458.320 0.140 ;
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.995000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 506.980 0.000 507.120 0.140 ;
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.995000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 555.780 0.000 555.920 0.140 ;
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.995000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 604.580 0.000 604.720 0.140 ;
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.995000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 653.380 0.000 653.520 0.140 ;
        END 
    END wmask[7] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 256.160 0.000 256.480 0.320 ;
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 250.040 0.000 250.360 0.320 ;
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 243.920 0.000 244.240 0.320 ;
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 237.800 0.000 238.120 0.320 ;
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 231.680 0.000 232.000 0.320 ;
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 225.560 0.000 225.880 0.320 ;
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 219.440 0.000 219.760 0.320 ;
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 213.320 0.000 213.640 0.320 ;
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 207.880 0.000 208.200 0.320 ;
        END 
    END addr[8] 
    PIN addr[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 201.760 0.000 202.080 0.320 ;
        END 
    END addr[9] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 268.400 0.000 268.720 0.320 ;
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.791100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 262.280 0.000 262.600 0.320 ;
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 41.850000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 271.800 0.000 272.120 0.320 ;
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 45.756000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 272.480 0.000 272.800 0.320 ;
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 311.560 6.240 ;
                RECT 313.280 5.920 317.680 6.240 ;
                RECT 319.400 5.920 323.800 6.240 ;
                RECT 325.520 5.920 329.920 6.240 ;
                RECT 331.640 5.920 336.040 6.240 ;
                RECT 337.760 5.920 342.160 6.240 ;
                RECT 343.880 5.920 348.280 6.240 ;
                RECT 350.000 5.920 354.400 6.240 ;
                RECT 356.120 5.920 360.520 6.240 ;
                RECT 362.240 5.920 366.640 6.240 ;
                RECT 368.360 5.920 372.760 6.240 ;
                RECT 374.480 5.920 378.880 6.240 ;
                RECT 380.600 5.920 385.000 6.240 ;
                RECT 386.720 5.920 391.120 6.240 ;
                RECT 392.840 5.920 397.240 6.240 ;
                RECT 398.960 5.920 403.360 6.240 ;
                RECT 405.080 5.920 409.480 6.240 ;
                RECT 411.200 5.920 415.600 6.240 ;
                RECT 417.320 5.920 421.720 6.240 ;
                RECT 423.440 5.920 427.840 6.240 ;
                RECT 429.560 5.920 433.960 6.240 ;
                RECT 435.680 5.920 440.080 6.240 ;
                RECT 441.800 5.920 446.200 6.240 ;
                RECT 447.920 5.920 452.320 6.240 ;
                RECT 453.360 5.920 458.440 6.240 ;
                RECT 459.480 5.920 464.560 6.240 ;
                RECT 465.600 5.920 470.680 6.240 ;
                RECT 471.720 5.920 476.800 6.240 ;
                RECT 477.840 5.920 482.920 6.240 ;
                RECT 483.960 5.920 489.040 6.240 ;
                RECT 490.080 5.920 495.160 6.240 ;
                RECT 496.200 5.920 501.280 6.240 ;
                RECT 502.320 5.920 506.720 6.240 ;
                RECT 508.440 5.920 512.840 6.240 ;
                RECT 514.560 5.920 518.960 6.240 ;
                RECT 520.680 5.920 525.080 6.240 ;
                RECT 526.800 5.920 531.200 6.240 ;
                RECT 532.920 5.920 537.320 6.240 ;
                RECT 539.040 5.920 543.440 6.240 ;
                RECT 545.160 5.920 549.560 6.240 ;
                RECT 551.280 5.920 555.680 6.240 ;
                RECT 557.400 5.920 561.800 6.240 ;
                RECT 563.520 5.920 567.920 6.240 ;
                RECT 569.640 5.920 574.040 6.240 ;
                RECT 575.760 5.920 580.160 6.240 ;
                RECT 581.880 5.920 586.280 6.240 ;
                RECT 588.000 5.920 592.400 6.240 ;
                RECT 594.120 5.920 598.520 6.240 ;
                RECT 600.240 5.920 604.640 6.240 ;
                RECT 606.360 5.920 610.760 6.240 ;
                RECT 612.480 5.920 616.880 6.240 ;
                RECT 618.600 5.920 623.000 6.240 ;
                RECT 624.720 5.920 629.120 6.240 ;
                RECT 630.840 5.920 635.240 6.240 ;
                RECT 636.960 5.920 641.360 6.240 ;
                RECT 643.080 5.920 647.480 6.240 ;
                RECT 649.200 5.920 653.600 6.240 ;
                RECT 655.320 5.920 659.720 6.240 ;
                RECT 660.760 5.920 665.840 6.240 ;
                RECT 666.880 5.920 671.960 6.240 ;
                RECT 673.000 5.920 678.080 6.240 ;
                RECT 679.120 5.920 684.200 6.240 ;
                RECT 685.240 5.920 690.320 6.240 ;
                RECT 691.360 5.920 696.440 6.240 ;
                RECT 697.480 5.920 715.800 6.240 ;
                RECT 0.160 7.280 715.800 7.600 ;
                RECT 0.160 8.640 715.800 8.960 ;
                RECT 0.160 10.000 271.440 10.320 ;
                RECT 307.840 10.000 715.800 10.320 ;
                RECT 0.160 11.360 715.800 11.680 ;
                RECT 0.160 12.720 197.320 13.040 ;
                RECT 273.160 12.720 715.800 13.040 ;
                RECT 0.160 14.080 715.800 14.400 ;
                RECT 0.160 15.440 715.800 15.760 ;
                RECT 0.160 16.800 715.800 17.120 ;
                RECT 0.160 18.160 197.320 18.480 ;
                RECT 272.480 18.160 715.800 18.480 ;
                RECT 0.160 19.520 310.880 19.840 ;
                RECT 653.960 19.520 715.800 19.840 ;
                RECT 0.160 20.880 301.360 21.200 ;
                RECT 706.320 20.880 715.800 21.200 ;
                RECT 0.160 22.240 301.360 22.560 ;
                RECT 706.320 22.240 715.800 22.560 ;
                RECT 0.160 23.600 301.360 23.920 ;
                RECT 706.320 23.600 715.800 23.920 ;
                RECT 0.160 24.960 301.360 25.280 ;
                RECT 706.320 24.960 715.800 25.280 ;
                RECT 0.160 26.320 301.360 26.640 ;
                RECT 706.320 26.320 715.800 26.640 ;
                RECT 0.160 27.680 301.360 28.000 ;
                RECT 706.320 27.680 715.800 28.000 ;
                RECT 0.160 29.040 301.360 29.360 ;
                RECT 706.320 29.040 715.800 29.360 ;
                RECT 0.160 30.400 301.360 30.720 ;
                RECT 706.320 30.400 715.800 30.720 ;
                RECT 0.160 31.760 301.360 32.080 ;
                RECT 706.320 31.760 715.800 32.080 ;
                RECT 0.160 33.120 301.360 33.440 ;
                RECT 706.320 33.120 715.800 33.440 ;
                RECT 0.160 34.480 301.360 34.800 ;
                RECT 706.320 34.480 715.800 34.800 ;
                RECT 0.160 35.840 301.360 36.160 ;
                RECT 706.320 35.840 715.800 36.160 ;
                RECT 0.160 37.200 145.640 37.520 ;
                RECT 250.040 37.200 300.680 37.520 ;
                RECT 706.320 37.200 715.800 37.520 ;
                RECT 0.160 38.560 144.280 38.880 ;
                RECT 256.160 38.560 301.360 38.880 ;
                RECT 706.320 38.560 715.800 38.880 ;
                RECT 0.160 39.920 125.240 40.240 ;
                RECT 273.160 39.920 301.360 40.240 ;
                RECT 706.320 39.920 715.800 40.240 ;
                RECT 0.160 41.280 123.880 41.600 ;
                RECT 269.080 41.280 301.360 41.600 ;
                RECT 706.320 41.280 715.800 41.600 ;
                RECT 0.160 42.640 301.360 42.960 ;
                RECT 706.320 42.640 715.800 42.960 ;
                RECT 0.160 44.000 265.320 44.320 ;
                RECT 271.120 44.000 301.360 44.320 ;
                RECT 706.320 44.000 715.800 44.320 ;
                RECT 0.160 45.360 265.320 45.680 ;
                RECT 271.120 45.360 301.360 45.680 ;
                RECT 706.320 45.360 715.800 45.680 ;
                RECT 0.160 46.720 265.320 47.040 ;
                RECT 706.320 46.720 715.800 47.040 ;
                RECT 0.160 48.080 265.320 48.400 ;
                RECT 706.320 48.080 715.800 48.400 ;
                RECT 0.160 49.440 265.320 49.760 ;
                RECT 271.120 49.440 301.360 49.760 ;
                RECT 706.320 49.440 715.800 49.760 ;
                RECT 0.160 50.800 301.360 51.120 ;
                RECT 706.320 50.800 715.800 51.120 ;
                RECT 0.160 52.160 301.360 52.480 ;
                RECT 706.320 52.160 715.800 52.480 ;
                RECT 0.160 53.520 301.360 53.840 ;
                RECT 706.320 53.520 715.800 53.840 ;
                RECT 0.160 54.880 301.360 55.200 ;
                RECT 706.320 54.880 715.800 55.200 ;
                RECT 0.160 56.240 144.280 56.560 ;
                RECT 150.080 56.240 155.840 56.560 ;
                RECT 269.760 56.240 301.360 56.560 ;
                RECT 706.320 56.240 715.800 56.560 ;
                RECT 0.160 57.600 145.640 57.920 ;
                RECT 149.400 57.600 155.840 57.920 ;
                RECT 285.400 57.600 301.360 57.920 ;
                RECT 706.320 57.600 715.800 57.920 ;
                RECT 0.160 58.960 155.840 59.280 ;
                RECT 285.400 58.960 301.360 59.280 ;
                RECT 706.320 58.960 715.800 59.280 ;
                RECT 0.160 60.320 155.840 60.640 ;
                RECT 282.680 60.320 301.360 60.640 ;
                RECT 706.320 60.320 715.800 60.640 ;
                RECT 0.160 61.680 155.840 62.000 ;
                RECT 285.400 61.680 301.360 62.000 ;
                RECT 706.320 61.680 715.800 62.000 ;
                RECT 0.160 63.040 155.840 63.360 ;
                RECT 285.400 63.040 301.360 63.360 ;
                RECT 706.320 63.040 715.800 63.360 ;
                RECT 0.160 64.400 155.840 64.720 ;
                RECT 269.760 64.400 301.360 64.720 ;
                RECT 706.320 64.400 715.800 64.720 ;
                RECT 0.160 65.760 155.840 66.080 ;
                RECT 285.400 65.760 301.360 66.080 ;
                RECT 706.320 65.760 715.800 66.080 ;
                RECT 0.160 67.120 155.840 67.440 ;
                RECT 282.680 67.120 301.360 67.440 ;
                RECT 706.320 67.120 715.800 67.440 ;
                RECT 0.160 68.480 155.840 68.800 ;
                RECT 285.400 68.480 301.360 68.800 ;
                RECT 706.320 68.480 715.800 68.800 ;
                RECT 0.160 69.840 155.840 70.160 ;
                RECT 285.400 69.840 301.360 70.160 ;
                RECT 706.320 69.840 715.800 70.160 ;
                RECT 0.160 71.200 155.840 71.520 ;
                RECT 285.400 71.200 301.360 71.520 ;
                RECT 706.320 71.200 715.800 71.520 ;
                RECT 0.160 72.560 155.840 72.880 ;
                RECT 282.680 72.560 301.360 72.880 ;
                RECT 706.320 72.560 715.800 72.880 ;
                RECT 0.160 73.920 155.840 74.240 ;
                RECT 269.760 73.920 301.360 74.240 ;
                RECT 706.320 73.920 715.800 74.240 ;
                RECT 0.160 75.280 155.840 75.600 ;
                RECT 285.400 75.280 301.360 75.600 ;
                RECT 706.320 75.280 715.800 75.600 ;
                RECT 0.160 76.640 155.840 76.960 ;
                RECT 290.840 76.640 301.360 76.960 ;
                RECT 706.320 76.640 715.800 76.960 ;
                RECT 0.160 78.000 155.840 78.320 ;
                RECT 290.840 78.000 301.360 78.320 ;
                RECT 706.320 78.000 715.800 78.320 ;
                RECT 0.160 79.360 155.840 79.680 ;
                RECT 288.120 79.360 301.360 79.680 ;
                RECT 706.320 79.360 715.800 79.680 ;
                RECT 0.160 80.720 155.840 81.040 ;
                RECT 290.840 80.720 301.360 81.040 ;
                RECT 706.320 80.720 715.800 81.040 ;
                RECT 0.160 82.080 155.840 82.400 ;
                RECT 269.760 82.080 301.360 82.400 ;
                RECT 706.320 82.080 715.800 82.400 ;
                RECT 0.160 83.440 155.840 83.760 ;
                RECT 290.840 83.440 301.360 83.760 ;
                RECT 706.320 83.440 715.800 83.760 ;
                RECT 0.160 84.800 155.840 85.120 ;
                RECT 290.840 84.800 301.360 85.120 ;
                RECT 706.320 84.800 715.800 85.120 ;
                RECT 0.160 86.160 155.840 86.480 ;
                RECT 288.120 86.160 301.360 86.480 ;
                RECT 706.320 86.160 715.800 86.480 ;
                RECT 0.160 87.520 155.840 87.840 ;
                RECT 290.840 87.520 301.360 87.840 ;
                RECT 706.320 87.520 715.800 87.840 ;
                RECT 0.160 88.880 155.840 89.200 ;
                RECT 290.840 88.880 301.360 89.200 ;
                RECT 706.320 88.880 715.800 89.200 ;
                RECT 0.160 90.240 155.840 90.560 ;
                RECT 269.760 90.240 301.360 90.560 ;
                RECT 706.320 90.240 715.800 90.560 ;
                RECT 0.160 91.600 155.840 91.920 ;
                RECT 290.840 91.600 301.360 91.920 ;
                RECT 706.320 91.600 715.800 91.920 ;
                RECT 0.160 92.960 155.840 93.280 ;
                RECT 288.120 92.960 301.360 93.280 ;
                RECT 706.320 92.960 715.800 93.280 ;
                RECT 0.160 94.320 155.840 94.640 ;
                RECT 290.840 94.320 301.360 94.640 ;
                RECT 706.320 94.320 715.800 94.640 ;
                RECT 0.160 95.680 155.840 96.000 ;
                RECT 296.280 95.680 301.360 96.000 ;
                RECT 706.320 95.680 715.800 96.000 ;
                RECT 0.160 97.040 155.840 97.360 ;
                RECT 296.280 97.040 301.360 97.360 ;
                RECT 706.320 97.040 715.800 97.360 ;
                RECT 0.160 98.400 155.840 98.720 ;
                RECT 293.560 98.400 301.360 98.720 ;
                RECT 706.320 98.400 715.800 98.720 ;
                RECT 0.160 99.760 155.840 100.080 ;
                RECT 269.760 99.760 301.360 100.080 ;
                RECT 706.320 99.760 715.800 100.080 ;
                RECT 0.160 101.120 155.840 101.440 ;
                RECT 293.560 101.120 301.360 101.440 ;
                RECT 706.320 101.120 715.800 101.440 ;
                RECT 0.160 102.480 155.840 102.800 ;
                RECT 296.280 102.480 301.360 102.800 ;
                RECT 706.320 102.480 715.800 102.800 ;
                RECT 0.160 103.840 155.840 104.160 ;
                RECT 296.280 103.840 301.360 104.160 ;
                RECT 706.320 103.840 715.800 104.160 ;
                RECT 0.160 105.200 155.840 105.520 ;
                RECT 293.560 105.200 301.360 105.520 ;
                RECT 706.320 105.200 715.800 105.520 ;
                RECT 0.160 106.560 155.840 106.880 ;
                RECT 296.280 106.560 301.360 106.880 ;
                RECT 706.320 106.560 715.800 106.880 ;
                RECT 0.160 107.920 155.840 108.240 ;
                RECT 269.760 107.920 301.360 108.240 ;
                RECT 706.320 107.920 715.800 108.240 ;
                RECT 0.160 109.280 155.840 109.600 ;
                RECT 296.280 109.280 301.360 109.600 ;
                RECT 706.320 109.280 715.800 109.600 ;
                RECT 0.160 110.640 155.840 110.960 ;
                RECT 296.280 110.640 301.360 110.960 ;
                RECT 706.320 110.640 715.800 110.960 ;
                RECT 0.160 112.000 155.840 112.320 ;
                RECT 293.560 112.000 301.360 112.320 ;
                RECT 706.320 112.000 715.800 112.320 ;
                RECT 0.160 113.360 155.840 113.680 ;
                RECT 296.280 113.360 301.360 113.680 ;
                RECT 706.320 113.360 715.800 113.680 ;
                RECT 0.160 114.720 155.840 115.040 ;
                RECT 706.320 114.720 715.800 115.040 ;
                RECT 0.160 116.080 155.840 116.400 ;
                RECT 269.760 116.080 301.360 116.400 ;
                RECT 706.320 116.080 715.800 116.400 ;
                RECT 0.160 117.440 155.840 117.760 ;
                RECT 706.320 117.440 715.800 117.760 ;
                RECT 0.160 118.800 155.840 119.120 ;
                RECT 706.320 118.800 715.800 119.120 ;
                RECT 0.160 120.160 155.840 120.480 ;
                RECT 706.320 120.160 715.800 120.480 ;
                RECT 0.160 121.520 155.840 121.840 ;
                RECT 706.320 121.520 715.800 121.840 ;
                RECT 0.160 122.880 155.840 123.200 ;
                RECT 706.320 122.880 715.800 123.200 ;
                RECT 0.160 124.240 155.840 124.560 ;
                RECT 706.320 124.240 715.800 124.560 ;
                RECT 0.160 125.600 155.840 125.920 ;
                RECT 269.760 125.600 301.360 125.920 ;
                RECT 706.320 125.600 715.800 125.920 ;
                RECT 0.160 126.960 155.840 127.280 ;
                RECT 706.320 126.960 715.800 127.280 ;
                RECT 0.160 128.320 155.840 128.640 ;
                RECT 706.320 128.320 715.800 128.640 ;
                RECT 0.160 129.680 155.840 130.000 ;
                RECT 706.320 129.680 715.800 130.000 ;
                RECT 0.160 131.040 155.840 131.360 ;
                RECT 706.320 131.040 715.800 131.360 ;
                RECT 0.160 132.400 155.840 132.720 ;
                RECT 706.320 132.400 715.800 132.720 ;
                RECT 0.160 133.760 155.840 134.080 ;
                RECT 269.760 133.760 301.360 134.080 ;
                RECT 706.320 133.760 715.800 134.080 ;
                RECT 0.160 135.120 301.360 135.440 ;
                RECT 706.320 135.120 715.800 135.440 ;
                RECT 0.160 136.480 98.720 136.800 ;
                RECT 117.440 136.480 276.880 136.800 ;
                RECT 706.320 136.480 715.800 136.800 ;
                RECT 0.160 137.840 98.720 138.160 ;
                RECT 117.440 137.840 295.920 138.160 ;
                RECT 706.320 137.840 715.800 138.160 ;
                RECT 0.160 139.200 98.720 139.520 ;
                RECT 117.440 139.200 295.920 139.520 ;
                RECT 706.320 139.200 715.800 139.520 ;
                RECT 0.160 140.560 98.720 140.880 ;
                RECT 117.440 140.560 295.920 140.880 ;
                RECT 706.320 140.560 715.800 140.880 ;
                RECT 0.160 141.920 98.720 142.240 ;
                RECT 117.440 141.920 290.480 142.240 ;
                RECT 706.320 141.920 715.800 142.240 ;
                RECT 0.160 143.280 98.720 143.600 ;
                RECT 117.440 143.280 290.480 143.600 ;
                RECT 706.320 143.280 715.800 143.600 ;
                RECT 0.160 144.640 98.720 144.960 ;
                RECT 117.440 144.640 120.480 144.960 ;
                RECT 131.040 144.640 285.040 144.960 ;
                RECT 706.320 144.640 715.800 144.960 ;
                RECT 0.160 146.000 98.720 146.320 ;
                RECT 117.440 146.000 121.840 146.320 ;
                RECT 127.640 146.000 135.440 146.320 ;
                RECT 137.840 146.000 285.040 146.320 ;
                RECT 706.320 146.000 715.800 146.320 ;
                RECT 0.160 147.360 98.720 147.680 ;
                RECT 117.440 147.360 123.200 147.680 ;
                RECT 126.960 147.360 279.600 147.680 ;
                RECT 706.320 147.360 715.800 147.680 ;
                RECT 0.160 148.720 98.720 149.040 ;
                RECT 117.440 148.720 129.320 149.040 ;
                RECT 137.160 148.720 279.600 149.040 ;
                RECT 706.320 148.720 715.800 149.040 ;
                RECT 0.160 150.080 98.720 150.400 ;
                RECT 117.440 150.080 125.240 150.400 ;
                RECT 138.520 150.080 301.360 150.400 ;
                RECT 706.320 150.080 715.800 150.400 ;
                RECT 0.160 151.440 98.720 151.760 ;
                RECT 117.440 151.440 122.520 151.760 ;
                RECT 131.040 151.440 301.360 151.760 ;
                RECT 706.320 151.440 715.800 151.760 ;
                RECT 0.160 152.800 98.720 153.120 ;
                RECT 117.440 152.800 301.360 153.120 ;
                RECT 706.320 152.800 715.800 153.120 ;
                RECT 0.160 154.160 98.720 154.480 ;
                RECT 117.440 154.160 121.840 154.480 ;
                RECT 124.240 154.160 301.360 154.480 ;
                RECT 706.320 154.160 715.800 154.480 ;
                RECT 0.160 155.520 98.720 155.840 ;
                RECT 117.440 155.520 119.800 155.840 ;
                RECT 137.160 155.520 301.360 155.840 ;
                RECT 706.320 155.520 715.800 155.840 ;
                RECT 0.160 156.880 98.720 157.200 ;
                RECT 117.440 156.880 128.640 157.200 ;
                RECT 131.040 156.880 301.360 157.200 ;
                RECT 706.320 156.880 715.800 157.200 ;
                RECT 0.160 158.240 98.720 158.560 ;
                RECT 117.440 158.240 301.360 158.560 ;
                RECT 706.320 158.240 715.800 158.560 ;
                RECT 0.160 159.600 98.720 159.920 ;
                RECT 117.440 159.600 129.320 159.920 ;
                RECT 137.840 159.600 301.360 159.920 ;
                RECT 706.320 159.600 715.800 159.920 ;
                RECT 0.160 160.960 98.720 161.280 ;
                RECT 117.440 160.960 126.600 161.280 ;
                RECT 131.040 160.960 301.360 161.280 ;
                RECT 706.320 160.960 715.800 161.280 ;
                RECT 0.160 162.320 98.720 162.640 ;
                RECT 117.440 162.320 128.640 162.640 ;
                RECT 131.040 162.320 301.360 162.640 ;
                RECT 706.320 162.320 715.800 162.640 ;
                RECT 0.160 163.680 98.720 164.000 ;
                RECT 117.440 163.680 301.360 164.000 ;
                RECT 706.320 163.680 715.800 164.000 ;
                RECT 0.160 165.040 98.720 165.360 ;
                RECT 117.440 165.040 119.800 165.360 ;
                RECT 142.600 165.040 301.360 165.360 ;
                RECT 706.320 165.040 715.800 165.360 ;
                RECT 0.160 166.400 98.720 166.720 ;
                RECT 117.440 166.400 138.160 166.720 ;
                RECT 143.960 166.400 301.360 166.720 ;
                RECT 706.320 166.400 715.800 166.720 ;
                RECT 0.160 167.760 98.720 168.080 ;
                RECT 117.440 167.760 128.640 168.080 ;
                RECT 131.040 167.760 140.880 168.080 ;
                RECT 144.640 167.760 301.360 168.080 ;
                RECT 706.320 167.760 715.800 168.080 ;
                RECT 0.160 169.120 98.720 169.440 ;
                RECT 117.440 169.120 120.480 169.440 ;
                RECT 133.760 169.120 301.360 169.440 ;
                RECT 706.320 169.120 715.800 169.440 ;
                RECT 0.160 170.480 98.720 170.800 ;
                RECT 117.440 170.480 129.320 170.800 ;
                RECT 137.840 170.480 301.360 170.800 ;
                RECT 706.320 170.480 715.800 170.800 ;
                RECT 0.160 171.840 98.720 172.160 ;
                RECT 117.440 171.840 126.600 172.160 ;
                RECT 131.040 171.840 301.360 172.160 ;
                RECT 706.320 171.840 715.800 172.160 ;
                RECT 0.160 173.200 98.720 173.520 ;
                RECT 117.440 173.200 129.320 173.520 ;
                RECT 138.520 173.200 301.360 173.520 ;
                RECT 706.320 173.200 715.800 173.520 ;
                RECT 0.160 174.560 98.720 174.880 ;
                RECT 117.440 174.560 301.360 174.880 ;
                RECT 706.320 174.560 715.800 174.880 ;
                RECT 0.160 175.920 98.720 176.240 ;
                RECT 117.440 175.920 122.520 176.240 ;
                RECT 125.600 175.920 301.360 176.240 ;
                RECT 706.320 175.920 715.800 176.240 ;
                RECT 0.160 177.280 98.720 177.600 ;
                RECT 117.440 177.280 122.520 177.600 ;
                RECT 131.040 177.280 301.360 177.600 ;
                RECT 706.320 177.280 715.800 177.600 ;
                RECT 0.160 178.640 98.720 178.960 ;
                RECT 117.440 178.640 301.360 178.960 ;
                RECT 706.320 178.640 715.800 178.960 ;
                RECT 0.160 180.000 98.720 180.320 ;
                RECT 117.440 180.000 128.640 180.320 ;
                RECT 131.040 180.000 301.360 180.320 ;
                RECT 706.320 180.000 715.800 180.320 ;
                RECT 0.160 181.360 98.720 181.680 ;
                RECT 117.440 181.360 121.840 181.680 ;
                RECT 127.640 181.360 129.320 181.680 ;
                RECT 131.720 181.360 301.360 181.680 ;
                RECT 706.320 181.360 715.800 181.680 ;
                RECT 0.160 182.720 98.720 183.040 ;
                RECT 117.440 182.720 125.920 183.040 ;
                RECT 137.160 182.720 301.360 183.040 ;
                RECT 706.320 182.720 715.800 183.040 ;
                RECT 0.160 184.080 98.720 184.400 ;
                RECT 117.440 184.080 128.640 184.400 ;
                RECT 131.040 184.080 301.360 184.400 ;
                RECT 706.320 184.080 715.800 184.400 ;
                RECT 0.160 185.440 98.720 185.760 ;
                RECT 117.440 185.440 123.880 185.760 ;
                RECT 131.040 185.440 301.360 185.760 ;
                RECT 706.320 185.440 715.800 185.760 ;
                RECT 0.160 186.800 98.720 187.120 ;
                RECT 117.440 186.800 129.320 187.120 ;
                RECT 131.720 186.800 301.360 187.120 ;
                RECT 706.320 186.800 715.800 187.120 ;
                RECT 0.160 188.160 98.720 188.480 ;
                RECT 117.440 188.160 120.480 188.480 ;
                RECT 127.640 188.160 195.280 188.480 ;
                RECT 269.080 188.160 301.360 188.480 ;
                RECT 706.320 188.160 715.800 188.480 ;
                RECT 0.160 189.520 98.720 189.840 ;
                RECT 117.440 189.520 119.800 189.840 ;
                RECT 137.840 189.520 195.280 189.840 ;
                RECT 269.080 189.520 301.360 189.840 ;
                RECT 706.320 189.520 715.800 189.840 ;
                RECT 0.160 190.880 98.720 191.200 ;
                RECT 130.360 190.880 195.280 191.200 ;
                RECT 269.080 190.880 301.360 191.200 ;
                RECT 706.320 190.880 715.800 191.200 ;
                RECT 0.160 192.240 98.720 192.560 ;
                RECT 117.440 192.240 120.480 192.560 ;
                RECT 133.760 192.240 195.280 192.560 ;
                RECT 269.080 192.240 301.360 192.560 ;
                RECT 706.320 192.240 715.800 192.560 ;
                RECT 0.160 193.600 98.720 193.920 ;
                RECT 117.440 193.600 135.440 193.920 ;
                RECT 137.840 193.600 195.280 193.920 ;
                RECT 269.080 193.600 301.360 193.920 ;
                RECT 706.320 193.600 715.800 193.920 ;
                RECT 0.160 194.960 98.720 195.280 ;
                RECT 117.440 194.960 301.360 195.280 ;
                RECT 706.320 194.960 715.800 195.280 ;
                RECT 0.160 196.320 98.720 196.640 ;
                RECT 117.440 196.320 132.040 196.640 ;
                RECT 139.880 196.320 301.360 196.640 ;
                RECT 706.320 196.320 715.800 196.640 ;
                RECT 0.160 197.680 98.720 198.000 ;
                RECT 117.440 197.680 282.320 198.000 ;
                RECT 706.320 197.680 715.800 198.000 ;
                RECT 0.160 199.040 98.720 199.360 ;
                RECT 117.440 199.040 202.080 199.360 ;
                RECT 269.760 199.040 282.320 199.360 ;
                RECT 706.320 199.040 715.800 199.360 ;
                RECT 0.160 200.400 98.720 200.720 ;
                RECT 117.440 200.400 122.520 200.720 ;
                RECT 125.600 200.400 202.080 200.720 ;
                RECT 269.760 200.400 282.320 200.720 ;
                RECT 706.320 200.400 715.800 200.720 ;
                RECT 0.160 201.760 98.720 202.080 ;
                RECT 117.440 201.760 119.800 202.080 ;
                RECT 124.240 201.760 202.080 202.080 ;
                RECT 269.760 201.760 287.760 202.080 ;
                RECT 706.320 201.760 715.800 202.080 ;
                RECT 0.160 203.120 98.720 203.440 ;
                RECT 117.440 203.120 202.080 203.440 ;
                RECT 269.760 203.120 287.760 203.440 ;
                RECT 706.320 203.120 715.800 203.440 ;
                RECT 0.160 204.480 98.720 204.800 ;
                RECT 117.440 204.480 202.080 204.800 ;
                RECT 269.760 204.480 293.200 204.800 ;
                RECT 706.320 204.480 715.800 204.800 ;
                RECT 0.160 205.840 98.720 206.160 ;
                RECT 117.440 205.840 125.240 206.160 ;
                RECT 137.840 205.840 202.080 206.160 ;
                RECT 269.760 205.840 293.200 206.160 ;
                RECT 706.320 205.840 715.800 206.160 ;
                RECT 0.160 207.200 98.720 207.520 ;
                RECT 117.440 207.200 202.080 207.520 ;
                RECT 269.760 207.200 298.640 207.520 ;
                RECT 706.320 207.200 715.800 207.520 ;
                RECT 0.160 208.560 98.720 208.880 ;
                RECT 117.440 208.560 202.080 208.880 ;
                RECT 269.760 208.560 298.640 208.880 ;
                RECT 706.320 208.560 715.800 208.880 ;
                RECT 0.160 209.920 98.720 210.240 ;
                RECT 117.440 209.920 202.080 210.240 ;
                RECT 269.760 209.920 301.360 210.240 ;
                RECT 706.320 209.920 715.800 210.240 ;
                RECT 0.160 211.280 98.720 211.600 ;
                RECT 117.440 211.280 122.520 211.600 ;
                RECT 126.960 211.280 202.080 211.600 ;
                RECT 706.320 211.280 715.800 211.600 ;
                RECT 0.160 212.640 98.720 212.960 ;
                RECT 117.440 212.640 202.080 212.960 ;
                RECT 706.320 212.640 715.800 212.960 ;
                RECT 0.160 214.000 98.720 214.320 ;
                RECT 117.440 214.000 135.440 214.320 ;
                RECT 138.520 214.000 202.080 214.320 ;
                RECT 706.320 214.000 715.800 214.320 ;
                RECT 0.160 215.360 98.720 215.680 ;
                RECT 117.440 215.360 202.080 215.680 ;
                RECT 269.760 215.360 301.360 215.680 ;
                RECT 706.320 215.360 715.800 215.680 ;
                RECT 0.160 216.720 98.720 217.040 ;
                RECT 117.440 216.720 202.080 217.040 ;
                RECT 269.760 216.720 301.360 217.040 ;
                RECT 706.320 216.720 715.800 217.040 ;
                RECT 0.160 218.080 98.720 218.400 ;
                RECT 117.440 218.080 121.840 218.400 ;
                RECT 124.920 218.080 202.080 218.400 ;
                RECT 269.760 218.080 301.360 218.400 ;
                RECT 706.320 218.080 715.800 218.400 ;
                RECT 0.160 219.440 98.720 219.760 ;
                RECT 117.440 219.440 202.080 219.760 ;
                RECT 269.760 219.440 301.360 219.760 ;
                RECT 706.320 219.440 715.800 219.760 ;
                RECT 0.160 220.800 98.720 221.120 ;
                RECT 117.440 220.800 202.080 221.120 ;
                RECT 269.760 220.800 301.360 221.120 ;
                RECT 706.320 220.800 715.800 221.120 ;
                RECT 0.160 222.160 98.720 222.480 ;
                RECT 117.440 222.160 128.640 222.480 ;
                RECT 137.160 222.160 202.080 222.480 ;
                RECT 269.760 222.160 301.360 222.480 ;
                RECT 706.320 222.160 715.800 222.480 ;
                RECT 0.160 223.520 98.720 223.840 ;
                RECT 117.440 223.520 202.080 223.840 ;
                RECT 269.760 223.520 301.360 223.840 ;
                RECT 706.320 223.520 715.800 223.840 ;
                RECT 0.160 224.880 98.720 225.200 ;
                RECT 117.440 224.880 125.240 225.200 ;
                RECT 127.640 224.880 202.080 225.200 ;
                RECT 269.760 224.880 301.360 225.200 ;
                RECT 706.320 224.880 715.800 225.200 ;
                RECT 0.160 226.240 98.720 226.560 ;
                RECT 117.440 226.240 202.080 226.560 ;
                RECT 269.760 226.240 301.360 226.560 ;
                RECT 706.320 226.240 715.800 226.560 ;
                RECT 0.160 227.600 98.720 227.920 ;
                RECT 117.440 227.600 202.080 227.920 ;
                RECT 269.760 227.600 301.360 227.920 ;
                RECT 706.320 227.600 715.800 227.920 ;
                RECT 0.160 228.960 98.720 229.280 ;
                RECT 117.440 228.960 202.080 229.280 ;
                RECT 269.760 228.960 301.360 229.280 ;
                RECT 706.320 228.960 715.800 229.280 ;
                RECT 0.160 230.320 98.720 230.640 ;
                RECT 117.440 230.320 202.080 230.640 ;
                RECT 269.760 230.320 301.360 230.640 ;
                RECT 706.320 230.320 715.800 230.640 ;
                RECT 0.160 231.680 98.720 232.000 ;
                RECT 117.440 231.680 202.080 232.000 ;
                RECT 269.760 231.680 301.360 232.000 ;
                RECT 706.320 231.680 715.800 232.000 ;
                RECT 0.160 233.040 202.080 233.360 ;
                RECT 269.760 233.040 301.360 233.360 ;
                RECT 706.320 233.040 715.800 233.360 ;
                RECT 0.160 234.400 202.080 234.720 ;
                RECT 269.760 234.400 301.360 234.720 ;
                RECT 706.320 234.400 715.800 234.720 ;
                RECT 0.160 235.760 202.080 236.080 ;
                RECT 269.760 235.760 301.360 236.080 ;
                RECT 706.320 235.760 715.800 236.080 ;
                RECT 0.160 237.120 79.000 237.440 ;
                RECT 98.400 237.120 123.880 237.440 ;
                RECT 127.640 237.120 202.080 237.440 ;
                RECT 269.760 237.120 301.360 237.440 ;
                RECT 706.320 237.120 715.800 237.440 ;
                RECT 0.160 238.480 79.000 238.800 ;
                RECT 98.400 238.480 202.080 238.800 ;
                RECT 269.760 238.480 301.360 238.800 ;
                RECT 706.320 238.480 715.800 238.800 ;
                RECT 0.160 239.840 79.000 240.160 ;
                RECT 98.400 239.840 104.840 240.160 ;
                RECT 112.000 239.840 202.080 240.160 ;
                RECT 269.760 239.840 301.360 240.160 ;
                RECT 706.320 239.840 715.800 240.160 ;
                RECT 0.160 241.200 79.000 241.520 ;
                RECT 98.400 241.200 125.920 241.520 ;
                RECT 131.720 241.200 202.080 241.520 ;
                RECT 269.760 241.200 301.360 241.520 ;
                RECT 706.320 241.200 715.800 241.520 ;
                RECT 0.160 242.560 79.000 242.880 ;
                RECT 98.400 242.560 99.400 242.880 ;
                RECT 116.760 242.560 202.080 242.880 ;
                RECT 706.320 242.560 715.800 242.880 ;
                RECT 0.160 243.920 79.000 244.240 ;
                RECT 98.400 243.920 99.400 244.240 ;
                RECT 116.760 243.920 202.080 244.240 ;
                RECT 706.320 243.920 715.800 244.240 ;
                RECT 0.160 245.280 79.000 245.600 ;
                RECT 98.400 245.280 202.080 245.600 ;
                RECT 706.320 245.280 715.800 245.600 ;
                RECT 0.160 246.640 73.560 246.960 ;
                RECT 112.000 246.640 120.480 246.960 ;
                RECT 130.360 246.640 202.080 246.960 ;
                RECT 269.760 246.640 301.360 246.960 ;
                RECT 706.320 246.640 715.800 246.960 ;
                RECT 0.160 248.000 104.840 248.320 ;
                RECT 124.920 248.000 715.800 248.320 ;
                RECT 0.160 249.360 33.440 249.680 ;
                RECT 124.240 249.360 715.800 249.680 ;
                RECT 0.160 250.720 298.640 251.040 ;
                RECT 708.360 250.720 715.800 251.040 ;
                RECT 0.160 252.080 298.640 252.400 ;
                RECT 708.360 252.080 715.800 252.400 ;
                RECT 0.160 253.440 28.680 253.760 ;
                RECT 35.160 253.440 106.200 253.760 ;
                RECT 708.360 253.440 715.800 253.760 ;
                RECT 0.160 254.800 26.640 255.120 ;
                RECT 37.200 254.800 38.200 255.120 ;
                RECT 50.800 254.800 106.200 255.120 ;
                RECT 708.360 254.800 715.800 255.120 ;
                RECT 0.160 256.160 26.640 256.480 ;
                RECT 37.200 256.160 39.560 256.480 ;
                RECT 50.120 256.160 62.680 256.480 ;
                RECT 64.400 256.160 77.640 256.480 ;
                RECT 95.680 256.160 106.200 256.480 ;
                RECT 708.360 256.160 715.800 256.480 ;
                RECT 0.160 257.520 62.680 257.840 ;
                RECT 64.400 257.520 77.640 257.840 ;
                RECT 95.680 257.520 106.200 257.840 ;
                RECT 708.360 257.520 715.800 257.840 ;
                RECT 0.160 258.880 26.640 259.200 ;
                RECT 37.200 258.880 62.680 259.200 ;
                RECT 67.120 258.880 77.640 259.200 ;
                RECT 95.680 258.880 106.200 259.200 ;
                RECT 708.360 258.880 715.800 259.200 ;
                RECT 0.160 260.240 62.680 260.560 ;
                RECT 67.800 260.240 77.640 260.560 ;
                RECT 95.680 260.240 106.200 260.560 ;
                RECT 708.360 260.240 715.800 260.560 ;
                RECT 0.160 261.600 26.640 261.920 ;
                RECT 37.200 261.600 62.680 261.920 ;
                RECT 68.480 261.600 77.640 261.920 ;
                RECT 95.680 261.600 106.200 261.920 ;
                RECT 708.360 261.600 715.800 261.920 ;
                RECT 0.160 262.960 26.640 263.280 ;
                RECT 37.200 262.960 106.200 263.280 ;
                RECT 708.360 262.960 715.800 263.280 ;
                RECT 0.160 264.320 77.640 264.640 ;
                RECT 95.680 264.320 106.200 264.640 ;
                RECT 708.360 264.320 715.800 264.640 ;
                RECT 0.160 265.680 77.640 266.000 ;
                RECT 95.680 265.680 106.200 266.000 ;
                RECT 708.360 265.680 715.800 266.000 ;
                RECT 0.160 267.040 77.640 267.360 ;
                RECT 95.680 267.040 106.200 267.360 ;
                RECT 708.360 267.040 715.800 267.360 ;
                RECT 0.160 268.400 19.840 268.720 ;
                RECT 22.240 268.400 35.480 268.720 ;
                RECT 38.560 268.400 77.640 268.720 ;
                RECT 95.680 268.400 106.200 268.720 ;
                RECT 708.360 268.400 715.800 268.720 ;
                RECT 0.160 269.760 19.160 270.080 ;
                RECT 22.240 269.760 40.240 270.080 ;
                RECT 51.480 269.760 77.640 270.080 ;
                RECT 88.880 269.760 106.200 270.080 ;
                RECT 708.360 269.760 715.800 270.080 ;
                RECT 0.160 271.120 18.480 271.440 ;
                RECT 22.240 271.120 41.600 271.440 ;
                RECT 50.800 271.120 89.880 271.440 ;
                RECT 95.680 271.120 106.200 271.440 ;
                RECT 708.360 271.120 715.800 271.440 ;
                RECT 0.160 272.480 17.800 272.800 ;
                RECT 22.240 272.480 62.680 272.800 ;
                RECT 65.080 272.480 77.640 272.800 ;
                RECT 95.680 272.480 106.200 272.800 ;
                RECT 708.360 272.480 715.800 272.800 ;
                RECT 0.160 273.840 62.680 274.160 ;
                RECT 65.760 273.840 77.640 274.160 ;
                RECT 95.680 273.840 106.200 274.160 ;
                RECT 708.360 273.840 715.800 274.160 ;
                RECT 0.160 275.200 17.120 275.520 ;
                RECT 22.240 275.200 62.680 275.520 ;
                RECT 65.760 275.200 77.640 275.520 ;
                RECT 95.680 275.200 106.200 275.520 ;
                RECT 708.360 275.200 715.800 275.520 ;
                RECT 0.160 276.560 16.440 276.880 ;
                RECT 22.240 276.560 62.680 276.880 ;
                RECT 64.400 276.560 77.640 276.880 ;
                RECT 95.680 276.560 106.200 276.880 ;
                RECT 708.360 276.560 715.800 276.880 ;
                RECT 0.160 277.920 62.680 278.240 ;
                RECT 66.440 277.920 77.640 278.240 ;
                RECT 88.880 277.920 106.200 278.240 ;
                RECT 708.360 277.920 715.800 278.240 ;
                RECT 0.160 279.280 15.760 279.600 ;
                RECT 22.240 279.280 35.480 279.600 ;
                RECT 42.640 279.280 77.640 279.600 ;
                RECT 95.680 279.280 106.200 279.600 ;
                RECT 708.360 279.280 715.800 279.600 ;
                RECT 0.160 280.640 15.080 280.960 ;
                RECT 22.240 280.640 35.480 280.960 ;
                RECT 43.320 280.640 77.640 280.960 ;
                RECT 95.680 280.640 106.200 280.960 ;
                RECT 708.360 280.640 715.800 280.960 ;
                RECT 0.160 282.000 77.640 282.320 ;
                RECT 95.680 282.000 106.200 282.320 ;
                RECT 708.360 282.000 715.800 282.320 ;
                RECT 0.160 283.360 14.400 283.680 ;
                RECT 22.240 283.360 35.480 283.680 ;
                RECT 43.320 283.360 77.640 283.680 ;
                RECT 95.680 283.360 106.200 283.680 ;
                RECT 708.360 283.360 715.800 283.680 ;
                RECT 0.160 284.720 13.720 285.040 ;
                RECT 22.240 284.720 35.480 285.040 ;
                RECT 42.640 284.720 77.640 285.040 ;
                RECT 95.680 284.720 106.200 285.040 ;
                RECT 708.360 284.720 715.800 285.040 ;
                RECT 0.160 286.080 13.040 286.400 ;
                RECT 22.240 286.080 106.200 286.400 ;
                RECT 708.360 286.080 715.800 286.400 ;
                RECT 0.160 287.440 12.360 287.760 ;
                RECT 22.240 287.440 77.640 287.760 ;
                RECT 95.680 287.440 106.200 287.760 ;
                RECT 708.360 287.440 715.800 287.760 ;
                RECT 0.160 288.800 77.640 289.120 ;
                RECT 95.680 288.800 106.200 289.120 ;
                RECT 708.360 288.800 715.800 289.120 ;
                RECT 0.160 290.160 11.680 290.480 ;
                RECT 22.240 290.160 77.640 290.480 ;
                RECT 95.680 290.160 106.200 290.480 ;
                RECT 708.360 290.160 715.800 290.480 ;
                RECT 0.160 291.520 11.000 291.840 ;
                RECT 22.240 291.520 77.640 291.840 ;
                RECT 95.680 291.520 106.200 291.840 ;
                RECT 708.360 291.520 715.800 291.840 ;
                RECT 0.160 292.880 10.320 293.200 ;
                RECT 22.240 292.880 77.640 293.200 ;
                RECT 95.680 292.880 106.200 293.200 ;
                RECT 708.360 292.880 715.800 293.200 ;
                RECT 0.160 294.240 106.200 294.560 ;
                RECT 708.360 294.240 715.800 294.560 ;
                RECT 0.160 295.600 9.640 295.920 ;
                RECT 22.240 295.600 35.480 295.920 ;
                RECT 38.560 295.600 77.640 295.920 ;
                RECT 95.680 295.600 106.200 295.920 ;
                RECT 708.360 295.600 715.800 295.920 ;
                RECT 0.160 296.960 77.640 297.280 ;
                RECT 95.680 296.960 106.200 297.280 ;
                RECT 708.360 296.960 715.800 297.280 ;
                RECT 0.160 298.320 77.640 298.640 ;
                RECT 95.680 298.320 106.200 298.640 ;
                RECT 708.360 298.320 715.800 298.640 ;
                RECT 0.160 299.680 77.640 300.000 ;
                RECT 95.680 299.680 106.200 300.000 ;
                RECT 708.360 299.680 715.800 300.000 ;
                RECT 0.160 301.040 77.640 301.360 ;
                RECT 95.680 301.040 106.200 301.360 ;
                RECT 708.360 301.040 715.800 301.360 ;
                RECT 0.160 302.400 106.200 302.720 ;
                RECT 708.360 302.400 715.800 302.720 ;
                RECT 0.160 303.760 77.640 304.080 ;
                RECT 95.680 303.760 106.200 304.080 ;
                RECT 708.360 303.760 715.800 304.080 ;
                RECT 0.160 305.120 77.640 305.440 ;
                RECT 95.680 305.120 106.200 305.440 ;
                RECT 708.360 305.120 715.800 305.440 ;
                RECT 0.160 306.480 77.640 306.800 ;
                RECT 95.680 306.480 106.200 306.800 ;
                RECT 708.360 306.480 715.800 306.800 ;
                RECT 0.160 307.840 77.640 308.160 ;
                RECT 95.680 307.840 106.200 308.160 ;
                RECT 708.360 307.840 715.800 308.160 ;
                RECT 0.160 309.200 77.640 309.520 ;
                RECT 92.280 309.200 106.200 309.520 ;
                RECT 708.360 309.200 715.800 309.520 ;
                RECT 0.160 310.560 91.920 310.880 ;
                RECT 95.680 310.560 106.200 310.880 ;
                RECT 708.360 310.560 715.800 310.880 ;
                RECT 0.160 311.920 77.640 312.240 ;
                RECT 95.680 311.920 106.200 312.240 ;
                RECT 708.360 311.920 715.800 312.240 ;
                RECT 0.160 313.280 77.640 313.600 ;
                RECT 95.680 313.280 106.200 313.600 ;
                RECT 708.360 313.280 715.800 313.600 ;
                RECT 0.160 314.640 77.640 314.960 ;
                RECT 95.680 314.640 106.200 314.960 ;
                RECT 708.360 314.640 715.800 314.960 ;
                RECT 0.160 316.000 77.640 316.320 ;
                RECT 95.680 316.000 106.200 316.320 ;
                RECT 708.360 316.000 715.800 316.320 ;
                RECT 0.160 317.360 77.640 317.680 ;
                RECT 92.280 317.360 106.200 317.680 ;
                RECT 708.360 317.360 715.800 317.680 ;
                RECT 0.160 318.720 77.640 319.040 ;
                RECT 95.680 318.720 106.200 319.040 ;
                RECT 708.360 318.720 715.800 319.040 ;
                RECT 0.160 320.080 77.640 320.400 ;
                RECT 95.680 320.080 106.200 320.400 ;
                RECT 708.360 320.080 715.800 320.400 ;
                RECT 0.160 321.440 77.640 321.760 ;
                RECT 95.680 321.440 106.200 321.760 ;
                RECT 708.360 321.440 715.800 321.760 ;
                RECT 0.160 322.800 77.640 323.120 ;
                RECT 95.680 322.800 106.200 323.120 ;
                RECT 708.360 322.800 715.800 323.120 ;
                RECT 0.160 324.160 77.640 324.480 ;
                RECT 95.680 324.160 106.200 324.480 ;
                RECT 708.360 324.160 715.800 324.480 ;
                RECT 0.160 325.520 106.200 325.840 ;
                RECT 708.360 325.520 715.800 325.840 ;
                RECT 0.160 326.880 77.640 327.200 ;
                RECT 95.680 326.880 106.200 327.200 ;
                RECT 708.360 326.880 715.800 327.200 ;
                RECT 0.160 328.240 77.640 328.560 ;
                RECT 95.680 328.240 106.200 328.560 ;
                RECT 708.360 328.240 715.800 328.560 ;
                RECT 0.160 329.600 77.640 329.920 ;
                RECT 95.680 329.600 106.200 329.920 ;
                RECT 708.360 329.600 715.800 329.920 ;
                RECT 0.160 330.960 77.640 331.280 ;
                RECT 95.680 330.960 106.200 331.280 ;
                RECT 708.360 330.960 715.800 331.280 ;
                RECT 0.160 332.320 77.640 332.640 ;
                RECT 95.680 332.320 106.200 332.640 ;
                RECT 708.360 332.320 715.800 332.640 ;
                RECT 0.160 333.680 106.200 334.000 ;
                RECT 708.360 333.680 715.800 334.000 ;
                RECT 0.160 335.040 77.640 335.360 ;
                RECT 95.680 335.040 106.200 335.360 ;
                RECT 708.360 335.040 715.800 335.360 ;
                RECT 0.160 336.400 77.640 336.720 ;
                RECT 95.680 336.400 106.200 336.720 ;
                RECT 708.360 336.400 715.800 336.720 ;
                RECT 0.160 337.760 77.640 338.080 ;
                RECT 95.680 337.760 106.200 338.080 ;
                RECT 708.360 337.760 715.800 338.080 ;
                RECT 0.160 339.120 77.640 339.440 ;
                RECT 95.680 339.120 106.200 339.440 ;
                RECT 708.360 339.120 715.800 339.440 ;
                RECT 0.160 340.480 77.640 340.800 ;
                RECT 95.680 340.480 106.200 340.800 ;
                RECT 708.360 340.480 715.800 340.800 ;
                RECT 0.160 341.840 106.200 342.160 ;
                RECT 708.360 341.840 715.800 342.160 ;
                RECT 0.160 343.200 77.640 343.520 ;
                RECT 95.680 343.200 106.200 343.520 ;
                RECT 708.360 343.200 715.800 343.520 ;
                RECT 0.160 344.560 77.640 344.880 ;
                RECT 95.680 344.560 106.200 344.880 ;
                RECT 708.360 344.560 715.800 344.880 ;
                RECT 0.160 345.920 77.640 346.240 ;
                RECT 95.680 345.920 106.200 346.240 ;
                RECT 708.360 345.920 715.800 346.240 ;
                RECT 0.160 347.280 77.640 347.600 ;
                RECT 95.680 347.280 106.200 347.600 ;
                RECT 708.360 347.280 715.800 347.600 ;
                RECT 0.160 348.640 77.640 348.960 ;
                RECT 95.000 348.640 106.200 348.960 ;
                RECT 708.360 348.640 715.800 348.960 ;
                RECT 0.160 350.000 85.800 350.320 ;
                RECT 95.680 350.000 106.200 350.320 ;
                RECT 708.360 350.000 715.800 350.320 ;
                RECT 0.160 351.360 79.680 351.680 ;
                RECT 95.680 351.360 106.200 351.680 ;
                RECT 708.360 351.360 715.800 351.680 ;
                RECT 0.160 352.720 79.680 353.040 ;
                RECT 95.680 352.720 106.200 353.040 ;
                RECT 708.360 352.720 715.800 353.040 ;
                RECT 0.160 354.080 79.680 354.400 ;
                RECT 95.680 354.080 106.200 354.400 ;
                RECT 708.360 354.080 715.800 354.400 ;
                RECT 0.160 355.440 79.680 355.760 ;
                RECT 95.680 355.440 106.200 355.760 ;
                RECT 708.360 355.440 715.800 355.760 ;
                RECT 0.160 356.800 42.280 357.120 ;
                RECT 51.480 356.800 106.200 357.120 ;
                RECT 708.360 356.800 715.800 357.120 ;
                RECT 0.160 358.160 40.920 358.480 ;
                RECT 50.800 358.160 62.680 358.480 ;
                RECT 64.400 358.160 77.640 358.480 ;
                RECT 95.680 358.160 106.200 358.480 ;
                RECT 708.360 358.160 715.800 358.480 ;
                RECT 0.160 359.520 62.680 359.840 ;
                RECT 67.120 359.520 77.640 359.840 ;
                RECT 95.680 359.520 106.200 359.840 ;
                RECT 708.360 359.520 715.800 359.840 ;
                RECT 0.160 360.880 62.680 361.200 ;
                RECT 67.120 360.880 77.640 361.200 ;
                RECT 95.680 360.880 106.200 361.200 ;
                RECT 708.360 360.880 715.800 361.200 ;
                RECT 0.160 362.240 62.680 362.560 ;
                RECT 67.800 362.240 77.640 362.560 ;
                RECT 95.680 362.240 106.200 362.560 ;
                RECT 708.360 362.240 715.800 362.560 ;
                RECT 0.160 363.600 62.680 363.920 ;
                RECT 64.400 363.600 77.640 363.920 ;
                RECT 95.680 363.600 106.200 363.920 ;
                RECT 708.360 363.600 715.800 363.920 ;
                RECT 0.160 364.960 106.200 365.280 ;
                RECT 708.360 364.960 715.800 365.280 ;
                RECT 0.160 366.320 77.640 366.640 ;
                RECT 95.680 366.320 106.200 366.640 ;
                RECT 708.360 366.320 715.800 366.640 ;
                RECT 0.160 367.680 77.640 368.000 ;
                RECT 95.680 367.680 106.200 368.000 ;
                RECT 708.360 367.680 715.800 368.000 ;
                RECT 0.160 369.040 77.640 369.360 ;
                RECT 95.680 369.040 106.200 369.360 ;
                RECT 708.360 369.040 715.800 369.360 ;
                RECT 0.160 370.400 77.640 370.720 ;
                RECT 95.680 370.400 106.200 370.720 ;
                RECT 708.360 370.400 715.800 370.720 ;
                RECT 0.160 371.760 77.640 372.080 ;
                RECT 95.680 371.760 106.200 372.080 ;
                RECT 708.360 371.760 715.800 372.080 ;
                RECT 0.160 373.120 38.880 373.440 ;
                RECT 50.800 373.120 106.200 373.440 ;
                RECT 708.360 373.120 715.800 373.440 ;
                RECT 0.160 374.480 37.520 374.800 ;
                RECT 50.120 374.480 62.680 374.800 ;
                RECT 64.400 374.480 77.640 374.800 ;
                RECT 95.680 374.480 106.200 374.800 ;
                RECT 708.360 374.480 715.800 374.800 ;
                RECT 0.160 375.840 62.680 376.160 ;
                RECT 65.080 375.840 77.640 376.160 ;
                RECT 95.680 375.840 106.200 376.160 ;
                RECT 708.360 375.840 715.800 376.160 ;
                RECT 0.160 377.200 62.680 377.520 ;
                RECT 65.760 377.200 77.640 377.520 ;
                RECT 95.680 377.200 106.200 377.520 ;
                RECT 708.360 377.200 715.800 377.520 ;
                RECT 0.160 378.560 62.680 378.880 ;
                RECT 65.760 378.560 77.640 378.880 ;
                RECT 95.680 378.560 106.200 378.880 ;
                RECT 708.360 378.560 715.800 378.880 ;
                RECT 0.160 379.920 62.680 380.240 ;
                RECT 66.440 379.920 77.640 380.240 ;
                RECT 95.680 379.920 106.200 380.240 ;
                RECT 708.360 379.920 715.800 380.240 ;
                RECT 0.160 381.280 106.200 381.600 ;
                RECT 708.360 381.280 715.800 381.600 ;
                RECT 0.160 382.640 77.640 382.960 ;
                RECT 95.680 382.640 106.200 382.960 ;
                RECT 708.360 382.640 715.800 382.960 ;
                RECT 0.160 384.000 77.640 384.320 ;
                RECT 95.680 384.000 106.200 384.320 ;
                RECT 708.360 384.000 715.800 384.320 ;
                RECT 0.160 385.360 77.640 385.680 ;
                RECT 95.680 385.360 106.200 385.680 ;
                RECT 708.360 385.360 715.800 385.680 ;
                RECT 0.160 386.720 77.640 387.040 ;
                RECT 95.680 386.720 106.200 387.040 ;
                RECT 708.360 386.720 715.800 387.040 ;
                RECT 0.160 388.080 77.640 388.400 ;
                RECT 82.080 388.080 106.200 388.400 ;
                RECT 708.360 388.080 715.800 388.400 ;
                RECT 0.160 389.440 106.200 389.760 ;
                RECT 708.360 389.440 715.800 389.760 ;
                RECT 0.160 390.800 77.640 391.120 ;
                RECT 95.680 390.800 106.200 391.120 ;
                RECT 708.360 390.800 715.800 391.120 ;
                RECT 0.160 392.160 77.640 392.480 ;
                RECT 95.680 392.160 106.200 392.480 ;
                RECT 708.360 392.160 715.800 392.480 ;
                RECT 0.160 393.520 77.640 393.840 ;
                RECT 95.680 393.520 106.200 393.840 ;
                RECT 708.360 393.520 715.800 393.840 ;
                RECT 0.160 394.880 77.640 395.200 ;
                RECT 95.680 394.880 106.200 395.200 ;
                RECT 708.360 394.880 715.800 395.200 ;
                RECT 0.160 396.240 77.640 396.560 ;
                RECT 82.760 396.240 106.200 396.560 ;
                RECT 708.360 396.240 715.800 396.560 ;
                RECT 0.160 397.600 77.640 397.920 ;
                RECT 95.680 397.600 106.200 397.920 ;
                RECT 708.360 397.600 715.800 397.920 ;
                RECT 0.160 398.960 77.640 399.280 ;
                RECT 95.680 398.960 106.200 399.280 ;
                RECT 708.360 398.960 715.800 399.280 ;
                RECT 0.160 400.320 77.640 400.640 ;
                RECT 95.680 400.320 106.200 400.640 ;
                RECT 708.360 400.320 715.800 400.640 ;
                RECT 0.160 401.680 77.640 402.000 ;
                RECT 95.680 401.680 106.200 402.000 ;
                RECT 708.360 401.680 715.800 402.000 ;
                RECT 0.160 403.040 77.640 403.360 ;
                RECT 95.680 403.040 106.200 403.360 ;
                RECT 708.360 403.040 715.800 403.360 ;
                RECT 0.160 404.400 77.640 404.720 ;
                RECT 83.440 404.400 106.200 404.720 ;
                RECT 708.360 404.400 715.800 404.720 ;
                RECT 0.160 405.760 77.640 406.080 ;
                RECT 95.680 405.760 106.200 406.080 ;
                RECT 708.360 405.760 715.800 406.080 ;
                RECT 0.160 407.120 77.640 407.440 ;
                RECT 95.680 407.120 106.200 407.440 ;
                RECT 708.360 407.120 715.800 407.440 ;
                RECT 0.160 408.480 77.640 408.800 ;
                RECT 95.680 408.480 106.200 408.800 ;
                RECT 708.360 408.480 715.800 408.800 ;
                RECT 0.160 409.840 77.640 410.160 ;
                RECT 95.680 409.840 106.200 410.160 ;
                RECT 708.360 409.840 715.800 410.160 ;
                RECT 0.160 411.200 77.640 411.520 ;
                RECT 95.680 411.200 106.200 411.520 ;
                RECT 708.360 411.200 715.800 411.520 ;
                RECT 0.160 412.560 106.200 412.880 ;
                RECT 708.360 412.560 715.800 412.880 ;
                RECT 0.160 413.920 77.640 414.240 ;
                RECT 95.680 413.920 106.200 414.240 ;
                RECT 708.360 413.920 715.800 414.240 ;
                RECT 0.160 415.280 77.640 415.600 ;
                RECT 95.680 415.280 106.200 415.600 ;
                RECT 708.360 415.280 715.800 415.600 ;
                RECT 0.160 416.640 77.640 416.960 ;
                RECT 95.680 416.640 106.200 416.960 ;
                RECT 708.360 416.640 715.800 416.960 ;
                RECT 0.160 418.000 77.640 418.320 ;
                RECT 95.680 418.000 106.200 418.320 ;
                RECT 708.360 418.000 715.800 418.320 ;
                RECT 0.160 419.360 77.640 419.680 ;
                RECT 95.680 419.360 106.200 419.680 ;
                RECT 708.360 419.360 715.800 419.680 ;
                RECT 0.160 420.720 106.200 421.040 ;
                RECT 708.360 420.720 715.800 421.040 ;
                RECT 0.160 422.080 77.640 422.400 ;
                RECT 95.680 422.080 106.200 422.400 ;
                RECT 708.360 422.080 715.800 422.400 ;
                RECT 0.160 423.440 77.640 423.760 ;
                RECT 95.680 423.440 106.200 423.760 ;
                RECT 708.360 423.440 715.800 423.760 ;
                RECT 0.160 424.800 77.640 425.120 ;
                RECT 95.680 424.800 106.200 425.120 ;
                RECT 708.360 424.800 715.800 425.120 ;
                RECT 0.160 426.160 77.640 426.480 ;
                RECT 95.680 426.160 106.200 426.480 ;
                RECT 708.360 426.160 715.800 426.480 ;
                RECT 0.160 427.520 77.640 427.840 ;
                RECT 95.680 427.520 106.200 427.840 ;
                RECT 708.360 427.520 715.800 427.840 ;
                RECT 0.160 428.880 106.200 429.200 ;
                RECT 708.360 428.880 715.800 429.200 ;
                RECT 0.160 430.240 77.640 430.560 ;
                RECT 95.680 430.240 106.200 430.560 ;
                RECT 708.360 430.240 715.800 430.560 ;
                RECT 0.160 431.600 77.640 431.920 ;
                RECT 95.680 431.600 106.200 431.920 ;
                RECT 708.360 431.600 715.800 431.920 ;
                RECT 0.160 432.960 77.640 433.280 ;
                RECT 95.680 432.960 106.200 433.280 ;
                RECT 708.360 432.960 715.800 433.280 ;
                RECT 0.160 434.320 77.640 434.640 ;
                RECT 95.680 434.320 106.200 434.640 ;
                RECT 708.360 434.320 715.800 434.640 ;
                RECT 0.160 435.680 77.640 436.000 ;
                RECT 86.160 435.680 106.200 436.000 ;
                RECT 708.360 435.680 715.800 436.000 ;
                RECT 0.160 437.040 91.920 437.360 ;
                RECT 95.680 437.040 106.200 437.360 ;
                RECT 708.360 437.040 715.800 437.360 ;
                RECT 0.160 438.400 77.640 438.720 ;
                RECT 95.680 438.400 106.200 438.720 ;
                RECT 708.360 438.400 715.800 438.720 ;
                RECT 0.160 439.760 77.640 440.080 ;
                RECT 95.680 439.760 106.200 440.080 ;
                RECT 708.360 439.760 715.800 440.080 ;
                RECT 0.160 441.120 77.640 441.440 ;
                RECT 95.680 441.120 106.200 441.440 ;
                RECT 708.360 441.120 715.800 441.440 ;
                RECT 0.160 442.480 77.640 442.800 ;
                RECT 95.680 442.480 106.200 442.800 ;
                RECT 708.360 442.480 715.800 442.800 ;
                RECT 0.160 443.840 77.640 444.160 ;
                RECT 86.840 443.840 106.200 444.160 ;
                RECT 708.360 443.840 715.800 444.160 ;
                RECT 0.160 445.200 77.640 445.520 ;
                RECT 95.680 445.200 106.200 445.520 ;
                RECT 708.360 445.200 715.800 445.520 ;
                RECT 0.160 446.560 77.640 446.880 ;
                RECT 95.680 446.560 106.200 446.880 ;
                RECT 708.360 446.560 715.800 446.880 ;
                RECT 0.160 447.920 77.640 448.240 ;
                RECT 95.680 447.920 106.200 448.240 ;
                RECT 708.360 447.920 715.800 448.240 ;
                RECT 0.160 449.280 77.640 449.600 ;
                RECT 95.680 449.280 106.200 449.600 ;
                RECT 708.360 449.280 715.800 449.600 ;
                RECT 0.160 450.640 77.640 450.960 ;
                RECT 95.680 450.640 106.200 450.960 ;
                RECT 708.360 450.640 715.800 450.960 ;
                RECT 0.160 452.000 106.200 452.320 ;
                RECT 708.360 452.000 715.800 452.320 ;
                RECT 0.160 453.360 81.040 453.680 ;
                RECT 95.680 453.360 106.200 453.680 ;
                RECT 708.360 453.360 715.800 453.680 ;
                RECT 0.160 454.720 81.040 455.040 ;
                RECT 95.680 454.720 106.200 455.040 ;
                RECT 708.360 454.720 715.800 455.040 ;
                RECT 0.160 456.080 88.520 456.400 ;
                RECT 95.680 456.080 106.200 456.400 ;
                RECT 708.360 456.080 715.800 456.400 ;
                RECT 0.160 457.440 81.040 457.760 ;
                RECT 95.680 457.440 106.200 457.760 ;
                RECT 708.360 457.440 715.800 457.760 ;
                RECT 0.160 458.800 81.040 459.120 ;
                RECT 95.680 458.800 106.200 459.120 ;
                RECT 708.360 458.800 715.800 459.120 ;
                RECT 0.160 460.160 106.200 460.480 ;
                RECT 708.360 460.160 715.800 460.480 ;
                RECT 0.160 461.520 81.040 461.840 ;
                RECT 95.680 461.520 106.200 461.840 ;
                RECT 708.360 461.520 715.800 461.840 ;
                RECT 0.160 462.880 81.040 463.200 ;
                RECT 95.680 462.880 106.200 463.200 ;
                RECT 708.360 462.880 715.800 463.200 ;
                RECT 0.160 464.240 81.040 464.560 ;
                RECT 95.680 464.240 106.200 464.560 ;
                RECT 708.360 464.240 715.800 464.560 ;
                RECT 0.160 465.600 91.240 465.920 ;
                RECT 95.680 465.600 106.200 465.920 ;
                RECT 708.360 465.600 715.800 465.920 ;
                RECT 0.160 466.960 81.040 467.280 ;
                RECT 95.680 466.960 106.200 467.280 ;
                RECT 708.360 466.960 715.800 467.280 ;
                RECT 0.160 468.320 106.200 468.640 ;
                RECT 708.360 468.320 715.800 468.640 ;
                RECT 0.160 469.680 81.040 470.000 ;
                RECT 95.680 469.680 106.200 470.000 ;
                RECT 708.360 469.680 715.800 470.000 ;
                RECT 0.160 471.040 81.040 471.360 ;
                RECT 95.680 471.040 106.200 471.360 ;
                RECT 708.360 471.040 715.800 471.360 ;
                RECT 0.160 472.400 81.040 472.720 ;
                RECT 95.680 472.400 106.200 472.720 ;
                RECT 708.360 472.400 715.800 472.720 ;
                RECT 0.160 473.760 81.040 474.080 ;
                RECT 95.680 473.760 106.200 474.080 ;
                RECT 708.360 473.760 715.800 474.080 ;
                RECT 0.160 475.120 106.200 475.440 ;
                RECT 708.360 475.120 715.800 475.440 ;
                RECT 0.160 476.480 85.800 476.800 ;
                RECT 95.680 476.480 106.200 476.800 ;
                RECT 708.360 476.480 715.800 476.800 ;
                RECT 0.160 477.840 81.720 478.160 ;
                RECT 95.680 477.840 106.200 478.160 ;
                RECT 708.360 477.840 715.800 478.160 ;
                RECT 0.160 479.200 81.720 479.520 ;
                RECT 95.680 479.200 106.200 479.520 ;
                RECT 708.360 479.200 715.800 479.520 ;
                RECT 0.160 480.560 81.720 480.880 ;
                RECT 95.680 480.560 106.200 480.880 ;
                RECT 708.360 480.560 715.800 480.880 ;
                RECT 0.160 481.920 81.720 482.240 ;
                RECT 95.680 481.920 106.200 482.240 ;
                RECT 708.360 481.920 715.800 482.240 ;
                RECT 0.160 483.280 106.200 483.600 ;
                RECT 708.360 483.280 715.800 483.600 ;
                RECT 0.160 484.640 87.840 484.960 ;
                RECT 95.680 484.640 106.200 484.960 ;
                RECT 708.360 484.640 715.800 484.960 ;
                RECT 0.160 486.000 81.720 486.320 ;
                RECT 95.680 486.000 106.200 486.320 ;
                RECT 708.360 486.000 715.800 486.320 ;
                RECT 0.160 487.360 81.720 487.680 ;
                RECT 95.680 487.360 106.200 487.680 ;
                RECT 708.360 487.360 715.800 487.680 ;
                RECT 0.160 488.720 81.720 489.040 ;
                RECT 95.680 488.720 106.200 489.040 ;
                RECT 708.360 488.720 715.800 489.040 ;
                RECT 0.160 490.080 81.720 490.400 ;
                RECT 95.680 490.080 106.200 490.400 ;
                RECT 708.360 490.080 715.800 490.400 ;
                RECT 0.160 491.440 106.200 491.760 ;
                RECT 708.360 491.440 715.800 491.760 ;
                RECT 0.160 492.800 81.720 493.120 ;
                RECT 95.680 492.800 106.200 493.120 ;
                RECT 708.360 492.800 715.800 493.120 ;
                RECT 0.160 494.160 90.560 494.480 ;
                RECT 95.680 494.160 106.200 494.480 ;
                RECT 708.360 494.160 715.800 494.480 ;
                RECT 0.160 495.520 90.560 495.840 ;
                RECT 95.680 495.520 106.200 495.840 ;
                RECT 708.360 495.520 715.800 495.840 ;
                RECT 0.160 496.880 81.720 497.200 ;
                RECT 95.680 496.880 106.200 497.200 ;
                RECT 708.360 496.880 715.800 497.200 ;
                RECT 0.160 498.240 81.720 498.560 ;
                RECT 95.680 498.240 106.200 498.560 ;
                RECT 708.360 498.240 715.800 498.560 ;
                RECT 0.160 499.600 106.200 499.920 ;
                RECT 708.360 499.600 715.800 499.920 ;
                RECT 0.160 500.960 81.720 501.280 ;
                RECT 95.680 500.960 106.200 501.280 ;
                RECT 708.360 500.960 715.800 501.280 ;
                RECT 0.160 502.320 81.720 502.640 ;
                RECT 95.680 502.320 106.200 502.640 ;
                RECT 708.360 502.320 715.800 502.640 ;
                RECT 0.160 503.680 92.600 504.000 ;
                RECT 95.680 503.680 106.200 504.000 ;
                RECT 708.360 503.680 715.800 504.000 ;
                RECT 0.160 505.040 93.280 505.360 ;
                RECT 95.680 505.040 106.200 505.360 ;
                RECT 708.360 505.040 715.800 505.360 ;
                RECT 0.160 506.400 81.720 506.720 ;
                RECT 95.680 506.400 106.200 506.720 ;
                RECT 708.360 506.400 715.800 506.720 ;
                RECT 0.160 507.760 106.200 508.080 ;
                RECT 708.360 507.760 715.800 508.080 ;
                RECT 0.160 509.120 82.400 509.440 ;
                RECT 95.680 509.120 106.200 509.440 ;
                RECT 708.360 509.120 715.800 509.440 ;
                RECT 0.160 510.480 82.400 510.800 ;
                RECT 95.680 510.480 106.200 510.800 ;
                RECT 708.360 510.480 715.800 510.800 ;
                RECT 0.160 511.840 82.400 512.160 ;
                RECT 95.680 511.840 106.200 512.160 ;
                RECT 708.360 511.840 715.800 512.160 ;
                RECT 0.160 513.200 82.400 513.520 ;
                RECT 95.680 513.200 106.200 513.520 ;
                RECT 708.360 513.200 715.800 513.520 ;
                RECT 0.160 514.560 106.200 514.880 ;
                RECT 708.360 514.560 715.800 514.880 ;
                RECT 0.160 515.920 87.840 516.240 ;
                RECT 95.680 515.920 106.200 516.240 ;
                RECT 708.360 515.920 715.800 516.240 ;
                RECT 0.160 517.280 82.400 517.600 ;
                RECT 95.680 517.280 106.200 517.600 ;
                RECT 708.360 517.280 715.800 517.600 ;
                RECT 0.160 518.640 82.400 518.960 ;
                RECT 95.680 518.640 106.200 518.960 ;
                RECT 708.360 518.640 715.800 518.960 ;
                RECT 0.160 520.000 82.400 520.320 ;
                RECT 95.680 520.000 106.200 520.320 ;
                RECT 708.360 520.000 715.800 520.320 ;
                RECT 0.160 521.360 82.400 521.680 ;
                RECT 95.680 521.360 106.200 521.680 ;
                RECT 708.360 521.360 715.800 521.680 ;
                RECT 0.160 522.720 106.200 523.040 ;
                RECT 708.360 522.720 715.800 523.040 ;
                RECT 0.160 524.080 89.880 524.400 ;
                RECT 95.680 524.080 106.200 524.400 ;
                RECT 708.360 524.080 715.800 524.400 ;
                RECT 0.160 525.440 82.400 525.760 ;
                RECT 95.680 525.440 106.200 525.760 ;
                RECT 708.360 525.440 715.800 525.760 ;
                RECT 0.160 526.800 82.400 527.120 ;
                RECT 95.680 526.800 106.200 527.120 ;
                RECT 708.360 526.800 715.800 527.120 ;
                RECT 0.160 528.160 82.400 528.480 ;
                RECT 95.680 528.160 106.200 528.480 ;
                RECT 708.360 528.160 715.800 528.480 ;
                RECT 0.160 529.520 82.400 529.840 ;
                RECT 95.680 529.520 106.200 529.840 ;
                RECT 708.360 529.520 715.800 529.840 ;
                RECT 0.160 530.880 106.200 531.200 ;
                RECT 708.360 530.880 715.800 531.200 ;
                RECT 0.160 532.240 82.400 532.560 ;
                RECT 95.680 532.240 106.200 532.560 ;
                RECT 708.360 532.240 715.800 532.560 ;
                RECT 0.160 533.600 91.920 533.920 ;
                RECT 95.680 533.600 106.200 533.920 ;
                RECT 708.360 533.600 715.800 533.920 ;
                RECT 0.160 534.960 82.400 535.280 ;
                RECT 95.680 534.960 106.200 535.280 ;
                RECT 708.360 534.960 715.800 535.280 ;
                RECT 0.160 536.320 82.400 536.640 ;
                RECT 95.680 536.320 106.200 536.640 ;
                RECT 708.360 536.320 715.800 536.640 ;
                RECT 0.160 537.680 82.400 538.000 ;
                RECT 95.680 537.680 106.200 538.000 ;
                RECT 708.360 537.680 715.800 538.000 ;
                RECT 0.160 539.040 106.200 539.360 ;
                RECT 708.360 539.040 715.800 539.360 ;
                RECT 0.160 540.400 82.400 540.720 ;
                RECT 95.680 540.400 106.200 540.720 ;
                RECT 708.360 540.400 715.800 540.720 ;
                RECT 0.160 541.760 82.400 542.080 ;
                RECT 95.680 541.760 106.200 542.080 ;
                RECT 708.360 541.760 715.800 542.080 ;
                RECT 0.160 543.120 87.160 543.440 ;
                RECT 95.680 543.120 106.200 543.440 ;
                RECT 708.360 543.120 715.800 543.440 ;
                RECT 0.160 544.480 82.400 544.800 ;
                RECT 95.680 544.480 106.200 544.800 ;
                RECT 708.360 544.480 715.800 544.800 ;
                RECT 0.160 545.840 82.400 546.160 ;
                RECT 95.680 545.840 106.200 546.160 ;
                RECT 708.360 545.840 715.800 546.160 ;
                RECT 0.160 547.200 106.200 547.520 ;
                RECT 708.360 547.200 715.800 547.520 ;
                RECT 0.160 548.560 82.400 548.880 ;
                RECT 95.680 548.560 106.200 548.880 ;
                RECT 708.360 548.560 715.800 548.880 ;
                RECT 0.160 549.920 82.400 550.240 ;
                RECT 95.680 549.920 106.200 550.240 ;
                RECT 708.360 549.920 715.800 550.240 ;
                RECT 0.160 551.280 82.400 551.600 ;
                RECT 95.680 551.280 106.200 551.600 ;
                RECT 708.360 551.280 715.800 551.600 ;
                RECT 0.160 552.640 89.200 552.960 ;
                RECT 95.680 552.640 106.200 552.960 ;
                RECT 708.360 552.640 715.800 552.960 ;
                RECT 0.160 554.000 106.200 554.320 ;
                RECT 708.360 554.000 715.800 554.320 ;
                RECT 0.160 555.360 89.880 555.680 ;
                RECT 95.680 555.360 106.200 555.680 ;
                RECT 708.360 555.360 715.800 555.680 ;
                RECT 0.160 556.720 82.400 557.040 ;
                RECT 95.680 556.720 106.200 557.040 ;
                RECT 708.360 556.720 715.800 557.040 ;
                RECT 0.160 558.080 82.400 558.400 ;
                RECT 95.680 558.080 106.200 558.400 ;
                RECT 708.360 558.080 715.800 558.400 ;
                RECT 0.160 559.440 82.400 559.760 ;
                RECT 95.680 559.440 106.200 559.760 ;
                RECT 708.360 559.440 715.800 559.760 ;
                RECT 0.160 560.800 82.400 561.120 ;
                RECT 95.680 560.800 106.200 561.120 ;
                RECT 708.360 560.800 715.800 561.120 ;
                RECT 0.160 562.160 106.200 562.480 ;
                RECT 708.360 562.160 715.800 562.480 ;
                RECT 0.160 563.520 91.920 563.840 ;
                RECT 95.680 563.520 106.200 563.840 ;
                RECT 708.360 563.520 715.800 563.840 ;
                RECT 0.160 564.880 82.400 565.200 ;
                RECT 95.680 564.880 106.200 565.200 ;
                RECT 708.360 564.880 715.800 565.200 ;
                RECT 0.160 566.240 82.400 566.560 ;
                RECT 95.680 566.240 106.200 566.560 ;
                RECT 708.360 566.240 715.800 566.560 ;
                RECT 0.160 567.600 82.400 567.920 ;
                RECT 95.680 567.600 106.200 567.920 ;
                RECT 708.360 567.600 715.800 567.920 ;
                RECT 0.160 568.960 82.400 569.280 ;
                RECT 95.680 568.960 106.200 569.280 ;
                RECT 708.360 568.960 715.800 569.280 ;
                RECT 0.160 570.320 106.200 570.640 ;
                RECT 708.360 570.320 715.800 570.640 ;
                RECT 0.160 571.680 83.080 572.000 ;
                RECT 95.680 571.680 106.200 572.000 ;
                RECT 708.360 571.680 715.800 572.000 ;
                RECT 0.160 573.040 86.480 573.360 ;
                RECT 95.680 573.040 106.200 573.360 ;
                RECT 708.360 573.040 715.800 573.360 ;
                RECT 0.160 574.400 83.080 574.720 ;
                RECT 95.680 574.400 106.200 574.720 ;
                RECT 708.360 574.400 715.800 574.720 ;
                RECT 0.160 575.760 83.080 576.080 ;
                RECT 95.680 575.760 106.200 576.080 ;
                RECT 708.360 575.760 715.800 576.080 ;
                RECT 0.160 577.120 83.080 577.440 ;
                RECT 95.680 577.120 106.200 577.440 ;
                RECT 708.360 577.120 715.800 577.440 ;
                RECT 0.160 578.480 106.200 578.800 ;
                RECT 708.360 578.480 715.800 578.800 ;
                RECT 0.160 579.840 83.080 580.160 ;
                RECT 95.680 579.840 106.200 580.160 ;
                RECT 708.360 579.840 715.800 580.160 ;
                RECT 0.160 581.200 83.080 581.520 ;
                RECT 95.680 581.200 106.200 581.520 ;
                RECT 708.360 581.200 715.800 581.520 ;
                RECT 0.160 582.560 88.520 582.880 ;
                RECT 95.680 582.560 106.200 582.880 ;
                RECT 708.360 582.560 715.800 582.880 ;
                RECT 0.160 583.920 83.080 584.240 ;
                RECT 95.680 583.920 106.200 584.240 ;
                RECT 708.360 583.920 715.800 584.240 ;
                RECT 0.160 585.280 83.080 585.600 ;
                RECT 95.680 585.280 106.200 585.600 ;
                RECT 708.360 585.280 715.800 585.600 ;
                RECT 0.160 586.640 106.200 586.960 ;
                RECT 708.360 586.640 715.800 586.960 ;
                RECT 0.160 588.000 83.080 588.320 ;
                RECT 95.680 588.000 106.200 588.320 ;
                RECT 708.360 588.000 715.800 588.320 ;
                RECT 0.160 589.360 83.080 589.680 ;
                RECT 95.680 589.360 106.200 589.680 ;
                RECT 708.360 589.360 715.800 589.680 ;
                RECT 0.160 590.720 83.080 591.040 ;
                RECT 95.680 590.720 106.200 591.040 ;
                RECT 708.360 590.720 715.800 591.040 ;
                RECT 0.160 592.080 91.240 592.400 ;
                RECT 95.680 592.080 106.200 592.400 ;
                RECT 708.360 592.080 715.800 592.400 ;
                RECT 0.160 593.440 83.080 593.760 ;
                RECT 95.680 593.440 106.200 593.760 ;
                RECT 708.360 593.440 715.800 593.760 ;
                RECT 0.160 594.800 106.200 595.120 ;
                RECT 708.360 594.800 715.800 595.120 ;
                RECT 0.160 596.160 83.080 596.480 ;
                RECT 95.680 596.160 106.200 596.480 ;
                RECT 708.360 596.160 715.800 596.480 ;
                RECT 0.160 597.520 83.080 597.840 ;
                RECT 95.680 597.520 106.200 597.840 ;
                RECT 708.360 597.520 715.800 597.840 ;
                RECT 0.160 598.880 83.080 599.200 ;
                RECT 95.680 598.880 106.200 599.200 ;
                RECT 708.360 598.880 715.800 599.200 ;
                RECT 0.160 600.240 83.080 600.560 ;
                RECT 95.680 600.240 106.200 600.560 ;
                RECT 708.360 600.240 715.800 600.560 ;
                RECT 0.160 601.600 106.200 601.920 ;
                RECT 708.360 601.600 715.800 601.920 ;
                RECT 0.160 602.960 85.800 603.280 ;
                RECT 95.680 602.960 106.200 603.280 ;
                RECT 708.360 602.960 715.800 603.280 ;
                RECT 0.160 604.320 83.760 604.640 ;
                RECT 95.680 604.320 106.200 604.640 ;
                RECT 708.360 604.320 715.800 604.640 ;
                RECT 0.160 605.680 83.760 606.000 ;
                RECT 95.680 605.680 106.200 606.000 ;
                RECT 708.360 605.680 715.800 606.000 ;
                RECT 0.160 607.040 83.760 607.360 ;
                RECT 95.680 607.040 106.200 607.360 ;
                RECT 708.360 607.040 715.800 607.360 ;
                RECT 0.160 608.400 83.760 608.720 ;
                RECT 95.680 608.400 106.200 608.720 ;
                RECT 708.360 608.400 715.800 608.720 ;
                RECT 0.160 609.760 106.200 610.080 ;
                RECT 708.360 609.760 715.800 610.080 ;
                RECT 0.160 611.120 87.840 611.440 ;
                RECT 95.680 611.120 106.200 611.440 ;
                RECT 708.360 611.120 715.800 611.440 ;
                RECT 0.160 612.480 88.520 612.800 ;
                RECT 95.680 612.480 106.200 612.800 ;
                RECT 708.360 612.480 715.800 612.800 ;
                RECT 0.160 613.840 83.760 614.160 ;
                RECT 95.680 613.840 106.200 614.160 ;
                RECT 708.360 613.840 715.800 614.160 ;
                RECT 0.160 615.200 83.760 615.520 ;
                RECT 95.680 615.200 106.200 615.520 ;
                RECT 708.360 615.200 715.800 615.520 ;
                RECT 0.160 616.560 83.760 616.880 ;
                RECT 95.680 616.560 106.200 616.880 ;
                RECT 708.360 616.560 715.800 616.880 ;
                RECT 0.160 617.920 106.200 618.240 ;
                RECT 708.360 617.920 715.800 618.240 ;
                RECT 0.160 619.280 83.760 619.600 ;
                RECT 95.680 619.280 106.200 619.600 ;
                RECT 708.360 619.280 715.800 619.600 ;
                RECT 0.160 620.640 83.760 620.960 ;
                RECT 95.680 620.640 106.200 620.960 ;
                RECT 708.360 620.640 715.800 620.960 ;
                RECT 0.160 622.000 90.560 622.320 ;
                RECT 95.680 622.000 106.200 622.320 ;
                RECT 708.360 622.000 715.800 622.320 ;
                RECT 0.160 623.360 83.760 623.680 ;
                RECT 95.680 623.360 106.200 623.680 ;
                RECT 708.360 623.360 715.800 623.680 ;
                RECT 0.160 624.720 83.760 625.040 ;
                RECT 95.680 624.720 106.200 625.040 ;
                RECT 708.360 624.720 715.800 625.040 ;
                RECT 0.160 626.080 106.200 626.400 ;
                RECT 708.360 626.080 715.800 626.400 ;
                RECT 0.160 627.440 83.760 627.760 ;
                RECT 95.680 627.440 106.200 627.760 ;
                RECT 708.360 627.440 715.800 627.760 ;
                RECT 0.160 628.800 83.760 629.120 ;
                RECT 95.680 628.800 106.200 629.120 ;
                RECT 708.360 628.800 715.800 629.120 ;
                RECT 0.160 630.160 83.760 630.480 ;
                RECT 95.680 630.160 106.200 630.480 ;
                RECT 708.360 630.160 715.800 630.480 ;
                RECT 0.160 631.520 93.280 631.840 ;
                RECT 95.680 631.520 106.200 631.840 ;
                RECT 708.360 631.520 715.800 631.840 ;
                RECT 0.160 632.880 83.760 633.200 ;
                RECT 95.680 632.880 106.200 633.200 ;
                RECT 708.360 632.880 715.800 633.200 ;
                RECT 0.160 634.240 106.200 634.560 ;
                RECT 708.360 634.240 715.800 634.560 ;
                RECT 0.160 635.600 83.760 635.920 ;
                RECT 95.680 635.600 106.200 635.920 ;
                RECT 708.360 635.600 715.800 635.920 ;
                RECT 0.160 636.960 83.760 637.280 ;
                RECT 95.680 636.960 106.200 637.280 ;
                RECT 708.360 636.960 715.800 637.280 ;
                RECT 0.160 638.320 83.760 638.640 ;
                RECT 95.680 638.320 106.200 638.640 ;
                RECT 708.360 638.320 715.800 638.640 ;
                RECT 0.160 639.680 83.760 640.000 ;
                RECT 95.680 639.680 106.200 640.000 ;
                RECT 708.360 639.680 715.800 640.000 ;
                RECT 0.160 641.040 106.200 641.360 ;
                RECT 708.360 641.040 715.800 641.360 ;
                RECT 0.160 642.400 87.840 642.720 ;
                RECT 95.680 642.400 106.200 642.720 ;
                RECT 708.360 642.400 715.800 642.720 ;
                RECT 0.160 643.760 83.760 644.080 ;
                RECT 95.680 643.760 106.200 644.080 ;
                RECT 708.360 643.760 715.800 644.080 ;
                RECT 0.160 645.120 83.760 645.440 ;
                RECT 95.680 645.120 106.200 645.440 ;
                RECT 708.360 645.120 715.800 645.440 ;
                RECT 0.160 646.480 83.760 646.800 ;
                RECT 95.680 646.480 106.200 646.800 ;
                RECT 708.360 646.480 715.800 646.800 ;
                RECT 0.160 647.840 83.760 648.160 ;
                RECT 95.680 647.840 106.200 648.160 ;
                RECT 708.360 647.840 715.800 648.160 ;
                RECT 0.160 649.200 106.200 649.520 ;
                RECT 708.360 649.200 715.800 649.520 ;
                RECT 0.160 650.560 89.880 650.880 ;
                RECT 95.680 650.560 106.200 650.880 ;
                RECT 708.360 650.560 715.800 650.880 ;
                RECT 0.160 651.920 83.760 652.240 ;
                RECT 95.680 651.920 106.200 652.240 ;
                RECT 708.360 651.920 715.800 652.240 ;
                RECT 0.160 653.280 83.760 653.600 ;
                RECT 95.680 653.280 106.200 653.600 ;
                RECT 708.360 653.280 715.800 653.600 ;
                RECT 0.160 654.640 83.760 654.960 ;
                RECT 95.680 654.640 106.200 654.960 ;
                RECT 708.360 654.640 715.800 654.960 ;
                RECT 0.160 656.000 83.760 656.320 ;
                RECT 95.680 656.000 106.200 656.320 ;
                RECT 708.360 656.000 715.800 656.320 ;
                RECT 0.160 657.360 106.200 657.680 ;
                RECT 708.360 657.360 715.800 657.680 ;
                RECT 0.160 658.720 83.760 659.040 ;
                RECT 95.680 658.720 106.200 659.040 ;
                RECT 708.360 658.720 715.800 659.040 ;
                RECT 0.160 660.080 91.920 660.400 ;
                RECT 95.680 660.080 106.200 660.400 ;
                RECT 708.360 660.080 715.800 660.400 ;
                RECT 0.160 661.440 92.600 661.760 ;
                RECT 95.680 661.440 106.200 661.760 ;
                RECT 708.360 661.440 715.800 661.760 ;
                RECT 0.160 662.800 83.760 663.120 ;
                RECT 95.680 662.800 106.200 663.120 ;
                RECT 708.360 662.800 715.800 663.120 ;
                RECT 0.160 664.160 83.760 664.480 ;
                RECT 95.680 664.160 106.200 664.480 ;
                RECT 708.360 664.160 715.800 664.480 ;
                RECT 0.160 665.520 106.200 665.840 ;
                RECT 708.360 665.520 715.800 665.840 ;
                RECT 0.160 666.880 84.440 667.200 ;
                RECT 95.680 666.880 106.200 667.200 ;
                RECT 708.360 666.880 715.800 667.200 ;
                RECT 0.160 668.240 84.440 668.560 ;
                RECT 95.680 668.240 106.200 668.560 ;
                RECT 708.360 668.240 715.800 668.560 ;
                RECT 0.160 669.600 84.440 669.920 ;
                RECT 95.680 669.600 106.200 669.920 ;
                RECT 708.360 669.600 715.800 669.920 ;
                RECT 0.160 670.960 87.160 671.280 ;
                RECT 95.680 670.960 106.200 671.280 ;
                RECT 708.360 670.960 715.800 671.280 ;
                RECT 0.160 672.320 84.440 672.640 ;
                RECT 95.680 672.320 106.200 672.640 ;
                RECT 708.360 672.320 715.800 672.640 ;
                RECT 0.160 673.680 106.200 674.000 ;
                RECT 708.360 673.680 715.800 674.000 ;
                RECT 0.160 675.040 84.440 675.360 ;
                RECT 95.680 675.040 106.200 675.360 ;
                RECT 708.360 675.040 715.800 675.360 ;
                RECT 0.160 676.400 84.440 676.720 ;
                RECT 95.680 676.400 106.200 676.720 ;
                RECT 708.360 676.400 715.800 676.720 ;
                RECT 0.160 677.760 84.440 678.080 ;
                RECT 95.680 677.760 106.200 678.080 ;
                RECT 708.360 677.760 715.800 678.080 ;
                RECT 0.160 679.120 84.440 679.440 ;
                RECT 95.680 679.120 106.200 679.440 ;
                RECT 708.360 679.120 715.800 679.440 ;
                RECT 0.160 680.480 106.200 680.800 ;
                RECT 708.360 680.480 715.800 680.800 ;
                RECT 0.160 681.840 89.880 682.160 ;
                RECT 95.680 681.840 106.200 682.160 ;
                RECT 708.360 681.840 715.800 682.160 ;
                RECT 0.160 683.200 84.440 683.520 ;
                RECT 95.680 683.200 106.200 683.520 ;
                RECT 708.360 683.200 715.800 683.520 ;
                RECT 0.160 684.560 84.440 684.880 ;
                RECT 95.680 684.560 106.200 684.880 ;
                RECT 708.360 684.560 715.800 684.880 ;
                RECT 0.160 685.920 84.440 686.240 ;
                RECT 95.680 685.920 106.200 686.240 ;
                RECT 708.360 685.920 715.800 686.240 ;
                RECT 0.160 687.280 84.440 687.600 ;
                RECT 95.680 687.280 106.200 687.600 ;
                RECT 708.360 687.280 715.800 687.600 ;
                RECT 0.160 688.640 106.200 688.960 ;
                RECT 708.360 688.640 715.800 688.960 ;
                RECT 0.160 690.000 91.920 690.320 ;
                RECT 95.680 690.000 106.200 690.320 ;
                RECT 708.360 690.000 715.800 690.320 ;
                RECT 0.160 691.360 84.440 691.680 ;
                RECT 95.680 691.360 106.200 691.680 ;
                RECT 708.360 691.360 715.800 691.680 ;
                RECT 0.160 692.720 84.440 693.040 ;
                RECT 95.680 692.720 106.200 693.040 ;
                RECT 708.360 692.720 715.800 693.040 ;
                RECT 0.160 694.080 84.440 694.400 ;
                RECT 95.680 694.080 106.200 694.400 ;
                RECT 708.360 694.080 715.800 694.400 ;
                RECT 0.160 695.440 84.440 695.760 ;
                RECT 95.680 695.440 106.200 695.760 ;
                RECT 708.360 695.440 715.800 695.760 ;
                RECT 0.160 696.800 106.200 697.120 ;
                RECT 708.360 696.800 715.800 697.120 ;
                RECT 0.160 698.160 85.120 698.480 ;
                RECT 95.680 698.160 106.200 698.480 ;
                RECT 708.360 698.160 715.800 698.480 ;
                RECT 0.160 699.520 86.480 699.840 ;
                RECT 95.680 699.520 106.200 699.840 ;
                RECT 708.360 699.520 715.800 699.840 ;
                RECT 0.160 700.880 85.120 701.200 ;
                RECT 95.680 700.880 106.200 701.200 ;
                RECT 708.360 700.880 715.800 701.200 ;
                RECT 0.160 702.240 85.120 702.560 ;
                RECT 95.680 702.240 106.200 702.560 ;
                RECT 708.360 702.240 715.800 702.560 ;
                RECT 0.160 703.600 85.120 703.920 ;
                RECT 95.680 703.600 106.200 703.920 ;
                RECT 708.360 703.600 715.800 703.920 ;
                RECT 0.160 704.960 106.200 705.280 ;
                RECT 708.360 704.960 715.800 705.280 ;
                RECT 0.160 706.320 85.120 706.640 ;
                RECT 95.680 706.320 106.200 706.640 ;
                RECT 708.360 706.320 715.800 706.640 ;
                RECT 0.160 707.680 85.120 708.000 ;
                RECT 95.680 707.680 106.200 708.000 ;
                RECT 708.360 707.680 715.800 708.000 ;
                RECT 0.160 709.040 88.520 709.360 ;
                RECT 95.680 709.040 106.200 709.360 ;
                RECT 708.360 709.040 715.800 709.360 ;
                RECT 0.160 710.400 89.200 710.720 ;
                RECT 95.680 710.400 106.200 710.720 ;
                RECT 708.360 710.400 715.800 710.720 ;
                RECT 0.160 711.760 85.120 712.080 ;
                RECT 95.680 711.760 106.200 712.080 ;
                RECT 708.360 711.760 715.800 712.080 ;
                RECT 0.160 713.120 106.200 713.440 ;
                RECT 708.360 713.120 715.800 713.440 ;
                RECT 0.160 714.480 85.120 714.800 ;
                RECT 95.680 714.480 106.200 714.800 ;
                RECT 708.360 714.480 715.800 714.800 ;
                RECT 0.160 715.840 85.120 716.160 ;
                RECT 95.680 715.840 106.200 716.160 ;
                RECT 708.360 715.840 715.800 716.160 ;
                RECT 0.160 717.200 85.120 717.520 ;
                RECT 95.680 717.200 106.200 717.520 ;
                RECT 708.360 717.200 715.800 717.520 ;
                RECT 0.160 718.560 91.240 718.880 ;
                RECT 95.680 718.560 106.200 718.880 ;
                RECT 708.360 718.560 715.800 718.880 ;
                RECT 0.160 719.920 106.200 720.240 ;
                RECT 708.360 719.920 715.800 720.240 ;
                RECT 0.160 721.280 91.920 721.600 ;
                RECT 95.680 721.280 106.200 721.600 ;
                RECT 708.360 721.280 715.800 721.600 ;
                RECT 0.160 722.640 85.120 722.960 ;
                RECT 95.680 722.640 106.200 722.960 ;
                RECT 708.360 722.640 715.800 722.960 ;
                RECT 0.160 724.000 85.120 724.320 ;
                RECT 95.680 724.000 106.200 724.320 ;
                RECT 708.360 724.000 715.800 724.320 ;
                RECT 0.160 725.360 85.120 725.680 ;
                RECT 95.680 725.360 106.200 725.680 ;
                RECT 708.360 725.360 715.800 725.680 ;
                RECT 0.160 726.720 85.120 727.040 ;
                RECT 95.680 726.720 106.200 727.040 ;
                RECT 708.360 726.720 715.800 727.040 ;
                RECT 0.160 728.080 106.200 728.400 ;
                RECT 708.360 728.080 715.800 728.400 ;
                RECT 0.160 729.440 85.800 729.760 ;
                RECT 95.680 729.440 106.200 729.760 ;
                RECT 708.360 729.440 715.800 729.760 ;
                RECT 0.160 730.800 85.800 731.120 ;
                RECT 95.680 730.800 106.200 731.120 ;
                RECT 708.360 730.800 715.800 731.120 ;
                RECT 0.160 732.160 85.800 732.480 ;
                RECT 95.680 732.160 106.200 732.480 ;
                RECT 708.360 732.160 715.800 732.480 ;
                RECT 0.160 733.520 85.800 733.840 ;
                RECT 95.680 733.520 106.200 733.840 ;
                RECT 708.360 733.520 715.800 733.840 ;
                RECT 0.160 734.880 85.800 735.200 ;
                RECT 95.680 734.880 106.200 735.200 ;
                RECT 708.360 734.880 715.800 735.200 ;
                RECT 0.160 736.240 106.200 736.560 ;
                RECT 708.360 736.240 715.800 736.560 ;
                RECT 0.160 737.600 85.800 737.920 ;
                RECT 95.680 737.600 106.200 737.920 ;
                RECT 708.360 737.600 715.800 737.920 ;
                RECT 0.160 738.960 88.520 739.280 ;
                RECT 95.680 738.960 106.200 739.280 ;
                RECT 708.360 738.960 715.800 739.280 ;
                RECT 0.160 740.320 85.800 740.640 ;
                RECT 95.680 740.320 106.200 740.640 ;
                RECT 708.360 740.320 715.800 740.640 ;
                RECT 0.160 741.680 85.800 742.000 ;
                RECT 95.680 741.680 106.200 742.000 ;
                RECT 708.360 741.680 715.800 742.000 ;
                RECT 0.160 743.040 85.800 743.360 ;
                RECT 95.680 743.040 106.200 743.360 ;
                RECT 708.360 743.040 715.800 743.360 ;
                RECT 0.160 744.400 106.200 744.720 ;
                RECT 708.360 744.400 715.800 744.720 ;
                RECT 0.160 745.760 85.800 746.080 ;
                RECT 95.680 745.760 106.200 746.080 ;
                RECT 708.360 745.760 715.800 746.080 ;
                RECT 0.160 747.120 85.800 747.440 ;
                RECT 95.680 747.120 106.200 747.440 ;
                RECT 708.360 747.120 715.800 747.440 ;
                RECT 0.160 748.480 90.560 748.800 ;
                RECT 95.680 748.480 106.200 748.800 ;
                RECT 708.360 748.480 715.800 748.800 ;
                RECT 0.160 749.840 85.800 750.160 ;
                RECT 95.680 749.840 106.200 750.160 ;
                RECT 708.360 749.840 715.800 750.160 ;
                RECT 0.160 751.200 85.800 751.520 ;
                RECT 95.680 751.200 106.200 751.520 ;
                RECT 708.360 751.200 715.800 751.520 ;
                RECT 0.160 752.560 106.200 752.880 ;
                RECT 708.360 752.560 715.800 752.880 ;
                RECT 0.160 753.920 85.800 754.240 ;
                RECT 95.680 753.920 106.200 754.240 ;
                RECT 708.360 753.920 715.800 754.240 ;
                RECT 0.160 755.280 85.800 755.600 ;
                RECT 95.680 755.280 106.200 755.600 ;
                RECT 708.360 755.280 715.800 755.600 ;
                RECT 0.160 756.640 85.800 756.960 ;
                RECT 95.680 756.640 106.200 756.960 ;
                RECT 708.360 756.640 715.800 756.960 ;
                RECT 0.160 758.000 93.280 758.320 ;
                RECT 95.680 758.000 106.200 758.320 ;
                RECT 708.360 758.000 715.800 758.320 ;
                RECT 0.160 759.360 85.800 759.680 ;
                RECT 95.680 759.360 106.200 759.680 ;
                RECT 708.360 759.360 715.800 759.680 ;
                RECT 0.160 760.720 106.200 761.040 ;
                RECT 708.360 760.720 715.800 761.040 ;
                RECT 0.160 762.080 298.640 762.400 ;
                RECT 708.360 762.080 715.800 762.400 ;
                RECT 0.160 763.440 298.640 763.760 ;
                RECT 708.360 763.440 715.800 763.760 ;
                RECT 0.160 764.800 298.640 765.120 ;
                RECT 708.360 764.800 715.800 765.120 ;
                RECT 0.160 766.160 715.800 766.480 ;
                RECT 0.160 767.520 715.800 767.840 ;
                RECT 0.160 768.880 715.800 769.200 ;
                RECT 0.160 770.240 715.800 770.560 ;
                RECT 0.160 0.160 715.800 1.520 ;
                RECT 0.160 774.960 715.800 776.320 ;
                RECT 302.780 41.890 308.580 43.260 ;
                RECT 698.680 41.890 704.480 43.260 ;
                RECT 302.780 47.145 308.580 48.695 ;
                RECT 698.680 47.145 704.480 48.695 ;
                RECT 302.780 53.000 308.580 54.800 ;
                RECT 698.680 53.000 704.480 54.800 ;
                RECT 302.780 58.530 308.580 59.780 ;
                RECT 698.680 58.530 704.480 59.780 ;
                RECT 302.780 63.290 308.580 64.580 ;
                RECT 698.680 63.290 704.480 64.580 ;
                RECT 302.780 68.110 308.580 69.400 ;
                RECT 698.680 68.110 704.480 69.400 ;
                RECT 302.780 87.530 704.480 88.330 ;
                RECT 302.780 229.725 704.480 233.325 ;
                RECT 302.780 90.540 704.480 91.340 ;
                RECT 302.780 123.035 704.480 123.325 ;
                RECT 302.780 113.230 704.480 116.830 ;
                RECT 302.780 95.430 704.480 96.230 ;
                RECT 302.780 76.060 704.480 77.860 ;
                RECT 302.780 163.385 704.480 165.185 ;
                RECT 302.780 26.135 704.480 27.935 ;
                RECT 110.570 253.835 112.490 761.015 ;
                RECT 114.410 253.835 116.330 761.015 ;
                RECT 126.605 253.835 128.525 761.015 ;
                RECT 130.445 253.835 132.365 761.015 ;
                RECT 134.285 253.835 136.205 761.015 ;
                RECT 138.125 253.835 140.045 761.015 ;
                RECT 159.440 253.835 161.360 761.015 ;
                RECT 163.280 253.835 165.200 761.015 ;
                RECT 167.120 253.835 169.040 761.015 ;
                RECT 170.960 253.835 172.880 761.015 ;
                RECT 174.800 253.835 176.720 761.015 ;
                RECT 178.640 253.835 180.560 761.015 ;
                RECT 182.480 253.835 184.400 761.015 ;
                RECT 186.320 253.835 188.240 761.015 ;
                RECT 224.845 253.835 226.765 761.015 ;
                RECT 228.685 253.835 230.605 761.015 ;
                RECT 232.525 253.835 234.445 761.015 ;
                RECT 236.365 253.835 238.285 761.015 ;
                RECT 240.205 253.835 242.125 761.015 ;
                RECT 244.045 253.835 245.965 761.015 ;
                RECT 247.885 253.835 249.805 761.015 ;
                RECT 251.725 253.835 253.645 761.015 ;
                RECT 255.565 253.835 257.485 761.015 ;
                RECT 259.405 253.835 261.325 761.015 ;
                RECT 263.245 253.835 265.165 761.015 ;
                RECT 267.085 253.835 269.005 761.015 ;
                RECT 270.925 253.835 272.845 761.015 ;
                RECT 274.765 253.835 276.685 761.015 ;
                RECT 278.605 253.835 280.525 761.015 ;
                RECT 282.445 253.835 284.365 761.015 ;
                RECT 286.285 253.835 288.205 761.015 ;
                RECT 290.125 253.835 292.045 761.015 ;
                RECT 293.965 253.835 295.885 761.015 ;
                RECT 159.035 55.635 160.785 134.035 ;
                RECT 165.495 55.635 167.415 134.035 ;
                RECT 172.125 55.635 173.875 134.035 ;
                RECT 178.585 55.635 180.505 134.035 ;
                RECT 187.080 55.635 189.000 134.035 ;
                RECT 190.920 55.635 192.840 134.035 ;
                RECT 203.115 55.635 205.035 134.035 ;
                RECT 206.955 55.635 208.875 134.035 ;
                RECT 210.795 55.635 212.715 134.035 ;
                RECT 214.635 55.635 216.555 134.035 ;
                RECT 236.180 55.635 238.100 134.035 ;
                RECT 240.020 55.635 241.940 134.035 ;
                RECT 243.860 55.635 245.780 134.035 ;
                RECT 247.700 55.635 249.620 134.035 ;
                RECT 251.540 55.635 253.460 134.035 ;
                RECT 255.380 55.635 257.300 134.035 ;
                RECT 259.220 55.635 261.140 134.035 ;
                RECT 263.060 55.635 264.980 134.035 ;
                RECT 266.900 55.635 268.820 134.035 ;
                RECT 206.635 199.700 208.555 247.200 ;
                RECT 214.125 199.700 215.875 247.200 ;
                RECT 220.345 199.700 221.885 247.200 ;
                RECT 228.220 199.700 230.140 247.200 ;
                RECT 232.060 199.700 233.980 247.200 ;
                RECT 248.155 199.700 250.075 247.200 ;
                RECT 251.995 199.700 253.915 247.200 ;
                RECT 255.835 199.700 257.755 247.200 ;
                RECT 259.675 199.700 261.595 247.200 ;
                RECT 263.515 199.700 265.435 247.200 ;
                RECT 267.355 199.700 269.275 247.200 ;
                RECT 198.525 188.540 200.275 193.700 ;
                RECT 209.085 188.540 211.005 193.700 ;
                RECT 212.925 188.540 214.845 193.700 ;
                RECT 235.945 188.540 237.865 193.700 ;
                RECT 239.785 188.540 241.705 193.700 ;
                RECT 243.625 188.540 245.545 193.700 ;
                RECT 247.465 188.540 249.385 193.700 ;
                RECT 251.305 188.540 253.225 193.700 ;
                RECT 255.145 188.540 257.065 193.700 ;
                RECT 258.985 188.540 260.905 193.700 ;
                RECT 262.825 188.540 264.745 193.700 ;
                RECT 266.665 188.540 268.585 193.700 ;
                RECT 268.375 44.475 270.125 49.635 ;
                RECT 27.350 256.105 36.510 256.855 ;
                RECT 27.350 261.505 36.510 263.425 ;
                RECT 99.910 242.115 115.950 243.765 ;
                RECT 79.510 242.295 97.950 245.895 ;
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 311.560 5.560 ;
                RECT 313.280 5.240 317.680 5.560 ;
                RECT 319.400 5.240 323.800 5.560 ;
                RECT 325.520 5.240 329.920 5.560 ;
                RECT 331.640 5.240 336.040 5.560 ;
                RECT 337.760 5.240 342.160 5.560 ;
                RECT 343.880 5.240 348.280 5.560 ;
                RECT 350.000 5.240 354.400 5.560 ;
                RECT 356.120 5.240 360.520 5.560 ;
                RECT 362.240 5.240 366.640 5.560 ;
                RECT 368.360 5.240 372.760 5.560 ;
                RECT 374.480 5.240 378.880 5.560 ;
                RECT 380.600 5.240 385.000 5.560 ;
                RECT 386.720 5.240 391.120 5.560 ;
                RECT 392.840 5.240 397.240 5.560 ;
                RECT 398.960 5.240 403.360 5.560 ;
                RECT 405.080 5.240 409.480 5.560 ;
                RECT 411.200 5.240 415.600 5.560 ;
                RECT 417.320 5.240 421.720 5.560 ;
                RECT 423.440 5.240 427.840 5.560 ;
                RECT 429.560 5.240 433.960 5.560 ;
                RECT 435.680 5.240 440.080 5.560 ;
                RECT 441.800 5.240 446.200 5.560 ;
                RECT 447.920 5.240 452.320 5.560 ;
                RECT 453.360 5.240 458.440 5.560 ;
                RECT 459.480 5.240 464.560 5.560 ;
                RECT 465.600 5.240 470.680 5.560 ;
                RECT 471.720 5.240 476.800 5.560 ;
                RECT 477.840 5.240 482.920 5.560 ;
                RECT 483.960 5.240 489.040 5.560 ;
                RECT 490.080 5.240 495.160 5.560 ;
                RECT 496.200 5.240 501.280 5.560 ;
                RECT 502.320 5.240 506.720 5.560 ;
                RECT 508.440 5.240 512.840 5.560 ;
                RECT 514.560 5.240 518.960 5.560 ;
                RECT 520.680 5.240 525.080 5.560 ;
                RECT 526.800 5.240 531.200 5.560 ;
                RECT 532.920 5.240 537.320 5.560 ;
                RECT 539.040 5.240 543.440 5.560 ;
                RECT 545.160 5.240 549.560 5.560 ;
                RECT 551.280 5.240 555.680 5.560 ;
                RECT 557.400 5.240 561.800 5.560 ;
                RECT 563.520 5.240 567.920 5.560 ;
                RECT 569.640 5.240 574.040 5.560 ;
                RECT 575.760 5.240 580.160 5.560 ;
                RECT 581.880 5.240 586.280 5.560 ;
                RECT 588.000 5.240 592.400 5.560 ;
                RECT 594.120 5.240 598.520 5.560 ;
                RECT 600.240 5.240 604.640 5.560 ;
                RECT 606.360 5.240 610.760 5.560 ;
                RECT 612.480 5.240 616.880 5.560 ;
                RECT 618.600 5.240 623.000 5.560 ;
                RECT 624.720 5.240 629.120 5.560 ;
                RECT 630.840 5.240 635.240 5.560 ;
                RECT 636.960 5.240 641.360 5.560 ;
                RECT 643.080 5.240 647.480 5.560 ;
                RECT 649.200 5.240 653.600 5.560 ;
                RECT 655.320 5.240 659.720 5.560 ;
                RECT 660.760 5.240 665.840 5.560 ;
                RECT 666.880 5.240 671.960 5.560 ;
                RECT 673.000 5.240 678.080 5.560 ;
                RECT 679.120 5.240 684.200 5.560 ;
                RECT 685.240 5.240 690.320 5.560 ;
                RECT 691.360 5.240 696.440 5.560 ;
                RECT 697.480 5.240 713.080 5.560 ;
                RECT 2.880 6.600 713.080 6.920 ;
                RECT 2.880 7.960 713.080 8.280 ;
                RECT 2.880 9.320 272.120 9.640 ;
                RECT 307.160 9.320 713.080 9.640 ;
                RECT 2.880 10.680 713.080 11.000 ;
                RECT 2.880 12.040 713.080 12.360 ;
                RECT 2.880 13.400 197.320 13.720 ;
                RECT 273.160 13.400 713.080 13.720 ;
                RECT 2.880 14.760 713.080 15.080 ;
                RECT 2.880 16.120 713.080 16.440 ;
                RECT 2.880 17.480 197.320 17.800 ;
                RECT 272.480 17.480 713.080 17.800 ;
                RECT 2.880 18.840 713.080 19.160 ;
                RECT 2.880 20.200 301.360 20.520 ;
                RECT 706.320 20.200 713.080 20.520 ;
                RECT 2.880 21.560 301.360 21.880 ;
                RECT 706.320 21.560 713.080 21.880 ;
                RECT 2.880 22.920 301.360 23.240 ;
                RECT 706.320 22.920 713.080 23.240 ;
                RECT 2.880 24.280 301.360 24.600 ;
                RECT 706.320 24.280 713.080 24.600 ;
                RECT 2.880 25.640 301.360 25.960 ;
                RECT 706.320 25.640 713.080 25.960 ;
                RECT 2.880 27.000 301.360 27.320 ;
                RECT 706.320 27.000 713.080 27.320 ;
                RECT 2.880 28.360 301.360 28.680 ;
                RECT 706.320 28.360 713.080 28.680 ;
                RECT 2.880 29.720 301.360 30.040 ;
                RECT 706.320 29.720 713.080 30.040 ;
                RECT 2.880 31.080 301.360 31.400 ;
                RECT 706.320 31.080 713.080 31.400 ;
                RECT 2.880 32.440 301.360 32.760 ;
                RECT 706.320 32.440 713.080 32.760 ;
                RECT 2.880 33.800 301.360 34.120 ;
                RECT 706.320 33.800 713.080 34.120 ;
                RECT 2.880 35.160 301.360 35.480 ;
                RECT 706.320 35.160 713.080 35.480 ;
                RECT 2.880 36.520 146.320 36.840 ;
                RECT 251.400 36.520 301.360 36.840 ;
                RECT 706.320 36.520 713.080 36.840 ;
                RECT 2.880 37.880 144.960 38.200 ;
                RECT 257.520 37.880 300.680 38.200 ;
                RECT 706.320 37.880 713.080 38.200 ;
                RECT 2.880 39.240 122.520 39.560 ;
                RECT 272.480 39.240 301.360 39.560 ;
                RECT 706.320 39.240 713.080 39.560 ;
                RECT 2.880 40.600 123.200 40.920 ;
                RECT 262.960 40.600 301.360 40.920 ;
                RECT 706.320 40.600 713.080 40.920 ;
                RECT 2.880 41.960 301.360 42.280 ;
                RECT 706.320 41.960 713.080 42.280 ;
                RECT 2.880 43.320 301.360 43.640 ;
                RECT 706.320 43.320 713.080 43.640 ;
                RECT 2.880 44.680 265.320 45.000 ;
                RECT 271.120 44.680 301.360 45.000 ;
                RECT 706.320 44.680 713.080 45.000 ;
                RECT 2.880 46.040 265.320 46.360 ;
                RECT 706.320 46.040 713.080 46.360 ;
                RECT 2.880 47.400 265.320 47.720 ;
                RECT 706.320 47.400 713.080 47.720 ;
                RECT 2.880 48.760 142.920 49.080 ;
                RECT 262.280 48.760 265.320 49.080 ;
                RECT 271.120 48.760 301.360 49.080 ;
                RECT 706.320 48.760 713.080 49.080 ;
                RECT 2.880 50.120 301.360 50.440 ;
                RECT 706.320 50.120 713.080 50.440 ;
                RECT 2.880 51.480 301.360 51.800 ;
                RECT 706.320 51.480 713.080 51.800 ;
                RECT 2.880 52.840 301.360 53.160 ;
                RECT 706.320 52.840 713.080 53.160 ;
                RECT 2.880 54.200 301.360 54.520 ;
                RECT 706.320 54.200 713.080 54.520 ;
                RECT 2.880 55.560 155.840 55.880 ;
                RECT 269.760 55.560 301.360 55.880 ;
                RECT 706.320 55.560 713.080 55.880 ;
                RECT 2.880 56.920 144.960 57.240 ;
                RECT 150.080 56.920 155.840 57.240 ;
                RECT 285.400 56.920 301.360 57.240 ;
                RECT 706.320 56.920 713.080 57.240 ;
                RECT 2.880 58.280 146.320 58.600 ;
                RECT 148.720 58.280 155.840 58.600 ;
                RECT 282.680 58.280 301.360 58.600 ;
                RECT 706.320 58.280 713.080 58.600 ;
                RECT 2.880 59.640 155.840 59.960 ;
                RECT 285.400 59.640 301.360 59.960 ;
                RECT 706.320 59.640 713.080 59.960 ;
                RECT 2.880 61.000 155.840 61.320 ;
                RECT 285.400 61.000 301.360 61.320 ;
                RECT 706.320 61.000 713.080 61.320 ;
                RECT 2.880 62.360 155.840 62.680 ;
                RECT 282.680 62.360 301.360 62.680 ;
                RECT 706.320 62.360 713.080 62.680 ;
                RECT 2.880 63.720 155.840 64.040 ;
                RECT 285.400 63.720 301.360 64.040 ;
                RECT 706.320 63.720 713.080 64.040 ;
                RECT 2.880 65.080 155.840 65.400 ;
                RECT 269.760 65.080 301.360 65.400 ;
                RECT 706.320 65.080 713.080 65.400 ;
                RECT 2.880 66.440 155.840 66.760 ;
                RECT 285.400 66.440 301.360 66.760 ;
                RECT 706.320 66.440 713.080 66.760 ;
                RECT 2.880 67.800 155.840 68.120 ;
                RECT 285.400 67.800 301.360 68.120 ;
                RECT 706.320 67.800 713.080 68.120 ;
                RECT 2.880 69.160 155.840 69.480 ;
                RECT 269.760 69.160 301.360 69.480 ;
                RECT 706.320 69.160 713.080 69.480 ;
                RECT 2.880 70.520 155.840 70.840 ;
                RECT 282.680 70.520 301.360 70.840 ;
                RECT 706.320 70.520 713.080 70.840 ;
                RECT 2.880 71.880 155.840 72.200 ;
                RECT 285.400 71.880 301.360 72.200 ;
                RECT 706.320 71.880 713.080 72.200 ;
                RECT 2.880 73.240 155.840 73.560 ;
                RECT 269.760 73.240 301.360 73.560 ;
                RECT 706.320 73.240 713.080 73.560 ;
                RECT 2.880 74.600 155.840 74.920 ;
                RECT 285.400 74.600 301.360 74.920 ;
                RECT 706.320 74.600 713.080 74.920 ;
                RECT 2.880 75.960 155.840 76.280 ;
                RECT 290.840 75.960 301.360 76.280 ;
                RECT 706.320 75.960 713.080 76.280 ;
                RECT 2.880 77.320 155.840 77.640 ;
                RECT 288.120 77.320 301.360 77.640 ;
                RECT 706.320 77.320 713.080 77.640 ;
                RECT 2.880 78.680 155.840 79.000 ;
                RECT 290.840 78.680 301.360 79.000 ;
                RECT 706.320 78.680 713.080 79.000 ;
                RECT 2.880 80.040 155.840 80.360 ;
                RECT 290.840 80.040 301.360 80.360 ;
                RECT 706.320 80.040 713.080 80.360 ;
                RECT 2.880 81.400 155.840 81.720 ;
                RECT 288.120 81.400 301.360 81.720 ;
                RECT 706.320 81.400 713.080 81.720 ;
                RECT 2.880 82.760 155.840 83.080 ;
                RECT 290.840 82.760 301.360 83.080 ;
                RECT 706.320 82.760 713.080 83.080 ;
                RECT 2.880 84.120 155.840 84.440 ;
                RECT 288.120 84.120 301.360 84.440 ;
                RECT 706.320 84.120 713.080 84.440 ;
                RECT 2.880 85.480 155.840 85.800 ;
                RECT 290.840 85.480 301.360 85.800 ;
                RECT 706.320 85.480 713.080 85.800 ;
                RECT 2.880 86.840 155.840 87.160 ;
                RECT 290.840 86.840 301.360 87.160 ;
                RECT 706.320 86.840 713.080 87.160 ;
                RECT 2.880 88.200 155.840 88.520 ;
                RECT 288.120 88.200 301.360 88.520 ;
                RECT 706.320 88.200 713.080 88.520 ;
                RECT 2.880 89.560 155.840 89.880 ;
                RECT 290.840 89.560 301.360 89.880 ;
                RECT 706.320 89.560 713.080 89.880 ;
                RECT 2.880 90.920 155.840 91.240 ;
                RECT 269.760 90.920 301.360 91.240 ;
                RECT 706.320 90.920 713.080 91.240 ;
                RECT 2.880 92.280 155.840 92.600 ;
                RECT 290.840 92.280 301.360 92.600 ;
                RECT 706.320 92.280 713.080 92.600 ;
                RECT 2.880 93.640 155.840 93.960 ;
                RECT 290.840 93.640 301.360 93.960 ;
                RECT 706.320 93.640 713.080 93.960 ;
                RECT 2.880 95.000 155.840 95.320 ;
                RECT 269.760 95.000 301.360 95.320 ;
                RECT 706.320 95.000 713.080 95.320 ;
                RECT 2.880 96.360 155.840 96.680 ;
                RECT 293.560 96.360 301.360 96.680 ;
                RECT 706.320 96.360 713.080 96.680 ;
                RECT 2.880 97.720 155.840 98.040 ;
                RECT 296.280 97.720 301.360 98.040 ;
                RECT 706.320 97.720 713.080 98.040 ;
                RECT 2.880 99.080 155.840 99.400 ;
                RECT 269.760 99.080 301.360 99.400 ;
                RECT 706.320 99.080 713.080 99.400 ;
                RECT 2.880 100.440 155.840 100.760 ;
                RECT 296.280 100.440 301.360 100.760 ;
                RECT 706.320 100.440 713.080 100.760 ;
                RECT 2.880 101.800 155.840 102.120 ;
                RECT 296.280 101.800 301.360 102.120 ;
                RECT 706.320 101.800 713.080 102.120 ;
                RECT 2.880 103.160 155.840 103.480 ;
                RECT 293.560 103.160 301.360 103.480 ;
                RECT 706.320 103.160 713.080 103.480 ;
                RECT 2.880 104.520 155.840 104.840 ;
                RECT 296.280 104.520 301.360 104.840 ;
                RECT 706.320 104.520 713.080 104.840 ;
                RECT 2.880 105.880 155.840 106.200 ;
                RECT 296.280 105.880 301.360 106.200 ;
                RECT 706.320 105.880 713.080 106.200 ;
                RECT 2.880 107.240 155.840 107.560 ;
                RECT 293.560 107.240 301.360 107.560 ;
                RECT 706.320 107.240 713.080 107.560 ;
                RECT 2.880 108.600 155.840 108.920 ;
                RECT 296.280 108.600 301.360 108.920 ;
                RECT 706.320 108.600 713.080 108.920 ;
                RECT 2.880 109.960 155.840 110.280 ;
                RECT 293.560 109.960 301.360 110.280 ;
                RECT 706.320 109.960 713.080 110.280 ;
                RECT 2.880 111.320 155.840 111.640 ;
                RECT 296.280 111.320 301.360 111.640 ;
                RECT 706.320 111.320 713.080 111.640 ;
                RECT 2.880 112.680 155.840 113.000 ;
                RECT 296.280 112.680 301.360 113.000 ;
                RECT 706.320 112.680 713.080 113.000 ;
                RECT 2.880 114.040 155.840 114.360 ;
                RECT 269.760 114.040 301.360 114.360 ;
                RECT 706.320 114.040 713.080 114.360 ;
                RECT 2.880 115.400 155.840 115.720 ;
                RECT 706.320 115.400 713.080 115.720 ;
                RECT 2.880 116.760 155.840 117.080 ;
                RECT 269.760 116.760 301.360 117.080 ;
                RECT 706.320 116.760 713.080 117.080 ;
                RECT 2.880 118.120 155.840 118.440 ;
                RECT 706.320 118.120 713.080 118.440 ;
                RECT 2.880 119.480 155.840 119.800 ;
                RECT 706.320 119.480 713.080 119.800 ;
                RECT 2.880 120.840 155.840 121.160 ;
                RECT 706.320 120.840 713.080 121.160 ;
                RECT 2.880 122.200 155.840 122.520 ;
                RECT 706.320 122.200 713.080 122.520 ;
                RECT 2.880 123.560 155.840 123.880 ;
                RECT 706.320 123.560 713.080 123.880 ;
                RECT 2.880 124.920 155.840 125.240 ;
                RECT 269.760 124.920 301.360 125.240 ;
                RECT 706.320 124.920 713.080 125.240 ;
                RECT 2.880 126.280 155.840 126.600 ;
                RECT 706.320 126.280 713.080 126.600 ;
                RECT 2.880 127.640 155.840 127.960 ;
                RECT 706.320 127.640 713.080 127.960 ;
                RECT 2.880 129.000 155.840 129.320 ;
                RECT 706.320 129.000 713.080 129.320 ;
                RECT 2.880 130.360 155.840 130.680 ;
                RECT 706.320 130.360 713.080 130.680 ;
                RECT 2.880 131.720 155.840 132.040 ;
                RECT 706.320 131.720 713.080 132.040 ;
                RECT 2.880 133.080 155.840 133.400 ;
                RECT 706.320 133.080 713.080 133.400 ;
                RECT 2.880 134.440 301.360 134.760 ;
                RECT 706.320 134.440 713.080 134.760 ;
                RECT 2.880 135.800 98.720 136.120 ;
                RECT 117.440 135.800 301.360 136.120 ;
                RECT 706.320 135.800 713.080 136.120 ;
                RECT 2.880 137.160 98.720 137.480 ;
                RECT 117.440 137.160 276.880 137.480 ;
                RECT 706.320 137.160 713.080 137.480 ;
                RECT 2.880 138.520 98.720 138.840 ;
                RECT 117.440 138.520 295.920 138.840 ;
                RECT 706.320 138.520 713.080 138.840 ;
                RECT 2.880 139.880 98.720 140.200 ;
                RECT 117.440 139.880 295.920 140.200 ;
                RECT 706.320 139.880 713.080 140.200 ;
                RECT 2.880 141.240 98.720 141.560 ;
                RECT 117.440 141.240 290.480 141.560 ;
                RECT 706.320 141.240 713.080 141.560 ;
                RECT 2.880 142.600 98.720 142.920 ;
                RECT 117.440 142.600 290.480 142.920 ;
                RECT 706.320 142.600 713.080 142.920 ;
                RECT 2.880 143.960 98.720 144.280 ;
                RECT 117.440 143.960 120.480 144.280 ;
                RECT 131.040 143.960 285.040 144.280 ;
                RECT 706.320 143.960 713.080 144.280 ;
                RECT 2.880 145.320 98.720 145.640 ;
                RECT 117.440 145.320 121.840 145.640 ;
                RECT 125.600 145.320 285.040 145.640 ;
                RECT 706.320 145.320 713.080 145.640 ;
                RECT 2.880 146.680 98.720 147.000 ;
                RECT 117.440 146.680 123.200 147.000 ;
                RECT 127.640 146.680 135.440 147.000 ;
                RECT 137.840 146.680 279.600 147.000 ;
                RECT 706.320 146.680 713.080 147.000 ;
                RECT 2.880 148.040 98.720 148.360 ;
                RECT 117.440 148.040 279.600 148.360 ;
                RECT 706.320 148.040 713.080 148.360 ;
                RECT 2.880 149.400 98.720 149.720 ;
                RECT 117.440 149.400 129.320 149.720 ;
                RECT 138.520 149.400 279.600 149.720 ;
                RECT 706.320 149.400 713.080 149.720 ;
                RECT 2.880 150.760 98.720 151.080 ;
                RECT 117.440 150.760 122.520 151.080 ;
                RECT 131.040 150.760 301.360 151.080 ;
                RECT 706.320 150.760 713.080 151.080 ;
                RECT 2.880 152.120 98.720 152.440 ;
                RECT 117.440 152.120 125.920 152.440 ;
                RECT 131.040 152.120 301.360 152.440 ;
                RECT 706.320 152.120 713.080 152.440 ;
                RECT 2.880 153.480 98.720 153.800 ;
                RECT 117.440 153.480 301.360 153.800 ;
                RECT 706.320 153.480 713.080 153.800 ;
                RECT 2.880 154.840 98.720 155.160 ;
                RECT 117.440 154.840 119.800 155.160 ;
                RECT 131.040 154.840 301.360 155.160 ;
                RECT 706.320 154.840 713.080 155.160 ;
                RECT 2.880 156.200 98.720 156.520 ;
                RECT 117.440 156.200 129.320 156.520 ;
                RECT 137.160 156.200 301.360 156.520 ;
                RECT 706.320 156.200 713.080 156.520 ;
                RECT 2.880 157.560 98.720 157.880 ;
                RECT 117.440 157.560 128.640 157.880 ;
                RECT 131.040 157.560 301.360 157.880 ;
                RECT 706.320 157.560 713.080 157.880 ;
                RECT 2.880 158.920 98.720 159.240 ;
                RECT 117.440 158.920 301.360 159.240 ;
                RECT 706.320 158.920 713.080 159.240 ;
                RECT 2.880 160.280 98.720 160.600 ;
                RECT 117.440 160.280 129.320 160.600 ;
                RECT 137.840 160.280 301.360 160.600 ;
                RECT 706.320 160.280 713.080 160.600 ;
                RECT 2.880 161.640 98.720 161.960 ;
                RECT 117.440 161.640 126.600 161.960 ;
                RECT 131.040 161.640 301.360 161.960 ;
                RECT 706.320 161.640 713.080 161.960 ;
                RECT 2.880 163.000 98.720 163.320 ;
                RECT 117.440 163.000 128.640 163.320 ;
                RECT 131.040 163.000 301.360 163.320 ;
                RECT 706.320 163.000 713.080 163.320 ;
                RECT 2.880 164.360 98.720 164.680 ;
                RECT 117.440 164.360 132.040 164.680 ;
                RECT 142.600 164.360 301.360 164.680 ;
                RECT 706.320 164.360 713.080 164.680 ;
                RECT 2.880 165.720 98.720 166.040 ;
                RECT 117.440 165.720 119.800 166.040 ;
                RECT 137.840 165.720 301.360 166.040 ;
                RECT 706.320 165.720 713.080 166.040 ;
                RECT 2.880 167.080 98.720 167.400 ;
                RECT 117.440 167.080 128.640 167.400 ;
                RECT 131.040 167.080 138.160 167.400 ;
                RECT 143.960 167.080 301.360 167.400 ;
                RECT 706.320 167.080 713.080 167.400 ;
                RECT 2.880 168.440 98.720 168.760 ;
                RECT 117.440 168.440 140.880 168.760 ;
                RECT 144.640 168.440 301.360 168.760 ;
                RECT 706.320 168.440 713.080 168.760 ;
                RECT 2.880 169.800 98.720 170.120 ;
                RECT 117.440 169.800 120.480 170.120 ;
                RECT 133.760 169.800 301.360 170.120 ;
                RECT 706.320 169.800 713.080 170.120 ;
                RECT 2.880 171.160 98.720 171.480 ;
                RECT 117.440 171.160 129.320 171.480 ;
                RECT 137.840 171.160 301.360 171.480 ;
                RECT 706.320 171.160 713.080 171.480 ;
                RECT 2.880 172.520 98.720 172.840 ;
                RECT 117.440 172.520 126.600 172.840 ;
                RECT 138.520 172.520 301.360 172.840 ;
                RECT 706.320 172.520 713.080 172.840 ;
                RECT 2.880 173.880 98.720 174.200 ;
                RECT 117.440 173.880 301.360 174.200 ;
                RECT 706.320 173.880 713.080 174.200 ;
                RECT 2.880 175.240 98.720 175.560 ;
                RECT 117.440 175.240 122.520 175.560 ;
                RECT 125.600 175.240 301.360 175.560 ;
                RECT 706.320 175.240 713.080 175.560 ;
                RECT 2.880 176.600 98.720 176.920 ;
                RECT 117.440 176.600 122.520 176.920 ;
                RECT 131.040 176.600 301.360 176.920 ;
                RECT 706.320 176.600 713.080 176.920 ;
                RECT 2.880 177.960 98.720 178.280 ;
                RECT 117.440 177.960 125.240 178.280 ;
                RECT 128.320 177.960 301.360 178.280 ;
                RECT 706.320 177.960 713.080 178.280 ;
                RECT 2.880 179.320 98.720 179.640 ;
                RECT 117.440 179.320 301.360 179.640 ;
                RECT 706.320 179.320 713.080 179.640 ;
                RECT 2.880 180.680 98.720 181.000 ;
                RECT 117.440 180.680 128.640 181.000 ;
                RECT 131.040 180.680 301.360 181.000 ;
                RECT 706.320 180.680 713.080 181.000 ;
                RECT 2.880 182.040 98.720 182.360 ;
                RECT 117.440 182.040 121.840 182.360 ;
                RECT 137.160 182.040 301.360 182.360 ;
                RECT 706.320 182.040 713.080 182.360 ;
                RECT 2.880 183.400 98.720 183.720 ;
                RECT 117.440 183.400 128.640 183.720 ;
                RECT 131.040 183.400 301.360 183.720 ;
                RECT 706.320 183.400 713.080 183.720 ;
                RECT 2.880 184.760 98.720 185.080 ;
                RECT 117.440 184.760 301.360 185.080 ;
                RECT 706.320 184.760 713.080 185.080 ;
                RECT 2.880 186.120 98.720 186.440 ;
                RECT 117.440 186.120 123.880 186.440 ;
                RECT 131.040 186.120 301.360 186.440 ;
                RECT 706.320 186.120 713.080 186.440 ;
                RECT 2.880 187.480 98.720 187.800 ;
                RECT 117.440 187.480 120.480 187.800 ;
                RECT 131.720 187.480 301.360 187.800 ;
                RECT 706.320 187.480 713.080 187.800 ;
                RECT 2.880 188.840 98.720 189.160 ;
                RECT 117.440 188.840 143.600 189.160 ;
                RECT 269.080 188.840 301.360 189.160 ;
                RECT 706.320 188.840 713.080 189.160 ;
                RECT 2.880 190.200 98.720 190.520 ;
                RECT 117.440 190.200 119.800 190.520 ;
                RECT 137.840 190.200 195.280 190.520 ;
                RECT 269.080 190.200 301.360 190.520 ;
                RECT 706.320 190.200 713.080 190.520 ;
                RECT 2.880 191.560 98.720 191.880 ;
                RECT 130.360 191.560 195.280 191.880 ;
                RECT 269.080 191.560 301.360 191.880 ;
                RECT 706.320 191.560 713.080 191.880 ;
                RECT 2.880 192.920 98.720 193.240 ;
                RECT 117.440 192.920 120.480 193.240 ;
                RECT 133.760 192.920 195.280 193.240 ;
                RECT 269.080 192.920 301.360 193.240 ;
                RECT 706.320 192.920 713.080 193.240 ;
                RECT 2.880 194.280 98.720 194.600 ;
                RECT 117.440 194.280 135.440 194.600 ;
                RECT 137.840 194.280 301.360 194.600 ;
                RECT 706.320 194.280 713.080 194.600 ;
                RECT 2.880 195.640 98.720 195.960 ;
                RECT 117.440 195.640 301.360 195.960 ;
                RECT 706.320 195.640 713.080 195.960 ;
                RECT 2.880 197.000 98.720 197.320 ;
                RECT 117.440 197.000 132.040 197.320 ;
                RECT 139.880 197.000 301.360 197.320 ;
                RECT 706.320 197.000 713.080 197.320 ;
                RECT 2.880 198.360 98.720 198.680 ;
                RECT 117.440 198.360 282.320 198.680 ;
                RECT 706.320 198.360 713.080 198.680 ;
                RECT 2.880 199.720 98.720 200.040 ;
                RECT 117.440 199.720 202.080 200.040 ;
                RECT 269.760 199.720 282.320 200.040 ;
                RECT 706.320 199.720 713.080 200.040 ;
                RECT 2.880 201.080 98.720 201.400 ;
                RECT 117.440 201.080 122.520 201.400 ;
                RECT 125.600 201.080 202.080 201.400 ;
                RECT 269.760 201.080 287.760 201.400 ;
                RECT 706.320 201.080 713.080 201.400 ;
                RECT 2.880 202.440 98.720 202.760 ;
                RECT 117.440 202.440 119.800 202.760 ;
                RECT 124.240 202.440 202.080 202.760 ;
                RECT 269.760 202.440 287.760 202.760 ;
                RECT 706.320 202.440 713.080 202.760 ;
                RECT 2.880 203.800 98.720 204.120 ;
                RECT 117.440 203.800 202.080 204.120 ;
                RECT 269.760 203.800 287.760 204.120 ;
                RECT 706.320 203.800 713.080 204.120 ;
                RECT 2.880 205.160 98.720 205.480 ;
                RECT 117.440 205.160 125.240 205.480 ;
                RECT 137.840 205.160 202.080 205.480 ;
                RECT 269.760 205.160 293.200 205.480 ;
                RECT 706.320 205.160 713.080 205.480 ;
                RECT 2.880 206.520 98.720 206.840 ;
                RECT 117.440 206.520 202.080 206.840 ;
                RECT 269.760 206.520 293.200 206.840 ;
                RECT 706.320 206.520 713.080 206.840 ;
                RECT 2.880 207.880 98.720 208.200 ;
                RECT 117.440 207.880 202.080 208.200 ;
                RECT 269.760 207.880 298.640 208.200 ;
                RECT 706.320 207.880 713.080 208.200 ;
                RECT 2.880 209.240 98.720 209.560 ;
                RECT 117.440 209.240 202.080 209.560 ;
                RECT 269.760 209.240 298.640 209.560 ;
                RECT 706.320 209.240 713.080 209.560 ;
                RECT 2.880 210.600 98.720 210.920 ;
                RECT 117.440 210.600 122.520 210.920 ;
                RECT 126.960 210.600 202.080 210.920 ;
                RECT 706.320 210.600 713.080 210.920 ;
                RECT 2.880 211.960 98.720 212.280 ;
                RECT 117.440 211.960 202.080 212.280 ;
                RECT 706.320 211.960 713.080 212.280 ;
                RECT 2.880 213.320 98.720 213.640 ;
                RECT 117.440 213.320 135.440 213.640 ;
                RECT 138.520 213.320 202.080 213.640 ;
                RECT 706.320 213.320 713.080 213.640 ;
                RECT 2.880 214.680 98.720 215.000 ;
                RECT 117.440 214.680 202.080 215.000 ;
                RECT 706.320 214.680 713.080 215.000 ;
                RECT 2.880 216.040 98.720 216.360 ;
                RECT 117.440 216.040 202.080 216.360 ;
                RECT 269.760 216.040 301.360 216.360 ;
                RECT 706.320 216.040 713.080 216.360 ;
                RECT 2.880 217.400 98.720 217.720 ;
                RECT 117.440 217.400 121.840 217.720 ;
                RECT 124.920 217.400 202.080 217.720 ;
                RECT 269.760 217.400 301.360 217.720 ;
                RECT 706.320 217.400 713.080 217.720 ;
                RECT 2.880 218.760 98.720 219.080 ;
                RECT 117.440 218.760 202.080 219.080 ;
                RECT 269.760 218.760 301.360 219.080 ;
                RECT 706.320 218.760 713.080 219.080 ;
                RECT 2.880 220.120 98.720 220.440 ;
                RECT 117.440 220.120 202.080 220.440 ;
                RECT 269.760 220.120 301.360 220.440 ;
                RECT 706.320 220.120 713.080 220.440 ;
                RECT 2.880 221.480 98.720 221.800 ;
                RECT 117.440 221.480 202.080 221.800 ;
                RECT 269.760 221.480 301.360 221.800 ;
                RECT 706.320 221.480 713.080 221.800 ;
                RECT 2.880 222.840 98.720 223.160 ;
                RECT 117.440 222.840 128.640 223.160 ;
                RECT 137.160 222.840 202.080 223.160 ;
                RECT 269.760 222.840 301.360 223.160 ;
                RECT 706.320 222.840 713.080 223.160 ;
                RECT 2.880 224.200 98.720 224.520 ;
                RECT 117.440 224.200 202.080 224.520 ;
                RECT 269.760 224.200 301.360 224.520 ;
                RECT 706.320 224.200 713.080 224.520 ;
                RECT 2.880 225.560 98.720 225.880 ;
                RECT 117.440 225.560 125.240 225.880 ;
                RECT 127.640 225.560 202.080 225.880 ;
                RECT 269.760 225.560 301.360 225.880 ;
                RECT 706.320 225.560 713.080 225.880 ;
                RECT 2.880 226.920 98.720 227.240 ;
                RECT 117.440 226.920 202.080 227.240 ;
                RECT 269.760 226.920 301.360 227.240 ;
                RECT 706.320 226.920 713.080 227.240 ;
                RECT 2.880 228.280 98.720 228.600 ;
                RECT 117.440 228.280 202.080 228.600 ;
                RECT 269.760 228.280 301.360 228.600 ;
                RECT 706.320 228.280 713.080 228.600 ;
                RECT 2.880 229.640 98.720 229.960 ;
                RECT 117.440 229.640 202.080 229.960 ;
                RECT 269.760 229.640 301.360 229.960 ;
                RECT 706.320 229.640 713.080 229.960 ;
                RECT 2.880 231.000 98.720 231.320 ;
                RECT 117.440 231.000 202.080 231.320 ;
                RECT 269.760 231.000 301.360 231.320 ;
                RECT 706.320 231.000 713.080 231.320 ;
                RECT 2.880 232.360 98.720 232.680 ;
                RECT 117.440 232.360 202.080 232.680 ;
                RECT 269.760 232.360 301.360 232.680 ;
                RECT 706.320 232.360 713.080 232.680 ;
                RECT 2.880 233.720 202.080 234.040 ;
                RECT 269.760 233.720 301.360 234.040 ;
                RECT 706.320 233.720 713.080 234.040 ;
                RECT 2.880 235.080 202.080 235.400 ;
                RECT 269.760 235.080 301.360 235.400 ;
                RECT 706.320 235.080 713.080 235.400 ;
                RECT 2.880 236.440 79.000 236.760 ;
                RECT 98.400 236.440 123.880 236.760 ;
                RECT 127.640 236.440 202.080 236.760 ;
                RECT 269.760 236.440 301.360 236.760 ;
                RECT 706.320 236.440 713.080 236.760 ;
                RECT 2.880 237.800 79.000 238.120 ;
                RECT 98.400 237.800 202.080 238.120 ;
                RECT 269.760 237.800 301.360 238.120 ;
                RECT 706.320 237.800 713.080 238.120 ;
                RECT 2.880 239.160 79.000 239.480 ;
                RECT 98.400 239.160 202.080 239.480 ;
                RECT 269.760 239.160 301.360 239.480 ;
                RECT 706.320 239.160 713.080 239.480 ;
                RECT 2.880 240.520 79.000 240.840 ;
                RECT 98.400 240.520 104.840 240.840 ;
                RECT 112.000 240.520 125.920 240.840 ;
                RECT 131.720 240.520 202.080 240.840 ;
                RECT 269.760 240.520 301.360 240.840 ;
                RECT 706.320 240.520 713.080 240.840 ;
                RECT 2.880 241.880 79.000 242.200 ;
                RECT 98.400 241.880 99.400 242.200 ;
                RECT 116.760 241.880 202.080 242.200 ;
                RECT 706.320 241.880 713.080 242.200 ;
                RECT 2.880 243.240 79.000 243.560 ;
                RECT 98.400 243.240 99.400 243.560 ;
                RECT 116.760 243.240 202.080 243.560 ;
                RECT 706.320 243.240 713.080 243.560 ;
                RECT 2.880 244.600 79.000 244.920 ;
                RECT 98.400 244.600 202.080 244.920 ;
                RECT 706.320 244.600 713.080 244.920 ;
                RECT 2.880 245.960 79.000 246.280 ;
                RECT 98.400 245.960 104.840 246.280 ;
                RECT 112.000 245.960 120.480 246.280 ;
                RECT 130.360 245.960 202.080 246.280 ;
                RECT 706.320 245.960 713.080 246.280 ;
                RECT 2.880 247.320 73.560 247.640 ;
                RECT 111.320 247.320 202.080 247.640 ;
                RECT 269.760 247.320 713.080 247.640 ;
                RECT 2.880 248.680 110.960 249.000 ;
                RECT 199.040 248.680 713.080 249.000 ;
                RECT 2.880 250.040 298.640 250.360 ;
                RECT 708.360 250.040 713.080 250.360 ;
                RECT 2.880 251.400 298.640 251.720 ;
                RECT 708.360 251.400 713.080 251.720 ;
                RECT 2.880 252.760 298.640 253.080 ;
                RECT 708.360 252.760 713.080 253.080 ;
                RECT 2.880 254.120 28.680 254.440 ;
                RECT 35.160 254.120 37.520 254.440 ;
                RECT 51.480 254.120 106.200 254.440 ;
                RECT 708.360 254.120 713.080 254.440 ;
                RECT 2.880 255.480 26.640 255.800 ;
                RECT 50.800 255.480 62.680 255.800 ;
                RECT 64.400 255.480 77.640 255.800 ;
                RECT 95.680 255.480 106.200 255.800 ;
                RECT 708.360 255.480 713.080 255.800 ;
                RECT 2.880 256.840 26.640 257.160 ;
                RECT 37.200 256.840 62.680 257.160 ;
                RECT 67.120 256.840 77.640 257.160 ;
                RECT 95.680 256.840 106.200 257.160 ;
                RECT 708.360 256.840 713.080 257.160 ;
                RECT 2.880 258.200 26.640 258.520 ;
                RECT 37.200 258.200 62.680 258.520 ;
                RECT 67.120 258.200 77.640 258.520 ;
                RECT 95.680 258.200 106.200 258.520 ;
                RECT 708.360 258.200 713.080 258.520 ;
                RECT 2.880 259.560 26.640 259.880 ;
                RECT 37.200 259.560 62.680 259.880 ;
                RECT 67.800 259.560 77.640 259.880 ;
                RECT 95.680 259.560 106.200 259.880 ;
                RECT 708.360 259.560 713.080 259.880 ;
                RECT 2.880 260.920 26.640 261.240 ;
                RECT 37.200 260.920 62.680 261.240 ;
                RECT 64.400 260.920 77.640 261.240 ;
                RECT 95.680 260.920 106.200 261.240 ;
                RECT 708.360 260.920 713.080 261.240 ;
                RECT 2.880 262.280 26.640 262.600 ;
                RECT 37.200 262.280 106.200 262.600 ;
                RECT 708.360 262.280 713.080 262.600 ;
                RECT 2.880 263.640 26.640 263.960 ;
                RECT 37.200 263.640 77.640 263.960 ;
                RECT 95.680 263.640 106.200 263.960 ;
                RECT 708.360 263.640 713.080 263.960 ;
                RECT 2.880 265.000 77.640 265.320 ;
                RECT 95.680 265.000 106.200 265.320 ;
                RECT 708.360 265.000 713.080 265.320 ;
                RECT 2.880 266.360 77.640 266.680 ;
                RECT 95.680 266.360 106.200 266.680 ;
                RECT 708.360 266.360 713.080 266.680 ;
                RECT 2.880 267.720 19.840 268.040 ;
                RECT 22.240 267.720 77.640 268.040 ;
                RECT 95.680 267.720 106.200 268.040 ;
                RECT 708.360 267.720 713.080 268.040 ;
                RECT 2.880 269.080 77.640 269.400 ;
                RECT 95.680 269.080 106.200 269.400 ;
                RECT 708.360 269.080 713.080 269.400 ;
                RECT 2.880 270.440 19.160 270.760 ;
                RECT 22.240 270.440 35.480 270.760 ;
                RECT 50.800 270.440 106.200 270.760 ;
                RECT 708.360 270.440 713.080 270.760 ;
                RECT 2.880 271.800 18.480 272.120 ;
                RECT 22.240 271.800 35.480 272.120 ;
                RECT 50.120 271.800 62.680 272.120 ;
                RECT 64.400 271.800 77.640 272.120 ;
                RECT 95.680 271.800 106.200 272.120 ;
                RECT 708.360 271.800 713.080 272.120 ;
                RECT 2.880 273.160 17.800 273.480 ;
                RECT 22.240 273.160 35.480 273.480 ;
                RECT 40.600 273.160 62.680 273.480 ;
                RECT 65.080 273.160 77.640 273.480 ;
                RECT 95.680 273.160 106.200 273.480 ;
                RECT 708.360 273.160 713.080 273.480 ;
                RECT 2.880 274.520 62.680 274.840 ;
                RECT 65.760 274.520 77.640 274.840 ;
                RECT 95.680 274.520 106.200 274.840 ;
                RECT 708.360 274.520 713.080 274.840 ;
                RECT 2.880 275.880 17.120 276.200 ;
                RECT 22.240 275.880 35.480 276.200 ;
                RECT 41.280 275.880 62.680 276.200 ;
                RECT 65.760 275.880 77.640 276.200 ;
                RECT 95.680 275.880 106.200 276.200 ;
                RECT 708.360 275.880 713.080 276.200 ;
                RECT 2.880 277.240 16.440 277.560 ;
                RECT 22.240 277.240 35.480 277.560 ;
                RECT 41.960 277.240 62.680 277.560 ;
                RECT 66.440 277.240 77.640 277.560 ;
                RECT 95.680 277.240 106.200 277.560 ;
                RECT 708.360 277.240 713.080 277.560 ;
                RECT 2.880 278.600 15.760 278.920 ;
                RECT 22.240 278.600 106.200 278.920 ;
                RECT 708.360 278.600 713.080 278.920 ;
                RECT 2.880 279.960 15.080 280.280 ;
                RECT 22.240 279.960 77.640 280.280 ;
                RECT 95.680 279.960 106.200 280.280 ;
                RECT 708.360 279.960 713.080 280.280 ;
                RECT 2.880 281.320 77.640 281.640 ;
                RECT 95.680 281.320 106.200 281.640 ;
                RECT 708.360 281.320 713.080 281.640 ;
                RECT 2.880 282.680 14.400 283.000 ;
                RECT 22.240 282.680 77.640 283.000 ;
                RECT 95.680 282.680 106.200 283.000 ;
                RECT 708.360 282.680 713.080 283.000 ;
                RECT 2.880 284.040 13.720 284.360 ;
                RECT 22.240 284.040 77.640 284.360 ;
                RECT 95.680 284.040 106.200 284.360 ;
                RECT 708.360 284.040 713.080 284.360 ;
                RECT 2.880 285.400 77.640 285.720 ;
                RECT 90.240 285.400 106.200 285.720 ;
                RECT 708.360 285.400 713.080 285.720 ;
                RECT 2.880 286.760 13.040 287.080 ;
                RECT 22.240 286.760 35.480 287.080 ;
                RECT 41.960 286.760 85.800 287.080 ;
                RECT 95.680 286.760 106.200 287.080 ;
                RECT 708.360 286.760 713.080 287.080 ;
                RECT 2.880 288.120 12.360 288.440 ;
                RECT 22.240 288.120 35.480 288.440 ;
                RECT 41.280 288.120 77.640 288.440 ;
                RECT 95.680 288.120 106.200 288.440 ;
                RECT 708.360 288.120 713.080 288.440 ;
                RECT 2.880 289.480 77.640 289.800 ;
                RECT 95.680 289.480 106.200 289.800 ;
                RECT 708.360 289.480 713.080 289.800 ;
                RECT 2.880 290.840 11.680 291.160 ;
                RECT 22.240 290.840 35.480 291.160 ;
                RECT 40.600 290.840 77.640 291.160 ;
                RECT 95.680 290.840 106.200 291.160 ;
                RECT 708.360 290.840 713.080 291.160 ;
                RECT 2.880 292.200 11.000 292.520 ;
                RECT 22.240 292.200 35.480 292.520 ;
                RECT 39.920 292.200 77.640 292.520 ;
                RECT 95.680 292.200 106.200 292.520 ;
                RECT 708.360 292.200 713.080 292.520 ;
                RECT 2.880 293.560 10.320 293.880 ;
                RECT 22.240 293.560 35.480 293.880 ;
                RECT 39.240 293.560 77.640 293.880 ;
                RECT 90.240 293.560 106.200 293.880 ;
                RECT 708.360 293.560 713.080 293.880 ;
                RECT 2.880 294.920 9.640 295.240 ;
                RECT 22.240 294.920 77.640 295.240 ;
                RECT 95.680 294.920 106.200 295.240 ;
                RECT 708.360 294.920 713.080 295.240 ;
                RECT 2.880 296.280 77.640 296.600 ;
                RECT 95.680 296.280 106.200 296.600 ;
                RECT 708.360 296.280 713.080 296.600 ;
                RECT 2.880 297.640 77.640 297.960 ;
                RECT 95.680 297.640 106.200 297.960 ;
                RECT 708.360 297.640 713.080 297.960 ;
                RECT 2.880 299.000 77.640 299.320 ;
                RECT 95.680 299.000 106.200 299.320 ;
                RECT 708.360 299.000 713.080 299.320 ;
                RECT 2.880 300.360 77.640 300.680 ;
                RECT 95.680 300.360 106.200 300.680 ;
                RECT 708.360 300.360 713.080 300.680 ;
                RECT 2.880 301.720 77.640 302.040 ;
                RECT 90.920 301.720 106.200 302.040 ;
                RECT 708.360 301.720 713.080 302.040 ;
                RECT 2.880 303.080 77.640 303.400 ;
                RECT 95.680 303.080 106.200 303.400 ;
                RECT 708.360 303.080 713.080 303.400 ;
                RECT 2.880 304.440 77.640 304.760 ;
                RECT 95.680 304.440 106.200 304.760 ;
                RECT 708.360 304.440 713.080 304.760 ;
                RECT 2.880 305.800 77.640 306.120 ;
                RECT 95.680 305.800 106.200 306.120 ;
                RECT 708.360 305.800 713.080 306.120 ;
                RECT 2.880 307.160 77.640 307.480 ;
                RECT 95.680 307.160 106.200 307.480 ;
                RECT 708.360 307.160 713.080 307.480 ;
                RECT 2.880 308.520 77.640 308.840 ;
                RECT 95.680 308.520 106.200 308.840 ;
                RECT 708.360 308.520 713.080 308.840 ;
                RECT 2.880 309.880 106.200 310.200 ;
                RECT 708.360 309.880 713.080 310.200 ;
                RECT 2.880 311.240 77.640 311.560 ;
                RECT 95.680 311.240 106.200 311.560 ;
                RECT 708.360 311.240 713.080 311.560 ;
                RECT 2.880 312.600 77.640 312.920 ;
                RECT 95.680 312.600 106.200 312.920 ;
                RECT 708.360 312.600 713.080 312.920 ;
                RECT 2.880 313.960 77.640 314.280 ;
                RECT 95.680 313.960 106.200 314.280 ;
                RECT 708.360 313.960 713.080 314.280 ;
                RECT 2.880 315.320 77.640 315.640 ;
                RECT 95.680 315.320 106.200 315.640 ;
                RECT 708.360 315.320 713.080 315.640 ;
                RECT 2.880 316.680 77.640 317.000 ;
                RECT 95.680 316.680 106.200 317.000 ;
                RECT 708.360 316.680 713.080 317.000 ;
                RECT 2.880 318.040 106.200 318.360 ;
                RECT 708.360 318.040 713.080 318.360 ;
                RECT 2.880 319.400 77.640 319.720 ;
                RECT 95.680 319.400 106.200 319.720 ;
                RECT 708.360 319.400 713.080 319.720 ;
                RECT 2.880 320.760 77.640 321.080 ;
                RECT 95.680 320.760 106.200 321.080 ;
                RECT 708.360 320.760 713.080 321.080 ;
                RECT 2.880 322.120 77.640 322.440 ;
                RECT 95.680 322.120 106.200 322.440 ;
                RECT 708.360 322.120 713.080 322.440 ;
                RECT 2.880 323.480 77.640 323.800 ;
                RECT 95.680 323.480 106.200 323.800 ;
                RECT 708.360 323.480 713.080 323.800 ;
                RECT 2.880 324.840 77.640 325.160 ;
                RECT 95.680 324.840 106.200 325.160 ;
                RECT 708.360 324.840 713.080 325.160 ;
                RECT 2.880 326.200 106.200 326.520 ;
                RECT 708.360 326.200 713.080 326.520 ;
                RECT 2.880 327.560 77.640 327.880 ;
                RECT 95.680 327.560 106.200 327.880 ;
                RECT 708.360 327.560 713.080 327.880 ;
                RECT 2.880 328.920 77.640 329.240 ;
                RECT 95.680 328.920 106.200 329.240 ;
                RECT 708.360 328.920 713.080 329.240 ;
                RECT 2.880 330.280 77.640 330.600 ;
                RECT 95.680 330.280 106.200 330.600 ;
                RECT 708.360 330.280 713.080 330.600 ;
                RECT 2.880 331.640 77.640 331.960 ;
                RECT 95.680 331.640 106.200 331.960 ;
                RECT 708.360 331.640 713.080 331.960 ;
                RECT 2.880 333.000 77.640 333.320 ;
                RECT 93.640 333.000 106.200 333.320 ;
                RECT 708.360 333.000 713.080 333.320 ;
                RECT 2.880 334.360 89.880 334.680 ;
                RECT 95.680 334.360 106.200 334.680 ;
                RECT 708.360 334.360 713.080 334.680 ;
                RECT 2.880 335.720 77.640 336.040 ;
                RECT 95.680 335.720 106.200 336.040 ;
                RECT 708.360 335.720 713.080 336.040 ;
                RECT 2.880 337.080 77.640 337.400 ;
                RECT 95.680 337.080 106.200 337.400 ;
                RECT 708.360 337.080 713.080 337.400 ;
                RECT 2.880 338.440 77.640 338.760 ;
                RECT 95.680 338.440 106.200 338.760 ;
                RECT 708.360 338.440 713.080 338.760 ;
                RECT 2.880 339.800 77.640 340.120 ;
                RECT 95.680 339.800 106.200 340.120 ;
                RECT 708.360 339.800 713.080 340.120 ;
                RECT 2.880 341.160 77.640 341.480 ;
                RECT 94.320 341.160 106.200 341.480 ;
                RECT 708.360 341.160 713.080 341.480 ;
                RECT 2.880 342.520 77.640 342.840 ;
                RECT 95.680 342.520 106.200 342.840 ;
                RECT 708.360 342.520 713.080 342.840 ;
                RECT 2.880 343.880 77.640 344.200 ;
                RECT 95.680 343.880 106.200 344.200 ;
                RECT 708.360 343.880 713.080 344.200 ;
                RECT 2.880 345.240 77.640 345.560 ;
                RECT 95.680 345.240 106.200 345.560 ;
                RECT 708.360 345.240 713.080 345.560 ;
                RECT 2.880 346.600 77.640 346.920 ;
                RECT 95.680 346.600 106.200 346.920 ;
                RECT 708.360 346.600 713.080 346.920 ;
                RECT 2.880 347.960 77.640 348.280 ;
                RECT 95.680 347.960 106.200 348.280 ;
                RECT 708.360 347.960 713.080 348.280 ;
                RECT 2.880 349.320 106.200 349.640 ;
                RECT 708.360 349.320 713.080 349.640 ;
                RECT 2.880 350.680 79.680 351.000 ;
                RECT 95.680 350.680 106.200 351.000 ;
                RECT 708.360 350.680 713.080 351.000 ;
                RECT 2.880 352.040 79.680 352.360 ;
                RECT 95.680 352.040 106.200 352.360 ;
                RECT 708.360 352.040 713.080 352.360 ;
                RECT 2.880 353.400 87.160 353.720 ;
                RECT 95.680 353.400 106.200 353.720 ;
                RECT 708.360 353.400 713.080 353.720 ;
                RECT 2.880 354.760 79.680 355.080 ;
                RECT 95.680 354.760 106.200 355.080 ;
                RECT 708.360 354.760 713.080 355.080 ;
                RECT 2.880 356.120 79.680 356.440 ;
                RECT 95.680 356.120 106.200 356.440 ;
                RECT 708.360 356.120 713.080 356.440 ;
                RECT 2.880 357.480 41.600 357.800 ;
                RECT 50.800 357.480 106.200 357.800 ;
                RECT 708.360 357.480 713.080 357.800 ;
                RECT 2.880 358.840 40.240 359.160 ;
                RECT 50.120 358.840 62.680 359.160 ;
                RECT 64.400 358.840 77.640 359.160 ;
                RECT 95.680 358.840 106.200 359.160 ;
                RECT 708.360 358.840 713.080 359.160 ;
                RECT 2.880 360.200 62.680 360.520 ;
                RECT 67.120 360.200 77.640 360.520 ;
                RECT 95.680 360.200 106.200 360.520 ;
                RECT 708.360 360.200 713.080 360.520 ;
                RECT 2.880 361.560 62.680 361.880 ;
                RECT 67.120 361.560 77.640 361.880 ;
                RECT 95.680 361.560 106.200 361.880 ;
                RECT 708.360 361.560 713.080 361.880 ;
                RECT 2.880 362.920 62.680 363.240 ;
                RECT 67.800 362.920 77.640 363.240 ;
                RECT 95.680 362.920 106.200 363.240 ;
                RECT 708.360 362.920 713.080 363.240 ;
                RECT 2.880 364.280 62.680 364.600 ;
                RECT 68.480 364.280 77.640 364.600 ;
                RECT 95.680 364.280 106.200 364.600 ;
                RECT 708.360 364.280 713.080 364.600 ;
                RECT 2.880 365.640 106.200 365.960 ;
                RECT 708.360 365.640 713.080 365.960 ;
                RECT 2.880 367.000 77.640 367.320 ;
                RECT 95.680 367.000 106.200 367.320 ;
                RECT 708.360 367.000 713.080 367.320 ;
                RECT 2.880 368.360 77.640 368.680 ;
                RECT 95.680 368.360 106.200 368.680 ;
                RECT 708.360 368.360 713.080 368.680 ;
                RECT 2.880 369.720 77.640 370.040 ;
                RECT 95.680 369.720 106.200 370.040 ;
                RECT 708.360 369.720 713.080 370.040 ;
                RECT 2.880 371.080 77.640 371.400 ;
                RECT 95.680 371.080 106.200 371.400 ;
                RECT 708.360 371.080 713.080 371.400 ;
                RECT 2.880 372.440 39.560 372.760 ;
                RECT 51.480 372.440 77.640 372.760 ;
                RECT 80.720 372.440 106.200 372.760 ;
                RECT 708.360 372.440 713.080 372.760 ;
                RECT 2.880 373.800 38.200 374.120 ;
                RECT 50.800 373.800 91.920 374.120 ;
                RECT 95.680 373.800 106.200 374.120 ;
                RECT 708.360 373.800 713.080 374.120 ;
                RECT 2.880 375.160 62.680 375.480 ;
                RECT 65.080 375.160 77.640 375.480 ;
                RECT 95.680 375.160 106.200 375.480 ;
                RECT 708.360 375.160 713.080 375.480 ;
                RECT 2.880 376.520 62.680 376.840 ;
                RECT 65.760 376.520 77.640 376.840 ;
                RECT 95.680 376.520 106.200 376.840 ;
                RECT 708.360 376.520 713.080 376.840 ;
                RECT 2.880 377.880 62.680 378.200 ;
                RECT 65.760 377.880 77.640 378.200 ;
                RECT 95.680 377.880 106.200 378.200 ;
                RECT 708.360 377.880 713.080 378.200 ;
                RECT 2.880 379.240 62.680 379.560 ;
                RECT 64.400 379.240 77.640 379.560 ;
                RECT 95.680 379.240 106.200 379.560 ;
                RECT 708.360 379.240 713.080 379.560 ;
                RECT 2.880 380.600 62.680 380.920 ;
                RECT 66.440 380.600 77.640 380.920 ;
                RECT 81.400 380.600 106.200 380.920 ;
                RECT 708.360 380.600 713.080 380.920 ;
                RECT 2.880 381.960 77.640 382.280 ;
                RECT 95.680 381.960 106.200 382.280 ;
                RECT 708.360 381.960 713.080 382.280 ;
                RECT 2.880 383.320 77.640 383.640 ;
                RECT 95.680 383.320 106.200 383.640 ;
                RECT 708.360 383.320 713.080 383.640 ;
                RECT 2.880 384.680 77.640 385.000 ;
                RECT 95.680 384.680 106.200 385.000 ;
                RECT 708.360 384.680 713.080 385.000 ;
                RECT 2.880 386.040 77.640 386.360 ;
                RECT 95.680 386.040 106.200 386.360 ;
                RECT 708.360 386.040 713.080 386.360 ;
                RECT 2.880 387.400 77.640 387.720 ;
                RECT 95.680 387.400 106.200 387.720 ;
                RECT 708.360 387.400 713.080 387.720 ;
                RECT 2.880 388.760 106.200 389.080 ;
                RECT 708.360 388.760 713.080 389.080 ;
                RECT 2.880 390.120 77.640 390.440 ;
                RECT 95.680 390.120 106.200 390.440 ;
                RECT 708.360 390.120 713.080 390.440 ;
                RECT 2.880 391.480 77.640 391.800 ;
                RECT 95.680 391.480 106.200 391.800 ;
                RECT 708.360 391.480 713.080 391.800 ;
                RECT 2.880 392.840 77.640 393.160 ;
                RECT 95.680 392.840 106.200 393.160 ;
                RECT 708.360 392.840 713.080 393.160 ;
                RECT 2.880 394.200 77.640 394.520 ;
                RECT 95.680 394.200 106.200 394.520 ;
                RECT 708.360 394.200 713.080 394.520 ;
                RECT 2.880 395.560 77.640 395.880 ;
                RECT 95.680 395.560 106.200 395.880 ;
                RECT 708.360 395.560 713.080 395.880 ;
                RECT 2.880 396.920 106.200 397.240 ;
                RECT 708.360 396.920 713.080 397.240 ;
                RECT 2.880 398.280 77.640 398.600 ;
                RECT 95.680 398.280 106.200 398.600 ;
                RECT 708.360 398.280 713.080 398.600 ;
                RECT 2.880 399.640 77.640 399.960 ;
                RECT 95.680 399.640 106.200 399.960 ;
                RECT 708.360 399.640 713.080 399.960 ;
                RECT 2.880 401.000 77.640 401.320 ;
                RECT 95.680 401.000 106.200 401.320 ;
                RECT 708.360 401.000 713.080 401.320 ;
                RECT 2.880 402.360 77.640 402.680 ;
                RECT 95.680 402.360 106.200 402.680 ;
                RECT 708.360 402.360 713.080 402.680 ;
                RECT 2.880 403.720 77.640 404.040 ;
                RECT 95.680 403.720 106.200 404.040 ;
                RECT 708.360 403.720 713.080 404.040 ;
                RECT 2.880 405.080 106.200 405.400 ;
                RECT 708.360 405.080 713.080 405.400 ;
                RECT 2.880 406.440 77.640 406.760 ;
                RECT 95.680 406.440 106.200 406.760 ;
                RECT 708.360 406.440 713.080 406.760 ;
                RECT 2.880 407.800 77.640 408.120 ;
                RECT 95.680 407.800 106.200 408.120 ;
                RECT 708.360 407.800 713.080 408.120 ;
                RECT 2.880 409.160 77.640 409.480 ;
                RECT 95.680 409.160 106.200 409.480 ;
                RECT 708.360 409.160 713.080 409.480 ;
                RECT 2.880 410.520 77.640 410.840 ;
                RECT 95.680 410.520 106.200 410.840 ;
                RECT 708.360 410.520 713.080 410.840 ;
                RECT 2.880 411.880 77.640 412.200 ;
                RECT 84.120 411.880 106.200 412.200 ;
                RECT 708.360 411.880 713.080 412.200 ;
                RECT 2.880 413.240 85.800 413.560 ;
                RECT 95.680 413.240 106.200 413.560 ;
                RECT 708.360 413.240 713.080 413.560 ;
                RECT 2.880 414.600 77.640 414.920 ;
                RECT 95.680 414.600 106.200 414.920 ;
                RECT 708.360 414.600 713.080 414.920 ;
                RECT 2.880 415.960 77.640 416.280 ;
                RECT 95.680 415.960 106.200 416.280 ;
                RECT 708.360 415.960 713.080 416.280 ;
                RECT 2.880 417.320 77.640 417.640 ;
                RECT 95.680 417.320 106.200 417.640 ;
                RECT 708.360 417.320 713.080 417.640 ;
                RECT 2.880 418.680 77.640 419.000 ;
                RECT 95.680 418.680 106.200 419.000 ;
                RECT 708.360 418.680 713.080 419.000 ;
                RECT 2.880 420.040 77.640 420.360 ;
                RECT 84.800 420.040 106.200 420.360 ;
                RECT 708.360 420.040 713.080 420.360 ;
                RECT 2.880 421.400 77.640 421.720 ;
                RECT 95.680 421.400 106.200 421.720 ;
                RECT 708.360 421.400 713.080 421.720 ;
                RECT 2.880 422.760 77.640 423.080 ;
                RECT 95.680 422.760 106.200 423.080 ;
                RECT 708.360 422.760 713.080 423.080 ;
                RECT 2.880 424.120 77.640 424.440 ;
                RECT 95.680 424.120 106.200 424.440 ;
                RECT 708.360 424.120 713.080 424.440 ;
                RECT 2.880 425.480 77.640 425.800 ;
                RECT 95.680 425.480 106.200 425.800 ;
                RECT 708.360 425.480 713.080 425.800 ;
                RECT 2.880 426.840 77.640 427.160 ;
                RECT 95.680 426.840 106.200 427.160 ;
                RECT 708.360 426.840 713.080 427.160 ;
                RECT 2.880 428.200 106.200 428.520 ;
                RECT 708.360 428.200 713.080 428.520 ;
                RECT 2.880 429.560 77.640 429.880 ;
                RECT 95.680 429.560 106.200 429.880 ;
                RECT 708.360 429.560 713.080 429.880 ;
                RECT 2.880 430.920 77.640 431.240 ;
                RECT 95.680 430.920 106.200 431.240 ;
                RECT 708.360 430.920 713.080 431.240 ;
                RECT 2.880 432.280 77.640 432.600 ;
                RECT 95.680 432.280 106.200 432.600 ;
                RECT 708.360 432.280 713.080 432.600 ;
                RECT 2.880 433.640 77.640 433.960 ;
                RECT 95.680 433.640 106.200 433.960 ;
                RECT 708.360 433.640 713.080 433.960 ;
                RECT 2.880 435.000 77.640 435.320 ;
                RECT 95.680 435.000 106.200 435.320 ;
                RECT 708.360 435.000 713.080 435.320 ;
                RECT 2.880 436.360 106.200 436.680 ;
                RECT 708.360 436.360 713.080 436.680 ;
                RECT 2.880 437.720 77.640 438.040 ;
                RECT 95.680 437.720 106.200 438.040 ;
                RECT 708.360 437.720 713.080 438.040 ;
                RECT 2.880 439.080 77.640 439.400 ;
                RECT 95.680 439.080 106.200 439.400 ;
                RECT 708.360 439.080 713.080 439.400 ;
                RECT 2.880 440.440 77.640 440.760 ;
                RECT 95.680 440.440 106.200 440.760 ;
                RECT 708.360 440.440 713.080 440.760 ;
                RECT 2.880 441.800 77.640 442.120 ;
                RECT 95.680 441.800 106.200 442.120 ;
                RECT 708.360 441.800 713.080 442.120 ;
                RECT 2.880 443.160 77.640 443.480 ;
                RECT 95.680 443.160 106.200 443.480 ;
                RECT 708.360 443.160 713.080 443.480 ;
                RECT 2.880 444.520 106.200 444.840 ;
                RECT 708.360 444.520 713.080 444.840 ;
                RECT 2.880 445.880 77.640 446.200 ;
                RECT 95.680 445.880 106.200 446.200 ;
                RECT 708.360 445.880 713.080 446.200 ;
                RECT 2.880 447.240 77.640 447.560 ;
                RECT 95.680 447.240 106.200 447.560 ;
                RECT 708.360 447.240 713.080 447.560 ;
                RECT 2.880 448.600 77.640 448.920 ;
                RECT 95.680 448.600 106.200 448.920 ;
                RECT 708.360 448.600 713.080 448.920 ;
                RECT 2.880 449.960 77.640 450.280 ;
                RECT 95.680 449.960 106.200 450.280 ;
                RECT 708.360 449.960 713.080 450.280 ;
                RECT 2.880 451.320 77.640 451.640 ;
                RECT 86.840 451.320 106.200 451.640 ;
                RECT 708.360 451.320 713.080 451.640 ;
                RECT 2.880 452.680 87.840 453.000 ;
                RECT 95.680 452.680 106.200 453.000 ;
                RECT 708.360 452.680 713.080 453.000 ;
                RECT 2.880 454.040 81.040 454.360 ;
                RECT 95.680 454.040 106.200 454.360 ;
                RECT 708.360 454.040 713.080 454.360 ;
                RECT 2.880 455.400 81.040 455.720 ;
                RECT 95.680 455.400 106.200 455.720 ;
                RECT 708.360 455.400 713.080 455.720 ;
                RECT 2.880 456.760 81.040 457.080 ;
                RECT 95.680 456.760 106.200 457.080 ;
                RECT 708.360 456.760 713.080 457.080 ;
                RECT 2.880 458.120 81.040 458.440 ;
                RECT 95.680 458.120 106.200 458.440 ;
                RECT 708.360 458.120 713.080 458.440 ;
                RECT 2.880 459.480 106.200 459.800 ;
                RECT 708.360 459.480 713.080 459.800 ;
                RECT 2.880 460.840 89.880 461.160 ;
                RECT 95.680 460.840 106.200 461.160 ;
                RECT 708.360 460.840 713.080 461.160 ;
                RECT 2.880 462.200 81.040 462.520 ;
                RECT 95.680 462.200 106.200 462.520 ;
                RECT 708.360 462.200 713.080 462.520 ;
                RECT 2.880 463.560 81.040 463.880 ;
                RECT 95.680 463.560 106.200 463.880 ;
                RECT 708.360 463.560 713.080 463.880 ;
                RECT 2.880 464.920 81.040 465.240 ;
                RECT 95.680 464.920 106.200 465.240 ;
                RECT 708.360 464.920 713.080 465.240 ;
                RECT 2.880 466.280 81.040 466.600 ;
                RECT 95.680 466.280 106.200 466.600 ;
                RECT 708.360 466.280 713.080 466.600 ;
                RECT 2.880 467.640 106.200 467.960 ;
                RECT 708.360 467.640 713.080 467.960 ;
                RECT 2.880 469.000 81.040 469.320 ;
                RECT 95.680 469.000 106.200 469.320 ;
                RECT 708.360 469.000 713.080 469.320 ;
                RECT 2.880 470.360 91.920 470.680 ;
                RECT 95.680 470.360 106.200 470.680 ;
                RECT 708.360 470.360 713.080 470.680 ;
                RECT 2.880 471.720 81.040 472.040 ;
                RECT 95.680 471.720 106.200 472.040 ;
                RECT 708.360 471.720 713.080 472.040 ;
                RECT 2.880 473.080 81.040 473.400 ;
                RECT 95.680 473.080 106.200 473.400 ;
                RECT 708.360 473.080 713.080 473.400 ;
                RECT 2.880 474.440 81.040 474.760 ;
                RECT 95.680 474.440 106.200 474.760 ;
                RECT 708.360 474.440 713.080 474.760 ;
                RECT 2.880 475.800 106.200 476.120 ;
                RECT 708.360 475.800 713.080 476.120 ;
                RECT 2.880 477.160 81.720 477.480 ;
                RECT 95.680 477.160 106.200 477.480 ;
                RECT 708.360 477.160 713.080 477.480 ;
                RECT 2.880 478.520 81.720 478.840 ;
                RECT 95.680 478.520 106.200 478.840 ;
                RECT 708.360 478.520 713.080 478.840 ;
                RECT 2.880 479.880 87.160 480.200 ;
                RECT 95.680 479.880 106.200 480.200 ;
                RECT 708.360 479.880 713.080 480.200 ;
                RECT 2.880 481.240 81.720 481.560 ;
                RECT 95.680 481.240 106.200 481.560 ;
                RECT 708.360 481.240 713.080 481.560 ;
                RECT 2.880 482.600 81.720 482.920 ;
                RECT 95.680 482.600 106.200 482.920 ;
                RECT 708.360 482.600 713.080 482.920 ;
                RECT 2.880 483.960 106.200 484.280 ;
                RECT 708.360 483.960 713.080 484.280 ;
                RECT 2.880 485.320 81.720 485.640 ;
                RECT 95.680 485.320 106.200 485.640 ;
                RECT 708.360 485.320 713.080 485.640 ;
                RECT 2.880 486.680 81.720 487.000 ;
                RECT 95.680 486.680 106.200 487.000 ;
                RECT 708.360 486.680 713.080 487.000 ;
                RECT 2.880 488.040 81.720 488.360 ;
                RECT 95.680 488.040 106.200 488.360 ;
                RECT 708.360 488.040 713.080 488.360 ;
                RECT 2.880 489.400 89.200 489.720 ;
                RECT 95.680 489.400 106.200 489.720 ;
                RECT 708.360 489.400 713.080 489.720 ;
                RECT 2.880 490.760 81.720 491.080 ;
                RECT 95.680 490.760 106.200 491.080 ;
                RECT 708.360 490.760 713.080 491.080 ;
                RECT 2.880 492.120 106.200 492.440 ;
                RECT 708.360 492.120 713.080 492.440 ;
                RECT 2.880 493.480 81.720 493.800 ;
                RECT 95.680 493.480 106.200 493.800 ;
                RECT 708.360 493.480 713.080 493.800 ;
                RECT 2.880 494.840 81.720 495.160 ;
                RECT 95.680 494.840 106.200 495.160 ;
                RECT 708.360 494.840 713.080 495.160 ;
                RECT 2.880 496.200 81.720 496.520 ;
                RECT 95.680 496.200 106.200 496.520 ;
                RECT 708.360 496.200 713.080 496.520 ;
                RECT 2.880 497.560 81.720 497.880 ;
                RECT 95.680 497.560 106.200 497.880 ;
                RECT 708.360 497.560 713.080 497.880 ;
                RECT 2.880 498.920 106.200 499.240 ;
                RECT 708.360 498.920 713.080 499.240 ;
                RECT 2.880 500.280 91.920 500.600 ;
                RECT 95.680 500.280 106.200 500.600 ;
                RECT 708.360 500.280 713.080 500.600 ;
                RECT 2.880 501.640 81.720 501.960 ;
                RECT 95.680 501.640 106.200 501.960 ;
                RECT 708.360 501.640 713.080 501.960 ;
                RECT 2.880 503.000 81.720 503.320 ;
                RECT 95.680 503.000 106.200 503.320 ;
                RECT 708.360 503.000 713.080 503.320 ;
                RECT 2.880 504.360 81.720 504.680 ;
                RECT 95.680 504.360 106.200 504.680 ;
                RECT 708.360 504.360 713.080 504.680 ;
                RECT 2.880 505.720 81.720 506.040 ;
                RECT 95.680 505.720 106.200 506.040 ;
                RECT 708.360 505.720 713.080 506.040 ;
                RECT 2.880 507.080 106.200 507.400 ;
                RECT 708.360 507.080 713.080 507.400 ;
                RECT 2.880 508.440 82.400 508.760 ;
                RECT 95.680 508.440 106.200 508.760 ;
                RECT 708.360 508.440 713.080 508.760 ;
                RECT 2.880 509.800 86.480 510.120 ;
                RECT 95.680 509.800 106.200 510.120 ;
                RECT 708.360 509.800 713.080 510.120 ;
                RECT 2.880 511.160 82.400 511.480 ;
                RECT 95.680 511.160 106.200 511.480 ;
                RECT 708.360 511.160 713.080 511.480 ;
                RECT 2.880 512.520 82.400 512.840 ;
                RECT 95.680 512.520 106.200 512.840 ;
                RECT 708.360 512.520 713.080 512.840 ;
                RECT 2.880 513.880 82.400 514.200 ;
                RECT 95.680 513.880 106.200 514.200 ;
                RECT 708.360 513.880 713.080 514.200 ;
                RECT 2.880 515.240 106.200 515.560 ;
                RECT 708.360 515.240 713.080 515.560 ;
                RECT 2.880 516.600 82.400 516.920 ;
                RECT 95.680 516.600 106.200 516.920 ;
                RECT 708.360 516.600 713.080 516.920 ;
                RECT 2.880 517.960 82.400 518.280 ;
                RECT 95.680 517.960 106.200 518.280 ;
                RECT 708.360 517.960 713.080 518.280 ;
                RECT 2.880 519.320 88.520 519.640 ;
                RECT 95.680 519.320 106.200 519.640 ;
                RECT 708.360 519.320 713.080 519.640 ;
                RECT 2.880 520.680 82.400 521.000 ;
                RECT 95.680 520.680 106.200 521.000 ;
                RECT 708.360 520.680 713.080 521.000 ;
                RECT 2.880 522.040 82.400 522.360 ;
                RECT 95.680 522.040 106.200 522.360 ;
                RECT 708.360 522.040 713.080 522.360 ;
                RECT 2.880 523.400 106.200 523.720 ;
                RECT 708.360 523.400 713.080 523.720 ;
                RECT 2.880 524.760 82.400 525.080 ;
                RECT 95.680 524.760 106.200 525.080 ;
                RECT 708.360 524.760 713.080 525.080 ;
                RECT 2.880 526.120 82.400 526.440 ;
                RECT 95.680 526.120 106.200 526.440 ;
                RECT 708.360 526.120 713.080 526.440 ;
                RECT 2.880 527.480 82.400 527.800 ;
                RECT 95.680 527.480 106.200 527.800 ;
                RECT 708.360 527.480 713.080 527.800 ;
                RECT 2.880 528.840 91.240 529.160 ;
                RECT 95.680 528.840 106.200 529.160 ;
                RECT 708.360 528.840 713.080 529.160 ;
                RECT 2.880 530.200 82.400 530.520 ;
                RECT 95.680 530.200 106.200 530.520 ;
                RECT 708.360 530.200 713.080 530.520 ;
                RECT 2.880 531.560 106.200 531.880 ;
                RECT 708.360 531.560 713.080 531.880 ;
                RECT 2.880 532.920 82.400 533.240 ;
                RECT 95.680 532.920 106.200 533.240 ;
                RECT 708.360 532.920 713.080 533.240 ;
                RECT 2.880 534.280 82.400 534.600 ;
                RECT 95.680 534.280 106.200 534.600 ;
                RECT 708.360 534.280 713.080 534.600 ;
                RECT 2.880 535.640 82.400 535.960 ;
                RECT 95.680 535.640 106.200 535.960 ;
                RECT 708.360 535.640 713.080 535.960 ;
                RECT 2.880 537.000 82.400 537.320 ;
                RECT 95.680 537.000 106.200 537.320 ;
                RECT 708.360 537.000 713.080 537.320 ;
                RECT 2.880 538.360 106.200 538.680 ;
                RECT 708.360 538.360 713.080 538.680 ;
                RECT 2.880 539.720 85.800 540.040 ;
                RECT 95.680 539.720 106.200 540.040 ;
                RECT 708.360 539.720 713.080 540.040 ;
                RECT 2.880 541.080 82.400 541.400 ;
                RECT 95.680 541.080 106.200 541.400 ;
                RECT 708.360 541.080 713.080 541.400 ;
                RECT 2.880 542.440 82.400 542.760 ;
                RECT 95.680 542.440 106.200 542.760 ;
                RECT 708.360 542.440 713.080 542.760 ;
                RECT 2.880 543.800 82.400 544.120 ;
                RECT 95.680 543.800 106.200 544.120 ;
                RECT 708.360 543.800 713.080 544.120 ;
                RECT 2.880 545.160 82.400 545.480 ;
                RECT 95.680 545.160 106.200 545.480 ;
                RECT 708.360 545.160 713.080 545.480 ;
                RECT 2.880 546.520 106.200 546.840 ;
                RECT 708.360 546.520 713.080 546.840 ;
                RECT 2.880 547.880 87.840 548.200 ;
                RECT 95.680 547.880 106.200 548.200 ;
                RECT 708.360 547.880 713.080 548.200 ;
                RECT 2.880 549.240 88.520 549.560 ;
                RECT 95.680 549.240 106.200 549.560 ;
                RECT 708.360 549.240 713.080 549.560 ;
                RECT 2.880 550.600 82.400 550.920 ;
                RECT 95.680 550.600 106.200 550.920 ;
                RECT 708.360 550.600 713.080 550.920 ;
                RECT 2.880 551.960 82.400 552.280 ;
                RECT 95.680 551.960 106.200 552.280 ;
                RECT 708.360 551.960 713.080 552.280 ;
                RECT 2.880 553.320 82.400 553.640 ;
                RECT 95.680 553.320 106.200 553.640 ;
                RECT 708.360 553.320 713.080 553.640 ;
                RECT 2.880 554.680 106.200 555.000 ;
                RECT 708.360 554.680 713.080 555.000 ;
                RECT 2.880 556.040 82.400 556.360 ;
                RECT 95.680 556.040 106.200 556.360 ;
                RECT 708.360 556.040 713.080 556.360 ;
                RECT 2.880 557.400 90.560 557.720 ;
                RECT 95.680 557.400 106.200 557.720 ;
                RECT 708.360 557.400 713.080 557.720 ;
                RECT 2.880 558.760 90.560 559.080 ;
                RECT 95.680 558.760 106.200 559.080 ;
                RECT 708.360 558.760 713.080 559.080 ;
                RECT 2.880 560.120 82.400 560.440 ;
                RECT 95.680 560.120 106.200 560.440 ;
                RECT 708.360 560.120 713.080 560.440 ;
                RECT 2.880 561.480 82.400 561.800 ;
                RECT 95.680 561.480 106.200 561.800 ;
                RECT 708.360 561.480 713.080 561.800 ;
                RECT 2.880 562.840 106.200 563.160 ;
                RECT 708.360 562.840 713.080 563.160 ;
                RECT 2.880 564.200 82.400 564.520 ;
                RECT 95.680 564.200 106.200 564.520 ;
                RECT 708.360 564.200 713.080 564.520 ;
                RECT 2.880 565.560 82.400 565.880 ;
                RECT 95.680 565.560 106.200 565.880 ;
                RECT 708.360 565.560 713.080 565.880 ;
                RECT 2.880 566.920 82.400 567.240 ;
                RECT 95.680 566.920 106.200 567.240 ;
                RECT 708.360 566.920 713.080 567.240 ;
                RECT 2.880 568.280 93.280 568.600 ;
                RECT 95.680 568.280 106.200 568.600 ;
                RECT 708.360 568.280 713.080 568.600 ;
                RECT 2.880 569.640 82.400 569.960 ;
                RECT 95.680 569.640 106.200 569.960 ;
                RECT 708.360 569.640 713.080 569.960 ;
                RECT 2.880 571.000 106.200 571.320 ;
                RECT 708.360 571.000 713.080 571.320 ;
                RECT 2.880 572.360 83.080 572.680 ;
                RECT 95.680 572.360 106.200 572.680 ;
                RECT 708.360 572.360 713.080 572.680 ;
                RECT 2.880 573.720 83.080 574.040 ;
                RECT 95.680 573.720 106.200 574.040 ;
                RECT 708.360 573.720 713.080 574.040 ;
                RECT 2.880 575.080 83.080 575.400 ;
                RECT 95.680 575.080 106.200 575.400 ;
                RECT 708.360 575.080 713.080 575.400 ;
                RECT 2.880 576.440 83.080 576.760 ;
                RECT 95.680 576.440 106.200 576.760 ;
                RECT 708.360 576.440 713.080 576.760 ;
                RECT 2.880 577.800 106.200 578.120 ;
                RECT 708.360 577.800 713.080 578.120 ;
                RECT 2.880 579.160 87.840 579.480 ;
                RECT 95.680 579.160 106.200 579.480 ;
                RECT 708.360 579.160 713.080 579.480 ;
                RECT 2.880 580.520 83.080 580.840 ;
                RECT 95.680 580.520 106.200 580.840 ;
                RECT 708.360 580.520 713.080 580.840 ;
                RECT 2.880 581.880 83.080 582.200 ;
                RECT 95.680 581.880 106.200 582.200 ;
                RECT 708.360 581.880 713.080 582.200 ;
                RECT 2.880 583.240 83.080 583.560 ;
                RECT 95.680 583.240 106.200 583.560 ;
                RECT 708.360 583.240 713.080 583.560 ;
                RECT 2.880 584.600 83.080 584.920 ;
                RECT 95.680 584.600 106.200 584.920 ;
                RECT 708.360 584.600 713.080 584.920 ;
                RECT 2.880 585.960 106.200 586.280 ;
                RECT 708.360 585.960 713.080 586.280 ;
                RECT 2.880 587.320 89.880 587.640 ;
                RECT 95.680 587.320 106.200 587.640 ;
                RECT 708.360 587.320 713.080 587.640 ;
                RECT 2.880 588.680 83.080 589.000 ;
                RECT 95.680 588.680 106.200 589.000 ;
                RECT 708.360 588.680 713.080 589.000 ;
                RECT 2.880 590.040 83.080 590.360 ;
                RECT 95.680 590.040 106.200 590.360 ;
                RECT 708.360 590.040 713.080 590.360 ;
                RECT 2.880 591.400 83.080 591.720 ;
                RECT 95.680 591.400 106.200 591.720 ;
                RECT 708.360 591.400 713.080 591.720 ;
                RECT 2.880 592.760 83.080 593.080 ;
                RECT 95.680 592.760 106.200 593.080 ;
                RECT 708.360 592.760 713.080 593.080 ;
                RECT 2.880 594.120 106.200 594.440 ;
                RECT 708.360 594.120 713.080 594.440 ;
                RECT 2.880 595.480 83.080 595.800 ;
                RECT 95.680 595.480 106.200 595.800 ;
                RECT 708.360 595.480 713.080 595.800 ;
                RECT 2.880 596.840 91.920 597.160 ;
                RECT 95.680 596.840 106.200 597.160 ;
                RECT 708.360 596.840 713.080 597.160 ;
                RECT 2.880 598.200 83.080 598.520 ;
                RECT 95.680 598.200 106.200 598.520 ;
                RECT 708.360 598.200 713.080 598.520 ;
                RECT 2.880 599.560 83.080 599.880 ;
                RECT 95.680 599.560 106.200 599.880 ;
                RECT 708.360 599.560 713.080 599.880 ;
                RECT 2.880 600.920 83.080 601.240 ;
                RECT 95.680 600.920 106.200 601.240 ;
                RECT 708.360 600.920 713.080 601.240 ;
                RECT 2.880 602.280 106.200 602.600 ;
                RECT 708.360 602.280 713.080 602.600 ;
                RECT 2.880 603.640 83.760 603.960 ;
                RECT 95.680 603.640 106.200 603.960 ;
                RECT 708.360 603.640 713.080 603.960 ;
                RECT 2.880 605.000 83.760 605.320 ;
                RECT 95.680 605.000 106.200 605.320 ;
                RECT 708.360 605.000 713.080 605.320 ;
                RECT 2.880 606.360 87.160 606.680 ;
                RECT 95.680 606.360 106.200 606.680 ;
                RECT 708.360 606.360 713.080 606.680 ;
                RECT 2.880 607.720 87.160 608.040 ;
                RECT 95.680 607.720 106.200 608.040 ;
                RECT 708.360 607.720 713.080 608.040 ;
                RECT 2.880 609.080 83.760 609.400 ;
                RECT 95.680 609.080 106.200 609.400 ;
                RECT 708.360 609.080 713.080 609.400 ;
                RECT 2.880 610.440 106.200 610.760 ;
                RECT 708.360 610.440 713.080 610.760 ;
                RECT 2.880 611.800 83.760 612.120 ;
                RECT 95.680 611.800 106.200 612.120 ;
                RECT 708.360 611.800 713.080 612.120 ;
                RECT 2.880 613.160 83.760 613.480 ;
                RECT 95.680 613.160 106.200 613.480 ;
                RECT 708.360 613.160 713.080 613.480 ;
                RECT 2.880 614.520 83.760 614.840 ;
                RECT 95.680 614.520 106.200 614.840 ;
                RECT 708.360 614.520 713.080 614.840 ;
                RECT 2.880 615.880 83.760 616.200 ;
                RECT 95.680 615.880 106.200 616.200 ;
                RECT 708.360 615.880 713.080 616.200 ;
                RECT 2.880 617.240 106.200 617.560 ;
                RECT 708.360 617.240 713.080 617.560 ;
                RECT 2.880 618.600 89.880 618.920 ;
                RECT 95.680 618.600 106.200 618.920 ;
                RECT 708.360 618.600 713.080 618.920 ;
                RECT 2.880 619.960 83.760 620.280 ;
                RECT 95.680 619.960 106.200 620.280 ;
                RECT 708.360 619.960 713.080 620.280 ;
                RECT 2.880 621.320 83.760 621.640 ;
                RECT 95.680 621.320 106.200 621.640 ;
                RECT 708.360 621.320 713.080 621.640 ;
                RECT 2.880 622.680 83.760 623.000 ;
                RECT 95.680 622.680 106.200 623.000 ;
                RECT 708.360 622.680 713.080 623.000 ;
                RECT 2.880 624.040 83.760 624.360 ;
                RECT 95.680 624.040 106.200 624.360 ;
                RECT 708.360 624.040 713.080 624.360 ;
                RECT 2.880 625.400 106.200 625.720 ;
                RECT 708.360 625.400 713.080 625.720 ;
                RECT 2.880 626.760 91.920 627.080 ;
                RECT 95.680 626.760 106.200 627.080 ;
                RECT 708.360 626.760 713.080 627.080 ;
                RECT 2.880 628.120 83.760 628.440 ;
                RECT 95.680 628.120 106.200 628.440 ;
                RECT 708.360 628.120 713.080 628.440 ;
                RECT 2.880 629.480 83.760 629.800 ;
                RECT 95.680 629.480 106.200 629.800 ;
                RECT 708.360 629.480 713.080 629.800 ;
                RECT 2.880 630.840 83.760 631.160 ;
                RECT 95.680 630.840 106.200 631.160 ;
                RECT 708.360 630.840 713.080 631.160 ;
                RECT 2.880 632.200 83.760 632.520 ;
                RECT 95.680 632.200 106.200 632.520 ;
                RECT 708.360 632.200 713.080 632.520 ;
                RECT 2.880 633.560 106.200 633.880 ;
                RECT 708.360 633.560 713.080 633.880 ;
                RECT 2.880 634.920 83.760 635.240 ;
                RECT 95.680 634.920 106.200 635.240 ;
                RECT 708.360 634.920 713.080 635.240 ;
                RECT 2.880 636.280 86.480 636.600 ;
                RECT 95.680 636.280 106.200 636.600 ;
                RECT 708.360 636.280 713.080 636.600 ;
                RECT 2.880 637.640 83.760 637.960 ;
                RECT 95.680 637.640 106.200 637.960 ;
                RECT 708.360 637.640 713.080 637.960 ;
                RECT 2.880 639.000 83.760 639.320 ;
                RECT 95.680 639.000 106.200 639.320 ;
                RECT 708.360 639.000 713.080 639.320 ;
                RECT 2.880 640.360 83.760 640.680 ;
                RECT 95.680 640.360 106.200 640.680 ;
                RECT 708.360 640.360 713.080 640.680 ;
                RECT 2.880 641.720 106.200 642.040 ;
                RECT 708.360 641.720 713.080 642.040 ;
                RECT 2.880 643.080 83.760 643.400 ;
                RECT 95.680 643.080 106.200 643.400 ;
                RECT 708.360 643.080 713.080 643.400 ;
                RECT 2.880 644.440 83.760 644.760 ;
                RECT 95.680 644.440 106.200 644.760 ;
                RECT 708.360 644.440 713.080 644.760 ;
                RECT 2.880 645.800 88.520 646.120 ;
                RECT 95.680 645.800 106.200 646.120 ;
                RECT 708.360 645.800 713.080 646.120 ;
                RECT 2.880 647.160 83.760 647.480 ;
                RECT 95.680 647.160 106.200 647.480 ;
                RECT 708.360 647.160 713.080 647.480 ;
                RECT 2.880 648.520 83.760 648.840 ;
                RECT 95.680 648.520 106.200 648.840 ;
                RECT 708.360 648.520 713.080 648.840 ;
                RECT 2.880 649.880 106.200 650.200 ;
                RECT 708.360 649.880 713.080 650.200 ;
                RECT 2.880 651.240 83.760 651.560 ;
                RECT 95.680 651.240 106.200 651.560 ;
                RECT 708.360 651.240 713.080 651.560 ;
                RECT 2.880 652.600 83.760 652.920 ;
                RECT 95.680 652.600 106.200 652.920 ;
                RECT 708.360 652.600 713.080 652.920 ;
                RECT 2.880 653.960 83.760 654.280 ;
                RECT 95.680 653.960 106.200 654.280 ;
                RECT 708.360 653.960 713.080 654.280 ;
                RECT 2.880 655.320 91.240 655.640 ;
                RECT 95.680 655.320 106.200 655.640 ;
                RECT 708.360 655.320 713.080 655.640 ;
                RECT 2.880 656.680 106.200 657.000 ;
                RECT 708.360 656.680 713.080 657.000 ;
                RECT 2.880 658.040 106.200 658.360 ;
                RECT 708.360 658.040 713.080 658.360 ;
                RECT 2.880 659.400 83.760 659.720 ;
                RECT 95.680 659.400 106.200 659.720 ;
                RECT 708.360 659.400 713.080 659.720 ;
                RECT 2.880 660.760 83.760 661.080 ;
                RECT 95.680 660.760 106.200 661.080 ;
                RECT 708.360 660.760 713.080 661.080 ;
                RECT 2.880 662.120 83.760 662.440 ;
                RECT 95.680 662.120 106.200 662.440 ;
                RECT 708.360 662.120 713.080 662.440 ;
                RECT 2.880 663.480 83.760 663.800 ;
                RECT 95.680 663.480 106.200 663.800 ;
                RECT 708.360 663.480 713.080 663.800 ;
                RECT 2.880 664.840 106.200 665.160 ;
                RECT 708.360 664.840 713.080 665.160 ;
                RECT 2.880 666.200 85.800 666.520 ;
                RECT 95.680 666.200 106.200 666.520 ;
                RECT 708.360 666.200 713.080 666.520 ;
                RECT 2.880 667.560 84.440 667.880 ;
                RECT 95.680 667.560 106.200 667.880 ;
                RECT 708.360 667.560 713.080 667.880 ;
                RECT 2.880 668.920 84.440 669.240 ;
                RECT 95.680 668.920 106.200 669.240 ;
                RECT 708.360 668.920 713.080 669.240 ;
                RECT 2.880 670.280 84.440 670.600 ;
                RECT 95.680 670.280 106.200 670.600 ;
                RECT 708.360 670.280 713.080 670.600 ;
                RECT 2.880 671.640 84.440 671.960 ;
                RECT 95.680 671.640 106.200 671.960 ;
                RECT 708.360 671.640 713.080 671.960 ;
                RECT 2.880 673.000 106.200 673.320 ;
                RECT 708.360 673.000 713.080 673.320 ;
                RECT 2.880 674.360 84.440 674.680 ;
                RECT 95.680 674.360 106.200 674.680 ;
                RECT 708.360 674.360 713.080 674.680 ;
                RECT 2.880 675.720 88.520 676.040 ;
                RECT 95.680 675.720 106.200 676.040 ;
                RECT 708.360 675.720 713.080 676.040 ;
                RECT 2.880 677.080 84.440 677.400 ;
                RECT 95.680 677.080 106.200 677.400 ;
                RECT 708.360 677.080 713.080 677.400 ;
                RECT 2.880 678.440 84.440 678.760 ;
                RECT 95.680 678.440 106.200 678.760 ;
                RECT 708.360 678.440 713.080 678.760 ;
                RECT 2.880 679.800 84.440 680.120 ;
                RECT 95.680 679.800 106.200 680.120 ;
                RECT 708.360 679.800 713.080 680.120 ;
                RECT 2.880 681.160 106.200 681.480 ;
                RECT 708.360 681.160 713.080 681.480 ;
                RECT 2.880 682.520 84.440 682.840 ;
                RECT 95.680 682.520 106.200 682.840 ;
                RECT 708.360 682.520 713.080 682.840 ;
                RECT 2.880 683.880 84.440 684.200 ;
                RECT 95.680 683.880 106.200 684.200 ;
                RECT 708.360 683.880 713.080 684.200 ;
                RECT 2.880 685.240 90.560 685.560 ;
                RECT 95.680 685.240 106.200 685.560 ;
                RECT 708.360 685.240 713.080 685.560 ;
                RECT 2.880 686.600 84.440 686.920 ;
                RECT 95.680 686.600 106.200 686.920 ;
                RECT 708.360 686.600 713.080 686.920 ;
                RECT 2.880 687.960 84.440 688.280 ;
                RECT 95.680 687.960 106.200 688.280 ;
                RECT 708.360 687.960 713.080 688.280 ;
                RECT 2.880 689.320 106.200 689.640 ;
                RECT 708.360 689.320 713.080 689.640 ;
                RECT 2.880 690.680 84.440 691.000 ;
                RECT 95.680 690.680 106.200 691.000 ;
                RECT 708.360 690.680 713.080 691.000 ;
                RECT 2.880 692.040 84.440 692.360 ;
                RECT 95.680 692.040 106.200 692.360 ;
                RECT 708.360 692.040 713.080 692.360 ;
                RECT 2.880 693.400 84.440 693.720 ;
                RECT 95.680 693.400 106.200 693.720 ;
                RECT 708.360 693.400 713.080 693.720 ;
                RECT 2.880 694.760 93.280 695.080 ;
                RECT 95.680 694.760 106.200 695.080 ;
                RECT 708.360 694.760 713.080 695.080 ;
                RECT 2.880 696.120 84.440 696.440 ;
                RECT 95.680 696.120 106.200 696.440 ;
                RECT 708.360 696.120 713.080 696.440 ;
                RECT 2.880 697.480 106.200 697.800 ;
                RECT 708.360 697.480 713.080 697.800 ;
                RECT 2.880 698.840 85.120 699.160 ;
                RECT 95.680 698.840 106.200 699.160 ;
                RECT 708.360 698.840 713.080 699.160 ;
                RECT 2.880 700.200 85.120 700.520 ;
                RECT 95.680 700.200 106.200 700.520 ;
                RECT 708.360 700.200 713.080 700.520 ;
                RECT 2.880 701.560 85.120 701.880 ;
                RECT 95.680 701.560 106.200 701.880 ;
                RECT 708.360 701.560 713.080 701.880 ;
                RECT 2.880 702.920 85.120 703.240 ;
                RECT 95.680 702.920 106.200 703.240 ;
                RECT 708.360 702.920 713.080 703.240 ;
                RECT 2.880 704.280 106.200 704.600 ;
                RECT 708.360 704.280 713.080 704.600 ;
                RECT 2.880 705.640 87.840 705.960 ;
                RECT 95.680 705.640 106.200 705.960 ;
                RECT 708.360 705.640 713.080 705.960 ;
                RECT 2.880 707.000 85.120 707.320 ;
                RECT 95.680 707.000 106.200 707.320 ;
                RECT 708.360 707.000 713.080 707.320 ;
                RECT 2.880 708.360 85.120 708.680 ;
                RECT 95.680 708.360 106.200 708.680 ;
                RECT 708.360 708.360 713.080 708.680 ;
                RECT 2.880 709.720 85.120 710.040 ;
                RECT 95.680 709.720 106.200 710.040 ;
                RECT 708.360 709.720 713.080 710.040 ;
                RECT 2.880 711.080 85.120 711.400 ;
                RECT 95.680 711.080 106.200 711.400 ;
                RECT 708.360 711.080 713.080 711.400 ;
                RECT 2.880 712.440 106.200 712.760 ;
                RECT 708.360 712.440 713.080 712.760 ;
                RECT 2.880 713.800 89.880 714.120 ;
                RECT 95.680 713.800 106.200 714.120 ;
                RECT 708.360 713.800 713.080 714.120 ;
                RECT 2.880 715.160 90.560 715.480 ;
                RECT 95.680 715.160 106.200 715.480 ;
                RECT 708.360 715.160 713.080 715.480 ;
                RECT 2.880 716.520 85.120 716.840 ;
                RECT 95.680 716.520 106.200 716.840 ;
                RECT 708.360 716.520 713.080 716.840 ;
                RECT 2.880 717.880 85.120 718.200 ;
                RECT 95.680 717.880 106.200 718.200 ;
                RECT 708.360 717.880 713.080 718.200 ;
                RECT 2.880 719.240 85.120 719.560 ;
                RECT 95.680 719.240 106.200 719.560 ;
                RECT 708.360 719.240 713.080 719.560 ;
                RECT 2.880 720.600 106.200 720.920 ;
                RECT 708.360 720.600 713.080 720.920 ;
                RECT 2.880 721.960 85.120 722.280 ;
                RECT 95.680 721.960 106.200 722.280 ;
                RECT 708.360 721.960 713.080 722.280 ;
                RECT 2.880 723.320 85.120 723.640 ;
                RECT 95.680 723.320 106.200 723.640 ;
                RECT 708.360 723.320 713.080 723.640 ;
                RECT 2.880 724.680 92.600 725.000 ;
                RECT 95.680 724.680 106.200 725.000 ;
                RECT 708.360 724.680 713.080 725.000 ;
                RECT 2.880 726.040 85.120 726.360 ;
                RECT 95.680 726.040 106.200 726.360 ;
                RECT 708.360 726.040 713.080 726.360 ;
                RECT 2.880 727.400 85.120 727.720 ;
                RECT 95.680 727.400 106.200 727.720 ;
                RECT 708.360 727.400 713.080 727.720 ;
                RECT 2.880 728.760 106.200 729.080 ;
                RECT 708.360 728.760 713.080 729.080 ;
                RECT 2.880 730.120 85.800 730.440 ;
                RECT 95.680 730.120 106.200 730.440 ;
                RECT 708.360 730.120 713.080 730.440 ;
                RECT 2.880 731.480 85.800 731.800 ;
                RECT 95.680 731.480 106.200 731.800 ;
                RECT 708.360 731.480 713.080 731.800 ;
                RECT 2.880 732.840 85.800 733.160 ;
                RECT 95.680 732.840 106.200 733.160 ;
                RECT 708.360 732.840 713.080 733.160 ;
                RECT 2.880 734.200 87.160 734.520 ;
                RECT 95.680 734.200 106.200 734.520 ;
                RECT 708.360 734.200 713.080 734.520 ;
                RECT 2.880 735.560 85.800 735.880 ;
                RECT 95.680 735.560 106.200 735.880 ;
                RECT 708.360 735.560 713.080 735.880 ;
                RECT 2.880 736.920 106.200 737.240 ;
                RECT 708.360 736.920 713.080 737.240 ;
                RECT 2.880 738.280 85.800 738.600 ;
                RECT 95.680 738.280 106.200 738.600 ;
                RECT 708.360 738.280 713.080 738.600 ;
                RECT 2.880 739.640 85.800 739.960 ;
                RECT 95.680 739.640 106.200 739.960 ;
                RECT 708.360 739.640 713.080 739.960 ;
                RECT 2.880 741.000 85.800 741.320 ;
                RECT 95.680 741.000 106.200 741.320 ;
                RECT 708.360 741.000 713.080 741.320 ;
                RECT 2.880 742.360 85.800 742.680 ;
                RECT 95.680 742.360 106.200 742.680 ;
                RECT 708.360 742.360 713.080 742.680 ;
                RECT 2.880 743.720 106.200 744.040 ;
                RECT 708.360 743.720 713.080 744.040 ;
                RECT 2.880 745.080 89.880 745.400 ;
                RECT 95.680 745.080 106.200 745.400 ;
                RECT 708.360 745.080 713.080 745.400 ;
                RECT 2.880 746.440 85.800 746.760 ;
                RECT 95.680 746.440 106.200 746.760 ;
                RECT 708.360 746.440 713.080 746.760 ;
                RECT 2.880 747.800 85.800 748.120 ;
                RECT 95.680 747.800 106.200 748.120 ;
                RECT 708.360 747.800 713.080 748.120 ;
                RECT 2.880 749.160 85.800 749.480 ;
                RECT 95.680 749.160 106.200 749.480 ;
                RECT 708.360 749.160 713.080 749.480 ;
                RECT 2.880 750.520 85.800 750.840 ;
                RECT 95.680 750.520 106.200 750.840 ;
                RECT 708.360 750.520 713.080 750.840 ;
                RECT 2.880 751.880 106.200 752.200 ;
                RECT 708.360 751.880 713.080 752.200 ;
                RECT 2.880 753.240 91.920 753.560 ;
                RECT 95.680 753.240 106.200 753.560 ;
                RECT 708.360 753.240 713.080 753.560 ;
                RECT 2.880 754.600 85.800 754.920 ;
                RECT 95.680 754.600 106.200 754.920 ;
                RECT 708.360 754.600 713.080 754.920 ;
                RECT 2.880 755.960 85.800 756.280 ;
                RECT 95.680 755.960 106.200 756.280 ;
                RECT 708.360 755.960 713.080 756.280 ;
                RECT 2.880 757.320 85.800 757.640 ;
                RECT 95.680 757.320 106.200 757.640 ;
                RECT 708.360 757.320 713.080 757.640 ;
                RECT 2.880 758.680 85.800 759.000 ;
                RECT 95.680 758.680 106.200 759.000 ;
                RECT 708.360 758.680 713.080 759.000 ;
                RECT 2.880 760.040 106.200 760.360 ;
                RECT 708.360 760.040 713.080 760.360 ;
                RECT 2.880 761.400 298.640 761.720 ;
                RECT 708.360 761.400 713.080 761.720 ;
                RECT 2.880 762.760 298.640 763.080 ;
                RECT 708.360 762.760 713.080 763.080 ;
                RECT 2.880 764.120 298.640 764.440 ;
                RECT 708.360 764.120 713.080 764.440 ;
                RECT 2.880 765.480 713.080 765.800 ;
                RECT 2.880 766.840 713.080 767.160 ;
                RECT 2.880 768.200 713.080 768.520 ;
                RECT 2.880 769.560 713.080 769.880 ;
                RECT 2.880 770.920 713.080 771.240 ;
                RECT 2.880 2.880 713.080 4.240 ;
                RECT 2.880 772.240 713.080 773.600 ;
                RECT 302.780 39.245 308.580 40.365 ;
                RECT 698.680 39.245 704.480 40.365 ;
                RECT 302.780 45.065 308.580 45.755 ;
                RECT 698.680 45.065 704.480 45.755 ;
                RECT 302.780 50.640 308.580 51.430 ;
                RECT 698.680 50.640 704.480 51.430 ;
                RECT 302.780 56.760 308.580 57.340 ;
                RECT 698.680 56.760 704.480 57.340 ;
                RECT 302.780 61.480 308.580 62.070 ;
                RECT 698.680 61.480 704.480 62.070 ;
                RECT 302.780 66.300 308.580 66.890 ;
                RECT 698.680 66.300 704.480 66.890 ;
                RECT 302.780 88.850 704.480 89.650 ;
                RECT 302.780 91.860 704.480 92.660 ;
                RECT 302.780 102.860 704.480 106.460 ;
                RECT 302.780 135.595 704.480 135.885 ;
                RECT 302.780 79.800 704.480 81.600 ;
                RECT 302.780 187.490 704.480 189.290 ;
                RECT 302.780 93.540 704.480 94.340 ;
                RECT 302.780 96.750 704.480 97.550 ;
                RECT 302.780 29.875 704.480 31.675 ;
                RECT 106.640 253.835 108.390 761.015 ;
                RECT 120.625 253.835 122.545 761.015 ;
                RECT 144.400 253.835 146.320 761.015 ;
                RECT 148.240 253.835 150.160 761.015 ;
                RECT 152.080 253.835 154.000 761.015 ;
                RECT 194.650 253.835 196.570 761.015 ;
                RECT 198.490 253.835 200.410 761.015 ;
                RECT 202.330 253.835 204.250 761.015 ;
                RECT 206.170 253.835 208.090 761.015 ;
                RECT 210.010 253.835 211.930 761.015 ;
                RECT 213.850 253.835 215.770 761.015 ;
                RECT 217.690 253.835 219.610 761.015 ;
                RECT 156.540 55.635 157.430 134.035 ;
                RECT 162.870 55.635 163.760 134.035 ;
                RECT 169.630 55.635 170.520 134.035 ;
                RECT 175.960 55.635 176.850 134.035 ;
                RECT 183.150 55.635 184.900 134.035 ;
                RECT 197.135 55.635 199.055 134.035 ;
                RECT 221.340 55.635 223.260 134.035 ;
                RECT 225.180 55.635 227.100 134.035 ;
                RECT 229.020 55.635 230.940 134.035 ;
                RECT 202.505 199.700 203.825 247.200 ;
                RECT 211.630 199.700 212.520 247.200 ;
                RECT 217.960 199.700 218.850 247.200 ;
                RECT 224.290 199.700 226.040 247.200 ;
                RECT 238.075 199.700 239.995 247.200 ;
                RECT 241.915 199.700 243.835 247.200 ;
                RECT 196.030 188.540 196.920 193.700 ;
                RECT 203.135 188.540 205.055 193.700 ;
                RECT 220.890 188.540 222.810 193.700 ;
                RECT 224.730 188.540 226.650 193.700 ;
                RECT 228.570 188.540 230.490 193.700 ;
                RECT 265.880 44.475 266.770 49.635 ;
                RECT 27.350 254.900 36.510 255.270 ;
                RECT 27.350 258.340 36.510 259.450 ;
                RECT 79.510 236.660 97.950 237.330 ;
                RECT 79.510 237.890 97.950 240.940 ;
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 715.960 776.480 ;
        LAYER met2 ;
            RECT 0.000 0.000 715.960 776.480 ;
    END 
END sram22_1024x64m4w8 
END LIBRARY 

