VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram22_1024x32m8w32
  CLASS BLOCK ;
  ORIGIN 89.065 244.085 ;
  FOREIGN sram22_1024x32m8w32 -89.065 -244.085 ;
  SIZE 458.29 BY 492.25 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 361.595 246.76 361.925 247.89 ;
        RECT 361.595 241.915 361.925 242.245 ;
        RECT 361.595 240.555 361.925 240.885 ;
        RECT 361.595 239.195 361.925 239.525 ;
        RECT 361.595 237.835 361.925 238.165 ;
        RECT 361.595 236.475 361.925 236.805 ;
        RECT 361.595 235.115 361.925 235.445 ;
        RECT 361.595 233.755 361.925 234.085 ;
        RECT 361.595 232.395 361.925 232.725 ;
        RECT 361.595 231.035 361.925 231.365 ;
        RECT 361.595 229.675 361.925 230.005 ;
        RECT 361.595 228.315 361.925 228.645 ;
        RECT 361.595 226.955 361.925 227.285 ;
        RECT 361.595 225.595 361.925 225.925 ;
        RECT 361.595 224.235 361.925 224.565 ;
        RECT 361.595 222.875 361.925 223.205 ;
        RECT 361.595 221.515 361.925 221.845 ;
        RECT 361.595 220.155 361.925 220.485 ;
        RECT 361.595 218.795 361.925 219.125 ;
        RECT 361.595 217.435 361.925 217.765 ;
        RECT 361.595 216.075 361.925 216.405 ;
        RECT 361.595 214.715 361.925 215.045 ;
        RECT 361.595 213.355 361.925 213.685 ;
        RECT 361.595 211.995 361.925 212.325 ;
        RECT 361.595 210.635 361.925 210.965 ;
        RECT 361.595 209.275 361.925 209.605 ;
        RECT 361.595 207.915 361.925 208.245 ;
        RECT 361.595 206.555 361.925 206.885 ;
        RECT 361.595 205.195 361.925 205.525 ;
        RECT 361.595 203.835 361.925 204.165 ;
        RECT 361.595 202.475 361.925 202.805 ;
        RECT 361.595 201.115 361.925 201.445 ;
        RECT 361.595 199.755 361.925 200.085 ;
        RECT 361.595 198.395 361.925 198.725 ;
        RECT 361.595 197.035 361.925 197.365 ;
        RECT 361.595 195.675 361.925 196.005 ;
        RECT 361.595 194.315 361.925 194.645 ;
        RECT 361.595 192.955 361.925 193.285 ;
        RECT 361.595 191.595 361.925 191.925 ;
        RECT 361.595 190.235 361.925 190.565 ;
        RECT 361.595 188.875 361.925 189.205 ;
        RECT 361.595 187.515 361.925 187.845 ;
        RECT 361.595 186.155 361.925 186.485 ;
        RECT 361.595 184.795 361.925 185.125 ;
        RECT 361.595 183.435 361.925 183.765 ;
        RECT 361.595 182.075 361.925 182.405 ;
        RECT 361.595 180.715 361.925 181.045 ;
        RECT 361.595 179.355 361.925 179.685 ;
        RECT 361.595 177.995 361.925 178.325 ;
        RECT 361.595 176.635 361.925 176.965 ;
        RECT 361.595 175.275 361.925 175.605 ;
        RECT 361.595 173.915 361.925 174.245 ;
        RECT 361.595 172.555 361.925 172.885 ;
        RECT 361.595 171.195 361.925 171.525 ;
        RECT 361.595 169.835 361.925 170.165 ;
        RECT 361.595 168.475 361.925 168.805 ;
        RECT 361.595 167.115 361.925 167.445 ;
        RECT 361.595 165.755 361.925 166.085 ;
        RECT 361.595 164.395 361.925 164.725 ;
        RECT 361.595 163.035 361.925 163.365 ;
        RECT 361.595 161.675 361.925 162.005 ;
        RECT 361.595 160.315 361.925 160.645 ;
        RECT 361.595 158.955 361.925 159.285 ;
        RECT 361.595 157.595 361.925 157.925 ;
        RECT 361.595 156.235 361.925 156.565 ;
        RECT 361.595 154.875 361.925 155.205 ;
        RECT 361.595 153.515 361.925 153.845 ;
        RECT 361.595 152.155 361.925 152.485 ;
        RECT 361.595 150.795 361.925 151.125 ;
        RECT 361.595 149.435 361.925 149.765 ;
        RECT 361.595 148.075 361.925 148.405 ;
        RECT 361.595 146.715 361.925 147.045 ;
        RECT 361.595 145.355 361.925 145.685 ;
        RECT 361.595 143.995 361.925 144.325 ;
        RECT 361.595 142.635 361.925 142.965 ;
        RECT 361.595 141.275 361.925 141.605 ;
        RECT 361.595 139.915 361.925 140.245 ;
        RECT 361.595 138.555 361.925 138.885 ;
        RECT 361.595 137.195 361.925 137.525 ;
        RECT 361.595 135.835 361.925 136.165 ;
        RECT 361.595 134.475 361.925 134.805 ;
        RECT 361.595 133.115 361.925 133.445 ;
        RECT 361.595 131.755 361.925 132.085 ;
        RECT 361.595 130.395 361.925 130.725 ;
        RECT 361.595 129.035 361.925 129.365 ;
        RECT 361.595 127.675 361.925 128.005 ;
        RECT 361.595 126.315 361.925 126.645 ;
        RECT 361.595 124.955 361.925 125.285 ;
        RECT 361.595 123.595 361.925 123.925 ;
        RECT 361.595 122.235 361.925 122.565 ;
        RECT 361.595 120.875 361.925 121.205 ;
        RECT 361.595 119.515 361.925 119.845 ;
        RECT 361.595 118.155 361.925 118.485 ;
        RECT 361.595 116.795 361.925 117.125 ;
        RECT 361.595 115.435 361.925 115.765 ;
        RECT 361.595 114.075 361.925 114.405 ;
        RECT 361.595 112.715 361.925 113.045 ;
        RECT 361.595 111.355 361.925 111.685 ;
        RECT 361.595 109.995 361.925 110.325 ;
        RECT 361.595 108.635 361.925 108.965 ;
        RECT 361.595 107.275 361.925 107.605 ;
        RECT 361.595 105.915 361.925 106.245 ;
        RECT 361.595 104.555 361.925 104.885 ;
        RECT 361.595 103.195 361.925 103.525 ;
        RECT 361.595 101.835 361.925 102.165 ;
        RECT 361.595 100.475 361.925 100.805 ;
        RECT 361.595 99.115 361.925 99.445 ;
        RECT 361.595 97.755 361.925 98.085 ;
        RECT 361.595 96.395 361.925 96.725 ;
        RECT 361.595 95.035 361.925 95.365 ;
        RECT 361.595 93.675 361.925 94.005 ;
        RECT 361.595 92.315 361.925 92.645 ;
        RECT 361.595 90.955 361.925 91.285 ;
        RECT 361.595 89.595 361.925 89.925 ;
        RECT 361.595 88.235 361.925 88.565 ;
        RECT 361.595 86.875 361.925 87.205 ;
        RECT 361.595 85.515 361.925 85.845 ;
        RECT 361.595 84.155 361.925 84.485 ;
        RECT 361.595 82.795 361.925 83.125 ;
        RECT 361.595 81.435 361.925 81.765 ;
        RECT 361.595 80.075 361.925 80.405 ;
        RECT 361.595 78.715 361.925 79.045 ;
        RECT 361.595 77.355 361.925 77.685 ;
        RECT 361.595 75.995 361.925 76.325 ;
        RECT 361.595 74.635 361.925 74.965 ;
        RECT 361.595 73.275 361.925 73.605 ;
        RECT 361.595 71.915 361.925 72.245 ;
        RECT 361.595 70.555 361.925 70.885 ;
        RECT 361.595 69.195 361.925 69.525 ;
        RECT 361.595 67.835 361.925 68.165 ;
        RECT 361.595 66.475 361.925 66.805 ;
        RECT 361.595 65.115 361.925 65.445 ;
        RECT 361.595 63.755 361.925 64.085 ;
        RECT 361.595 62.395 361.925 62.725 ;
        RECT 361.595 61.035 361.925 61.365 ;
        RECT 361.595 59.675 361.925 60.005 ;
        RECT 361.595 58.315 361.925 58.645 ;
        RECT 361.595 56.955 361.925 57.285 ;
        RECT 361.595 55.595 361.925 55.925 ;
        RECT 361.595 54.235 361.925 54.565 ;
        RECT 361.595 52.875 361.925 53.205 ;
        RECT 361.595 51.515 361.925 51.845 ;
        RECT 361.595 50.155 361.925 50.485 ;
        RECT 361.595 48.795 361.925 49.125 ;
        RECT 361.595 47.435 361.925 47.765 ;
        RECT 361.595 46.075 361.925 46.405 ;
        RECT 361.595 44.715 361.925 45.045 ;
        RECT 361.595 43.355 361.925 43.685 ;
        RECT 361.595 41.995 361.925 42.325 ;
        RECT 361.595 40.635 361.925 40.965 ;
        RECT 361.595 39.275 361.925 39.605 ;
        RECT 361.595 37.915 361.925 38.245 ;
        RECT 361.595 36.555 361.925 36.885 ;
        RECT 361.595 35.195 361.925 35.525 ;
        RECT 361.595 33.835 361.925 34.165 ;
        RECT 361.595 32.475 361.925 32.805 ;
        RECT 361.595 31.115 361.925 31.445 ;
        RECT 361.595 29.755 361.925 30.085 ;
        RECT 361.595 28.395 361.925 28.725 ;
        RECT 361.595 27.035 361.925 27.365 ;
        RECT 361.595 25.675 361.925 26.005 ;
        RECT 361.595 24.315 361.925 24.645 ;
        RECT 361.595 22.955 361.925 23.285 ;
        RECT 361.595 21.595 361.925 21.925 ;
        RECT 361.595 20.235 361.925 20.565 ;
        RECT 361.595 18.875 361.925 19.205 ;
        RECT 361.595 17.515 361.925 17.845 ;
        RECT 361.595 16.155 361.925 16.485 ;
        RECT 361.595 14.795 361.925 15.125 ;
        RECT 361.595 13.435 361.925 13.765 ;
        RECT 361.595 12.075 361.925 12.405 ;
        RECT 361.595 10.715 361.925 11.045 ;
        RECT 361.595 9.355 361.925 9.685 ;
        RECT 361.595 7.995 361.925 8.325 ;
        RECT 361.595 6.635 361.925 6.965 ;
        RECT 361.595 5.275 361.925 5.605 ;
        RECT 361.595 3.915 361.925 4.245 ;
        RECT 361.595 2.555 361.925 2.885 ;
        RECT 361.595 1.195 361.925 1.525 ;
        RECT 361.595 -0.165 361.925 0.165 ;
        RECT 361.595 -1.525 361.925 -1.195 ;
        RECT 361.595 -2.885 361.925 -2.555 ;
        RECT 361.595 -4.245 361.925 -3.915 ;
        RECT 361.595 -5.605 361.925 -5.275 ;
        RECT 361.595 -6.965 361.925 -6.635 ;
        RECT 361.595 -8.325 361.925 -7.995 ;
        RECT 361.595 -9.685 361.925 -9.355 ;
        RECT 361.595 -11.045 361.925 -10.715 ;
        RECT 361.595 -12.405 361.925 -12.075 ;
        RECT 361.595 -13.765 361.925 -13.435 ;
        RECT 361.595 -15.125 361.925 -14.795 ;
        RECT 361.595 -16.485 361.925 -16.155 ;
        RECT 361.595 -17.845 361.925 -17.515 ;
        RECT 361.595 -19.205 361.925 -18.875 ;
        RECT 361.595 -20.565 361.925 -20.235 ;
        RECT 361.595 -21.925 361.925 -21.595 ;
        RECT 361.595 -23.285 361.925 -22.955 ;
        RECT 361.595 -24.645 361.925 -24.315 ;
        RECT 361.595 -26.005 361.925 -25.675 ;
        RECT 361.595 -27.365 361.925 -27.035 ;
        RECT 361.595 -28.725 361.925 -28.395 ;
        RECT 361.595 -30.085 361.925 -29.755 ;
        RECT 361.595 -31.445 361.925 -31.115 ;
        RECT 361.595 -32.805 361.925 -32.475 ;
        RECT 361.595 -34.165 361.925 -33.835 ;
        RECT 361.595 -35.525 361.925 -35.195 ;
        RECT 361.595 -36.885 361.925 -36.555 ;
        RECT 361.595 -38.245 361.925 -37.915 ;
        RECT 361.595 -39.605 361.925 -39.275 ;
        RECT 361.595 -40.965 361.925 -40.635 ;
        RECT 361.595 -42.325 361.925 -41.995 ;
        RECT 361.595 -43.685 361.925 -43.355 ;
        RECT 361.595 -45.045 361.925 -44.715 ;
        RECT 361.595 -46.405 361.925 -46.075 ;
        RECT 361.595 -47.765 361.925 -47.435 ;
        RECT 361.595 -49.125 361.925 -48.795 ;
        RECT 361.595 -50.485 361.925 -50.155 ;
        RECT 361.595 -51.845 361.925 -51.515 ;
        RECT 361.595 -53.205 361.925 -52.875 ;
        RECT 361.595 -54.565 361.925 -54.235 ;
        RECT 361.595 -55.925 361.925 -55.595 ;
        RECT 361.595 -57.285 361.925 -56.955 ;
        RECT 361.595 -58.645 361.925 -58.315 ;
        RECT 361.595 -60.005 361.925 -59.675 ;
        RECT 361.595 -61.365 361.925 -61.035 ;
        RECT 361.595 -62.725 361.925 -62.395 ;
        RECT 361.595 -64.085 361.925 -63.755 ;
        RECT 361.595 -65.445 361.925 -65.115 ;
        RECT 361.595 -66.805 361.925 -66.475 ;
        RECT 361.595 -68.165 361.925 -67.835 ;
        RECT 361.595 -69.525 361.925 -69.195 ;
        RECT 361.595 -70.885 361.925 -70.555 ;
        RECT 361.595 -72.245 361.925 -71.915 ;
        RECT 361.595 -73.605 361.925 -73.275 ;
        RECT 361.595 -74.965 361.925 -74.635 ;
        RECT 361.595 -76.325 361.925 -75.995 ;
        RECT 361.595 -77.685 361.925 -77.355 ;
        RECT 361.595 -79.045 361.925 -78.715 ;
        RECT 361.595 -80.405 361.925 -80.075 ;
        RECT 361.595 -81.765 361.925 -81.435 ;
        RECT 361.595 -83.125 361.925 -82.795 ;
        RECT 361.595 -84.485 361.925 -84.155 ;
        RECT 361.595 -85.845 361.925 -85.515 ;
        RECT 361.595 -87.205 361.925 -86.875 ;
        RECT 361.595 -88.565 361.925 -88.235 ;
        RECT 361.595 -89.925 361.925 -89.595 ;
        RECT 361.595 -91.285 361.925 -90.955 ;
        RECT 361.595 -92.645 361.925 -92.315 ;
        RECT 361.595 -94.005 361.925 -93.675 ;
        RECT 361.595 -95.365 361.925 -95.035 ;
        RECT 361.595 -96.725 361.925 -96.395 ;
        RECT 361.595 -98.085 361.925 -97.755 ;
        RECT 361.595 -99.445 361.925 -99.115 ;
        RECT 361.595 -100.805 361.925 -100.475 ;
        RECT 361.595 -102.165 361.925 -101.835 ;
        RECT 361.595 -103.525 361.925 -103.195 ;
        RECT 361.595 -104.885 361.925 -104.555 ;
        RECT 361.595 -106.245 361.925 -105.915 ;
        RECT 361.595 -107.605 361.925 -107.275 ;
        RECT 361.595 -108.965 361.925 -108.635 ;
        RECT 361.595 -110.325 361.925 -109.995 ;
        RECT 361.595 -111.685 361.925 -111.355 ;
        RECT 361.595 -113.045 361.925 -112.715 ;
        RECT 361.595 -114.405 361.925 -114.075 ;
        RECT 361.595 -115.765 361.925 -115.435 ;
        RECT 361.595 -117.125 361.925 -116.795 ;
        RECT 361.595 -118.485 361.925 -118.155 ;
        RECT 361.595 -119.845 361.925 -119.515 ;
        RECT 361.595 -121.205 361.925 -120.875 ;
        RECT 361.595 -122.565 361.925 -122.235 ;
        RECT 361.595 -123.925 361.925 -123.595 ;
        RECT 361.595 -125.285 361.925 -124.955 ;
        RECT 361.595 -126.645 361.925 -126.315 ;
        RECT 361.595 -128.005 361.925 -127.675 ;
        RECT 361.595 -129.365 361.925 -129.035 ;
        RECT 361.595 -130.725 361.925 -130.395 ;
        RECT 361.595 -132.085 361.925 -131.755 ;
        RECT 361.595 -133.445 361.925 -133.115 ;
        RECT 361.595 -134.805 361.925 -134.475 ;
        RECT 361.595 -136.165 361.925 -135.835 ;
        RECT 361.595 -137.525 361.925 -137.195 ;
        RECT 361.595 -138.885 361.925 -138.555 ;
        RECT 361.595 -140.245 361.925 -139.915 ;
        RECT 361.595 -141.605 361.925 -141.275 ;
        RECT 361.595 -142.965 361.925 -142.635 ;
        RECT 361.595 -144.325 361.925 -143.995 ;
        RECT 361.595 -145.685 361.925 -145.355 ;
        RECT 361.595 -147.045 361.925 -146.715 ;
        RECT 361.595 -148.405 361.925 -148.075 ;
        RECT 361.595 -149.765 361.925 -149.435 ;
        RECT 361.595 -151.125 361.925 -150.795 ;
        RECT 361.595 -152.485 361.925 -152.155 ;
        RECT 361.595 -153.845 361.925 -153.515 ;
        RECT 361.595 -155.205 361.925 -154.875 ;
        RECT 361.595 -156.565 361.925 -156.235 ;
        RECT 361.595 -157.925 361.925 -157.595 ;
        RECT 361.595 -159.285 361.925 -158.955 ;
        RECT 361.595 -160.645 361.925 -160.315 ;
        RECT 361.595 -162.005 361.925 -161.675 ;
        RECT 361.595 -163.365 361.925 -163.035 ;
        RECT 361.595 -164.725 361.925 -164.395 ;
        RECT 361.595 -166.085 361.925 -165.755 ;
        RECT 361.595 -167.445 361.925 -167.115 ;
        RECT 361.595 -168.805 361.925 -168.475 ;
        RECT 361.595 -170.165 361.925 -169.835 ;
        RECT 361.595 -171.525 361.925 -171.195 ;
        RECT 361.595 -172.885 361.925 -172.555 ;
        RECT 361.595 -174.245 361.925 -173.915 ;
        RECT 361.595 -175.605 361.925 -175.275 ;
        RECT 361.595 -176.965 361.925 -176.635 ;
        RECT 361.595 -178.325 361.925 -177.995 ;
        RECT 361.595 -179.685 361.925 -179.355 ;
        RECT 361.595 -181.045 361.925 -180.715 ;
        RECT 361.595 -182.405 361.925 -182.075 ;
        RECT 361.595 -183.765 361.925 -183.435 ;
        RECT 361.595 -185.125 361.925 -184.795 ;
        RECT 361.595 -186.485 361.925 -186.155 ;
        RECT 361.595 -187.845 361.925 -187.515 ;
        RECT 361.595 -189.205 361.925 -188.875 ;
        RECT 361.595 -190.565 361.925 -190.235 ;
        RECT 361.595 -191.925 361.925 -191.595 ;
        RECT 361.595 -193.285 361.925 -192.955 ;
        RECT 361.595 -194.645 361.925 -194.315 ;
        RECT 361.595 -196.005 361.925 -195.675 ;
        RECT 361.595 -197.365 361.925 -197.035 ;
        RECT 361.595 -198.725 361.925 -198.395 ;
        RECT 361.595 -200.085 361.925 -199.755 ;
        RECT 361.595 -201.445 361.925 -201.115 ;
        RECT 361.595 -202.805 361.925 -202.475 ;
        RECT 361.595 -204.165 361.925 -203.835 ;
        RECT 361.595 -205.525 361.925 -205.195 ;
        RECT 361.595 -206.885 361.925 -206.555 ;
        RECT 361.595 -208.245 361.925 -207.915 ;
        RECT 361.595 -209.605 361.925 -209.275 ;
        RECT 361.595 -210.965 361.925 -210.635 ;
        RECT 361.595 -212.325 361.925 -211.995 ;
        RECT 361.595 -213.685 361.925 -213.355 ;
        RECT 361.595 -215.045 361.925 -214.715 ;
        RECT 361.595 -216.405 361.925 -216.075 ;
        RECT 361.595 -217.765 361.925 -217.435 ;
        RECT 361.595 -219.125 361.925 -218.795 ;
        RECT 361.595 -220.485 361.925 -220.155 ;
        RECT 361.595 -221.845 361.925 -221.515 ;
        RECT 361.595 -223.205 361.925 -222.875 ;
        RECT 361.595 -224.565 361.925 -224.235 ;
        RECT 361.595 -225.925 361.925 -225.595 ;
        RECT 361.595 -227.285 361.925 -226.955 ;
        RECT 361.595 -228.645 361.925 -228.315 ;
        RECT 361.595 -230.005 361.925 -229.675 ;
        RECT 361.595 -231.365 361.925 -231.035 ;
        RECT 361.595 -232.725 361.925 -232.395 ;
        RECT 361.595 -234.085 361.925 -233.755 ;
        RECT 361.595 -235.445 361.925 -235.115 ;
        RECT 361.595 -236.805 361.925 -236.475 ;
        RECT 361.595 -238.165 361.925 -237.835 ;
        RECT 361.595 -243.81 361.925 -242.68 ;
        RECT 361.6 -243.925 361.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.955 246.76 363.285 247.89 ;
        RECT 362.955 241.915 363.285 242.245 ;
        RECT 362.955 240.555 363.285 240.885 ;
        RECT 362.955 239.195 363.285 239.525 ;
        RECT 362.955 237.835 363.285 238.165 ;
        RECT 362.955 236.475 363.285 236.805 ;
        RECT 362.955 235.115 363.285 235.445 ;
        RECT 362.955 233.755 363.285 234.085 ;
        RECT 362.955 232.395 363.285 232.725 ;
        RECT 362.955 231.035 363.285 231.365 ;
        RECT 362.955 229.675 363.285 230.005 ;
        RECT 362.955 228.315 363.285 228.645 ;
        RECT 362.955 226.955 363.285 227.285 ;
        RECT 362.955 225.595 363.285 225.925 ;
        RECT 362.955 224.235 363.285 224.565 ;
        RECT 362.955 222.875 363.285 223.205 ;
        RECT 362.955 221.515 363.285 221.845 ;
        RECT 362.955 220.155 363.285 220.485 ;
        RECT 362.955 218.795 363.285 219.125 ;
        RECT 362.955 217.435 363.285 217.765 ;
        RECT 362.955 216.075 363.285 216.405 ;
        RECT 362.955 214.715 363.285 215.045 ;
        RECT 362.955 213.355 363.285 213.685 ;
        RECT 362.955 211.995 363.285 212.325 ;
        RECT 362.955 210.635 363.285 210.965 ;
        RECT 362.955 209.275 363.285 209.605 ;
        RECT 362.955 207.915 363.285 208.245 ;
        RECT 362.955 206.555 363.285 206.885 ;
        RECT 362.955 205.195 363.285 205.525 ;
        RECT 362.955 203.835 363.285 204.165 ;
        RECT 362.955 202.475 363.285 202.805 ;
        RECT 362.955 201.115 363.285 201.445 ;
        RECT 362.955 199.755 363.285 200.085 ;
        RECT 362.955 198.395 363.285 198.725 ;
        RECT 362.955 197.035 363.285 197.365 ;
        RECT 362.955 195.675 363.285 196.005 ;
        RECT 362.955 194.315 363.285 194.645 ;
        RECT 362.955 192.955 363.285 193.285 ;
        RECT 362.955 191.595 363.285 191.925 ;
        RECT 362.955 190.235 363.285 190.565 ;
        RECT 362.955 188.875 363.285 189.205 ;
        RECT 362.955 187.515 363.285 187.845 ;
        RECT 362.955 186.155 363.285 186.485 ;
        RECT 362.955 184.795 363.285 185.125 ;
        RECT 362.955 183.435 363.285 183.765 ;
        RECT 362.955 182.075 363.285 182.405 ;
        RECT 362.955 180.715 363.285 181.045 ;
        RECT 362.955 179.355 363.285 179.685 ;
        RECT 362.955 177.995 363.285 178.325 ;
        RECT 362.955 176.635 363.285 176.965 ;
        RECT 362.955 175.275 363.285 175.605 ;
        RECT 362.955 173.915 363.285 174.245 ;
        RECT 362.955 172.555 363.285 172.885 ;
        RECT 362.955 171.195 363.285 171.525 ;
        RECT 362.955 169.835 363.285 170.165 ;
        RECT 362.955 168.475 363.285 168.805 ;
        RECT 362.955 167.115 363.285 167.445 ;
        RECT 362.955 165.755 363.285 166.085 ;
        RECT 362.955 164.395 363.285 164.725 ;
        RECT 362.955 163.035 363.285 163.365 ;
        RECT 362.955 161.675 363.285 162.005 ;
        RECT 362.955 160.315 363.285 160.645 ;
        RECT 362.955 158.955 363.285 159.285 ;
        RECT 362.955 157.595 363.285 157.925 ;
        RECT 362.955 156.235 363.285 156.565 ;
        RECT 362.955 154.875 363.285 155.205 ;
        RECT 362.955 153.515 363.285 153.845 ;
        RECT 362.955 152.155 363.285 152.485 ;
        RECT 362.955 150.795 363.285 151.125 ;
        RECT 362.955 149.435 363.285 149.765 ;
        RECT 362.955 148.075 363.285 148.405 ;
        RECT 362.955 146.715 363.285 147.045 ;
        RECT 362.955 145.355 363.285 145.685 ;
        RECT 362.955 143.995 363.285 144.325 ;
        RECT 362.955 142.635 363.285 142.965 ;
        RECT 362.955 141.275 363.285 141.605 ;
        RECT 362.955 139.915 363.285 140.245 ;
        RECT 362.955 138.555 363.285 138.885 ;
        RECT 362.955 137.195 363.285 137.525 ;
        RECT 362.955 135.835 363.285 136.165 ;
        RECT 362.955 134.475 363.285 134.805 ;
        RECT 362.955 133.115 363.285 133.445 ;
        RECT 362.955 131.755 363.285 132.085 ;
        RECT 362.955 130.395 363.285 130.725 ;
        RECT 362.955 129.035 363.285 129.365 ;
        RECT 362.955 127.675 363.285 128.005 ;
        RECT 362.955 126.315 363.285 126.645 ;
        RECT 362.955 124.955 363.285 125.285 ;
        RECT 362.955 123.595 363.285 123.925 ;
        RECT 362.955 122.235 363.285 122.565 ;
        RECT 362.955 120.875 363.285 121.205 ;
        RECT 362.955 119.515 363.285 119.845 ;
        RECT 362.955 118.155 363.285 118.485 ;
        RECT 362.955 116.795 363.285 117.125 ;
        RECT 362.955 115.435 363.285 115.765 ;
        RECT 362.955 114.075 363.285 114.405 ;
        RECT 362.955 112.715 363.285 113.045 ;
        RECT 362.955 111.355 363.285 111.685 ;
        RECT 362.955 109.995 363.285 110.325 ;
        RECT 362.955 108.635 363.285 108.965 ;
        RECT 362.955 107.275 363.285 107.605 ;
        RECT 362.955 105.915 363.285 106.245 ;
        RECT 362.955 104.555 363.285 104.885 ;
        RECT 362.955 103.195 363.285 103.525 ;
        RECT 362.955 101.835 363.285 102.165 ;
        RECT 362.955 100.475 363.285 100.805 ;
        RECT 362.955 99.115 363.285 99.445 ;
        RECT 362.955 97.755 363.285 98.085 ;
        RECT 362.955 96.395 363.285 96.725 ;
        RECT 362.955 95.035 363.285 95.365 ;
        RECT 362.955 93.675 363.285 94.005 ;
        RECT 362.955 92.315 363.285 92.645 ;
        RECT 362.955 90.955 363.285 91.285 ;
        RECT 362.955 89.595 363.285 89.925 ;
        RECT 362.955 88.235 363.285 88.565 ;
        RECT 362.955 86.875 363.285 87.205 ;
        RECT 362.955 85.515 363.285 85.845 ;
        RECT 362.955 84.155 363.285 84.485 ;
        RECT 362.955 82.795 363.285 83.125 ;
        RECT 362.955 81.435 363.285 81.765 ;
        RECT 362.955 80.075 363.285 80.405 ;
        RECT 362.955 78.715 363.285 79.045 ;
        RECT 362.955 77.355 363.285 77.685 ;
        RECT 362.955 75.995 363.285 76.325 ;
        RECT 362.955 74.635 363.285 74.965 ;
        RECT 362.955 73.275 363.285 73.605 ;
        RECT 362.955 71.915 363.285 72.245 ;
        RECT 362.955 70.555 363.285 70.885 ;
        RECT 362.955 69.195 363.285 69.525 ;
        RECT 362.955 67.835 363.285 68.165 ;
        RECT 362.955 66.475 363.285 66.805 ;
        RECT 362.955 65.115 363.285 65.445 ;
        RECT 362.955 63.755 363.285 64.085 ;
        RECT 362.955 62.395 363.285 62.725 ;
        RECT 362.955 61.035 363.285 61.365 ;
        RECT 362.955 59.675 363.285 60.005 ;
        RECT 362.955 58.315 363.285 58.645 ;
        RECT 362.955 56.955 363.285 57.285 ;
        RECT 362.955 55.595 363.285 55.925 ;
        RECT 362.955 54.235 363.285 54.565 ;
        RECT 362.955 52.875 363.285 53.205 ;
        RECT 362.955 51.515 363.285 51.845 ;
        RECT 362.955 50.155 363.285 50.485 ;
        RECT 362.955 48.795 363.285 49.125 ;
        RECT 362.955 47.435 363.285 47.765 ;
        RECT 362.955 46.075 363.285 46.405 ;
        RECT 362.955 44.715 363.285 45.045 ;
        RECT 362.955 43.355 363.285 43.685 ;
        RECT 362.955 41.995 363.285 42.325 ;
        RECT 362.955 40.635 363.285 40.965 ;
        RECT 362.955 39.275 363.285 39.605 ;
        RECT 362.955 37.915 363.285 38.245 ;
        RECT 362.955 36.555 363.285 36.885 ;
        RECT 362.955 35.195 363.285 35.525 ;
        RECT 362.955 33.835 363.285 34.165 ;
        RECT 362.955 32.475 363.285 32.805 ;
        RECT 362.955 31.115 363.285 31.445 ;
        RECT 362.955 29.755 363.285 30.085 ;
        RECT 362.955 28.395 363.285 28.725 ;
        RECT 362.955 27.035 363.285 27.365 ;
        RECT 362.955 25.675 363.285 26.005 ;
        RECT 362.955 24.315 363.285 24.645 ;
        RECT 362.955 22.955 363.285 23.285 ;
        RECT 362.955 21.595 363.285 21.925 ;
        RECT 362.955 20.235 363.285 20.565 ;
        RECT 362.955 18.875 363.285 19.205 ;
        RECT 362.955 17.515 363.285 17.845 ;
        RECT 362.955 16.155 363.285 16.485 ;
        RECT 362.955 14.795 363.285 15.125 ;
        RECT 362.955 13.435 363.285 13.765 ;
        RECT 362.955 12.075 363.285 12.405 ;
        RECT 362.955 10.715 363.285 11.045 ;
        RECT 362.955 9.355 363.285 9.685 ;
        RECT 362.955 7.995 363.285 8.325 ;
        RECT 362.955 6.635 363.285 6.965 ;
        RECT 362.955 5.275 363.285 5.605 ;
        RECT 362.955 3.915 363.285 4.245 ;
        RECT 362.955 2.555 363.285 2.885 ;
        RECT 362.955 1.195 363.285 1.525 ;
        RECT 362.955 -0.165 363.285 0.165 ;
        RECT 362.955 -1.525 363.285 -1.195 ;
        RECT 362.955 -2.885 363.285 -2.555 ;
        RECT 362.955 -4.245 363.285 -3.915 ;
        RECT 362.955 -5.605 363.285 -5.275 ;
        RECT 362.955 -6.965 363.285 -6.635 ;
        RECT 362.955 -8.325 363.285 -7.995 ;
        RECT 362.955 -9.685 363.285 -9.355 ;
        RECT 362.955 -11.045 363.285 -10.715 ;
        RECT 362.955 -12.405 363.285 -12.075 ;
        RECT 362.955 -13.765 363.285 -13.435 ;
        RECT 362.955 -15.125 363.285 -14.795 ;
        RECT 362.955 -16.485 363.285 -16.155 ;
        RECT 362.955 -17.845 363.285 -17.515 ;
        RECT 362.955 -19.205 363.285 -18.875 ;
        RECT 362.955 -20.565 363.285 -20.235 ;
        RECT 362.955 -21.925 363.285 -21.595 ;
        RECT 362.955 -23.285 363.285 -22.955 ;
        RECT 362.955 -24.645 363.285 -24.315 ;
        RECT 362.955 -26.005 363.285 -25.675 ;
        RECT 362.955 -27.365 363.285 -27.035 ;
        RECT 362.955 -28.725 363.285 -28.395 ;
        RECT 362.955 -30.085 363.285 -29.755 ;
        RECT 362.955 -31.445 363.285 -31.115 ;
        RECT 362.955 -32.805 363.285 -32.475 ;
        RECT 362.955 -34.165 363.285 -33.835 ;
        RECT 362.955 -35.525 363.285 -35.195 ;
        RECT 362.955 -36.885 363.285 -36.555 ;
        RECT 362.955 -38.245 363.285 -37.915 ;
        RECT 362.955 -39.605 363.285 -39.275 ;
        RECT 362.955 -40.965 363.285 -40.635 ;
        RECT 362.955 -42.325 363.285 -41.995 ;
        RECT 362.955 -43.685 363.285 -43.355 ;
        RECT 362.955 -45.045 363.285 -44.715 ;
        RECT 362.955 -46.405 363.285 -46.075 ;
        RECT 362.955 -47.765 363.285 -47.435 ;
        RECT 362.955 -49.125 363.285 -48.795 ;
        RECT 362.955 -50.485 363.285 -50.155 ;
        RECT 362.955 -51.845 363.285 -51.515 ;
        RECT 362.955 -53.205 363.285 -52.875 ;
        RECT 362.955 -54.565 363.285 -54.235 ;
        RECT 362.955 -55.925 363.285 -55.595 ;
        RECT 362.955 -57.285 363.285 -56.955 ;
        RECT 362.955 -58.645 363.285 -58.315 ;
        RECT 362.955 -60.005 363.285 -59.675 ;
        RECT 362.955 -61.365 363.285 -61.035 ;
        RECT 362.955 -62.725 363.285 -62.395 ;
        RECT 362.955 -64.085 363.285 -63.755 ;
        RECT 362.955 -65.445 363.285 -65.115 ;
        RECT 362.955 -66.805 363.285 -66.475 ;
        RECT 362.955 -68.165 363.285 -67.835 ;
        RECT 362.955 -69.525 363.285 -69.195 ;
        RECT 362.955 -70.885 363.285 -70.555 ;
        RECT 362.955 -72.245 363.285 -71.915 ;
        RECT 362.955 -73.605 363.285 -73.275 ;
        RECT 362.955 -74.965 363.285 -74.635 ;
        RECT 362.955 -76.325 363.285 -75.995 ;
        RECT 362.955 -77.685 363.285 -77.355 ;
        RECT 362.955 -79.045 363.285 -78.715 ;
        RECT 362.955 -80.405 363.285 -80.075 ;
        RECT 362.955 -81.765 363.285 -81.435 ;
        RECT 362.955 -83.125 363.285 -82.795 ;
        RECT 362.955 -84.485 363.285 -84.155 ;
        RECT 362.955 -85.845 363.285 -85.515 ;
        RECT 362.955 -87.205 363.285 -86.875 ;
        RECT 362.955 -88.565 363.285 -88.235 ;
        RECT 362.955 -89.925 363.285 -89.595 ;
        RECT 362.955 -91.285 363.285 -90.955 ;
        RECT 362.955 -92.645 363.285 -92.315 ;
        RECT 362.955 -94.005 363.285 -93.675 ;
        RECT 362.955 -95.365 363.285 -95.035 ;
        RECT 362.955 -96.725 363.285 -96.395 ;
        RECT 362.955 -98.085 363.285 -97.755 ;
        RECT 362.955 -99.445 363.285 -99.115 ;
        RECT 362.955 -100.805 363.285 -100.475 ;
        RECT 362.955 -102.165 363.285 -101.835 ;
        RECT 362.955 -103.525 363.285 -103.195 ;
        RECT 362.955 -104.885 363.285 -104.555 ;
        RECT 362.955 -106.245 363.285 -105.915 ;
        RECT 362.955 -107.605 363.285 -107.275 ;
        RECT 362.955 -108.965 363.285 -108.635 ;
        RECT 362.955 -110.325 363.285 -109.995 ;
        RECT 362.955 -111.685 363.285 -111.355 ;
        RECT 362.955 -113.045 363.285 -112.715 ;
        RECT 362.955 -114.405 363.285 -114.075 ;
        RECT 362.955 -115.765 363.285 -115.435 ;
        RECT 362.955 -117.125 363.285 -116.795 ;
        RECT 362.955 -118.485 363.285 -118.155 ;
        RECT 362.955 -119.845 363.285 -119.515 ;
        RECT 362.955 -121.205 363.285 -120.875 ;
        RECT 362.955 -122.565 363.285 -122.235 ;
        RECT 362.955 -123.925 363.285 -123.595 ;
        RECT 362.955 -125.285 363.285 -124.955 ;
        RECT 362.955 -126.645 363.285 -126.315 ;
        RECT 362.955 -128.005 363.285 -127.675 ;
        RECT 362.955 -129.365 363.285 -129.035 ;
        RECT 362.955 -130.725 363.285 -130.395 ;
        RECT 362.955 -132.085 363.285 -131.755 ;
        RECT 362.955 -133.445 363.285 -133.115 ;
        RECT 362.955 -134.805 363.285 -134.475 ;
        RECT 362.955 -136.165 363.285 -135.835 ;
        RECT 362.955 -137.525 363.285 -137.195 ;
        RECT 362.955 -138.885 363.285 -138.555 ;
        RECT 362.955 -140.245 363.285 -139.915 ;
        RECT 362.955 -141.605 363.285 -141.275 ;
        RECT 362.955 -142.965 363.285 -142.635 ;
        RECT 362.955 -144.325 363.285 -143.995 ;
        RECT 362.955 -145.685 363.285 -145.355 ;
        RECT 362.955 -147.045 363.285 -146.715 ;
        RECT 362.955 -148.405 363.285 -148.075 ;
        RECT 362.955 -149.765 363.285 -149.435 ;
        RECT 362.955 -151.125 363.285 -150.795 ;
        RECT 362.955 -152.485 363.285 -152.155 ;
        RECT 362.955 -153.845 363.285 -153.515 ;
        RECT 362.955 -155.205 363.285 -154.875 ;
        RECT 362.955 -156.565 363.285 -156.235 ;
        RECT 362.955 -157.925 363.285 -157.595 ;
        RECT 362.955 -159.285 363.285 -158.955 ;
        RECT 362.955 -160.645 363.285 -160.315 ;
        RECT 362.955 -162.005 363.285 -161.675 ;
        RECT 362.955 -163.365 363.285 -163.035 ;
        RECT 362.955 -164.725 363.285 -164.395 ;
        RECT 362.955 -166.085 363.285 -165.755 ;
        RECT 362.955 -167.445 363.285 -167.115 ;
        RECT 362.955 -168.805 363.285 -168.475 ;
        RECT 362.955 -170.165 363.285 -169.835 ;
        RECT 362.955 -171.525 363.285 -171.195 ;
        RECT 362.955 -172.885 363.285 -172.555 ;
        RECT 362.955 -174.245 363.285 -173.915 ;
        RECT 362.955 -175.605 363.285 -175.275 ;
        RECT 362.955 -176.965 363.285 -176.635 ;
        RECT 362.955 -178.325 363.285 -177.995 ;
        RECT 362.955 -179.685 363.285 -179.355 ;
        RECT 362.955 -181.045 363.285 -180.715 ;
        RECT 362.955 -182.405 363.285 -182.075 ;
        RECT 362.955 -183.765 363.285 -183.435 ;
        RECT 362.955 -185.125 363.285 -184.795 ;
        RECT 362.955 -186.485 363.285 -186.155 ;
        RECT 362.955 -187.845 363.285 -187.515 ;
        RECT 362.955 -189.205 363.285 -188.875 ;
        RECT 362.955 -190.565 363.285 -190.235 ;
        RECT 362.955 -191.925 363.285 -191.595 ;
        RECT 362.955 -193.285 363.285 -192.955 ;
        RECT 362.955 -194.645 363.285 -194.315 ;
        RECT 362.955 -196.005 363.285 -195.675 ;
        RECT 362.955 -197.365 363.285 -197.035 ;
        RECT 362.955 -198.725 363.285 -198.395 ;
        RECT 362.955 -200.085 363.285 -199.755 ;
        RECT 362.955 -201.445 363.285 -201.115 ;
        RECT 362.955 -202.805 363.285 -202.475 ;
        RECT 362.955 -204.165 363.285 -203.835 ;
        RECT 362.955 -205.525 363.285 -205.195 ;
        RECT 362.955 -206.885 363.285 -206.555 ;
        RECT 362.955 -208.245 363.285 -207.915 ;
        RECT 362.955 -209.605 363.285 -209.275 ;
        RECT 362.955 -210.965 363.285 -210.635 ;
        RECT 362.955 -212.325 363.285 -211.995 ;
        RECT 362.955 -213.685 363.285 -213.355 ;
        RECT 362.955 -215.045 363.285 -214.715 ;
        RECT 362.955 -216.405 363.285 -216.075 ;
        RECT 362.955 -217.765 363.285 -217.435 ;
        RECT 362.955 -219.125 363.285 -218.795 ;
        RECT 362.955 -220.485 363.285 -220.155 ;
        RECT 362.955 -221.845 363.285 -221.515 ;
        RECT 362.955 -223.205 363.285 -222.875 ;
        RECT 362.955 -224.565 363.285 -224.235 ;
        RECT 362.955 -225.925 363.285 -225.595 ;
        RECT 362.955 -227.285 363.285 -226.955 ;
        RECT 362.955 -228.645 363.285 -228.315 ;
        RECT 362.955 -230.005 363.285 -229.675 ;
        RECT 362.955 -231.365 363.285 -231.035 ;
        RECT 362.955 -232.725 363.285 -232.395 ;
        RECT 362.955 -234.085 363.285 -233.755 ;
        RECT 362.955 -235.445 363.285 -235.115 ;
        RECT 362.955 -236.805 363.285 -236.475 ;
        RECT 362.955 -238.165 363.285 -237.835 ;
        RECT 362.955 -243.81 363.285 -242.68 ;
        RECT 362.96 -243.925 363.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.515 246.76 357.845 247.89 ;
        RECT 357.515 241.915 357.845 242.245 ;
        RECT 357.515 240.555 357.845 240.885 ;
        RECT 357.515 239.195 357.845 239.525 ;
        RECT 357.515 237.835 357.845 238.165 ;
        RECT 357.515 235.17 357.845 235.5 ;
        RECT 357.515 232.995 357.845 233.325 ;
        RECT 357.515 231.415 357.845 231.745 ;
        RECT 357.515 230.565 357.845 230.895 ;
        RECT 357.515 228.255 357.845 228.585 ;
        RECT 357.515 227.405 357.845 227.735 ;
        RECT 357.515 225.095 357.845 225.425 ;
        RECT 357.515 224.245 357.845 224.575 ;
        RECT 357.515 221.935 357.845 222.265 ;
        RECT 357.515 221.085 357.845 221.415 ;
        RECT 357.515 218.775 357.845 219.105 ;
        RECT 357.515 217.195 357.845 217.525 ;
        RECT 357.515 216.345 357.845 216.675 ;
        RECT 357.515 214.035 357.845 214.365 ;
        RECT 357.515 213.185 357.845 213.515 ;
        RECT 357.515 210.875 357.845 211.205 ;
        RECT 357.515 210.025 357.845 210.355 ;
        RECT 357.515 207.715 357.845 208.045 ;
        RECT 357.515 206.865 357.845 207.195 ;
        RECT 357.515 204.555 357.845 204.885 ;
        RECT 357.515 202.975 357.845 203.305 ;
        RECT 357.515 202.125 357.845 202.455 ;
        RECT 357.515 199.815 357.845 200.145 ;
        RECT 357.515 198.965 357.845 199.295 ;
        RECT 357.515 196.655 357.845 196.985 ;
        RECT 357.515 195.805 357.845 196.135 ;
        RECT 357.515 193.495 357.845 193.825 ;
        RECT 357.515 192.645 357.845 192.975 ;
        RECT 357.515 190.335 357.845 190.665 ;
        RECT 357.515 188.755 357.845 189.085 ;
        RECT 357.515 187.905 357.845 188.235 ;
        RECT 357.515 185.595 357.845 185.925 ;
        RECT 357.515 184.745 357.845 185.075 ;
        RECT 357.515 182.435 357.845 182.765 ;
        RECT 357.515 181.585 357.845 181.915 ;
        RECT 357.515 179.275 357.845 179.605 ;
        RECT 357.515 178.425 357.845 178.755 ;
        RECT 357.515 176.115 357.845 176.445 ;
        RECT 357.515 174.535 357.845 174.865 ;
        RECT 357.515 173.685 357.845 174.015 ;
        RECT 357.515 171.375 357.845 171.705 ;
        RECT 357.515 170.525 357.845 170.855 ;
        RECT 357.515 168.215 357.845 168.545 ;
        RECT 357.515 167.365 357.845 167.695 ;
        RECT 357.515 165.055 357.845 165.385 ;
        RECT 357.515 164.205 357.845 164.535 ;
        RECT 357.515 161.895 357.845 162.225 ;
        RECT 357.515 160.315 357.845 160.645 ;
        RECT 357.515 159.465 357.845 159.795 ;
        RECT 357.515 157.155 357.845 157.485 ;
        RECT 357.515 156.305 357.845 156.635 ;
        RECT 357.515 153.995 357.845 154.325 ;
        RECT 357.515 153.145 357.845 153.475 ;
        RECT 357.515 150.835 357.845 151.165 ;
        RECT 357.515 149.985 357.845 150.315 ;
        RECT 357.515 147.675 357.845 148.005 ;
        RECT 357.515 146.095 357.845 146.425 ;
        RECT 357.515 145.245 357.845 145.575 ;
        RECT 357.515 142.935 357.845 143.265 ;
        RECT 357.515 142.085 357.845 142.415 ;
        RECT 357.515 139.775 357.845 140.105 ;
        RECT 357.515 138.925 357.845 139.255 ;
        RECT 357.515 136.615 357.845 136.945 ;
        RECT 357.515 135.765 357.845 136.095 ;
        RECT 357.515 133.455 357.845 133.785 ;
        RECT 357.515 131.875 357.845 132.205 ;
        RECT 357.515 131.025 357.845 131.355 ;
        RECT 357.515 128.715 357.845 129.045 ;
        RECT 357.515 127.865 357.845 128.195 ;
        RECT 357.515 125.555 357.845 125.885 ;
        RECT 357.515 124.705 357.845 125.035 ;
        RECT 357.515 122.395 357.845 122.725 ;
        RECT 357.515 121.545 357.845 121.875 ;
        RECT 357.515 119.235 357.845 119.565 ;
        RECT 357.515 117.655 357.845 117.985 ;
        RECT 357.515 116.805 357.845 117.135 ;
        RECT 357.515 114.495 357.845 114.825 ;
        RECT 357.515 113.645 357.845 113.975 ;
        RECT 357.515 111.335 357.845 111.665 ;
        RECT 357.515 110.485 357.845 110.815 ;
        RECT 357.515 108.175 357.845 108.505 ;
        RECT 357.515 107.325 357.845 107.655 ;
        RECT 357.515 105.015 357.845 105.345 ;
        RECT 357.515 103.435 357.845 103.765 ;
        RECT 357.515 102.585 357.845 102.915 ;
        RECT 357.515 100.275 357.845 100.605 ;
        RECT 357.515 99.425 357.845 99.755 ;
        RECT 357.515 97.115 357.845 97.445 ;
        RECT 357.515 96.265 357.845 96.595 ;
        RECT 357.515 93.955 357.845 94.285 ;
        RECT 357.515 93.105 357.845 93.435 ;
        RECT 357.515 90.795 357.845 91.125 ;
        RECT 357.515 89.215 357.845 89.545 ;
        RECT 357.515 88.365 357.845 88.695 ;
        RECT 357.515 86.055 357.845 86.385 ;
        RECT 357.515 85.205 357.845 85.535 ;
        RECT 357.515 82.895 357.845 83.225 ;
        RECT 357.515 82.045 357.845 82.375 ;
        RECT 357.515 79.735 357.845 80.065 ;
        RECT 357.515 78.885 357.845 79.215 ;
        RECT 357.515 76.575 357.845 76.905 ;
        RECT 357.515 74.995 357.845 75.325 ;
        RECT 357.515 74.145 357.845 74.475 ;
        RECT 357.515 71.835 357.845 72.165 ;
        RECT 357.515 70.985 357.845 71.315 ;
        RECT 357.515 68.675 357.845 69.005 ;
        RECT 357.515 67.825 357.845 68.155 ;
        RECT 357.515 65.515 357.845 65.845 ;
        RECT 357.515 64.665 357.845 64.995 ;
        RECT 357.515 62.355 357.845 62.685 ;
        RECT 357.515 60.775 357.845 61.105 ;
        RECT 357.515 59.925 357.845 60.255 ;
        RECT 357.515 57.615 357.845 57.945 ;
        RECT 357.515 56.765 357.845 57.095 ;
        RECT 357.515 54.455 357.845 54.785 ;
        RECT 357.515 53.605 357.845 53.935 ;
        RECT 357.515 51.295 357.845 51.625 ;
        RECT 357.515 50.445 357.845 50.775 ;
        RECT 357.515 48.135 357.845 48.465 ;
        RECT 357.515 46.555 357.845 46.885 ;
        RECT 357.515 45.705 357.845 46.035 ;
        RECT 357.515 43.395 357.845 43.725 ;
        RECT 357.515 42.545 357.845 42.875 ;
        RECT 357.515 40.235 357.845 40.565 ;
        RECT 357.515 39.385 357.845 39.715 ;
        RECT 357.515 37.075 357.845 37.405 ;
        RECT 357.515 36.225 357.845 36.555 ;
        RECT 357.515 33.915 357.845 34.245 ;
        RECT 357.515 32.335 357.845 32.665 ;
        RECT 357.515 31.485 357.845 31.815 ;
        RECT 357.515 29.175 357.845 29.505 ;
        RECT 357.515 28.325 357.845 28.655 ;
        RECT 357.515 26.015 357.845 26.345 ;
        RECT 357.515 25.165 357.845 25.495 ;
        RECT 357.515 22.855 357.845 23.185 ;
        RECT 357.515 22.005 357.845 22.335 ;
        RECT 357.515 19.695 357.845 20.025 ;
        RECT 357.515 18.115 357.845 18.445 ;
        RECT 357.515 17.265 357.845 17.595 ;
        RECT 357.515 14.955 357.845 15.285 ;
        RECT 357.515 14.105 357.845 14.435 ;
        RECT 357.515 11.795 357.845 12.125 ;
        RECT 357.515 10.945 357.845 11.275 ;
        RECT 357.515 8.635 357.845 8.965 ;
        RECT 357.515 7.785 357.845 8.115 ;
        RECT 357.515 5.475 357.845 5.805 ;
        RECT 357.515 3.895 357.845 4.225 ;
        RECT 357.515 3.045 357.845 3.375 ;
        RECT 357.515 0.87 357.845 1.2 ;
        RECT 357.515 -1.525 357.845 -1.195 ;
        RECT 357.515 -2.885 357.845 -2.555 ;
        RECT 357.515 -4.245 357.845 -3.915 ;
        RECT 357.515 -5.605 357.845 -5.275 ;
        RECT 357.515 -6.965 357.845 -6.635 ;
        RECT 357.515 -8.325 357.845 -7.995 ;
        RECT 357.515 -9.685 357.845 -9.355 ;
        RECT 357.515 -11.045 357.845 -10.715 ;
        RECT 357.515 -12.405 357.845 -12.075 ;
        RECT 357.515 -13.765 357.845 -13.435 ;
        RECT 357.515 -15.125 357.845 -14.795 ;
        RECT 357.515 -16.485 357.845 -16.155 ;
        RECT 357.515 -17.845 357.845 -17.515 ;
        RECT 357.515 -19.205 357.845 -18.875 ;
        RECT 357.515 -20.565 357.845 -20.235 ;
        RECT 357.515 -21.925 357.845 -21.595 ;
        RECT 357.515 -23.285 357.845 -22.955 ;
        RECT 357.515 -24.645 357.845 -24.315 ;
        RECT 357.515 -26.005 357.845 -25.675 ;
        RECT 357.515 -27.365 357.845 -27.035 ;
        RECT 357.515 -28.725 357.845 -28.395 ;
        RECT 357.515 -30.085 357.845 -29.755 ;
        RECT 357.515 -31.445 357.845 -31.115 ;
        RECT 357.515 -32.805 357.845 -32.475 ;
        RECT 357.515 -34.165 357.845 -33.835 ;
        RECT 357.515 -35.525 357.845 -35.195 ;
        RECT 357.515 -36.885 357.845 -36.555 ;
        RECT 357.515 -38.245 357.845 -37.915 ;
        RECT 357.515 -39.605 357.845 -39.275 ;
        RECT 357.515 -40.965 357.845 -40.635 ;
        RECT 357.515 -42.325 357.845 -41.995 ;
        RECT 357.515 -43.685 357.845 -43.355 ;
        RECT 357.515 -45.045 357.845 -44.715 ;
        RECT 357.515 -46.405 357.845 -46.075 ;
        RECT 357.515 -47.765 357.845 -47.435 ;
        RECT 357.515 -49.125 357.845 -48.795 ;
        RECT 357.515 -50.485 357.845 -50.155 ;
        RECT 357.515 -51.845 357.845 -51.515 ;
        RECT 357.515 -53.205 357.845 -52.875 ;
        RECT 357.515 -54.565 357.845 -54.235 ;
        RECT 357.515 -55.925 357.845 -55.595 ;
        RECT 357.515 -57.285 357.845 -56.955 ;
        RECT 357.515 -58.645 357.845 -58.315 ;
        RECT 357.515 -60.005 357.845 -59.675 ;
        RECT 357.515 -61.365 357.845 -61.035 ;
        RECT 357.515 -62.725 357.845 -62.395 ;
        RECT 357.515 -64.085 357.845 -63.755 ;
        RECT 357.515 -65.445 357.845 -65.115 ;
        RECT 357.515 -66.805 357.845 -66.475 ;
        RECT 357.515 -68.165 357.845 -67.835 ;
        RECT 357.515 -69.525 357.845 -69.195 ;
        RECT 357.515 -70.885 357.845 -70.555 ;
        RECT 357.515 -72.245 357.845 -71.915 ;
        RECT 357.515 -73.605 357.845 -73.275 ;
        RECT 357.515 -74.965 357.845 -74.635 ;
        RECT 357.515 -76.325 357.845 -75.995 ;
        RECT 357.515 -77.685 357.845 -77.355 ;
        RECT 357.515 -79.045 357.845 -78.715 ;
        RECT 357.515 -80.405 357.845 -80.075 ;
        RECT 357.515 -81.765 357.845 -81.435 ;
        RECT 357.515 -83.125 357.845 -82.795 ;
        RECT 357.515 -84.485 357.845 -84.155 ;
        RECT 357.515 -85.845 357.845 -85.515 ;
        RECT 357.515 -87.205 357.845 -86.875 ;
        RECT 357.515 -88.565 357.845 -88.235 ;
        RECT 357.515 -89.925 357.845 -89.595 ;
        RECT 357.515 -91.285 357.845 -90.955 ;
        RECT 357.515 -92.645 357.845 -92.315 ;
        RECT 357.515 -94.005 357.845 -93.675 ;
        RECT 357.515 -95.365 357.845 -95.035 ;
        RECT 357.515 -96.725 357.845 -96.395 ;
        RECT 357.515 -98.085 357.845 -97.755 ;
        RECT 357.515 -99.445 357.845 -99.115 ;
        RECT 357.515 -100.805 357.845 -100.475 ;
        RECT 357.515 -102.165 357.845 -101.835 ;
        RECT 357.515 -103.525 357.845 -103.195 ;
        RECT 357.515 -104.885 357.845 -104.555 ;
        RECT 357.515 -106.245 357.845 -105.915 ;
        RECT 357.515 -107.605 357.845 -107.275 ;
        RECT 357.515 -108.965 357.845 -108.635 ;
        RECT 357.515 -110.325 357.845 -109.995 ;
        RECT 357.515 -111.685 357.845 -111.355 ;
        RECT 357.515 -113.045 357.845 -112.715 ;
        RECT 357.515 -114.405 357.845 -114.075 ;
        RECT 357.515 -115.765 357.845 -115.435 ;
        RECT 357.515 -117.125 357.845 -116.795 ;
        RECT 357.515 -118.485 357.845 -118.155 ;
        RECT 357.515 -119.845 357.845 -119.515 ;
        RECT 357.515 -121.205 357.845 -120.875 ;
        RECT 357.515 -122.565 357.845 -122.235 ;
        RECT 357.515 -123.925 357.845 -123.595 ;
        RECT 357.515 -125.285 357.845 -124.955 ;
        RECT 357.515 -126.645 357.845 -126.315 ;
        RECT 357.515 -128.005 357.845 -127.675 ;
        RECT 357.515 -129.365 357.845 -129.035 ;
        RECT 357.515 -130.725 357.845 -130.395 ;
        RECT 357.515 -132.085 357.845 -131.755 ;
        RECT 357.515 -133.445 357.845 -133.115 ;
        RECT 357.515 -134.805 357.845 -134.475 ;
        RECT 357.515 -136.165 357.845 -135.835 ;
        RECT 357.515 -137.525 357.845 -137.195 ;
        RECT 357.515 -138.885 357.845 -138.555 ;
        RECT 357.515 -140.245 357.845 -139.915 ;
        RECT 357.515 -141.605 357.845 -141.275 ;
        RECT 357.515 -142.965 357.845 -142.635 ;
        RECT 357.515 -144.325 357.845 -143.995 ;
        RECT 357.515 -145.685 357.845 -145.355 ;
        RECT 357.515 -147.045 357.845 -146.715 ;
        RECT 357.515 -148.405 357.845 -148.075 ;
        RECT 357.515 -149.765 357.845 -149.435 ;
        RECT 357.515 -151.125 357.845 -150.795 ;
        RECT 357.515 -152.485 357.845 -152.155 ;
        RECT 357.515 -153.845 357.845 -153.515 ;
        RECT 357.515 -155.205 357.845 -154.875 ;
        RECT 357.515 -156.565 357.845 -156.235 ;
        RECT 357.515 -157.925 357.845 -157.595 ;
        RECT 357.515 -159.285 357.845 -158.955 ;
        RECT 357.515 -160.645 357.845 -160.315 ;
        RECT 357.515 -162.005 357.845 -161.675 ;
        RECT 357.515 -163.365 357.845 -163.035 ;
        RECT 357.515 -164.725 357.845 -164.395 ;
        RECT 357.515 -166.085 357.845 -165.755 ;
        RECT 357.515 -167.445 357.845 -167.115 ;
        RECT 357.515 -168.805 357.845 -168.475 ;
        RECT 357.515 -170.165 357.845 -169.835 ;
        RECT 357.515 -171.525 357.845 -171.195 ;
        RECT 357.515 -172.885 357.845 -172.555 ;
        RECT 357.515 -174.245 357.845 -173.915 ;
        RECT 357.515 -175.605 357.845 -175.275 ;
        RECT 357.515 -176.965 357.845 -176.635 ;
        RECT 357.515 -178.325 357.845 -177.995 ;
        RECT 357.515 -179.685 357.845 -179.355 ;
        RECT 357.515 -181.045 357.845 -180.715 ;
        RECT 357.515 -182.405 357.845 -182.075 ;
        RECT 357.515 -183.765 357.845 -183.435 ;
        RECT 357.515 -185.125 357.845 -184.795 ;
        RECT 357.515 -186.485 357.845 -186.155 ;
        RECT 357.515 -187.845 357.845 -187.515 ;
        RECT 357.515 -189.205 357.845 -188.875 ;
        RECT 357.515 -190.565 357.845 -190.235 ;
        RECT 357.515 -191.925 357.845 -191.595 ;
        RECT 357.515 -193.285 357.845 -192.955 ;
        RECT 357.515 -194.645 357.845 -194.315 ;
        RECT 357.515 -196.005 357.845 -195.675 ;
        RECT 357.515 -197.365 357.845 -197.035 ;
        RECT 357.515 -198.725 357.845 -198.395 ;
        RECT 357.515 -200.085 357.845 -199.755 ;
        RECT 357.515 -201.445 357.845 -201.115 ;
        RECT 357.515 -202.805 357.845 -202.475 ;
        RECT 357.515 -204.165 357.845 -203.835 ;
        RECT 357.515 -205.525 357.845 -205.195 ;
        RECT 357.515 -206.885 357.845 -206.555 ;
        RECT 357.515 -208.245 357.845 -207.915 ;
        RECT 357.515 -209.605 357.845 -209.275 ;
        RECT 357.515 -210.965 357.845 -210.635 ;
        RECT 357.515 -212.325 357.845 -211.995 ;
        RECT 357.515 -213.685 357.845 -213.355 ;
        RECT 357.515 -215.045 357.845 -214.715 ;
        RECT 357.515 -216.405 357.845 -216.075 ;
        RECT 357.515 -217.765 357.845 -217.435 ;
        RECT 357.515 -219.125 357.845 -218.795 ;
        RECT 357.515 -220.485 357.845 -220.155 ;
        RECT 357.515 -221.845 357.845 -221.515 ;
        RECT 357.515 -223.205 357.845 -222.875 ;
        RECT 357.515 -224.565 357.845 -224.235 ;
        RECT 357.515 -225.925 357.845 -225.595 ;
        RECT 357.515 -227.285 357.845 -226.955 ;
        RECT 357.515 -228.645 357.845 -228.315 ;
        RECT 357.515 -230.005 357.845 -229.675 ;
        RECT 357.515 -231.365 357.845 -231.035 ;
        RECT 357.515 -232.725 357.845 -232.395 ;
        RECT 357.515 -234.085 357.845 -233.755 ;
        RECT 357.515 -235.445 357.845 -235.115 ;
        RECT 357.515 -236.805 357.845 -236.475 ;
        RECT 357.515 -238.165 357.845 -237.835 ;
        RECT 357.515 -243.81 357.845 -242.68 ;
        RECT 357.52 -243.925 357.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.875 246.76 359.205 247.89 ;
        RECT 358.875 241.915 359.205 242.245 ;
        RECT 358.875 240.555 359.205 240.885 ;
        RECT 358.875 239.195 359.205 239.525 ;
        RECT 358.875 237.835 359.205 238.165 ;
        RECT 358.875 235.17 359.205 235.5 ;
        RECT 358.875 232.995 359.205 233.325 ;
        RECT 358.875 231.415 359.205 231.745 ;
        RECT 358.875 230.565 359.205 230.895 ;
        RECT 358.875 228.255 359.205 228.585 ;
        RECT 358.875 227.405 359.205 227.735 ;
        RECT 358.875 225.095 359.205 225.425 ;
        RECT 358.875 224.245 359.205 224.575 ;
        RECT 358.875 221.935 359.205 222.265 ;
        RECT 358.875 221.085 359.205 221.415 ;
        RECT 358.875 218.775 359.205 219.105 ;
        RECT 358.875 217.195 359.205 217.525 ;
        RECT 358.875 216.345 359.205 216.675 ;
        RECT 358.875 214.035 359.205 214.365 ;
        RECT 358.875 213.185 359.205 213.515 ;
        RECT 358.875 210.875 359.205 211.205 ;
        RECT 358.875 210.025 359.205 210.355 ;
        RECT 358.875 207.715 359.205 208.045 ;
        RECT 358.875 206.865 359.205 207.195 ;
        RECT 358.875 204.555 359.205 204.885 ;
        RECT 358.875 202.975 359.205 203.305 ;
        RECT 358.875 202.125 359.205 202.455 ;
        RECT 358.875 199.815 359.205 200.145 ;
        RECT 358.875 198.965 359.205 199.295 ;
        RECT 358.875 196.655 359.205 196.985 ;
        RECT 358.875 195.805 359.205 196.135 ;
        RECT 358.875 193.495 359.205 193.825 ;
        RECT 358.875 192.645 359.205 192.975 ;
        RECT 358.875 190.335 359.205 190.665 ;
        RECT 358.875 188.755 359.205 189.085 ;
        RECT 358.875 187.905 359.205 188.235 ;
        RECT 358.875 185.595 359.205 185.925 ;
        RECT 358.875 184.745 359.205 185.075 ;
        RECT 358.875 182.435 359.205 182.765 ;
        RECT 358.875 181.585 359.205 181.915 ;
        RECT 358.875 179.275 359.205 179.605 ;
        RECT 358.875 178.425 359.205 178.755 ;
        RECT 358.875 176.115 359.205 176.445 ;
        RECT 358.875 174.535 359.205 174.865 ;
        RECT 358.875 173.685 359.205 174.015 ;
        RECT 358.875 171.375 359.205 171.705 ;
        RECT 358.875 170.525 359.205 170.855 ;
        RECT 358.875 168.215 359.205 168.545 ;
        RECT 358.875 167.365 359.205 167.695 ;
        RECT 358.875 165.055 359.205 165.385 ;
        RECT 358.875 164.205 359.205 164.535 ;
        RECT 358.875 161.895 359.205 162.225 ;
        RECT 358.875 160.315 359.205 160.645 ;
        RECT 358.875 159.465 359.205 159.795 ;
        RECT 358.875 157.155 359.205 157.485 ;
        RECT 358.875 156.305 359.205 156.635 ;
        RECT 358.875 153.995 359.205 154.325 ;
        RECT 358.875 153.145 359.205 153.475 ;
        RECT 358.875 150.835 359.205 151.165 ;
        RECT 358.875 149.985 359.205 150.315 ;
        RECT 358.875 147.675 359.205 148.005 ;
        RECT 358.875 146.095 359.205 146.425 ;
        RECT 358.875 145.245 359.205 145.575 ;
        RECT 358.875 142.935 359.205 143.265 ;
        RECT 358.875 142.085 359.205 142.415 ;
        RECT 358.875 139.775 359.205 140.105 ;
        RECT 358.875 138.925 359.205 139.255 ;
        RECT 358.875 136.615 359.205 136.945 ;
        RECT 358.875 135.765 359.205 136.095 ;
        RECT 358.875 133.455 359.205 133.785 ;
        RECT 358.875 131.875 359.205 132.205 ;
        RECT 358.875 131.025 359.205 131.355 ;
        RECT 358.875 128.715 359.205 129.045 ;
        RECT 358.875 127.865 359.205 128.195 ;
        RECT 358.875 125.555 359.205 125.885 ;
        RECT 358.875 124.705 359.205 125.035 ;
        RECT 358.875 122.395 359.205 122.725 ;
        RECT 358.875 121.545 359.205 121.875 ;
        RECT 358.875 119.235 359.205 119.565 ;
        RECT 358.875 117.655 359.205 117.985 ;
        RECT 358.875 116.805 359.205 117.135 ;
        RECT 358.875 114.495 359.205 114.825 ;
        RECT 358.875 113.645 359.205 113.975 ;
        RECT 358.875 111.335 359.205 111.665 ;
        RECT 358.875 110.485 359.205 110.815 ;
        RECT 358.875 108.175 359.205 108.505 ;
        RECT 358.875 107.325 359.205 107.655 ;
        RECT 358.875 105.015 359.205 105.345 ;
        RECT 358.875 103.435 359.205 103.765 ;
        RECT 358.875 102.585 359.205 102.915 ;
        RECT 358.875 100.275 359.205 100.605 ;
        RECT 358.875 99.425 359.205 99.755 ;
        RECT 358.875 97.115 359.205 97.445 ;
        RECT 358.875 96.265 359.205 96.595 ;
        RECT 358.875 93.955 359.205 94.285 ;
        RECT 358.875 93.105 359.205 93.435 ;
        RECT 358.875 90.795 359.205 91.125 ;
        RECT 358.875 89.215 359.205 89.545 ;
        RECT 358.875 88.365 359.205 88.695 ;
        RECT 358.875 86.055 359.205 86.385 ;
        RECT 358.875 85.205 359.205 85.535 ;
        RECT 358.875 82.895 359.205 83.225 ;
        RECT 358.875 82.045 359.205 82.375 ;
        RECT 358.875 79.735 359.205 80.065 ;
        RECT 358.875 78.885 359.205 79.215 ;
        RECT 358.875 76.575 359.205 76.905 ;
        RECT 358.875 74.995 359.205 75.325 ;
        RECT 358.875 74.145 359.205 74.475 ;
        RECT 358.875 71.835 359.205 72.165 ;
        RECT 358.875 70.985 359.205 71.315 ;
        RECT 358.875 68.675 359.205 69.005 ;
        RECT 358.875 67.825 359.205 68.155 ;
        RECT 358.875 65.515 359.205 65.845 ;
        RECT 358.875 64.665 359.205 64.995 ;
        RECT 358.875 62.355 359.205 62.685 ;
        RECT 358.875 60.775 359.205 61.105 ;
        RECT 358.875 59.925 359.205 60.255 ;
        RECT 358.875 57.615 359.205 57.945 ;
        RECT 358.875 56.765 359.205 57.095 ;
        RECT 358.875 54.455 359.205 54.785 ;
        RECT 358.875 53.605 359.205 53.935 ;
        RECT 358.875 51.295 359.205 51.625 ;
        RECT 358.875 50.445 359.205 50.775 ;
        RECT 358.875 48.135 359.205 48.465 ;
        RECT 358.875 46.555 359.205 46.885 ;
        RECT 358.875 45.705 359.205 46.035 ;
        RECT 358.875 43.395 359.205 43.725 ;
        RECT 358.875 42.545 359.205 42.875 ;
        RECT 358.875 40.235 359.205 40.565 ;
        RECT 358.875 39.385 359.205 39.715 ;
        RECT 358.875 37.075 359.205 37.405 ;
        RECT 358.875 36.225 359.205 36.555 ;
        RECT 358.875 33.915 359.205 34.245 ;
        RECT 358.875 32.335 359.205 32.665 ;
        RECT 358.875 31.485 359.205 31.815 ;
        RECT 358.875 29.175 359.205 29.505 ;
        RECT 358.875 28.325 359.205 28.655 ;
        RECT 358.875 26.015 359.205 26.345 ;
        RECT 358.875 25.165 359.205 25.495 ;
        RECT 358.875 22.855 359.205 23.185 ;
        RECT 358.875 22.005 359.205 22.335 ;
        RECT 358.875 19.695 359.205 20.025 ;
        RECT 358.875 18.115 359.205 18.445 ;
        RECT 358.875 17.265 359.205 17.595 ;
        RECT 358.875 14.955 359.205 15.285 ;
        RECT 358.875 14.105 359.205 14.435 ;
        RECT 358.875 11.795 359.205 12.125 ;
        RECT 358.875 10.945 359.205 11.275 ;
        RECT 358.875 8.635 359.205 8.965 ;
        RECT 358.875 7.785 359.205 8.115 ;
        RECT 358.875 5.475 359.205 5.805 ;
        RECT 358.875 3.895 359.205 4.225 ;
        RECT 358.875 3.045 359.205 3.375 ;
        RECT 358.875 0.87 359.205 1.2 ;
        RECT 358.875 -1.525 359.205 -1.195 ;
        RECT 358.875 -2.885 359.205 -2.555 ;
        RECT 358.875 -4.245 359.205 -3.915 ;
        RECT 358.875 -5.605 359.205 -5.275 ;
        RECT 358.875 -6.965 359.205 -6.635 ;
        RECT 358.875 -8.325 359.205 -7.995 ;
        RECT 358.875 -9.685 359.205 -9.355 ;
        RECT 358.875 -11.045 359.205 -10.715 ;
        RECT 358.875 -12.405 359.205 -12.075 ;
        RECT 358.875 -13.765 359.205 -13.435 ;
        RECT 358.875 -15.125 359.205 -14.795 ;
        RECT 358.875 -16.485 359.205 -16.155 ;
        RECT 358.875 -17.845 359.205 -17.515 ;
        RECT 358.875 -19.205 359.205 -18.875 ;
        RECT 358.875 -20.565 359.205 -20.235 ;
        RECT 358.875 -21.925 359.205 -21.595 ;
        RECT 358.875 -23.285 359.205 -22.955 ;
        RECT 358.875 -24.645 359.205 -24.315 ;
        RECT 358.875 -26.005 359.205 -25.675 ;
        RECT 358.875 -27.365 359.205 -27.035 ;
        RECT 358.875 -28.725 359.205 -28.395 ;
        RECT 358.875 -30.085 359.205 -29.755 ;
        RECT 358.875 -31.445 359.205 -31.115 ;
        RECT 358.875 -32.805 359.205 -32.475 ;
        RECT 358.875 -34.165 359.205 -33.835 ;
        RECT 358.875 -35.525 359.205 -35.195 ;
        RECT 358.875 -36.885 359.205 -36.555 ;
        RECT 358.875 -38.245 359.205 -37.915 ;
        RECT 358.875 -39.605 359.205 -39.275 ;
        RECT 358.875 -40.965 359.205 -40.635 ;
        RECT 358.875 -42.325 359.205 -41.995 ;
        RECT 358.875 -43.685 359.205 -43.355 ;
        RECT 358.875 -45.045 359.205 -44.715 ;
        RECT 358.875 -46.405 359.205 -46.075 ;
        RECT 358.875 -47.765 359.205 -47.435 ;
        RECT 358.875 -49.125 359.205 -48.795 ;
        RECT 358.875 -50.485 359.205 -50.155 ;
        RECT 358.875 -51.845 359.205 -51.515 ;
        RECT 358.875 -53.205 359.205 -52.875 ;
        RECT 358.875 -54.565 359.205 -54.235 ;
        RECT 358.875 -55.925 359.205 -55.595 ;
        RECT 358.875 -57.285 359.205 -56.955 ;
        RECT 358.875 -58.645 359.205 -58.315 ;
        RECT 358.875 -60.005 359.205 -59.675 ;
        RECT 358.875 -61.365 359.205 -61.035 ;
        RECT 358.875 -62.725 359.205 -62.395 ;
        RECT 358.875 -64.085 359.205 -63.755 ;
        RECT 358.875 -65.445 359.205 -65.115 ;
        RECT 358.875 -66.805 359.205 -66.475 ;
        RECT 358.875 -68.165 359.205 -67.835 ;
        RECT 358.875 -69.525 359.205 -69.195 ;
        RECT 358.875 -70.885 359.205 -70.555 ;
        RECT 358.875 -72.245 359.205 -71.915 ;
        RECT 358.875 -73.605 359.205 -73.275 ;
        RECT 358.875 -74.965 359.205 -74.635 ;
        RECT 358.875 -76.325 359.205 -75.995 ;
        RECT 358.875 -77.685 359.205 -77.355 ;
        RECT 358.875 -79.045 359.205 -78.715 ;
        RECT 358.875 -80.405 359.205 -80.075 ;
        RECT 358.875 -81.765 359.205 -81.435 ;
        RECT 358.875 -83.125 359.205 -82.795 ;
        RECT 358.875 -84.485 359.205 -84.155 ;
        RECT 358.875 -85.845 359.205 -85.515 ;
        RECT 358.875 -87.205 359.205 -86.875 ;
        RECT 358.875 -88.565 359.205 -88.235 ;
        RECT 358.875 -89.925 359.205 -89.595 ;
        RECT 358.875 -91.285 359.205 -90.955 ;
        RECT 358.875 -92.645 359.205 -92.315 ;
        RECT 358.875 -94.005 359.205 -93.675 ;
        RECT 358.875 -95.365 359.205 -95.035 ;
        RECT 358.875 -96.725 359.205 -96.395 ;
        RECT 358.875 -98.085 359.205 -97.755 ;
        RECT 358.875 -99.445 359.205 -99.115 ;
        RECT 358.875 -100.805 359.205 -100.475 ;
        RECT 358.875 -102.165 359.205 -101.835 ;
        RECT 358.875 -103.525 359.205 -103.195 ;
        RECT 358.875 -104.885 359.205 -104.555 ;
        RECT 358.875 -106.245 359.205 -105.915 ;
        RECT 358.875 -107.605 359.205 -107.275 ;
        RECT 358.875 -108.965 359.205 -108.635 ;
        RECT 358.875 -110.325 359.205 -109.995 ;
        RECT 358.875 -111.685 359.205 -111.355 ;
        RECT 358.875 -113.045 359.205 -112.715 ;
        RECT 358.875 -114.405 359.205 -114.075 ;
        RECT 358.875 -115.765 359.205 -115.435 ;
        RECT 358.875 -117.125 359.205 -116.795 ;
        RECT 358.875 -118.485 359.205 -118.155 ;
        RECT 358.875 -119.845 359.205 -119.515 ;
        RECT 358.875 -121.205 359.205 -120.875 ;
        RECT 358.875 -122.565 359.205 -122.235 ;
        RECT 358.875 -123.925 359.205 -123.595 ;
        RECT 358.875 -125.285 359.205 -124.955 ;
        RECT 358.875 -126.645 359.205 -126.315 ;
        RECT 358.875 -128.005 359.205 -127.675 ;
        RECT 358.875 -129.365 359.205 -129.035 ;
        RECT 358.875 -130.725 359.205 -130.395 ;
        RECT 358.875 -132.085 359.205 -131.755 ;
        RECT 358.875 -133.445 359.205 -133.115 ;
        RECT 358.875 -134.805 359.205 -134.475 ;
        RECT 358.875 -136.165 359.205 -135.835 ;
        RECT 358.875 -137.525 359.205 -137.195 ;
        RECT 358.875 -138.885 359.205 -138.555 ;
        RECT 358.875 -140.245 359.205 -139.915 ;
        RECT 358.875 -141.605 359.205 -141.275 ;
        RECT 358.875 -142.965 359.205 -142.635 ;
        RECT 358.875 -144.325 359.205 -143.995 ;
        RECT 358.875 -145.685 359.205 -145.355 ;
        RECT 358.875 -147.045 359.205 -146.715 ;
        RECT 358.875 -148.405 359.205 -148.075 ;
        RECT 358.875 -149.765 359.205 -149.435 ;
        RECT 358.875 -151.125 359.205 -150.795 ;
        RECT 358.875 -152.485 359.205 -152.155 ;
        RECT 358.875 -153.845 359.205 -153.515 ;
        RECT 358.875 -155.205 359.205 -154.875 ;
        RECT 358.875 -156.565 359.205 -156.235 ;
        RECT 358.875 -157.925 359.205 -157.595 ;
        RECT 358.875 -159.285 359.205 -158.955 ;
        RECT 358.875 -160.645 359.205 -160.315 ;
        RECT 358.875 -162.005 359.205 -161.675 ;
        RECT 358.875 -163.365 359.205 -163.035 ;
        RECT 358.875 -164.725 359.205 -164.395 ;
        RECT 358.875 -166.085 359.205 -165.755 ;
        RECT 358.875 -167.445 359.205 -167.115 ;
        RECT 358.875 -168.805 359.205 -168.475 ;
        RECT 358.875 -170.165 359.205 -169.835 ;
        RECT 358.875 -171.525 359.205 -171.195 ;
        RECT 358.875 -172.885 359.205 -172.555 ;
        RECT 358.875 -174.245 359.205 -173.915 ;
        RECT 358.875 -175.605 359.205 -175.275 ;
        RECT 358.875 -176.965 359.205 -176.635 ;
        RECT 358.875 -178.325 359.205 -177.995 ;
        RECT 358.875 -179.685 359.205 -179.355 ;
        RECT 358.875 -181.045 359.205 -180.715 ;
        RECT 358.875 -182.405 359.205 -182.075 ;
        RECT 358.875 -183.765 359.205 -183.435 ;
        RECT 358.875 -185.125 359.205 -184.795 ;
        RECT 358.875 -186.485 359.205 -186.155 ;
        RECT 358.875 -187.845 359.205 -187.515 ;
        RECT 358.875 -189.205 359.205 -188.875 ;
        RECT 358.875 -190.565 359.205 -190.235 ;
        RECT 358.875 -191.925 359.205 -191.595 ;
        RECT 358.875 -193.285 359.205 -192.955 ;
        RECT 358.875 -194.645 359.205 -194.315 ;
        RECT 358.875 -196.005 359.205 -195.675 ;
        RECT 358.875 -197.365 359.205 -197.035 ;
        RECT 358.875 -198.725 359.205 -198.395 ;
        RECT 358.875 -200.085 359.205 -199.755 ;
        RECT 358.875 -201.445 359.205 -201.115 ;
        RECT 358.875 -202.805 359.205 -202.475 ;
        RECT 358.875 -204.165 359.205 -203.835 ;
        RECT 358.875 -205.525 359.205 -205.195 ;
        RECT 358.875 -206.885 359.205 -206.555 ;
        RECT 358.875 -208.245 359.205 -207.915 ;
        RECT 358.875 -209.605 359.205 -209.275 ;
        RECT 358.875 -210.965 359.205 -210.635 ;
        RECT 358.875 -212.325 359.205 -211.995 ;
        RECT 358.875 -213.685 359.205 -213.355 ;
        RECT 358.875 -215.045 359.205 -214.715 ;
        RECT 358.875 -216.405 359.205 -216.075 ;
        RECT 358.875 -217.765 359.205 -217.435 ;
        RECT 358.875 -219.125 359.205 -218.795 ;
        RECT 358.875 -220.485 359.205 -220.155 ;
        RECT 358.875 -221.845 359.205 -221.515 ;
        RECT 358.875 -223.205 359.205 -222.875 ;
        RECT 358.875 -224.565 359.205 -224.235 ;
        RECT 358.875 -225.925 359.205 -225.595 ;
        RECT 358.875 -227.285 359.205 -226.955 ;
        RECT 358.875 -228.645 359.205 -228.315 ;
        RECT 358.875 -230.005 359.205 -229.675 ;
        RECT 358.875 -231.365 359.205 -231.035 ;
        RECT 358.875 -232.725 359.205 -232.395 ;
        RECT 358.875 -234.085 359.205 -233.755 ;
        RECT 358.875 -235.445 359.205 -235.115 ;
        RECT 358.875 -236.805 359.205 -236.475 ;
        RECT 358.875 -238.165 359.205 -237.835 ;
        RECT 358.875 -243.81 359.205 -242.68 ;
        RECT 358.88 -243.925 359.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 -181.045 360.565 -180.715 ;
        RECT 360.235 -182.405 360.565 -182.075 ;
        RECT 360.235 -183.765 360.565 -183.435 ;
        RECT 360.235 -185.125 360.565 -184.795 ;
        RECT 360.235 -186.485 360.565 -186.155 ;
        RECT 360.235 -187.845 360.565 -187.515 ;
        RECT 360.235 -189.205 360.565 -188.875 ;
        RECT 360.235 -190.565 360.565 -190.235 ;
        RECT 360.235 -191.925 360.565 -191.595 ;
        RECT 360.235 -193.285 360.565 -192.955 ;
        RECT 360.235 -194.645 360.565 -194.315 ;
        RECT 360.235 -196.005 360.565 -195.675 ;
        RECT 360.235 -197.365 360.565 -197.035 ;
        RECT 360.235 -198.725 360.565 -198.395 ;
        RECT 360.235 -200.085 360.565 -199.755 ;
        RECT 360.235 -201.445 360.565 -201.115 ;
        RECT 360.235 -202.805 360.565 -202.475 ;
        RECT 360.235 -204.165 360.565 -203.835 ;
        RECT 360.235 -205.525 360.565 -205.195 ;
        RECT 360.235 -206.885 360.565 -206.555 ;
        RECT 360.235 -208.245 360.565 -207.915 ;
        RECT 360.235 -209.605 360.565 -209.275 ;
        RECT 360.235 -210.965 360.565 -210.635 ;
        RECT 360.235 -212.325 360.565 -211.995 ;
        RECT 360.235 -213.685 360.565 -213.355 ;
        RECT 360.235 -215.045 360.565 -214.715 ;
        RECT 360.235 -216.405 360.565 -216.075 ;
        RECT 360.235 -217.765 360.565 -217.435 ;
        RECT 360.235 -219.125 360.565 -218.795 ;
        RECT 360.235 -220.485 360.565 -220.155 ;
        RECT 360.235 -221.845 360.565 -221.515 ;
        RECT 360.235 -223.205 360.565 -222.875 ;
        RECT 360.235 -224.565 360.565 -224.235 ;
        RECT 360.235 -225.925 360.565 -225.595 ;
        RECT 360.235 -227.285 360.565 -226.955 ;
        RECT 360.235 -228.645 360.565 -228.315 ;
        RECT 360.235 -230.005 360.565 -229.675 ;
        RECT 360.235 -231.365 360.565 -231.035 ;
        RECT 360.235 -232.725 360.565 -232.395 ;
        RECT 360.235 -234.085 360.565 -233.755 ;
        RECT 360.235 -235.445 360.565 -235.115 ;
        RECT 360.235 -236.805 360.565 -236.475 ;
        RECT 360.235 -238.165 360.565 -237.835 ;
        RECT 360.235 -243.81 360.565 -242.68 ;
        RECT 360.24 -243.925 360.56 248.005 ;
        RECT 360.235 246.76 360.565 247.89 ;
        RECT 360.235 241.915 360.565 242.245 ;
        RECT 360.235 240.555 360.565 240.885 ;
        RECT 360.235 239.195 360.565 239.525 ;
        RECT 360.235 237.835 360.565 238.165 ;
        RECT 360.235 235.17 360.565 235.5 ;
        RECT 360.235 232.995 360.565 233.325 ;
        RECT 360.235 231.415 360.565 231.745 ;
        RECT 360.235 230.565 360.565 230.895 ;
        RECT 360.235 228.255 360.565 228.585 ;
        RECT 360.235 227.405 360.565 227.735 ;
        RECT 360.235 225.095 360.565 225.425 ;
        RECT 360.235 224.245 360.565 224.575 ;
        RECT 360.235 221.935 360.565 222.265 ;
        RECT 360.235 221.085 360.565 221.415 ;
        RECT 360.235 218.775 360.565 219.105 ;
        RECT 360.235 217.195 360.565 217.525 ;
        RECT 360.235 216.345 360.565 216.675 ;
        RECT 360.235 214.035 360.565 214.365 ;
        RECT 360.235 213.185 360.565 213.515 ;
        RECT 360.235 210.875 360.565 211.205 ;
        RECT 360.235 210.025 360.565 210.355 ;
        RECT 360.235 207.715 360.565 208.045 ;
        RECT 360.235 206.865 360.565 207.195 ;
        RECT 360.235 204.555 360.565 204.885 ;
        RECT 360.235 202.975 360.565 203.305 ;
        RECT 360.235 202.125 360.565 202.455 ;
        RECT 360.235 199.815 360.565 200.145 ;
        RECT 360.235 198.965 360.565 199.295 ;
        RECT 360.235 196.655 360.565 196.985 ;
        RECT 360.235 195.805 360.565 196.135 ;
        RECT 360.235 193.495 360.565 193.825 ;
        RECT 360.235 192.645 360.565 192.975 ;
        RECT 360.235 190.335 360.565 190.665 ;
        RECT 360.235 188.755 360.565 189.085 ;
        RECT 360.235 187.905 360.565 188.235 ;
        RECT 360.235 185.595 360.565 185.925 ;
        RECT 360.235 184.745 360.565 185.075 ;
        RECT 360.235 182.435 360.565 182.765 ;
        RECT 360.235 181.585 360.565 181.915 ;
        RECT 360.235 179.275 360.565 179.605 ;
        RECT 360.235 178.425 360.565 178.755 ;
        RECT 360.235 176.115 360.565 176.445 ;
        RECT 360.235 174.535 360.565 174.865 ;
        RECT 360.235 173.685 360.565 174.015 ;
        RECT 360.235 171.375 360.565 171.705 ;
        RECT 360.235 170.525 360.565 170.855 ;
        RECT 360.235 168.215 360.565 168.545 ;
        RECT 360.235 167.365 360.565 167.695 ;
        RECT 360.235 165.055 360.565 165.385 ;
        RECT 360.235 164.205 360.565 164.535 ;
        RECT 360.235 161.895 360.565 162.225 ;
        RECT 360.235 160.315 360.565 160.645 ;
        RECT 360.235 159.465 360.565 159.795 ;
        RECT 360.235 157.155 360.565 157.485 ;
        RECT 360.235 156.305 360.565 156.635 ;
        RECT 360.235 153.995 360.565 154.325 ;
        RECT 360.235 153.145 360.565 153.475 ;
        RECT 360.235 150.835 360.565 151.165 ;
        RECT 360.235 149.985 360.565 150.315 ;
        RECT 360.235 147.675 360.565 148.005 ;
        RECT 360.235 146.095 360.565 146.425 ;
        RECT 360.235 145.245 360.565 145.575 ;
        RECT 360.235 142.935 360.565 143.265 ;
        RECT 360.235 142.085 360.565 142.415 ;
        RECT 360.235 139.775 360.565 140.105 ;
        RECT 360.235 138.925 360.565 139.255 ;
        RECT 360.235 136.615 360.565 136.945 ;
        RECT 360.235 135.765 360.565 136.095 ;
        RECT 360.235 133.455 360.565 133.785 ;
        RECT 360.235 131.875 360.565 132.205 ;
        RECT 360.235 131.025 360.565 131.355 ;
        RECT 360.235 128.715 360.565 129.045 ;
        RECT 360.235 127.865 360.565 128.195 ;
        RECT 360.235 125.555 360.565 125.885 ;
        RECT 360.235 124.705 360.565 125.035 ;
        RECT 360.235 122.395 360.565 122.725 ;
        RECT 360.235 121.545 360.565 121.875 ;
        RECT 360.235 119.235 360.565 119.565 ;
        RECT 360.235 117.655 360.565 117.985 ;
        RECT 360.235 116.805 360.565 117.135 ;
        RECT 360.235 114.495 360.565 114.825 ;
        RECT 360.235 113.645 360.565 113.975 ;
        RECT 360.235 111.335 360.565 111.665 ;
        RECT 360.235 110.485 360.565 110.815 ;
        RECT 360.235 108.175 360.565 108.505 ;
        RECT 360.235 107.325 360.565 107.655 ;
        RECT 360.235 105.015 360.565 105.345 ;
        RECT 360.235 103.435 360.565 103.765 ;
        RECT 360.235 102.585 360.565 102.915 ;
        RECT 360.235 100.275 360.565 100.605 ;
        RECT 360.235 99.425 360.565 99.755 ;
        RECT 360.235 97.115 360.565 97.445 ;
        RECT 360.235 96.265 360.565 96.595 ;
        RECT 360.235 93.955 360.565 94.285 ;
        RECT 360.235 93.105 360.565 93.435 ;
        RECT 360.235 90.795 360.565 91.125 ;
        RECT 360.235 89.215 360.565 89.545 ;
        RECT 360.235 88.365 360.565 88.695 ;
        RECT 360.235 86.055 360.565 86.385 ;
        RECT 360.235 85.205 360.565 85.535 ;
        RECT 360.235 82.895 360.565 83.225 ;
        RECT 360.235 82.045 360.565 82.375 ;
        RECT 360.235 79.735 360.565 80.065 ;
        RECT 360.235 78.885 360.565 79.215 ;
        RECT 360.235 76.575 360.565 76.905 ;
        RECT 360.235 74.995 360.565 75.325 ;
        RECT 360.235 74.145 360.565 74.475 ;
        RECT 360.235 71.835 360.565 72.165 ;
        RECT 360.235 70.985 360.565 71.315 ;
        RECT 360.235 68.675 360.565 69.005 ;
        RECT 360.235 67.825 360.565 68.155 ;
        RECT 360.235 65.515 360.565 65.845 ;
        RECT 360.235 64.665 360.565 64.995 ;
        RECT 360.235 62.355 360.565 62.685 ;
        RECT 360.235 60.775 360.565 61.105 ;
        RECT 360.235 59.925 360.565 60.255 ;
        RECT 360.235 57.615 360.565 57.945 ;
        RECT 360.235 56.765 360.565 57.095 ;
        RECT 360.235 54.455 360.565 54.785 ;
        RECT 360.235 53.605 360.565 53.935 ;
        RECT 360.235 51.295 360.565 51.625 ;
        RECT 360.235 50.445 360.565 50.775 ;
        RECT 360.235 48.135 360.565 48.465 ;
        RECT 360.235 46.555 360.565 46.885 ;
        RECT 360.235 45.705 360.565 46.035 ;
        RECT 360.235 43.395 360.565 43.725 ;
        RECT 360.235 42.545 360.565 42.875 ;
        RECT 360.235 40.235 360.565 40.565 ;
        RECT 360.235 39.385 360.565 39.715 ;
        RECT 360.235 37.075 360.565 37.405 ;
        RECT 360.235 36.225 360.565 36.555 ;
        RECT 360.235 33.915 360.565 34.245 ;
        RECT 360.235 32.335 360.565 32.665 ;
        RECT 360.235 31.485 360.565 31.815 ;
        RECT 360.235 29.175 360.565 29.505 ;
        RECT 360.235 28.325 360.565 28.655 ;
        RECT 360.235 26.015 360.565 26.345 ;
        RECT 360.235 25.165 360.565 25.495 ;
        RECT 360.235 22.855 360.565 23.185 ;
        RECT 360.235 22.005 360.565 22.335 ;
        RECT 360.235 19.695 360.565 20.025 ;
        RECT 360.235 18.115 360.565 18.445 ;
        RECT 360.235 17.265 360.565 17.595 ;
        RECT 360.235 14.955 360.565 15.285 ;
        RECT 360.235 14.105 360.565 14.435 ;
        RECT 360.235 11.795 360.565 12.125 ;
        RECT 360.235 10.945 360.565 11.275 ;
        RECT 360.235 8.635 360.565 8.965 ;
        RECT 360.235 7.785 360.565 8.115 ;
        RECT 360.235 5.475 360.565 5.805 ;
        RECT 360.235 3.895 360.565 4.225 ;
        RECT 360.235 3.045 360.565 3.375 ;
        RECT 360.235 0.87 360.565 1.2 ;
        RECT 360.235 -1.525 360.565 -1.195 ;
        RECT 360.235 -2.885 360.565 -2.555 ;
        RECT 360.235 -4.245 360.565 -3.915 ;
        RECT 360.235 -5.605 360.565 -5.275 ;
        RECT 360.235 -6.965 360.565 -6.635 ;
        RECT 360.235 -8.325 360.565 -7.995 ;
        RECT 360.235 -9.685 360.565 -9.355 ;
        RECT 360.235 -11.045 360.565 -10.715 ;
        RECT 360.235 -12.405 360.565 -12.075 ;
        RECT 360.235 -13.765 360.565 -13.435 ;
        RECT 360.235 -15.125 360.565 -14.795 ;
        RECT 360.235 -16.485 360.565 -16.155 ;
        RECT 360.235 -17.845 360.565 -17.515 ;
        RECT 360.235 -19.205 360.565 -18.875 ;
        RECT 360.235 -20.565 360.565 -20.235 ;
        RECT 360.235 -21.925 360.565 -21.595 ;
        RECT 360.235 -23.285 360.565 -22.955 ;
        RECT 360.235 -24.645 360.565 -24.315 ;
        RECT 360.235 -26.005 360.565 -25.675 ;
        RECT 360.235 -27.365 360.565 -27.035 ;
        RECT 360.235 -28.725 360.565 -28.395 ;
        RECT 360.235 -30.085 360.565 -29.755 ;
        RECT 360.235 -31.445 360.565 -31.115 ;
        RECT 360.235 -32.805 360.565 -32.475 ;
        RECT 360.235 -34.165 360.565 -33.835 ;
        RECT 360.235 -35.525 360.565 -35.195 ;
        RECT 360.235 -36.885 360.565 -36.555 ;
        RECT 360.235 -38.245 360.565 -37.915 ;
        RECT 360.235 -39.605 360.565 -39.275 ;
        RECT 360.235 -40.965 360.565 -40.635 ;
        RECT 360.235 -42.325 360.565 -41.995 ;
        RECT 360.235 -43.685 360.565 -43.355 ;
        RECT 360.235 -45.045 360.565 -44.715 ;
        RECT 360.235 -46.405 360.565 -46.075 ;
        RECT 360.235 -47.765 360.565 -47.435 ;
        RECT 360.235 -49.125 360.565 -48.795 ;
        RECT 360.235 -50.485 360.565 -50.155 ;
        RECT 360.235 -51.845 360.565 -51.515 ;
        RECT 360.235 -53.205 360.565 -52.875 ;
        RECT 360.235 -54.565 360.565 -54.235 ;
        RECT 360.235 -55.925 360.565 -55.595 ;
        RECT 360.235 -57.285 360.565 -56.955 ;
        RECT 360.235 -58.645 360.565 -58.315 ;
        RECT 360.235 -60.005 360.565 -59.675 ;
        RECT 360.235 -61.365 360.565 -61.035 ;
        RECT 360.235 -62.725 360.565 -62.395 ;
        RECT 360.235 -64.085 360.565 -63.755 ;
        RECT 360.235 -65.445 360.565 -65.115 ;
        RECT 360.235 -66.805 360.565 -66.475 ;
        RECT 360.235 -68.165 360.565 -67.835 ;
        RECT 360.235 -69.525 360.565 -69.195 ;
        RECT 360.235 -70.885 360.565 -70.555 ;
        RECT 360.235 -72.245 360.565 -71.915 ;
        RECT 360.235 -73.605 360.565 -73.275 ;
        RECT 360.235 -74.965 360.565 -74.635 ;
        RECT 360.235 -76.325 360.565 -75.995 ;
        RECT 360.235 -77.685 360.565 -77.355 ;
        RECT 360.235 -79.045 360.565 -78.715 ;
        RECT 360.235 -80.405 360.565 -80.075 ;
        RECT 360.235 -81.765 360.565 -81.435 ;
        RECT 360.235 -83.125 360.565 -82.795 ;
        RECT 360.235 -84.485 360.565 -84.155 ;
        RECT 360.235 -85.845 360.565 -85.515 ;
        RECT 360.235 -87.205 360.565 -86.875 ;
        RECT 360.235 -88.565 360.565 -88.235 ;
        RECT 360.235 -89.925 360.565 -89.595 ;
        RECT 360.235 -91.285 360.565 -90.955 ;
        RECT 360.235 -92.645 360.565 -92.315 ;
        RECT 360.235 -94.005 360.565 -93.675 ;
        RECT 360.235 -95.365 360.565 -95.035 ;
        RECT 360.235 -96.725 360.565 -96.395 ;
        RECT 360.235 -98.085 360.565 -97.755 ;
        RECT 360.235 -99.445 360.565 -99.115 ;
        RECT 360.235 -100.805 360.565 -100.475 ;
        RECT 360.235 -102.165 360.565 -101.835 ;
        RECT 360.235 -103.525 360.565 -103.195 ;
        RECT 360.235 -104.885 360.565 -104.555 ;
        RECT 360.235 -106.245 360.565 -105.915 ;
        RECT 360.235 -107.605 360.565 -107.275 ;
        RECT 360.235 -108.965 360.565 -108.635 ;
        RECT 360.235 -110.325 360.565 -109.995 ;
        RECT 360.235 -111.685 360.565 -111.355 ;
        RECT 360.235 -113.045 360.565 -112.715 ;
        RECT 360.235 -114.405 360.565 -114.075 ;
        RECT 360.235 -115.765 360.565 -115.435 ;
        RECT 360.235 -117.125 360.565 -116.795 ;
        RECT 360.235 -118.485 360.565 -118.155 ;
        RECT 360.235 -119.845 360.565 -119.515 ;
        RECT 360.235 -121.205 360.565 -120.875 ;
        RECT 360.235 -122.565 360.565 -122.235 ;
        RECT 360.235 -123.925 360.565 -123.595 ;
        RECT 360.235 -125.285 360.565 -124.955 ;
        RECT 360.235 -126.645 360.565 -126.315 ;
        RECT 360.235 -128.005 360.565 -127.675 ;
        RECT 360.235 -129.365 360.565 -129.035 ;
        RECT 360.235 -130.725 360.565 -130.395 ;
        RECT 360.235 -132.085 360.565 -131.755 ;
        RECT 360.235 -133.445 360.565 -133.115 ;
        RECT 360.235 -134.805 360.565 -134.475 ;
        RECT 360.235 -136.165 360.565 -135.835 ;
        RECT 360.235 -137.525 360.565 -137.195 ;
        RECT 360.235 -138.885 360.565 -138.555 ;
        RECT 360.235 -140.245 360.565 -139.915 ;
        RECT 360.235 -141.605 360.565 -141.275 ;
        RECT 360.235 -142.965 360.565 -142.635 ;
        RECT 360.235 -144.325 360.565 -143.995 ;
        RECT 360.235 -145.685 360.565 -145.355 ;
        RECT 360.235 -147.045 360.565 -146.715 ;
        RECT 360.235 -148.405 360.565 -148.075 ;
        RECT 360.235 -149.765 360.565 -149.435 ;
        RECT 360.235 -151.125 360.565 -150.795 ;
        RECT 360.235 -152.485 360.565 -152.155 ;
        RECT 360.235 -153.845 360.565 -153.515 ;
        RECT 360.235 -155.205 360.565 -154.875 ;
        RECT 360.235 -156.565 360.565 -156.235 ;
        RECT 360.235 -157.925 360.565 -157.595 ;
        RECT 360.235 -159.285 360.565 -158.955 ;
        RECT 360.235 -160.645 360.565 -160.315 ;
        RECT 360.235 -162.005 360.565 -161.675 ;
        RECT 360.235 -163.365 360.565 -163.035 ;
        RECT 360.235 -164.725 360.565 -164.395 ;
        RECT 360.235 -166.085 360.565 -165.755 ;
        RECT 360.235 -167.445 360.565 -167.115 ;
        RECT 360.235 -168.805 360.565 -168.475 ;
        RECT 360.235 -170.165 360.565 -169.835 ;
        RECT 360.235 -171.525 360.565 -171.195 ;
        RECT 360.235 -172.885 360.565 -172.555 ;
        RECT 360.235 -174.245 360.565 -173.915 ;
        RECT 360.235 -175.605 360.565 -175.275 ;
        RECT 360.235 -176.965 360.565 -176.635 ;
        RECT 360.235 -178.325 360.565 -177.995 ;
        RECT 360.235 -179.685 360.565 -179.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.56 -125.535 340.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 246.76 341.525 247.89 ;
        RECT 341.195 241.915 341.525 242.245 ;
        RECT 341.195 240.555 341.525 240.885 ;
        RECT 341.195 239.195 341.525 239.525 ;
        RECT 341.195 237.835 341.525 238.165 ;
        RECT 341.2 237.16 341.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 -126.645 341.525 -126.315 ;
        RECT 341.195 -128.005 341.525 -127.675 ;
        RECT 341.195 -129.365 341.525 -129.035 ;
        RECT 341.195 -130.725 341.525 -130.395 ;
        RECT 341.195 -132.085 341.525 -131.755 ;
        RECT 341.195 -133.445 341.525 -133.115 ;
        RECT 341.195 -134.805 341.525 -134.475 ;
        RECT 341.195 -136.165 341.525 -135.835 ;
        RECT 341.195 -137.525 341.525 -137.195 ;
        RECT 341.195 -138.885 341.525 -138.555 ;
        RECT 341.195 -140.245 341.525 -139.915 ;
        RECT 341.195 -141.605 341.525 -141.275 ;
        RECT 341.195 -142.965 341.525 -142.635 ;
        RECT 341.195 -144.325 341.525 -143.995 ;
        RECT 341.195 -145.685 341.525 -145.355 ;
        RECT 341.195 -147.045 341.525 -146.715 ;
        RECT 341.195 -148.405 341.525 -148.075 ;
        RECT 341.195 -149.765 341.525 -149.435 ;
        RECT 341.195 -151.125 341.525 -150.795 ;
        RECT 341.195 -152.485 341.525 -152.155 ;
        RECT 341.195 -153.845 341.525 -153.515 ;
        RECT 341.195 -155.205 341.525 -154.875 ;
        RECT 341.195 -156.565 341.525 -156.235 ;
        RECT 341.195 -157.925 341.525 -157.595 ;
        RECT 341.195 -159.285 341.525 -158.955 ;
        RECT 341.195 -160.645 341.525 -160.315 ;
        RECT 341.195 -162.005 341.525 -161.675 ;
        RECT 341.195 -163.365 341.525 -163.035 ;
        RECT 341.195 -164.725 341.525 -164.395 ;
        RECT 341.195 -166.085 341.525 -165.755 ;
        RECT 341.195 -167.445 341.525 -167.115 ;
        RECT 341.195 -168.805 341.525 -168.475 ;
        RECT 341.195 -170.165 341.525 -169.835 ;
        RECT 341.195 -171.525 341.525 -171.195 ;
        RECT 341.195 -172.885 341.525 -172.555 ;
        RECT 341.195 -174.245 341.525 -173.915 ;
        RECT 341.195 -175.605 341.525 -175.275 ;
        RECT 341.195 -176.965 341.525 -176.635 ;
        RECT 341.195 -178.325 341.525 -177.995 ;
        RECT 341.195 -179.685 341.525 -179.355 ;
        RECT 341.195 -181.045 341.525 -180.715 ;
        RECT 341.195 -182.405 341.525 -182.075 ;
        RECT 341.195 -183.765 341.525 -183.435 ;
        RECT 341.195 -185.125 341.525 -184.795 ;
        RECT 341.195 -186.485 341.525 -186.155 ;
        RECT 341.195 -187.845 341.525 -187.515 ;
        RECT 341.195 -189.205 341.525 -188.875 ;
        RECT 341.195 -190.565 341.525 -190.235 ;
        RECT 341.195 -191.925 341.525 -191.595 ;
        RECT 341.195 -193.285 341.525 -192.955 ;
        RECT 341.195 -194.645 341.525 -194.315 ;
        RECT 341.195 -196.005 341.525 -195.675 ;
        RECT 341.195 -197.365 341.525 -197.035 ;
        RECT 341.195 -198.725 341.525 -198.395 ;
        RECT 341.195 -200.085 341.525 -199.755 ;
        RECT 341.195 -201.445 341.525 -201.115 ;
        RECT 341.195 -202.805 341.525 -202.475 ;
        RECT 341.195 -204.165 341.525 -203.835 ;
        RECT 341.195 -205.525 341.525 -205.195 ;
        RECT 341.195 -206.885 341.525 -206.555 ;
        RECT 341.195 -208.245 341.525 -207.915 ;
        RECT 341.195 -209.605 341.525 -209.275 ;
        RECT 341.195 -210.965 341.525 -210.635 ;
        RECT 341.195 -212.325 341.525 -211.995 ;
        RECT 341.195 -213.685 341.525 -213.355 ;
        RECT 341.195 -215.045 341.525 -214.715 ;
        RECT 341.195 -216.405 341.525 -216.075 ;
        RECT 341.195 -217.765 341.525 -217.435 ;
        RECT 341.195 -219.125 341.525 -218.795 ;
        RECT 341.195 -220.485 341.525 -220.155 ;
        RECT 341.195 -221.845 341.525 -221.515 ;
        RECT 341.195 -223.205 341.525 -222.875 ;
        RECT 341.195 -224.565 341.525 -224.235 ;
        RECT 341.195 -225.925 341.525 -225.595 ;
        RECT 341.195 -227.285 341.525 -226.955 ;
        RECT 341.195 -228.645 341.525 -228.315 ;
        RECT 341.195 -230.005 341.525 -229.675 ;
        RECT 341.195 -231.365 341.525 -231.035 ;
        RECT 341.195 -232.725 341.525 -232.395 ;
        RECT 341.195 -234.085 341.525 -233.755 ;
        RECT 341.195 -235.445 341.525 -235.115 ;
        RECT 341.195 -236.805 341.525 -236.475 ;
        RECT 341.195 -238.165 341.525 -237.835 ;
        RECT 341.195 -243.81 341.525 -242.68 ;
        RECT 341.2 -243.925 341.52 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 246.76 342.885 247.89 ;
        RECT 342.555 241.915 342.885 242.245 ;
        RECT 342.555 240.555 342.885 240.885 ;
        RECT 342.555 239.195 342.885 239.525 ;
        RECT 342.555 237.835 342.885 238.165 ;
        RECT 342.56 237.16 342.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 -1.525 342.885 -1.195 ;
        RECT 342.555 -2.885 342.885 -2.555 ;
        RECT 342.56 -3.56 342.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 246.76 344.245 247.89 ;
        RECT 343.915 241.915 344.245 242.245 ;
        RECT 343.915 240.555 344.245 240.885 ;
        RECT 343.915 239.195 344.245 239.525 ;
        RECT 343.915 237.835 344.245 238.165 ;
        RECT 343.92 237.16 344.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 -1.525 344.245 -1.195 ;
        RECT 343.915 -2.885 344.245 -2.555 ;
        RECT 343.92 -3.56 344.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 246.76 345.605 247.89 ;
        RECT 345.275 241.915 345.605 242.245 ;
        RECT 345.275 240.555 345.605 240.885 ;
        RECT 345.275 239.195 345.605 239.525 ;
        RECT 345.275 237.835 345.605 238.165 ;
        RECT 345.28 237.16 345.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 -1.525 345.605 -1.195 ;
        RECT 345.275 -2.885 345.605 -2.555 ;
        RECT 345.28 -3.56 345.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 -122.565 345.605 -122.235 ;
        RECT 345.275 -123.925 345.605 -123.595 ;
        RECT 345.275 -125.285 345.605 -124.955 ;
        RECT 345.275 -126.645 345.605 -126.315 ;
        RECT 345.275 -128.005 345.605 -127.675 ;
        RECT 345.275 -129.365 345.605 -129.035 ;
        RECT 345.275 -130.725 345.605 -130.395 ;
        RECT 345.275 -132.085 345.605 -131.755 ;
        RECT 345.275 -133.445 345.605 -133.115 ;
        RECT 345.275 -134.805 345.605 -134.475 ;
        RECT 345.275 -136.165 345.605 -135.835 ;
        RECT 345.275 -137.525 345.605 -137.195 ;
        RECT 345.275 -138.885 345.605 -138.555 ;
        RECT 345.275 -140.245 345.605 -139.915 ;
        RECT 345.275 -141.605 345.605 -141.275 ;
        RECT 345.275 -142.965 345.605 -142.635 ;
        RECT 345.275 -144.325 345.605 -143.995 ;
        RECT 345.275 -145.685 345.605 -145.355 ;
        RECT 345.275 -147.045 345.605 -146.715 ;
        RECT 345.275 -148.405 345.605 -148.075 ;
        RECT 345.275 -149.765 345.605 -149.435 ;
        RECT 345.275 -151.125 345.605 -150.795 ;
        RECT 345.275 -152.485 345.605 -152.155 ;
        RECT 345.275 -153.845 345.605 -153.515 ;
        RECT 345.275 -155.205 345.605 -154.875 ;
        RECT 345.275 -156.565 345.605 -156.235 ;
        RECT 345.275 -157.925 345.605 -157.595 ;
        RECT 345.275 -159.285 345.605 -158.955 ;
        RECT 345.275 -160.645 345.605 -160.315 ;
        RECT 345.275 -162.005 345.605 -161.675 ;
        RECT 345.275 -163.365 345.605 -163.035 ;
        RECT 345.275 -164.725 345.605 -164.395 ;
        RECT 345.275 -166.085 345.605 -165.755 ;
        RECT 345.275 -167.445 345.605 -167.115 ;
        RECT 345.275 -168.805 345.605 -168.475 ;
        RECT 345.275 -170.165 345.605 -169.835 ;
        RECT 345.275 -171.525 345.605 -171.195 ;
        RECT 345.275 -172.885 345.605 -172.555 ;
        RECT 345.275 -174.245 345.605 -173.915 ;
        RECT 345.275 -175.605 345.605 -175.275 ;
        RECT 345.275 -176.965 345.605 -176.635 ;
        RECT 345.275 -178.325 345.605 -177.995 ;
        RECT 345.275 -179.685 345.605 -179.355 ;
        RECT 345.275 -181.045 345.605 -180.715 ;
        RECT 345.275 -182.405 345.605 -182.075 ;
        RECT 345.275 -183.765 345.605 -183.435 ;
        RECT 345.275 -185.125 345.605 -184.795 ;
        RECT 345.275 -186.485 345.605 -186.155 ;
        RECT 345.275 -187.845 345.605 -187.515 ;
        RECT 345.275 -189.205 345.605 -188.875 ;
        RECT 345.275 -190.565 345.605 -190.235 ;
        RECT 345.275 -191.925 345.605 -191.595 ;
        RECT 345.275 -193.285 345.605 -192.955 ;
        RECT 345.275 -194.645 345.605 -194.315 ;
        RECT 345.275 -196.005 345.605 -195.675 ;
        RECT 345.275 -197.365 345.605 -197.035 ;
        RECT 345.275 -198.725 345.605 -198.395 ;
        RECT 345.275 -200.085 345.605 -199.755 ;
        RECT 345.275 -201.445 345.605 -201.115 ;
        RECT 345.275 -202.805 345.605 -202.475 ;
        RECT 345.275 -204.165 345.605 -203.835 ;
        RECT 345.275 -205.525 345.605 -205.195 ;
        RECT 345.275 -206.885 345.605 -206.555 ;
        RECT 345.275 -208.245 345.605 -207.915 ;
        RECT 345.275 -209.605 345.605 -209.275 ;
        RECT 345.275 -210.965 345.605 -210.635 ;
        RECT 345.275 -212.325 345.605 -211.995 ;
        RECT 345.275 -213.685 345.605 -213.355 ;
        RECT 345.275 -215.045 345.605 -214.715 ;
        RECT 345.275 -216.405 345.605 -216.075 ;
        RECT 345.275 -217.765 345.605 -217.435 ;
        RECT 345.275 -219.125 345.605 -218.795 ;
        RECT 345.275 -220.485 345.605 -220.155 ;
        RECT 345.275 -221.845 345.605 -221.515 ;
        RECT 345.275 -223.205 345.605 -222.875 ;
        RECT 345.275 -224.565 345.605 -224.235 ;
        RECT 345.275 -225.925 345.605 -225.595 ;
        RECT 345.275 -227.285 345.605 -226.955 ;
        RECT 345.275 -228.645 345.605 -228.315 ;
        RECT 345.275 -230.005 345.605 -229.675 ;
        RECT 345.275 -231.365 345.605 -231.035 ;
        RECT 345.275 -232.725 345.605 -232.395 ;
        RECT 345.275 -234.085 345.605 -233.755 ;
        RECT 345.275 -235.445 345.605 -235.115 ;
        RECT 345.275 -236.805 345.605 -236.475 ;
        RECT 345.275 -238.165 345.605 -237.835 ;
        RECT 345.275 -243.81 345.605 -242.68 ;
        RECT 345.28 -243.925 345.6 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 246.76 346.965 247.89 ;
        RECT 346.635 241.915 346.965 242.245 ;
        RECT 346.635 240.555 346.965 240.885 ;
        RECT 346.635 239.195 346.965 239.525 ;
        RECT 346.635 237.835 346.965 238.165 ;
        RECT 346.64 237.16 346.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 -1.525 346.965 -1.195 ;
        RECT 346.635 -2.885 346.965 -2.555 ;
        RECT 346.64 -3.56 346.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 -122.565 346.965 -122.235 ;
        RECT 346.635 -123.925 346.965 -123.595 ;
        RECT 346.635 -125.285 346.965 -124.955 ;
        RECT 346.635 -126.645 346.965 -126.315 ;
        RECT 346.635 -128.005 346.965 -127.675 ;
        RECT 346.635 -129.365 346.965 -129.035 ;
        RECT 346.635 -130.725 346.965 -130.395 ;
        RECT 346.635 -132.085 346.965 -131.755 ;
        RECT 346.635 -133.445 346.965 -133.115 ;
        RECT 346.635 -134.805 346.965 -134.475 ;
        RECT 346.635 -136.165 346.965 -135.835 ;
        RECT 346.635 -137.525 346.965 -137.195 ;
        RECT 346.635 -138.885 346.965 -138.555 ;
        RECT 346.635 -140.245 346.965 -139.915 ;
        RECT 346.635 -141.605 346.965 -141.275 ;
        RECT 346.635 -142.965 346.965 -142.635 ;
        RECT 346.635 -144.325 346.965 -143.995 ;
        RECT 346.635 -145.685 346.965 -145.355 ;
        RECT 346.635 -147.045 346.965 -146.715 ;
        RECT 346.635 -148.405 346.965 -148.075 ;
        RECT 346.635 -149.765 346.965 -149.435 ;
        RECT 346.635 -151.125 346.965 -150.795 ;
        RECT 346.635 -152.485 346.965 -152.155 ;
        RECT 346.635 -153.845 346.965 -153.515 ;
        RECT 346.635 -155.205 346.965 -154.875 ;
        RECT 346.635 -156.565 346.965 -156.235 ;
        RECT 346.635 -157.925 346.965 -157.595 ;
        RECT 346.635 -159.285 346.965 -158.955 ;
        RECT 346.635 -160.645 346.965 -160.315 ;
        RECT 346.635 -162.005 346.965 -161.675 ;
        RECT 346.635 -163.365 346.965 -163.035 ;
        RECT 346.635 -164.725 346.965 -164.395 ;
        RECT 346.635 -166.085 346.965 -165.755 ;
        RECT 346.635 -167.445 346.965 -167.115 ;
        RECT 346.635 -168.805 346.965 -168.475 ;
        RECT 346.635 -170.165 346.965 -169.835 ;
        RECT 346.635 -171.525 346.965 -171.195 ;
        RECT 346.635 -172.885 346.965 -172.555 ;
        RECT 346.635 -174.245 346.965 -173.915 ;
        RECT 346.635 -175.605 346.965 -175.275 ;
        RECT 346.635 -176.965 346.965 -176.635 ;
        RECT 346.635 -178.325 346.965 -177.995 ;
        RECT 346.635 -179.685 346.965 -179.355 ;
        RECT 346.635 -181.045 346.965 -180.715 ;
        RECT 346.635 -182.405 346.965 -182.075 ;
        RECT 346.635 -183.765 346.965 -183.435 ;
        RECT 346.635 -185.125 346.965 -184.795 ;
        RECT 346.635 -186.485 346.965 -186.155 ;
        RECT 346.635 -187.845 346.965 -187.515 ;
        RECT 346.635 -189.205 346.965 -188.875 ;
        RECT 346.635 -190.565 346.965 -190.235 ;
        RECT 346.635 -191.925 346.965 -191.595 ;
        RECT 346.635 -193.285 346.965 -192.955 ;
        RECT 346.635 -194.645 346.965 -194.315 ;
        RECT 346.635 -196.005 346.965 -195.675 ;
        RECT 346.635 -197.365 346.965 -197.035 ;
        RECT 346.635 -198.725 346.965 -198.395 ;
        RECT 346.635 -200.085 346.965 -199.755 ;
        RECT 346.635 -201.445 346.965 -201.115 ;
        RECT 346.635 -202.805 346.965 -202.475 ;
        RECT 346.635 -204.165 346.965 -203.835 ;
        RECT 346.635 -205.525 346.965 -205.195 ;
        RECT 346.635 -206.885 346.965 -206.555 ;
        RECT 346.635 -208.245 346.965 -207.915 ;
        RECT 346.635 -209.605 346.965 -209.275 ;
        RECT 346.635 -210.965 346.965 -210.635 ;
        RECT 346.635 -212.325 346.965 -211.995 ;
        RECT 346.635 -213.685 346.965 -213.355 ;
        RECT 346.635 -215.045 346.965 -214.715 ;
        RECT 346.635 -216.405 346.965 -216.075 ;
        RECT 346.635 -217.765 346.965 -217.435 ;
        RECT 346.635 -219.125 346.965 -218.795 ;
        RECT 346.635 -220.485 346.965 -220.155 ;
        RECT 346.635 -221.845 346.965 -221.515 ;
        RECT 346.635 -223.205 346.965 -222.875 ;
        RECT 346.635 -224.565 346.965 -224.235 ;
        RECT 346.635 -225.925 346.965 -225.595 ;
        RECT 346.635 -227.285 346.965 -226.955 ;
        RECT 346.635 -228.645 346.965 -228.315 ;
        RECT 346.635 -230.005 346.965 -229.675 ;
        RECT 346.635 -231.365 346.965 -231.035 ;
        RECT 346.635 -232.725 346.965 -232.395 ;
        RECT 346.635 -234.085 346.965 -233.755 ;
        RECT 346.635 -235.445 346.965 -235.115 ;
        RECT 346.635 -236.805 346.965 -236.475 ;
        RECT 346.635 -238.165 346.965 -237.835 ;
        RECT 346.635 -243.81 346.965 -242.68 ;
        RECT 346.64 -243.925 346.96 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 246.76 348.325 247.89 ;
        RECT 347.995 241.915 348.325 242.245 ;
        RECT 347.995 240.555 348.325 240.885 ;
        RECT 347.995 239.195 348.325 239.525 ;
        RECT 347.995 237.835 348.325 238.165 ;
        RECT 348 237.16 348.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 -1.525 348.325 -1.195 ;
        RECT 347.995 -2.885 348.325 -2.555 ;
        RECT 348 -3.56 348.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 -122.565 348.325 -122.235 ;
        RECT 347.995 -123.925 348.325 -123.595 ;
        RECT 347.995 -125.285 348.325 -124.955 ;
        RECT 347.995 -126.645 348.325 -126.315 ;
        RECT 347.995 -128.005 348.325 -127.675 ;
        RECT 347.995 -129.365 348.325 -129.035 ;
        RECT 347.995 -130.725 348.325 -130.395 ;
        RECT 347.995 -132.085 348.325 -131.755 ;
        RECT 347.995 -133.445 348.325 -133.115 ;
        RECT 347.995 -134.805 348.325 -134.475 ;
        RECT 347.995 -136.165 348.325 -135.835 ;
        RECT 347.995 -137.525 348.325 -137.195 ;
        RECT 347.995 -138.885 348.325 -138.555 ;
        RECT 347.995 -140.245 348.325 -139.915 ;
        RECT 347.995 -141.605 348.325 -141.275 ;
        RECT 347.995 -142.965 348.325 -142.635 ;
        RECT 347.995 -144.325 348.325 -143.995 ;
        RECT 347.995 -145.685 348.325 -145.355 ;
        RECT 347.995 -147.045 348.325 -146.715 ;
        RECT 347.995 -148.405 348.325 -148.075 ;
        RECT 347.995 -149.765 348.325 -149.435 ;
        RECT 347.995 -151.125 348.325 -150.795 ;
        RECT 347.995 -152.485 348.325 -152.155 ;
        RECT 347.995 -153.845 348.325 -153.515 ;
        RECT 347.995 -155.205 348.325 -154.875 ;
        RECT 347.995 -156.565 348.325 -156.235 ;
        RECT 347.995 -157.925 348.325 -157.595 ;
        RECT 347.995 -159.285 348.325 -158.955 ;
        RECT 347.995 -160.645 348.325 -160.315 ;
        RECT 347.995 -162.005 348.325 -161.675 ;
        RECT 347.995 -163.365 348.325 -163.035 ;
        RECT 347.995 -164.725 348.325 -164.395 ;
        RECT 347.995 -166.085 348.325 -165.755 ;
        RECT 347.995 -167.445 348.325 -167.115 ;
        RECT 347.995 -168.805 348.325 -168.475 ;
        RECT 347.995 -170.165 348.325 -169.835 ;
        RECT 347.995 -171.525 348.325 -171.195 ;
        RECT 347.995 -172.885 348.325 -172.555 ;
        RECT 347.995 -174.245 348.325 -173.915 ;
        RECT 347.995 -175.605 348.325 -175.275 ;
        RECT 347.995 -176.965 348.325 -176.635 ;
        RECT 347.995 -178.325 348.325 -177.995 ;
        RECT 347.995 -179.685 348.325 -179.355 ;
        RECT 347.995 -181.045 348.325 -180.715 ;
        RECT 347.995 -182.405 348.325 -182.075 ;
        RECT 347.995 -183.765 348.325 -183.435 ;
        RECT 347.995 -185.125 348.325 -184.795 ;
        RECT 347.995 -186.485 348.325 -186.155 ;
        RECT 347.995 -187.845 348.325 -187.515 ;
        RECT 347.995 -189.205 348.325 -188.875 ;
        RECT 347.995 -190.565 348.325 -190.235 ;
        RECT 347.995 -191.925 348.325 -191.595 ;
        RECT 347.995 -193.285 348.325 -192.955 ;
        RECT 347.995 -194.645 348.325 -194.315 ;
        RECT 347.995 -196.005 348.325 -195.675 ;
        RECT 347.995 -197.365 348.325 -197.035 ;
        RECT 347.995 -198.725 348.325 -198.395 ;
        RECT 347.995 -200.085 348.325 -199.755 ;
        RECT 347.995 -201.445 348.325 -201.115 ;
        RECT 347.995 -202.805 348.325 -202.475 ;
        RECT 347.995 -204.165 348.325 -203.835 ;
        RECT 347.995 -205.525 348.325 -205.195 ;
        RECT 347.995 -206.885 348.325 -206.555 ;
        RECT 347.995 -208.245 348.325 -207.915 ;
        RECT 347.995 -209.605 348.325 -209.275 ;
        RECT 347.995 -210.965 348.325 -210.635 ;
        RECT 347.995 -212.325 348.325 -211.995 ;
        RECT 347.995 -213.685 348.325 -213.355 ;
        RECT 347.995 -215.045 348.325 -214.715 ;
        RECT 347.995 -216.405 348.325 -216.075 ;
        RECT 347.995 -217.765 348.325 -217.435 ;
        RECT 347.995 -219.125 348.325 -218.795 ;
        RECT 347.995 -220.485 348.325 -220.155 ;
        RECT 347.995 -221.845 348.325 -221.515 ;
        RECT 347.995 -223.205 348.325 -222.875 ;
        RECT 347.995 -224.565 348.325 -224.235 ;
        RECT 347.995 -225.925 348.325 -225.595 ;
        RECT 347.995 -227.285 348.325 -226.955 ;
        RECT 347.995 -228.645 348.325 -228.315 ;
        RECT 347.995 -230.005 348.325 -229.675 ;
        RECT 347.995 -231.365 348.325 -231.035 ;
        RECT 347.995 -232.725 348.325 -232.395 ;
        RECT 347.995 -234.085 348.325 -233.755 ;
        RECT 347.995 -235.445 348.325 -235.115 ;
        RECT 347.995 -236.805 348.325 -236.475 ;
        RECT 347.995 -238.165 348.325 -237.835 ;
        RECT 347.995 -243.81 348.325 -242.68 ;
        RECT 348 -243.925 348.32 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 246.76 349.685 247.89 ;
        RECT 349.355 241.915 349.685 242.245 ;
        RECT 349.355 240.555 349.685 240.885 ;
        RECT 349.355 239.195 349.685 239.525 ;
        RECT 349.355 237.835 349.685 238.165 ;
        RECT 349.36 237.16 349.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 -1.525 349.685 -1.195 ;
        RECT 349.355 -2.885 349.685 -2.555 ;
        RECT 349.36 -3.56 349.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 -122.565 349.685 -122.235 ;
        RECT 349.355 -123.925 349.685 -123.595 ;
        RECT 349.355 -125.285 349.685 -124.955 ;
        RECT 349.355 -126.645 349.685 -126.315 ;
        RECT 349.355 -128.005 349.685 -127.675 ;
        RECT 349.355 -129.365 349.685 -129.035 ;
        RECT 349.355 -130.725 349.685 -130.395 ;
        RECT 349.355 -132.085 349.685 -131.755 ;
        RECT 349.355 -133.445 349.685 -133.115 ;
        RECT 349.355 -134.805 349.685 -134.475 ;
        RECT 349.355 -136.165 349.685 -135.835 ;
        RECT 349.355 -137.525 349.685 -137.195 ;
        RECT 349.355 -138.885 349.685 -138.555 ;
        RECT 349.355 -140.245 349.685 -139.915 ;
        RECT 349.355 -141.605 349.685 -141.275 ;
        RECT 349.355 -142.965 349.685 -142.635 ;
        RECT 349.355 -144.325 349.685 -143.995 ;
        RECT 349.355 -145.685 349.685 -145.355 ;
        RECT 349.355 -147.045 349.685 -146.715 ;
        RECT 349.355 -148.405 349.685 -148.075 ;
        RECT 349.355 -149.765 349.685 -149.435 ;
        RECT 349.355 -151.125 349.685 -150.795 ;
        RECT 349.355 -152.485 349.685 -152.155 ;
        RECT 349.355 -153.845 349.685 -153.515 ;
        RECT 349.355 -155.205 349.685 -154.875 ;
        RECT 349.355 -156.565 349.685 -156.235 ;
        RECT 349.355 -157.925 349.685 -157.595 ;
        RECT 349.355 -159.285 349.685 -158.955 ;
        RECT 349.355 -160.645 349.685 -160.315 ;
        RECT 349.355 -162.005 349.685 -161.675 ;
        RECT 349.355 -163.365 349.685 -163.035 ;
        RECT 349.355 -164.725 349.685 -164.395 ;
        RECT 349.355 -166.085 349.685 -165.755 ;
        RECT 349.355 -167.445 349.685 -167.115 ;
        RECT 349.355 -168.805 349.685 -168.475 ;
        RECT 349.355 -170.165 349.685 -169.835 ;
        RECT 349.355 -171.525 349.685 -171.195 ;
        RECT 349.355 -172.885 349.685 -172.555 ;
        RECT 349.355 -174.245 349.685 -173.915 ;
        RECT 349.355 -175.605 349.685 -175.275 ;
        RECT 349.355 -176.965 349.685 -176.635 ;
        RECT 349.355 -178.325 349.685 -177.995 ;
        RECT 349.355 -179.685 349.685 -179.355 ;
        RECT 349.355 -181.045 349.685 -180.715 ;
        RECT 349.355 -182.405 349.685 -182.075 ;
        RECT 349.355 -183.765 349.685 -183.435 ;
        RECT 349.355 -185.125 349.685 -184.795 ;
        RECT 349.355 -186.485 349.685 -186.155 ;
        RECT 349.355 -187.845 349.685 -187.515 ;
        RECT 349.355 -189.205 349.685 -188.875 ;
        RECT 349.355 -190.565 349.685 -190.235 ;
        RECT 349.355 -191.925 349.685 -191.595 ;
        RECT 349.355 -193.285 349.685 -192.955 ;
        RECT 349.355 -194.645 349.685 -194.315 ;
        RECT 349.355 -196.005 349.685 -195.675 ;
        RECT 349.355 -197.365 349.685 -197.035 ;
        RECT 349.355 -198.725 349.685 -198.395 ;
        RECT 349.355 -200.085 349.685 -199.755 ;
        RECT 349.355 -201.445 349.685 -201.115 ;
        RECT 349.355 -202.805 349.685 -202.475 ;
        RECT 349.355 -204.165 349.685 -203.835 ;
        RECT 349.355 -205.525 349.685 -205.195 ;
        RECT 349.355 -206.885 349.685 -206.555 ;
        RECT 349.355 -208.245 349.685 -207.915 ;
        RECT 349.355 -209.605 349.685 -209.275 ;
        RECT 349.355 -210.965 349.685 -210.635 ;
        RECT 349.355 -212.325 349.685 -211.995 ;
        RECT 349.355 -213.685 349.685 -213.355 ;
        RECT 349.355 -215.045 349.685 -214.715 ;
        RECT 349.355 -216.405 349.685 -216.075 ;
        RECT 349.355 -217.765 349.685 -217.435 ;
        RECT 349.355 -219.125 349.685 -218.795 ;
        RECT 349.355 -220.485 349.685 -220.155 ;
        RECT 349.355 -221.845 349.685 -221.515 ;
        RECT 349.355 -223.205 349.685 -222.875 ;
        RECT 349.355 -224.565 349.685 -224.235 ;
        RECT 349.355 -225.925 349.685 -225.595 ;
        RECT 349.355 -227.285 349.685 -226.955 ;
        RECT 349.355 -228.645 349.685 -228.315 ;
        RECT 349.355 -230.005 349.685 -229.675 ;
        RECT 349.355 -231.365 349.685 -231.035 ;
        RECT 349.355 -232.725 349.685 -232.395 ;
        RECT 349.355 -234.085 349.685 -233.755 ;
        RECT 349.355 -235.445 349.685 -235.115 ;
        RECT 349.355 -236.805 349.685 -236.475 ;
        RECT 349.355 -238.165 349.685 -237.835 ;
        RECT 349.355 -243.81 349.685 -242.68 ;
        RECT 349.36 -243.925 349.68 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 246.76 351.045 247.89 ;
        RECT 350.715 241.915 351.045 242.245 ;
        RECT 350.715 240.555 351.045 240.885 ;
        RECT 350.715 239.195 351.045 239.525 ;
        RECT 350.715 237.835 351.045 238.165 ;
        RECT 350.72 237.16 351.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 -1.525 351.045 -1.195 ;
        RECT 350.715 -2.885 351.045 -2.555 ;
        RECT 350.72 -3.56 351.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 -122.565 351.045 -122.235 ;
        RECT 350.715 -123.925 351.045 -123.595 ;
        RECT 350.715 -125.285 351.045 -124.955 ;
        RECT 350.715 -126.645 351.045 -126.315 ;
        RECT 350.715 -128.005 351.045 -127.675 ;
        RECT 350.715 -129.365 351.045 -129.035 ;
        RECT 350.715 -130.725 351.045 -130.395 ;
        RECT 350.715 -132.085 351.045 -131.755 ;
        RECT 350.715 -133.445 351.045 -133.115 ;
        RECT 350.715 -134.805 351.045 -134.475 ;
        RECT 350.715 -136.165 351.045 -135.835 ;
        RECT 350.715 -137.525 351.045 -137.195 ;
        RECT 350.715 -138.885 351.045 -138.555 ;
        RECT 350.715 -140.245 351.045 -139.915 ;
        RECT 350.715 -141.605 351.045 -141.275 ;
        RECT 350.715 -142.965 351.045 -142.635 ;
        RECT 350.715 -144.325 351.045 -143.995 ;
        RECT 350.715 -145.685 351.045 -145.355 ;
        RECT 350.715 -147.045 351.045 -146.715 ;
        RECT 350.715 -148.405 351.045 -148.075 ;
        RECT 350.715 -149.765 351.045 -149.435 ;
        RECT 350.715 -151.125 351.045 -150.795 ;
        RECT 350.715 -152.485 351.045 -152.155 ;
        RECT 350.715 -153.845 351.045 -153.515 ;
        RECT 350.715 -155.205 351.045 -154.875 ;
        RECT 350.715 -156.565 351.045 -156.235 ;
        RECT 350.715 -157.925 351.045 -157.595 ;
        RECT 350.715 -159.285 351.045 -158.955 ;
        RECT 350.715 -160.645 351.045 -160.315 ;
        RECT 350.715 -162.005 351.045 -161.675 ;
        RECT 350.715 -163.365 351.045 -163.035 ;
        RECT 350.715 -164.725 351.045 -164.395 ;
        RECT 350.715 -166.085 351.045 -165.755 ;
        RECT 350.715 -167.445 351.045 -167.115 ;
        RECT 350.715 -168.805 351.045 -168.475 ;
        RECT 350.715 -170.165 351.045 -169.835 ;
        RECT 350.715 -171.525 351.045 -171.195 ;
        RECT 350.715 -172.885 351.045 -172.555 ;
        RECT 350.715 -174.245 351.045 -173.915 ;
        RECT 350.715 -175.605 351.045 -175.275 ;
        RECT 350.715 -176.965 351.045 -176.635 ;
        RECT 350.715 -178.325 351.045 -177.995 ;
        RECT 350.715 -179.685 351.045 -179.355 ;
        RECT 350.715 -181.045 351.045 -180.715 ;
        RECT 350.715 -182.405 351.045 -182.075 ;
        RECT 350.715 -183.765 351.045 -183.435 ;
        RECT 350.715 -185.125 351.045 -184.795 ;
        RECT 350.715 -186.485 351.045 -186.155 ;
        RECT 350.715 -187.845 351.045 -187.515 ;
        RECT 350.715 -189.205 351.045 -188.875 ;
        RECT 350.715 -190.565 351.045 -190.235 ;
        RECT 350.715 -191.925 351.045 -191.595 ;
        RECT 350.715 -193.285 351.045 -192.955 ;
        RECT 350.715 -194.645 351.045 -194.315 ;
        RECT 350.715 -196.005 351.045 -195.675 ;
        RECT 350.715 -197.365 351.045 -197.035 ;
        RECT 350.715 -198.725 351.045 -198.395 ;
        RECT 350.715 -200.085 351.045 -199.755 ;
        RECT 350.715 -201.445 351.045 -201.115 ;
        RECT 350.715 -202.805 351.045 -202.475 ;
        RECT 350.715 -204.165 351.045 -203.835 ;
        RECT 350.715 -205.525 351.045 -205.195 ;
        RECT 350.715 -206.885 351.045 -206.555 ;
        RECT 350.715 -208.245 351.045 -207.915 ;
        RECT 350.715 -209.605 351.045 -209.275 ;
        RECT 350.715 -210.965 351.045 -210.635 ;
        RECT 350.715 -212.325 351.045 -211.995 ;
        RECT 350.715 -213.685 351.045 -213.355 ;
        RECT 350.715 -215.045 351.045 -214.715 ;
        RECT 350.715 -216.405 351.045 -216.075 ;
        RECT 350.715 -217.765 351.045 -217.435 ;
        RECT 350.715 -219.125 351.045 -218.795 ;
        RECT 350.715 -220.485 351.045 -220.155 ;
        RECT 350.715 -221.845 351.045 -221.515 ;
        RECT 350.715 -223.205 351.045 -222.875 ;
        RECT 350.715 -224.565 351.045 -224.235 ;
        RECT 350.715 -225.925 351.045 -225.595 ;
        RECT 350.715 -227.285 351.045 -226.955 ;
        RECT 350.715 -228.645 351.045 -228.315 ;
        RECT 350.715 -230.005 351.045 -229.675 ;
        RECT 350.715 -231.365 351.045 -231.035 ;
        RECT 350.715 -232.725 351.045 -232.395 ;
        RECT 350.715 -234.085 351.045 -233.755 ;
        RECT 350.715 -235.445 351.045 -235.115 ;
        RECT 350.715 -236.805 351.045 -236.475 ;
        RECT 350.715 -238.165 351.045 -237.835 ;
        RECT 350.715 -243.81 351.045 -242.68 ;
        RECT 350.72 -243.925 351.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 246.76 352.405 247.89 ;
        RECT 352.075 241.915 352.405 242.245 ;
        RECT 352.075 240.555 352.405 240.885 ;
        RECT 352.075 239.195 352.405 239.525 ;
        RECT 352.075 237.835 352.405 238.165 ;
        RECT 352.08 237.16 352.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 -126.645 352.405 -126.315 ;
        RECT 352.075 -128.005 352.405 -127.675 ;
        RECT 352.075 -129.365 352.405 -129.035 ;
        RECT 352.075 -130.725 352.405 -130.395 ;
        RECT 352.075 -132.085 352.405 -131.755 ;
        RECT 352.075 -133.445 352.405 -133.115 ;
        RECT 352.075 -134.805 352.405 -134.475 ;
        RECT 352.075 -136.165 352.405 -135.835 ;
        RECT 352.075 -137.525 352.405 -137.195 ;
        RECT 352.075 -138.885 352.405 -138.555 ;
        RECT 352.075 -140.245 352.405 -139.915 ;
        RECT 352.075 -141.605 352.405 -141.275 ;
        RECT 352.075 -142.965 352.405 -142.635 ;
        RECT 352.075 -144.325 352.405 -143.995 ;
        RECT 352.075 -145.685 352.405 -145.355 ;
        RECT 352.075 -147.045 352.405 -146.715 ;
        RECT 352.075 -148.405 352.405 -148.075 ;
        RECT 352.075 -149.765 352.405 -149.435 ;
        RECT 352.075 -151.125 352.405 -150.795 ;
        RECT 352.075 -152.485 352.405 -152.155 ;
        RECT 352.075 -153.845 352.405 -153.515 ;
        RECT 352.075 -155.205 352.405 -154.875 ;
        RECT 352.075 -156.565 352.405 -156.235 ;
        RECT 352.075 -157.925 352.405 -157.595 ;
        RECT 352.075 -159.285 352.405 -158.955 ;
        RECT 352.075 -160.645 352.405 -160.315 ;
        RECT 352.075 -162.005 352.405 -161.675 ;
        RECT 352.075 -163.365 352.405 -163.035 ;
        RECT 352.075 -164.725 352.405 -164.395 ;
        RECT 352.075 -166.085 352.405 -165.755 ;
        RECT 352.075 -167.445 352.405 -167.115 ;
        RECT 352.075 -168.805 352.405 -168.475 ;
        RECT 352.075 -170.165 352.405 -169.835 ;
        RECT 352.075 -171.525 352.405 -171.195 ;
        RECT 352.075 -172.885 352.405 -172.555 ;
        RECT 352.075 -174.245 352.405 -173.915 ;
        RECT 352.075 -175.605 352.405 -175.275 ;
        RECT 352.075 -176.965 352.405 -176.635 ;
        RECT 352.075 -178.325 352.405 -177.995 ;
        RECT 352.075 -179.685 352.405 -179.355 ;
        RECT 352.075 -181.045 352.405 -180.715 ;
        RECT 352.075 -182.405 352.405 -182.075 ;
        RECT 352.075 -183.765 352.405 -183.435 ;
        RECT 352.075 -185.125 352.405 -184.795 ;
        RECT 352.075 -186.485 352.405 -186.155 ;
        RECT 352.075 -187.845 352.405 -187.515 ;
        RECT 352.075 -189.205 352.405 -188.875 ;
        RECT 352.075 -190.565 352.405 -190.235 ;
        RECT 352.075 -191.925 352.405 -191.595 ;
        RECT 352.075 -193.285 352.405 -192.955 ;
        RECT 352.075 -194.645 352.405 -194.315 ;
        RECT 352.075 -196.005 352.405 -195.675 ;
        RECT 352.075 -197.365 352.405 -197.035 ;
        RECT 352.075 -198.725 352.405 -198.395 ;
        RECT 352.075 -200.085 352.405 -199.755 ;
        RECT 352.075 -201.445 352.405 -201.115 ;
        RECT 352.075 -202.805 352.405 -202.475 ;
        RECT 352.075 -204.165 352.405 -203.835 ;
        RECT 352.075 -205.525 352.405 -205.195 ;
        RECT 352.075 -206.885 352.405 -206.555 ;
        RECT 352.075 -208.245 352.405 -207.915 ;
        RECT 352.075 -209.605 352.405 -209.275 ;
        RECT 352.075 -210.965 352.405 -210.635 ;
        RECT 352.075 -212.325 352.405 -211.995 ;
        RECT 352.075 -213.685 352.405 -213.355 ;
        RECT 352.075 -215.045 352.405 -214.715 ;
        RECT 352.075 -216.405 352.405 -216.075 ;
        RECT 352.075 -217.765 352.405 -217.435 ;
        RECT 352.075 -219.125 352.405 -218.795 ;
        RECT 352.075 -220.485 352.405 -220.155 ;
        RECT 352.075 -221.845 352.405 -221.515 ;
        RECT 352.075 -223.205 352.405 -222.875 ;
        RECT 352.075 -224.565 352.405 -224.235 ;
        RECT 352.075 -225.925 352.405 -225.595 ;
        RECT 352.075 -227.285 352.405 -226.955 ;
        RECT 352.075 -228.645 352.405 -228.315 ;
        RECT 352.075 -230.005 352.405 -229.675 ;
        RECT 352.075 -231.365 352.405 -231.035 ;
        RECT 352.075 -232.725 352.405 -232.395 ;
        RECT 352.075 -234.085 352.405 -233.755 ;
        RECT 352.075 -235.445 352.405 -235.115 ;
        RECT 352.075 -236.805 352.405 -236.475 ;
        RECT 352.075 -238.165 352.405 -237.835 ;
        RECT 352.075 -243.81 352.405 -242.68 ;
        RECT 352.08 -243.925 352.4 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.11 -125.535 352.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 246.76 353.765 247.89 ;
        RECT 353.435 241.915 353.765 242.245 ;
        RECT 353.435 240.555 353.765 240.885 ;
        RECT 353.435 239.195 353.765 239.525 ;
        RECT 353.435 237.835 353.765 238.165 ;
        RECT 353.44 237.16 353.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 -1.525 353.765 -1.195 ;
        RECT 353.435 -2.885 353.765 -2.555 ;
        RECT 353.44 -3.56 353.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 -122.565 353.765 -122.235 ;
        RECT 353.435 -123.925 353.765 -123.595 ;
        RECT 353.435 -125.285 353.765 -124.955 ;
        RECT 353.435 -126.645 353.765 -126.315 ;
        RECT 353.435 -128.005 353.765 -127.675 ;
        RECT 353.435 -129.365 353.765 -129.035 ;
        RECT 353.435 -130.725 353.765 -130.395 ;
        RECT 353.435 -132.085 353.765 -131.755 ;
        RECT 353.435 -133.445 353.765 -133.115 ;
        RECT 353.435 -134.805 353.765 -134.475 ;
        RECT 353.435 -136.165 353.765 -135.835 ;
        RECT 353.435 -137.525 353.765 -137.195 ;
        RECT 353.435 -138.885 353.765 -138.555 ;
        RECT 353.435 -140.245 353.765 -139.915 ;
        RECT 353.435 -141.605 353.765 -141.275 ;
        RECT 353.435 -142.965 353.765 -142.635 ;
        RECT 353.435 -144.325 353.765 -143.995 ;
        RECT 353.435 -145.685 353.765 -145.355 ;
        RECT 353.435 -147.045 353.765 -146.715 ;
        RECT 353.435 -148.405 353.765 -148.075 ;
        RECT 353.435 -149.765 353.765 -149.435 ;
        RECT 353.435 -151.125 353.765 -150.795 ;
        RECT 353.435 -152.485 353.765 -152.155 ;
        RECT 353.435 -153.845 353.765 -153.515 ;
        RECT 353.435 -155.205 353.765 -154.875 ;
        RECT 353.435 -156.565 353.765 -156.235 ;
        RECT 353.435 -157.925 353.765 -157.595 ;
        RECT 353.435 -159.285 353.765 -158.955 ;
        RECT 353.435 -160.645 353.765 -160.315 ;
        RECT 353.435 -162.005 353.765 -161.675 ;
        RECT 353.435 -163.365 353.765 -163.035 ;
        RECT 353.435 -164.725 353.765 -164.395 ;
        RECT 353.435 -166.085 353.765 -165.755 ;
        RECT 353.435 -167.445 353.765 -167.115 ;
        RECT 353.435 -168.805 353.765 -168.475 ;
        RECT 353.435 -170.165 353.765 -169.835 ;
        RECT 353.435 -171.525 353.765 -171.195 ;
        RECT 353.435 -172.885 353.765 -172.555 ;
        RECT 353.435 -174.245 353.765 -173.915 ;
        RECT 353.435 -175.605 353.765 -175.275 ;
        RECT 353.435 -176.965 353.765 -176.635 ;
        RECT 353.435 -178.325 353.765 -177.995 ;
        RECT 353.435 -179.685 353.765 -179.355 ;
        RECT 353.435 -181.045 353.765 -180.715 ;
        RECT 353.435 -182.405 353.765 -182.075 ;
        RECT 353.435 -183.765 353.765 -183.435 ;
        RECT 353.435 -185.125 353.765 -184.795 ;
        RECT 353.435 -186.485 353.765 -186.155 ;
        RECT 353.435 -187.845 353.765 -187.515 ;
        RECT 353.435 -189.205 353.765 -188.875 ;
        RECT 353.435 -190.565 353.765 -190.235 ;
        RECT 353.435 -191.925 353.765 -191.595 ;
        RECT 353.435 -193.285 353.765 -192.955 ;
        RECT 353.435 -194.645 353.765 -194.315 ;
        RECT 353.435 -196.005 353.765 -195.675 ;
        RECT 353.435 -197.365 353.765 -197.035 ;
        RECT 353.435 -198.725 353.765 -198.395 ;
        RECT 353.435 -200.085 353.765 -199.755 ;
        RECT 353.435 -201.445 353.765 -201.115 ;
        RECT 353.435 -202.805 353.765 -202.475 ;
        RECT 353.435 -204.165 353.765 -203.835 ;
        RECT 353.435 -205.525 353.765 -205.195 ;
        RECT 353.435 -206.885 353.765 -206.555 ;
        RECT 353.435 -208.245 353.765 -207.915 ;
        RECT 353.435 -209.605 353.765 -209.275 ;
        RECT 353.435 -210.965 353.765 -210.635 ;
        RECT 353.435 -212.325 353.765 -211.995 ;
        RECT 353.435 -213.685 353.765 -213.355 ;
        RECT 353.435 -215.045 353.765 -214.715 ;
        RECT 353.435 -216.405 353.765 -216.075 ;
        RECT 353.435 -217.765 353.765 -217.435 ;
        RECT 353.435 -219.125 353.765 -218.795 ;
        RECT 353.435 -220.485 353.765 -220.155 ;
        RECT 353.435 -221.845 353.765 -221.515 ;
        RECT 353.435 -223.205 353.765 -222.875 ;
        RECT 353.435 -224.565 353.765 -224.235 ;
        RECT 353.435 -225.925 353.765 -225.595 ;
        RECT 353.435 -227.285 353.765 -226.955 ;
        RECT 353.435 -228.645 353.765 -228.315 ;
        RECT 353.435 -230.005 353.765 -229.675 ;
        RECT 353.435 -231.365 353.765 -231.035 ;
        RECT 353.435 -232.725 353.765 -232.395 ;
        RECT 353.435 -234.085 353.765 -233.755 ;
        RECT 353.435 -235.445 353.765 -235.115 ;
        RECT 353.435 -236.805 353.765 -236.475 ;
        RECT 353.435 -238.165 353.765 -237.835 ;
        RECT 353.435 -243.81 353.765 -242.68 ;
        RECT 353.44 -243.925 353.76 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 246.76 355.125 247.89 ;
        RECT 354.795 241.915 355.125 242.245 ;
        RECT 354.795 240.555 355.125 240.885 ;
        RECT 354.795 239.195 355.125 239.525 ;
        RECT 354.795 237.835 355.125 238.165 ;
        RECT 354.8 237.16 355.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 -1.525 355.125 -1.195 ;
        RECT 354.795 -2.885 355.125 -2.555 ;
        RECT 354.8 -3.56 355.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 -122.565 355.125 -122.235 ;
        RECT 354.795 -123.925 355.125 -123.595 ;
        RECT 354.795 -125.285 355.125 -124.955 ;
        RECT 354.795 -126.645 355.125 -126.315 ;
        RECT 354.795 -128.005 355.125 -127.675 ;
        RECT 354.795 -129.365 355.125 -129.035 ;
        RECT 354.795 -130.725 355.125 -130.395 ;
        RECT 354.795 -132.085 355.125 -131.755 ;
        RECT 354.795 -133.445 355.125 -133.115 ;
        RECT 354.795 -134.805 355.125 -134.475 ;
        RECT 354.795 -136.165 355.125 -135.835 ;
        RECT 354.795 -137.525 355.125 -137.195 ;
        RECT 354.795 -138.885 355.125 -138.555 ;
        RECT 354.795 -140.245 355.125 -139.915 ;
        RECT 354.795 -141.605 355.125 -141.275 ;
        RECT 354.795 -142.965 355.125 -142.635 ;
        RECT 354.795 -144.325 355.125 -143.995 ;
        RECT 354.795 -145.685 355.125 -145.355 ;
        RECT 354.795 -147.045 355.125 -146.715 ;
        RECT 354.795 -148.405 355.125 -148.075 ;
        RECT 354.795 -149.765 355.125 -149.435 ;
        RECT 354.795 -151.125 355.125 -150.795 ;
        RECT 354.795 -152.485 355.125 -152.155 ;
        RECT 354.795 -153.845 355.125 -153.515 ;
        RECT 354.795 -155.205 355.125 -154.875 ;
        RECT 354.795 -156.565 355.125 -156.235 ;
        RECT 354.795 -157.925 355.125 -157.595 ;
        RECT 354.795 -159.285 355.125 -158.955 ;
        RECT 354.795 -160.645 355.125 -160.315 ;
        RECT 354.795 -162.005 355.125 -161.675 ;
        RECT 354.795 -163.365 355.125 -163.035 ;
        RECT 354.795 -164.725 355.125 -164.395 ;
        RECT 354.795 -166.085 355.125 -165.755 ;
        RECT 354.795 -167.445 355.125 -167.115 ;
        RECT 354.795 -168.805 355.125 -168.475 ;
        RECT 354.795 -170.165 355.125 -169.835 ;
        RECT 354.795 -171.525 355.125 -171.195 ;
        RECT 354.795 -172.885 355.125 -172.555 ;
        RECT 354.795 -174.245 355.125 -173.915 ;
        RECT 354.795 -175.605 355.125 -175.275 ;
        RECT 354.795 -176.965 355.125 -176.635 ;
        RECT 354.795 -178.325 355.125 -177.995 ;
        RECT 354.795 -179.685 355.125 -179.355 ;
        RECT 354.795 -181.045 355.125 -180.715 ;
        RECT 354.795 -182.405 355.125 -182.075 ;
        RECT 354.795 -183.765 355.125 -183.435 ;
        RECT 354.795 -185.125 355.125 -184.795 ;
        RECT 354.795 -186.485 355.125 -186.155 ;
        RECT 354.795 -187.845 355.125 -187.515 ;
        RECT 354.795 -189.205 355.125 -188.875 ;
        RECT 354.795 -190.565 355.125 -190.235 ;
        RECT 354.795 -191.925 355.125 -191.595 ;
        RECT 354.795 -193.285 355.125 -192.955 ;
        RECT 354.795 -194.645 355.125 -194.315 ;
        RECT 354.795 -196.005 355.125 -195.675 ;
        RECT 354.795 -197.365 355.125 -197.035 ;
        RECT 354.795 -198.725 355.125 -198.395 ;
        RECT 354.795 -200.085 355.125 -199.755 ;
        RECT 354.795 -201.445 355.125 -201.115 ;
        RECT 354.795 -202.805 355.125 -202.475 ;
        RECT 354.795 -204.165 355.125 -203.835 ;
        RECT 354.795 -205.525 355.125 -205.195 ;
        RECT 354.795 -206.885 355.125 -206.555 ;
        RECT 354.795 -208.245 355.125 -207.915 ;
        RECT 354.795 -209.605 355.125 -209.275 ;
        RECT 354.795 -210.965 355.125 -210.635 ;
        RECT 354.795 -212.325 355.125 -211.995 ;
        RECT 354.795 -213.685 355.125 -213.355 ;
        RECT 354.795 -215.045 355.125 -214.715 ;
        RECT 354.795 -216.405 355.125 -216.075 ;
        RECT 354.795 -217.765 355.125 -217.435 ;
        RECT 354.795 -219.125 355.125 -218.795 ;
        RECT 354.795 -220.485 355.125 -220.155 ;
        RECT 354.795 -221.845 355.125 -221.515 ;
        RECT 354.795 -223.205 355.125 -222.875 ;
        RECT 354.795 -224.565 355.125 -224.235 ;
        RECT 354.795 -225.925 355.125 -225.595 ;
        RECT 354.795 -227.285 355.125 -226.955 ;
        RECT 354.795 -228.645 355.125 -228.315 ;
        RECT 354.795 -230.005 355.125 -229.675 ;
        RECT 354.795 -231.365 355.125 -231.035 ;
        RECT 354.795 -232.725 355.125 -232.395 ;
        RECT 354.795 -234.085 355.125 -233.755 ;
        RECT 354.795 -235.445 355.125 -235.115 ;
        RECT 354.795 -236.805 355.125 -236.475 ;
        RECT 354.795 -238.165 355.125 -237.835 ;
        RECT 354.795 -243.81 355.125 -242.68 ;
        RECT 354.8 -243.925 355.12 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.155 -190.565 356.485 -190.235 ;
        RECT 356.155 -191.925 356.485 -191.595 ;
        RECT 356.155 -193.285 356.485 -192.955 ;
        RECT 356.155 -194.645 356.485 -194.315 ;
        RECT 356.155 -196.005 356.485 -195.675 ;
        RECT 356.155 -197.365 356.485 -197.035 ;
        RECT 356.155 -198.725 356.485 -198.395 ;
        RECT 356.155 -200.085 356.485 -199.755 ;
        RECT 356.155 -201.445 356.485 -201.115 ;
        RECT 356.155 -202.805 356.485 -202.475 ;
        RECT 356.155 -204.165 356.485 -203.835 ;
        RECT 356.155 -205.525 356.485 -205.195 ;
        RECT 356.155 -206.885 356.485 -206.555 ;
        RECT 356.155 -208.245 356.485 -207.915 ;
        RECT 356.155 -209.605 356.485 -209.275 ;
        RECT 356.155 -210.965 356.485 -210.635 ;
        RECT 356.155 -212.325 356.485 -211.995 ;
        RECT 356.155 -213.685 356.485 -213.355 ;
        RECT 356.155 -215.045 356.485 -214.715 ;
        RECT 356.155 -216.405 356.485 -216.075 ;
        RECT 356.155 -217.765 356.485 -217.435 ;
        RECT 356.155 -219.125 356.485 -218.795 ;
        RECT 356.155 -220.485 356.485 -220.155 ;
        RECT 356.155 -221.845 356.485 -221.515 ;
        RECT 356.155 -223.205 356.485 -222.875 ;
        RECT 356.155 -224.565 356.485 -224.235 ;
        RECT 356.155 -225.925 356.485 -225.595 ;
        RECT 356.155 -227.285 356.485 -226.955 ;
        RECT 356.155 -228.645 356.485 -228.315 ;
        RECT 356.155 -230.005 356.485 -229.675 ;
        RECT 356.155 -231.365 356.485 -231.035 ;
        RECT 356.155 -232.725 356.485 -232.395 ;
        RECT 356.155 -234.085 356.485 -233.755 ;
        RECT 356.155 -235.445 356.485 -235.115 ;
        RECT 356.155 -236.805 356.485 -236.475 ;
        RECT 356.155 -238.165 356.485 -237.835 ;
        RECT 356.155 -243.81 356.485 -242.68 ;
        RECT 356.16 -243.925 356.48 248.005 ;
        RECT 356.155 246.76 356.485 247.89 ;
        RECT 356.155 241.915 356.485 242.245 ;
        RECT 356.155 240.555 356.485 240.885 ;
        RECT 356.155 239.195 356.485 239.525 ;
        RECT 356.155 237.835 356.485 238.165 ;
        RECT 356.155 235.17 356.485 235.5 ;
        RECT 356.155 232.995 356.485 233.325 ;
        RECT 356.155 231.415 356.485 231.745 ;
        RECT 356.155 230.565 356.485 230.895 ;
        RECT 356.155 228.255 356.485 228.585 ;
        RECT 356.155 227.405 356.485 227.735 ;
        RECT 356.155 225.095 356.485 225.425 ;
        RECT 356.155 224.245 356.485 224.575 ;
        RECT 356.155 221.935 356.485 222.265 ;
        RECT 356.155 221.085 356.485 221.415 ;
        RECT 356.155 218.775 356.485 219.105 ;
        RECT 356.155 217.195 356.485 217.525 ;
        RECT 356.155 216.345 356.485 216.675 ;
        RECT 356.155 214.035 356.485 214.365 ;
        RECT 356.155 213.185 356.485 213.515 ;
        RECT 356.155 210.875 356.485 211.205 ;
        RECT 356.155 210.025 356.485 210.355 ;
        RECT 356.155 207.715 356.485 208.045 ;
        RECT 356.155 206.865 356.485 207.195 ;
        RECT 356.155 204.555 356.485 204.885 ;
        RECT 356.155 202.975 356.485 203.305 ;
        RECT 356.155 202.125 356.485 202.455 ;
        RECT 356.155 199.815 356.485 200.145 ;
        RECT 356.155 198.965 356.485 199.295 ;
        RECT 356.155 196.655 356.485 196.985 ;
        RECT 356.155 195.805 356.485 196.135 ;
        RECT 356.155 193.495 356.485 193.825 ;
        RECT 356.155 192.645 356.485 192.975 ;
        RECT 356.155 190.335 356.485 190.665 ;
        RECT 356.155 188.755 356.485 189.085 ;
        RECT 356.155 187.905 356.485 188.235 ;
        RECT 356.155 185.595 356.485 185.925 ;
        RECT 356.155 184.745 356.485 185.075 ;
        RECT 356.155 182.435 356.485 182.765 ;
        RECT 356.155 181.585 356.485 181.915 ;
        RECT 356.155 179.275 356.485 179.605 ;
        RECT 356.155 178.425 356.485 178.755 ;
        RECT 356.155 176.115 356.485 176.445 ;
        RECT 356.155 174.535 356.485 174.865 ;
        RECT 356.155 173.685 356.485 174.015 ;
        RECT 356.155 171.375 356.485 171.705 ;
        RECT 356.155 170.525 356.485 170.855 ;
        RECT 356.155 168.215 356.485 168.545 ;
        RECT 356.155 167.365 356.485 167.695 ;
        RECT 356.155 165.055 356.485 165.385 ;
        RECT 356.155 164.205 356.485 164.535 ;
        RECT 356.155 161.895 356.485 162.225 ;
        RECT 356.155 160.315 356.485 160.645 ;
        RECT 356.155 159.465 356.485 159.795 ;
        RECT 356.155 157.155 356.485 157.485 ;
        RECT 356.155 156.305 356.485 156.635 ;
        RECT 356.155 153.995 356.485 154.325 ;
        RECT 356.155 153.145 356.485 153.475 ;
        RECT 356.155 150.835 356.485 151.165 ;
        RECT 356.155 149.985 356.485 150.315 ;
        RECT 356.155 147.675 356.485 148.005 ;
        RECT 356.155 146.095 356.485 146.425 ;
        RECT 356.155 145.245 356.485 145.575 ;
        RECT 356.155 142.935 356.485 143.265 ;
        RECT 356.155 142.085 356.485 142.415 ;
        RECT 356.155 139.775 356.485 140.105 ;
        RECT 356.155 138.925 356.485 139.255 ;
        RECT 356.155 136.615 356.485 136.945 ;
        RECT 356.155 135.765 356.485 136.095 ;
        RECT 356.155 133.455 356.485 133.785 ;
        RECT 356.155 131.875 356.485 132.205 ;
        RECT 356.155 131.025 356.485 131.355 ;
        RECT 356.155 128.715 356.485 129.045 ;
        RECT 356.155 127.865 356.485 128.195 ;
        RECT 356.155 125.555 356.485 125.885 ;
        RECT 356.155 124.705 356.485 125.035 ;
        RECT 356.155 122.395 356.485 122.725 ;
        RECT 356.155 121.545 356.485 121.875 ;
        RECT 356.155 119.235 356.485 119.565 ;
        RECT 356.155 117.655 356.485 117.985 ;
        RECT 356.155 116.805 356.485 117.135 ;
        RECT 356.155 114.495 356.485 114.825 ;
        RECT 356.155 113.645 356.485 113.975 ;
        RECT 356.155 111.335 356.485 111.665 ;
        RECT 356.155 110.485 356.485 110.815 ;
        RECT 356.155 108.175 356.485 108.505 ;
        RECT 356.155 107.325 356.485 107.655 ;
        RECT 356.155 105.015 356.485 105.345 ;
        RECT 356.155 103.435 356.485 103.765 ;
        RECT 356.155 102.585 356.485 102.915 ;
        RECT 356.155 100.275 356.485 100.605 ;
        RECT 356.155 99.425 356.485 99.755 ;
        RECT 356.155 97.115 356.485 97.445 ;
        RECT 356.155 96.265 356.485 96.595 ;
        RECT 356.155 93.955 356.485 94.285 ;
        RECT 356.155 93.105 356.485 93.435 ;
        RECT 356.155 90.795 356.485 91.125 ;
        RECT 356.155 89.215 356.485 89.545 ;
        RECT 356.155 88.365 356.485 88.695 ;
        RECT 356.155 86.055 356.485 86.385 ;
        RECT 356.155 85.205 356.485 85.535 ;
        RECT 356.155 82.895 356.485 83.225 ;
        RECT 356.155 82.045 356.485 82.375 ;
        RECT 356.155 79.735 356.485 80.065 ;
        RECT 356.155 78.885 356.485 79.215 ;
        RECT 356.155 76.575 356.485 76.905 ;
        RECT 356.155 74.995 356.485 75.325 ;
        RECT 356.155 74.145 356.485 74.475 ;
        RECT 356.155 71.835 356.485 72.165 ;
        RECT 356.155 70.985 356.485 71.315 ;
        RECT 356.155 68.675 356.485 69.005 ;
        RECT 356.155 67.825 356.485 68.155 ;
        RECT 356.155 65.515 356.485 65.845 ;
        RECT 356.155 64.665 356.485 64.995 ;
        RECT 356.155 62.355 356.485 62.685 ;
        RECT 356.155 60.775 356.485 61.105 ;
        RECT 356.155 59.925 356.485 60.255 ;
        RECT 356.155 57.615 356.485 57.945 ;
        RECT 356.155 56.765 356.485 57.095 ;
        RECT 356.155 54.455 356.485 54.785 ;
        RECT 356.155 53.605 356.485 53.935 ;
        RECT 356.155 51.295 356.485 51.625 ;
        RECT 356.155 50.445 356.485 50.775 ;
        RECT 356.155 48.135 356.485 48.465 ;
        RECT 356.155 46.555 356.485 46.885 ;
        RECT 356.155 45.705 356.485 46.035 ;
        RECT 356.155 43.395 356.485 43.725 ;
        RECT 356.155 42.545 356.485 42.875 ;
        RECT 356.155 40.235 356.485 40.565 ;
        RECT 356.155 39.385 356.485 39.715 ;
        RECT 356.155 37.075 356.485 37.405 ;
        RECT 356.155 36.225 356.485 36.555 ;
        RECT 356.155 33.915 356.485 34.245 ;
        RECT 356.155 32.335 356.485 32.665 ;
        RECT 356.155 31.485 356.485 31.815 ;
        RECT 356.155 29.175 356.485 29.505 ;
        RECT 356.155 28.325 356.485 28.655 ;
        RECT 356.155 26.015 356.485 26.345 ;
        RECT 356.155 25.165 356.485 25.495 ;
        RECT 356.155 22.855 356.485 23.185 ;
        RECT 356.155 22.005 356.485 22.335 ;
        RECT 356.155 19.695 356.485 20.025 ;
        RECT 356.155 18.115 356.485 18.445 ;
        RECT 356.155 17.265 356.485 17.595 ;
        RECT 356.155 14.955 356.485 15.285 ;
        RECT 356.155 14.105 356.485 14.435 ;
        RECT 356.155 11.795 356.485 12.125 ;
        RECT 356.155 10.945 356.485 11.275 ;
        RECT 356.155 8.635 356.485 8.965 ;
        RECT 356.155 7.785 356.485 8.115 ;
        RECT 356.155 5.475 356.485 5.805 ;
        RECT 356.155 3.895 356.485 4.225 ;
        RECT 356.155 3.045 356.485 3.375 ;
        RECT 356.155 0.87 356.485 1.2 ;
        RECT 356.155 -1.525 356.485 -1.195 ;
        RECT 356.155 -2.885 356.485 -2.555 ;
        RECT 356.155 -4.245 356.485 -3.915 ;
        RECT 356.155 -5.605 356.485 -5.275 ;
        RECT 356.155 -6.965 356.485 -6.635 ;
        RECT 356.155 -8.325 356.485 -7.995 ;
        RECT 356.155 -9.685 356.485 -9.355 ;
        RECT 356.155 -11.045 356.485 -10.715 ;
        RECT 356.155 -12.405 356.485 -12.075 ;
        RECT 356.155 -13.765 356.485 -13.435 ;
        RECT 356.155 -15.125 356.485 -14.795 ;
        RECT 356.155 -16.485 356.485 -16.155 ;
        RECT 356.155 -17.845 356.485 -17.515 ;
        RECT 356.155 -19.205 356.485 -18.875 ;
        RECT 356.155 -20.565 356.485 -20.235 ;
        RECT 356.155 -21.925 356.485 -21.595 ;
        RECT 356.155 -23.285 356.485 -22.955 ;
        RECT 356.155 -24.645 356.485 -24.315 ;
        RECT 356.155 -26.005 356.485 -25.675 ;
        RECT 356.155 -27.365 356.485 -27.035 ;
        RECT 356.155 -28.725 356.485 -28.395 ;
        RECT 356.155 -30.085 356.485 -29.755 ;
        RECT 356.155 -31.445 356.485 -31.115 ;
        RECT 356.155 -32.805 356.485 -32.475 ;
        RECT 356.155 -34.165 356.485 -33.835 ;
        RECT 356.155 -35.525 356.485 -35.195 ;
        RECT 356.155 -36.885 356.485 -36.555 ;
        RECT 356.155 -38.245 356.485 -37.915 ;
        RECT 356.155 -39.605 356.485 -39.275 ;
        RECT 356.155 -40.965 356.485 -40.635 ;
        RECT 356.155 -42.325 356.485 -41.995 ;
        RECT 356.155 -43.685 356.485 -43.355 ;
        RECT 356.155 -45.045 356.485 -44.715 ;
        RECT 356.155 -46.405 356.485 -46.075 ;
        RECT 356.155 -47.765 356.485 -47.435 ;
        RECT 356.155 -49.125 356.485 -48.795 ;
        RECT 356.155 -50.485 356.485 -50.155 ;
        RECT 356.155 -51.845 356.485 -51.515 ;
        RECT 356.155 -53.205 356.485 -52.875 ;
        RECT 356.155 -54.565 356.485 -54.235 ;
        RECT 356.155 -55.925 356.485 -55.595 ;
        RECT 356.155 -57.285 356.485 -56.955 ;
        RECT 356.155 -58.645 356.485 -58.315 ;
        RECT 356.155 -60.005 356.485 -59.675 ;
        RECT 356.155 -61.365 356.485 -61.035 ;
        RECT 356.155 -62.725 356.485 -62.395 ;
        RECT 356.155 -64.085 356.485 -63.755 ;
        RECT 356.155 -65.445 356.485 -65.115 ;
        RECT 356.155 -66.805 356.485 -66.475 ;
        RECT 356.155 -68.165 356.485 -67.835 ;
        RECT 356.155 -69.525 356.485 -69.195 ;
        RECT 356.155 -70.885 356.485 -70.555 ;
        RECT 356.155 -72.245 356.485 -71.915 ;
        RECT 356.155 -73.605 356.485 -73.275 ;
        RECT 356.155 -74.965 356.485 -74.635 ;
        RECT 356.155 -76.325 356.485 -75.995 ;
        RECT 356.155 -77.685 356.485 -77.355 ;
        RECT 356.155 -79.045 356.485 -78.715 ;
        RECT 356.155 -80.405 356.485 -80.075 ;
        RECT 356.155 -81.765 356.485 -81.435 ;
        RECT 356.155 -83.125 356.485 -82.795 ;
        RECT 356.155 -84.485 356.485 -84.155 ;
        RECT 356.155 -85.845 356.485 -85.515 ;
        RECT 356.155 -87.205 356.485 -86.875 ;
        RECT 356.155 -88.565 356.485 -88.235 ;
        RECT 356.155 -89.925 356.485 -89.595 ;
        RECT 356.155 -91.285 356.485 -90.955 ;
        RECT 356.155 -92.645 356.485 -92.315 ;
        RECT 356.155 -94.005 356.485 -93.675 ;
        RECT 356.155 -95.365 356.485 -95.035 ;
        RECT 356.155 -96.725 356.485 -96.395 ;
        RECT 356.155 -98.085 356.485 -97.755 ;
        RECT 356.155 -99.445 356.485 -99.115 ;
        RECT 356.155 -100.805 356.485 -100.475 ;
        RECT 356.155 -102.165 356.485 -101.835 ;
        RECT 356.155 -103.525 356.485 -103.195 ;
        RECT 356.155 -104.885 356.485 -104.555 ;
        RECT 356.155 -106.245 356.485 -105.915 ;
        RECT 356.155 -107.605 356.485 -107.275 ;
        RECT 356.155 -108.965 356.485 -108.635 ;
        RECT 356.155 -110.325 356.485 -109.995 ;
        RECT 356.155 -111.685 356.485 -111.355 ;
        RECT 356.155 -113.045 356.485 -112.715 ;
        RECT 356.155 -114.405 356.485 -114.075 ;
        RECT 356.155 -115.765 356.485 -115.435 ;
        RECT 356.155 -117.125 356.485 -116.795 ;
        RECT 356.155 -118.485 356.485 -118.155 ;
        RECT 356.155 -119.845 356.485 -119.515 ;
        RECT 356.155 -121.205 356.485 -120.875 ;
        RECT 356.155 -122.565 356.485 -122.235 ;
        RECT 356.155 -123.925 356.485 -123.595 ;
        RECT 356.155 -125.285 356.485 -124.955 ;
        RECT 356.155 -126.645 356.485 -126.315 ;
        RECT 356.155 -128.005 356.485 -127.675 ;
        RECT 356.155 -129.365 356.485 -129.035 ;
        RECT 356.155 -130.725 356.485 -130.395 ;
        RECT 356.155 -132.085 356.485 -131.755 ;
        RECT 356.155 -133.445 356.485 -133.115 ;
        RECT 356.155 -134.805 356.485 -134.475 ;
        RECT 356.155 -136.165 356.485 -135.835 ;
        RECT 356.155 -137.525 356.485 -137.195 ;
        RECT 356.155 -138.885 356.485 -138.555 ;
        RECT 356.155 -140.245 356.485 -139.915 ;
        RECT 356.155 -141.605 356.485 -141.275 ;
        RECT 356.155 -142.965 356.485 -142.635 ;
        RECT 356.155 -144.325 356.485 -143.995 ;
        RECT 356.155 -145.685 356.485 -145.355 ;
        RECT 356.155 -147.045 356.485 -146.715 ;
        RECT 356.155 -148.405 356.485 -148.075 ;
        RECT 356.155 -149.765 356.485 -149.435 ;
        RECT 356.155 -151.125 356.485 -150.795 ;
        RECT 356.155 -152.485 356.485 -152.155 ;
        RECT 356.155 -153.845 356.485 -153.515 ;
        RECT 356.155 -155.205 356.485 -154.875 ;
        RECT 356.155 -156.565 356.485 -156.235 ;
        RECT 356.155 -157.925 356.485 -157.595 ;
        RECT 356.155 -159.285 356.485 -158.955 ;
        RECT 356.155 -160.645 356.485 -160.315 ;
        RECT 356.155 -162.005 356.485 -161.675 ;
        RECT 356.155 -163.365 356.485 -163.035 ;
        RECT 356.155 -164.725 356.485 -164.395 ;
        RECT 356.155 -166.085 356.485 -165.755 ;
        RECT 356.155 -167.445 356.485 -167.115 ;
        RECT 356.155 -168.805 356.485 -168.475 ;
        RECT 356.155 -170.165 356.485 -169.835 ;
        RECT 356.155 -171.525 356.485 -171.195 ;
        RECT 356.155 -172.885 356.485 -172.555 ;
        RECT 356.155 -174.245 356.485 -173.915 ;
        RECT 356.155 -175.605 356.485 -175.275 ;
        RECT 356.155 -176.965 356.485 -176.635 ;
        RECT 356.155 -178.325 356.485 -177.995 ;
        RECT 356.155 -179.685 356.485 -179.355 ;
        RECT 356.155 -181.045 356.485 -180.715 ;
        RECT 356.155 -182.405 356.485 -182.075 ;
        RECT 356.155 -183.765 356.485 -183.435 ;
        RECT 356.155 -185.125 356.485 -184.795 ;
        RECT 356.155 -186.485 356.485 -186.155 ;
        RECT 356.155 -187.845 356.485 -187.515 ;
        RECT 356.155 -189.205 356.485 -188.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 246.76 323.845 247.89 ;
        RECT 323.515 241.915 323.845 242.245 ;
        RECT 323.515 240.555 323.845 240.885 ;
        RECT 323.515 239.195 323.845 239.525 ;
        RECT 323.515 237.835 323.845 238.165 ;
        RECT 323.52 237.16 323.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 -1.525 323.845 -1.195 ;
        RECT 323.515 -2.885 323.845 -2.555 ;
        RECT 323.52 -3.56 323.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 -122.565 323.845 -122.235 ;
        RECT 323.515 -123.925 323.845 -123.595 ;
        RECT 323.515 -125.285 323.845 -124.955 ;
        RECT 323.515 -126.645 323.845 -126.315 ;
        RECT 323.515 -128.005 323.845 -127.675 ;
        RECT 323.515 -129.365 323.845 -129.035 ;
        RECT 323.515 -130.725 323.845 -130.395 ;
        RECT 323.515 -132.085 323.845 -131.755 ;
        RECT 323.515 -133.445 323.845 -133.115 ;
        RECT 323.515 -134.805 323.845 -134.475 ;
        RECT 323.515 -136.165 323.845 -135.835 ;
        RECT 323.515 -137.525 323.845 -137.195 ;
        RECT 323.515 -138.885 323.845 -138.555 ;
        RECT 323.515 -140.245 323.845 -139.915 ;
        RECT 323.515 -141.605 323.845 -141.275 ;
        RECT 323.515 -142.965 323.845 -142.635 ;
        RECT 323.515 -144.325 323.845 -143.995 ;
        RECT 323.515 -145.685 323.845 -145.355 ;
        RECT 323.515 -147.045 323.845 -146.715 ;
        RECT 323.515 -148.405 323.845 -148.075 ;
        RECT 323.515 -149.765 323.845 -149.435 ;
        RECT 323.515 -151.125 323.845 -150.795 ;
        RECT 323.515 -152.485 323.845 -152.155 ;
        RECT 323.515 -153.845 323.845 -153.515 ;
        RECT 323.515 -155.205 323.845 -154.875 ;
        RECT 323.515 -156.565 323.845 -156.235 ;
        RECT 323.515 -157.925 323.845 -157.595 ;
        RECT 323.515 -159.285 323.845 -158.955 ;
        RECT 323.515 -160.645 323.845 -160.315 ;
        RECT 323.515 -162.005 323.845 -161.675 ;
        RECT 323.515 -163.365 323.845 -163.035 ;
        RECT 323.515 -164.725 323.845 -164.395 ;
        RECT 323.515 -166.085 323.845 -165.755 ;
        RECT 323.515 -167.445 323.845 -167.115 ;
        RECT 323.515 -168.805 323.845 -168.475 ;
        RECT 323.515 -170.165 323.845 -169.835 ;
        RECT 323.515 -171.525 323.845 -171.195 ;
        RECT 323.515 -172.885 323.845 -172.555 ;
        RECT 323.515 -174.245 323.845 -173.915 ;
        RECT 323.515 -175.605 323.845 -175.275 ;
        RECT 323.515 -176.965 323.845 -176.635 ;
        RECT 323.515 -178.325 323.845 -177.995 ;
        RECT 323.515 -179.685 323.845 -179.355 ;
        RECT 323.515 -181.045 323.845 -180.715 ;
        RECT 323.515 -182.405 323.845 -182.075 ;
        RECT 323.515 -183.765 323.845 -183.435 ;
        RECT 323.515 -185.125 323.845 -184.795 ;
        RECT 323.515 -186.485 323.845 -186.155 ;
        RECT 323.515 -187.845 323.845 -187.515 ;
        RECT 323.515 -189.205 323.845 -188.875 ;
        RECT 323.515 -190.565 323.845 -190.235 ;
        RECT 323.515 -191.925 323.845 -191.595 ;
        RECT 323.515 -193.285 323.845 -192.955 ;
        RECT 323.515 -194.645 323.845 -194.315 ;
        RECT 323.515 -196.005 323.845 -195.675 ;
        RECT 323.515 -197.365 323.845 -197.035 ;
        RECT 323.515 -198.725 323.845 -198.395 ;
        RECT 323.515 -200.085 323.845 -199.755 ;
        RECT 323.515 -201.445 323.845 -201.115 ;
        RECT 323.515 -202.805 323.845 -202.475 ;
        RECT 323.515 -204.165 323.845 -203.835 ;
        RECT 323.515 -205.525 323.845 -205.195 ;
        RECT 323.515 -206.885 323.845 -206.555 ;
        RECT 323.515 -208.245 323.845 -207.915 ;
        RECT 323.515 -209.605 323.845 -209.275 ;
        RECT 323.515 -210.965 323.845 -210.635 ;
        RECT 323.515 -212.325 323.845 -211.995 ;
        RECT 323.515 -213.685 323.845 -213.355 ;
        RECT 323.515 -215.045 323.845 -214.715 ;
        RECT 323.515 -216.405 323.845 -216.075 ;
        RECT 323.515 -217.765 323.845 -217.435 ;
        RECT 323.515 -219.125 323.845 -218.795 ;
        RECT 323.515 -220.485 323.845 -220.155 ;
        RECT 323.515 -221.845 323.845 -221.515 ;
        RECT 323.515 -223.205 323.845 -222.875 ;
        RECT 323.515 -224.565 323.845 -224.235 ;
        RECT 323.515 -225.925 323.845 -225.595 ;
        RECT 323.515 -227.285 323.845 -226.955 ;
        RECT 323.515 -228.645 323.845 -228.315 ;
        RECT 323.515 -230.005 323.845 -229.675 ;
        RECT 323.515 -231.365 323.845 -231.035 ;
        RECT 323.515 -232.725 323.845 -232.395 ;
        RECT 323.515 -234.085 323.845 -233.755 ;
        RECT 323.515 -235.445 323.845 -235.115 ;
        RECT 323.515 -236.805 323.845 -236.475 ;
        RECT 323.515 -238.165 323.845 -237.835 ;
        RECT 323.515 -243.81 323.845 -242.68 ;
        RECT 323.52 -243.925 323.84 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 246.76 325.205 247.89 ;
        RECT 324.875 241.915 325.205 242.245 ;
        RECT 324.875 240.555 325.205 240.885 ;
        RECT 324.875 239.195 325.205 239.525 ;
        RECT 324.875 237.835 325.205 238.165 ;
        RECT 324.88 237.16 325.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 -1.525 325.205 -1.195 ;
        RECT 324.875 -2.885 325.205 -2.555 ;
        RECT 324.88 -3.56 325.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 -122.565 325.205 -122.235 ;
        RECT 324.875 -123.925 325.205 -123.595 ;
        RECT 324.875 -125.285 325.205 -124.955 ;
        RECT 324.875 -126.645 325.205 -126.315 ;
        RECT 324.875 -128.005 325.205 -127.675 ;
        RECT 324.875 -129.365 325.205 -129.035 ;
        RECT 324.875 -130.725 325.205 -130.395 ;
        RECT 324.875 -132.085 325.205 -131.755 ;
        RECT 324.875 -133.445 325.205 -133.115 ;
        RECT 324.875 -134.805 325.205 -134.475 ;
        RECT 324.875 -136.165 325.205 -135.835 ;
        RECT 324.875 -137.525 325.205 -137.195 ;
        RECT 324.875 -138.885 325.205 -138.555 ;
        RECT 324.875 -140.245 325.205 -139.915 ;
        RECT 324.875 -141.605 325.205 -141.275 ;
        RECT 324.875 -142.965 325.205 -142.635 ;
        RECT 324.875 -144.325 325.205 -143.995 ;
        RECT 324.875 -145.685 325.205 -145.355 ;
        RECT 324.875 -147.045 325.205 -146.715 ;
        RECT 324.875 -148.405 325.205 -148.075 ;
        RECT 324.875 -149.765 325.205 -149.435 ;
        RECT 324.875 -151.125 325.205 -150.795 ;
        RECT 324.875 -152.485 325.205 -152.155 ;
        RECT 324.875 -153.845 325.205 -153.515 ;
        RECT 324.875 -155.205 325.205 -154.875 ;
        RECT 324.875 -156.565 325.205 -156.235 ;
        RECT 324.875 -157.925 325.205 -157.595 ;
        RECT 324.875 -159.285 325.205 -158.955 ;
        RECT 324.875 -160.645 325.205 -160.315 ;
        RECT 324.875 -162.005 325.205 -161.675 ;
        RECT 324.875 -163.365 325.205 -163.035 ;
        RECT 324.875 -164.725 325.205 -164.395 ;
        RECT 324.875 -166.085 325.205 -165.755 ;
        RECT 324.875 -167.445 325.205 -167.115 ;
        RECT 324.875 -168.805 325.205 -168.475 ;
        RECT 324.875 -170.165 325.205 -169.835 ;
        RECT 324.875 -171.525 325.205 -171.195 ;
        RECT 324.875 -172.885 325.205 -172.555 ;
        RECT 324.875 -174.245 325.205 -173.915 ;
        RECT 324.875 -175.605 325.205 -175.275 ;
        RECT 324.875 -176.965 325.205 -176.635 ;
        RECT 324.875 -178.325 325.205 -177.995 ;
        RECT 324.875 -179.685 325.205 -179.355 ;
        RECT 324.875 -181.045 325.205 -180.715 ;
        RECT 324.875 -182.405 325.205 -182.075 ;
        RECT 324.875 -183.765 325.205 -183.435 ;
        RECT 324.875 -185.125 325.205 -184.795 ;
        RECT 324.875 -186.485 325.205 -186.155 ;
        RECT 324.875 -187.845 325.205 -187.515 ;
        RECT 324.875 -189.205 325.205 -188.875 ;
        RECT 324.875 -190.565 325.205 -190.235 ;
        RECT 324.875 -191.925 325.205 -191.595 ;
        RECT 324.875 -193.285 325.205 -192.955 ;
        RECT 324.875 -194.645 325.205 -194.315 ;
        RECT 324.875 -196.005 325.205 -195.675 ;
        RECT 324.875 -197.365 325.205 -197.035 ;
        RECT 324.875 -198.725 325.205 -198.395 ;
        RECT 324.875 -200.085 325.205 -199.755 ;
        RECT 324.875 -201.445 325.205 -201.115 ;
        RECT 324.875 -202.805 325.205 -202.475 ;
        RECT 324.875 -204.165 325.205 -203.835 ;
        RECT 324.875 -205.525 325.205 -205.195 ;
        RECT 324.875 -206.885 325.205 -206.555 ;
        RECT 324.875 -208.245 325.205 -207.915 ;
        RECT 324.875 -209.605 325.205 -209.275 ;
        RECT 324.875 -210.965 325.205 -210.635 ;
        RECT 324.875 -212.325 325.205 -211.995 ;
        RECT 324.875 -213.685 325.205 -213.355 ;
        RECT 324.875 -215.045 325.205 -214.715 ;
        RECT 324.875 -216.405 325.205 -216.075 ;
        RECT 324.875 -217.765 325.205 -217.435 ;
        RECT 324.875 -219.125 325.205 -218.795 ;
        RECT 324.875 -220.485 325.205 -220.155 ;
        RECT 324.875 -221.845 325.205 -221.515 ;
        RECT 324.875 -223.205 325.205 -222.875 ;
        RECT 324.875 -224.565 325.205 -224.235 ;
        RECT 324.875 -225.925 325.205 -225.595 ;
        RECT 324.875 -227.285 325.205 -226.955 ;
        RECT 324.875 -228.645 325.205 -228.315 ;
        RECT 324.875 -230.005 325.205 -229.675 ;
        RECT 324.875 -231.365 325.205 -231.035 ;
        RECT 324.875 -232.725 325.205 -232.395 ;
        RECT 324.875 -234.085 325.205 -233.755 ;
        RECT 324.875 -235.445 325.205 -235.115 ;
        RECT 324.875 -236.805 325.205 -236.475 ;
        RECT 324.875 -238.165 325.205 -237.835 ;
        RECT 324.875 -243.81 325.205 -242.68 ;
        RECT 324.88 -243.925 325.2 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 246.76 326.565 247.89 ;
        RECT 326.235 241.915 326.565 242.245 ;
        RECT 326.235 240.555 326.565 240.885 ;
        RECT 326.235 239.195 326.565 239.525 ;
        RECT 326.235 237.835 326.565 238.165 ;
        RECT 326.24 237.16 326.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 -1.525 326.565 -1.195 ;
        RECT 326.235 -2.885 326.565 -2.555 ;
        RECT 326.24 -3.56 326.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 -122.565 326.565 -122.235 ;
        RECT 326.235 -123.925 326.565 -123.595 ;
        RECT 326.235 -125.285 326.565 -124.955 ;
        RECT 326.235 -126.645 326.565 -126.315 ;
        RECT 326.235 -128.005 326.565 -127.675 ;
        RECT 326.235 -129.365 326.565 -129.035 ;
        RECT 326.235 -130.725 326.565 -130.395 ;
        RECT 326.235 -132.085 326.565 -131.755 ;
        RECT 326.235 -133.445 326.565 -133.115 ;
        RECT 326.235 -134.805 326.565 -134.475 ;
        RECT 326.235 -136.165 326.565 -135.835 ;
        RECT 326.235 -137.525 326.565 -137.195 ;
        RECT 326.235 -138.885 326.565 -138.555 ;
        RECT 326.235 -140.245 326.565 -139.915 ;
        RECT 326.235 -141.605 326.565 -141.275 ;
        RECT 326.235 -142.965 326.565 -142.635 ;
        RECT 326.235 -144.325 326.565 -143.995 ;
        RECT 326.235 -145.685 326.565 -145.355 ;
        RECT 326.235 -147.045 326.565 -146.715 ;
        RECT 326.235 -148.405 326.565 -148.075 ;
        RECT 326.235 -149.765 326.565 -149.435 ;
        RECT 326.235 -151.125 326.565 -150.795 ;
        RECT 326.235 -152.485 326.565 -152.155 ;
        RECT 326.235 -153.845 326.565 -153.515 ;
        RECT 326.235 -155.205 326.565 -154.875 ;
        RECT 326.235 -156.565 326.565 -156.235 ;
        RECT 326.235 -157.925 326.565 -157.595 ;
        RECT 326.235 -159.285 326.565 -158.955 ;
        RECT 326.235 -160.645 326.565 -160.315 ;
        RECT 326.235 -162.005 326.565 -161.675 ;
        RECT 326.235 -163.365 326.565 -163.035 ;
        RECT 326.235 -164.725 326.565 -164.395 ;
        RECT 326.235 -166.085 326.565 -165.755 ;
        RECT 326.235 -167.445 326.565 -167.115 ;
        RECT 326.235 -168.805 326.565 -168.475 ;
        RECT 326.235 -170.165 326.565 -169.835 ;
        RECT 326.235 -171.525 326.565 -171.195 ;
        RECT 326.235 -172.885 326.565 -172.555 ;
        RECT 326.235 -174.245 326.565 -173.915 ;
        RECT 326.235 -175.605 326.565 -175.275 ;
        RECT 326.235 -176.965 326.565 -176.635 ;
        RECT 326.235 -178.325 326.565 -177.995 ;
        RECT 326.235 -179.685 326.565 -179.355 ;
        RECT 326.235 -181.045 326.565 -180.715 ;
        RECT 326.235 -182.405 326.565 -182.075 ;
        RECT 326.235 -183.765 326.565 -183.435 ;
        RECT 326.235 -185.125 326.565 -184.795 ;
        RECT 326.235 -186.485 326.565 -186.155 ;
        RECT 326.235 -187.845 326.565 -187.515 ;
        RECT 326.235 -189.205 326.565 -188.875 ;
        RECT 326.235 -190.565 326.565 -190.235 ;
        RECT 326.235 -191.925 326.565 -191.595 ;
        RECT 326.235 -193.285 326.565 -192.955 ;
        RECT 326.235 -194.645 326.565 -194.315 ;
        RECT 326.235 -196.005 326.565 -195.675 ;
        RECT 326.235 -197.365 326.565 -197.035 ;
        RECT 326.235 -198.725 326.565 -198.395 ;
        RECT 326.235 -200.085 326.565 -199.755 ;
        RECT 326.235 -201.445 326.565 -201.115 ;
        RECT 326.235 -202.805 326.565 -202.475 ;
        RECT 326.235 -204.165 326.565 -203.835 ;
        RECT 326.235 -205.525 326.565 -205.195 ;
        RECT 326.235 -206.885 326.565 -206.555 ;
        RECT 326.235 -208.245 326.565 -207.915 ;
        RECT 326.235 -209.605 326.565 -209.275 ;
        RECT 326.235 -210.965 326.565 -210.635 ;
        RECT 326.235 -212.325 326.565 -211.995 ;
        RECT 326.235 -213.685 326.565 -213.355 ;
        RECT 326.235 -215.045 326.565 -214.715 ;
        RECT 326.235 -216.405 326.565 -216.075 ;
        RECT 326.235 -217.765 326.565 -217.435 ;
        RECT 326.235 -219.125 326.565 -218.795 ;
        RECT 326.235 -220.485 326.565 -220.155 ;
        RECT 326.235 -221.845 326.565 -221.515 ;
        RECT 326.235 -223.205 326.565 -222.875 ;
        RECT 326.235 -224.565 326.565 -224.235 ;
        RECT 326.235 -225.925 326.565 -225.595 ;
        RECT 326.235 -227.285 326.565 -226.955 ;
        RECT 326.235 -228.645 326.565 -228.315 ;
        RECT 326.235 -230.005 326.565 -229.675 ;
        RECT 326.235 -231.365 326.565 -231.035 ;
        RECT 326.235 -232.725 326.565 -232.395 ;
        RECT 326.235 -234.085 326.565 -233.755 ;
        RECT 326.235 -235.445 326.565 -235.115 ;
        RECT 326.235 -236.805 326.565 -236.475 ;
        RECT 326.235 -238.165 326.565 -237.835 ;
        RECT 326.235 -243.81 326.565 -242.68 ;
        RECT 326.24 -243.925 326.56 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 246.76 327.925 247.89 ;
        RECT 327.595 241.915 327.925 242.245 ;
        RECT 327.595 240.555 327.925 240.885 ;
        RECT 327.595 239.195 327.925 239.525 ;
        RECT 327.595 237.835 327.925 238.165 ;
        RECT 327.6 237.16 327.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 -1.525 327.925 -1.195 ;
        RECT 327.595 -2.885 327.925 -2.555 ;
        RECT 327.6 -3.56 327.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 -122.565 327.925 -122.235 ;
        RECT 327.595 -123.925 327.925 -123.595 ;
        RECT 327.595 -125.285 327.925 -124.955 ;
        RECT 327.595 -126.645 327.925 -126.315 ;
        RECT 327.595 -128.005 327.925 -127.675 ;
        RECT 327.595 -129.365 327.925 -129.035 ;
        RECT 327.595 -130.725 327.925 -130.395 ;
        RECT 327.595 -132.085 327.925 -131.755 ;
        RECT 327.595 -133.445 327.925 -133.115 ;
        RECT 327.595 -134.805 327.925 -134.475 ;
        RECT 327.595 -136.165 327.925 -135.835 ;
        RECT 327.595 -137.525 327.925 -137.195 ;
        RECT 327.595 -138.885 327.925 -138.555 ;
        RECT 327.595 -140.245 327.925 -139.915 ;
        RECT 327.595 -141.605 327.925 -141.275 ;
        RECT 327.595 -142.965 327.925 -142.635 ;
        RECT 327.595 -144.325 327.925 -143.995 ;
        RECT 327.595 -145.685 327.925 -145.355 ;
        RECT 327.595 -147.045 327.925 -146.715 ;
        RECT 327.595 -148.405 327.925 -148.075 ;
        RECT 327.595 -149.765 327.925 -149.435 ;
        RECT 327.595 -151.125 327.925 -150.795 ;
        RECT 327.595 -152.485 327.925 -152.155 ;
        RECT 327.595 -153.845 327.925 -153.515 ;
        RECT 327.595 -155.205 327.925 -154.875 ;
        RECT 327.595 -156.565 327.925 -156.235 ;
        RECT 327.595 -157.925 327.925 -157.595 ;
        RECT 327.595 -159.285 327.925 -158.955 ;
        RECT 327.595 -160.645 327.925 -160.315 ;
        RECT 327.595 -162.005 327.925 -161.675 ;
        RECT 327.595 -163.365 327.925 -163.035 ;
        RECT 327.595 -164.725 327.925 -164.395 ;
        RECT 327.595 -166.085 327.925 -165.755 ;
        RECT 327.595 -167.445 327.925 -167.115 ;
        RECT 327.595 -168.805 327.925 -168.475 ;
        RECT 327.595 -170.165 327.925 -169.835 ;
        RECT 327.595 -171.525 327.925 -171.195 ;
        RECT 327.595 -172.885 327.925 -172.555 ;
        RECT 327.595 -174.245 327.925 -173.915 ;
        RECT 327.595 -175.605 327.925 -175.275 ;
        RECT 327.595 -176.965 327.925 -176.635 ;
        RECT 327.595 -178.325 327.925 -177.995 ;
        RECT 327.595 -179.685 327.925 -179.355 ;
        RECT 327.595 -181.045 327.925 -180.715 ;
        RECT 327.595 -182.405 327.925 -182.075 ;
        RECT 327.595 -183.765 327.925 -183.435 ;
        RECT 327.595 -185.125 327.925 -184.795 ;
        RECT 327.595 -186.485 327.925 -186.155 ;
        RECT 327.595 -187.845 327.925 -187.515 ;
        RECT 327.595 -189.205 327.925 -188.875 ;
        RECT 327.595 -190.565 327.925 -190.235 ;
        RECT 327.595 -191.925 327.925 -191.595 ;
        RECT 327.595 -193.285 327.925 -192.955 ;
        RECT 327.595 -194.645 327.925 -194.315 ;
        RECT 327.595 -196.005 327.925 -195.675 ;
        RECT 327.595 -197.365 327.925 -197.035 ;
        RECT 327.595 -198.725 327.925 -198.395 ;
        RECT 327.595 -200.085 327.925 -199.755 ;
        RECT 327.595 -201.445 327.925 -201.115 ;
        RECT 327.595 -202.805 327.925 -202.475 ;
        RECT 327.595 -204.165 327.925 -203.835 ;
        RECT 327.595 -205.525 327.925 -205.195 ;
        RECT 327.595 -206.885 327.925 -206.555 ;
        RECT 327.595 -208.245 327.925 -207.915 ;
        RECT 327.595 -209.605 327.925 -209.275 ;
        RECT 327.595 -210.965 327.925 -210.635 ;
        RECT 327.595 -212.325 327.925 -211.995 ;
        RECT 327.595 -213.685 327.925 -213.355 ;
        RECT 327.595 -215.045 327.925 -214.715 ;
        RECT 327.595 -216.405 327.925 -216.075 ;
        RECT 327.595 -217.765 327.925 -217.435 ;
        RECT 327.595 -219.125 327.925 -218.795 ;
        RECT 327.595 -220.485 327.925 -220.155 ;
        RECT 327.595 -221.845 327.925 -221.515 ;
        RECT 327.595 -223.205 327.925 -222.875 ;
        RECT 327.595 -224.565 327.925 -224.235 ;
        RECT 327.595 -225.925 327.925 -225.595 ;
        RECT 327.595 -227.285 327.925 -226.955 ;
        RECT 327.595 -228.645 327.925 -228.315 ;
        RECT 327.595 -230.005 327.925 -229.675 ;
        RECT 327.595 -231.365 327.925 -231.035 ;
        RECT 327.595 -232.725 327.925 -232.395 ;
        RECT 327.595 -234.085 327.925 -233.755 ;
        RECT 327.595 -235.445 327.925 -235.115 ;
        RECT 327.595 -236.805 327.925 -236.475 ;
        RECT 327.595 -238.165 327.925 -237.835 ;
        RECT 327.595 -243.81 327.925 -242.68 ;
        RECT 327.6 -243.925 327.92 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 246.76 329.285 247.89 ;
        RECT 328.955 241.915 329.285 242.245 ;
        RECT 328.955 240.555 329.285 240.885 ;
        RECT 328.955 239.195 329.285 239.525 ;
        RECT 328.955 237.835 329.285 238.165 ;
        RECT 328.96 237.16 329.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 -1.525 329.285 -1.195 ;
        RECT 328.955 -2.885 329.285 -2.555 ;
        RECT 328.96 -3.56 329.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 -122.565 329.285 -122.235 ;
        RECT 328.955 -123.925 329.285 -123.595 ;
        RECT 328.955 -125.285 329.285 -124.955 ;
        RECT 328.955 -126.645 329.285 -126.315 ;
        RECT 328.955 -128.005 329.285 -127.675 ;
        RECT 328.955 -129.365 329.285 -129.035 ;
        RECT 328.955 -130.725 329.285 -130.395 ;
        RECT 328.955 -132.085 329.285 -131.755 ;
        RECT 328.955 -133.445 329.285 -133.115 ;
        RECT 328.955 -134.805 329.285 -134.475 ;
        RECT 328.955 -136.165 329.285 -135.835 ;
        RECT 328.955 -137.525 329.285 -137.195 ;
        RECT 328.955 -138.885 329.285 -138.555 ;
        RECT 328.955 -140.245 329.285 -139.915 ;
        RECT 328.955 -141.605 329.285 -141.275 ;
        RECT 328.955 -142.965 329.285 -142.635 ;
        RECT 328.955 -144.325 329.285 -143.995 ;
        RECT 328.955 -145.685 329.285 -145.355 ;
        RECT 328.955 -147.045 329.285 -146.715 ;
        RECT 328.955 -148.405 329.285 -148.075 ;
        RECT 328.955 -149.765 329.285 -149.435 ;
        RECT 328.955 -151.125 329.285 -150.795 ;
        RECT 328.955 -152.485 329.285 -152.155 ;
        RECT 328.955 -153.845 329.285 -153.515 ;
        RECT 328.955 -155.205 329.285 -154.875 ;
        RECT 328.955 -156.565 329.285 -156.235 ;
        RECT 328.955 -157.925 329.285 -157.595 ;
        RECT 328.955 -159.285 329.285 -158.955 ;
        RECT 328.955 -160.645 329.285 -160.315 ;
        RECT 328.955 -162.005 329.285 -161.675 ;
        RECT 328.955 -163.365 329.285 -163.035 ;
        RECT 328.955 -164.725 329.285 -164.395 ;
        RECT 328.955 -166.085 329.285 -165.755 ;
        RECT 328.955 -167.445 329.285 -167.115 ;
        RECT 328.955 -168.805 329.285 -168.475 ;
        RECT 328.955 -170.165 329.285 -169.835 ;
        RECT 328.955 -171.525 329.285 -171.195 ;
        RECT 328.955 -172.885 329.285 -172.555 ;
        RECT 328.955 -174.245 329.285 -173.915 ;
        RECT 328.955 -175.605 329.285 -175.275 ;
        RECT 328.955 -176.965 329.285 -176.635 ;
        RECT 328.955 -178.325 329.285 -177.995 ;
        RECT 328.955 -179.685 329.285 -179.355 ;
        RECT 328.955 -181.045 329.285 -180.715 ;
        RECT 328.955 -182.405 329.285 -182.075 ;
        RECT 328.955 -183.765 329.285 -183.435 ;
        RECT 328.955 -185.125 329.285 -184.795 ;
        RECT 328.955 -186.485 329.285 -186.155 ;
        RECT 328.955 -187.845 329.285 -187.515 ;
        RECT 328.955 -189.205 329.285 -188.875 ;
        RECT 328.955 -190.565 329.285 -190.235 ;
        RECT 328.955 -191.925 329.285 -191.595 ;
        RECT 328.955 -193.285 329.285 -192.955 ;
        RECT 328.955 -194.645 329.285 -194.315 ;
        RECT 328.955 -196.005 329.285 -195.675 ;
        RECT 328.955 -197.365 329.285 -197.035 ;
        RECT 328.955 -198.725 329.285 -198.395 ;
        RECT 328.955 -200.085 329.285 -199.755 ;
        RECT 328.955 -201.445 329.285 -201.115 ;
        RECT 328.955 -202.805 329.285 -202.475 ;
        RECT 328.955 -204.165 329.285 -203.835 ;
        RECT 328.955 -205.525 329.285 -205.195 ;
        RECT 328.955 -206.885 329.285 -206.555 ;
        RECT 328.955 -208.245 329.285 -207.915 ;
        RECT 328.955 -209.605 329.285 -209.275 ;
        RECT 328.955 -210.965 329.285 -210.635 ;
        RECT 328.955 -212.325 329.285 -211.995 ;
        RECT 328.955 -213.685 329.285 -213.355 ;
        RECT 328.955 -215.045 329.285 -214.715 ;
        RECT 328.955 -216.405 329.285 -216.075 ;
        RECT 328.955 -217.765 329.285 -217.435 ;
        RECT 328.955 -219.125 329.285 -218.795 ;
        RECT 328.955 -220.485 329.285 -220.155 ;
        RECT 328.955 -221.845 329.285 -221.515 ;
        RECT 328.955 -223.205 329.285 -222.875 ;
        RECT 328.955 -224.565 329.285 -224.235 ;
        RECT 328.955 -225.925 329.285 -225.595 ;
        RECT 328.955 -227.285 329.285 -226.955 ;
        RECT 328.955 -228.645 329.285 -228.315 ;
        RECT 328.955 -230.005 329.285 -229.675 ;
        RECT 328.955 -231.365 329.285 -231.035 ;
        RECT 328.955 -232.725 329.285 -232.395 ;
        RECT 328.955 -234.085 329.285 -233.755 ;
        RECT 328.955 -235.445 329.285 -235.115 ;
        RECT 328.955 -236.805 329.285 -236.475 ;
        RECT 328.955 -238.165 329.285 -237.835 ;
        RECT 328.955 -243.81 329.285 -242.68 ;
        RECT 328.96 -243.925 329.28 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.66 -125.535 329.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 246.76 330.645 247.89 ;
        RECT 330.315 241.915 330.645 242.245 ;
        RECT 330.315 240.555 330.645 240.885 ;
        RECT 330.315 239.195 330.645 239.525 ;
        RECT 330.315 237.835 330.645 238.165 ;
        RECT 330.32 237.16 330.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 -126.645 330.645 -126.315 ;
        RECT 330.315 -128.005 330.645 -127.675 ;
        RECT 330.315 -129.365 330.645 -129.035 ;
        RECT 330.315 -130.725 330.645 -130.395 ;
        RECT 330.315 -132.085 330.645 -131.755 ;
        RECT 330.315 -133.445 330.645 -133.115 ;
        RECT 330.315 -134.805 330.645 -134.475 ;
        RECT 330.315 -136.165 330.645 -135.835 ;
        RECT 330.315 -137.525 330.645 -137.195 ;
        RECT 330.315 -138.885 330.645 -138.555 ;
        RECT 330.315 -140.245 330.645 -139.915 ;
        RECT 330.315 -141.605 330.645 -141.275 ;
        RECT 330.315 -142.965 330.645 -142.635 ;
        RECT 330.315 -144.325 330.645 -143.995 ;
        RECT 330.315 -145.685 330.645 -145.355 ;
        RECT 330.315 -147.045 330.645 -146.715 ;
        RECT 330.315 -148.405 330.645 -148.075 ;
        RECT 330.315 -149.765 330.645 -149.435 ;
        RECT 330.315 -151.125 330.645 -150.795 ;
        RECT 330.315 -152.485 330.645 -152.155 ;
        RECT 330.315 -153.845 330.645 -153.515 ;
        RECT 330.315 -155.205 330.645 -154.875 ;
        RECT 330.315 -156.565 330.645 -156.235 ;
        RECT 330.315 -157.925 330.645 -157.595 ;
        RECT 330.315 -159.285 330.645 -158.955 ;
        RECT 330.315 -160.645 330.645 -160.315 ;
        RECT 330.315 -162.005 330.645 -161.675 ;
        RECT 330.315 -163.365 330.645 -163.035 ;
        RECT 330.315 -164.725 330.645 -164.395 ;
        RECT 330.315 -166.085 330.645 -165.755 ;
        RECT 330.315 -167.445 330.645 -167.115 ;
        RECT 330.315 -168.805 330.645 -168.475 ;
        RECT 330.315 -170.165 330.645 -169.835 ;
        RECT 330.315 -171.525 330.645 -171.195 ;
        RECT 330.315 -172.885 330.645 -172.555 ;
        RECT 330.315 -174.245 330.645 -173.915 ;
        RECT 330.315 -175.605 330.645 -175.275 ;
        RECT 330.315 -176.965 330.645 -176.635 ;
        RECT 330.315 -178.325 330.645 -177.995 ;
        RECT 330.315 -179.685 330.645 -179.355 ;
        RECT 330.315 -181.045 330.645 -180.715 ;
        RECT 330.315 -182.405 330.645 -182.075 ;
        RECT 330.315 -183.765 330.645 -183.435 ;
        RECT 330.315 -185.125 330.645 -184.795 ;
        RECT 330.315 -186.485 330.645 -186.155 ;
        RECT 330.315 -187.845 330.645 -187.515 ;
        RECT 330.315 -189.205 330.645 -188.875 ;
        RECT 330.315 -190.565 330.645 -190.235 ;
        RECT 330.315 -191.925 330.645 -191.595 ;
        RECT 330.315 -193.285 330.645 -192.955 ;
        RECT 330.315 -194.645 330.645 -194.315 ;
        RECT 330.315 -196.005 330.645 -195.675 ;
        RECT 330.315 -197.365 330.645 -197.035 ;
        RECT 330.315 -198.725 330.645 -198.395 ;
        RECT 330.315 -200.085 330.645 -199.755 ;
        RECT 330.315 -201.445 330.645 -201.115 ;
        RECT 330.315 -202.805 330.645 -202.475 ;
        RECT 330.315 -204.165 330.645 -203.835 ;
        RECT 330.315 -205.525 330.645 -205.195 ;
        RECT 330.315 -206.885 330.645 -206.555 ;
        RECT 330.315 -208.245 330.645 -207.915 ;
        RECT 330.315 -209.605 330.645 -209.275 ;
        RECT 330.315 -210.965 330.645 -210.635 ;
        RECT 330.315 -212.325 330.645 -211.995 ;
        RECT 330.315 -213.685 330.645 -213.355 ;
        RECT 330.315 -215.045 330.645 -214.715 ;
        RECT 330.315 -216.405 330.645 -216.075 ;
        RECT 330.315 -217.765 330.645 -217.435 ;
        RECT 330.315 -219.125 330.645 -218.795 ;
        RECT 330.315 -220.485 330.645 -220.155 ;
        RECT 330.315 -221.845 330.645 -221.515 ;
        RECT 330.315 -223.205 330.645 -222.875 ;
        RECT 330.315 -224.565 330.645 -224.235 ;
        RECT 330.315 -225.925 330.645 -225.595 ;
        RECT 330.315 -227.285 330.645 -226.955 ;
        RECT 330.315 -228.645 330.645 -228.315 ;
        RECT 330.315 -230.005 330.645 -229.675 ;
        RECT 330.315 -231.365 330.645 -231.035 ;
        RECT 330.315 -232.725 330.645 -232.395 ;
        RECT 330.315 -234.085 330.645 -233.755 ;
        RECT 330.315 -235.445 330.645 -235.115 ;
        RECT 330.315 -236.805 330.645 -236.475 ;
        RECT 330.315 -238.165 330.645 -237.835 ;
        RECT 330.315 -243.81 330.645 -242.68 ;
        RECT 330.32 -243.925 330.64 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 246.76 332.005 247.89 ;
        RECT 331.675 241.915 332.005 242.245 ;
        RECT 331.675 240.555 332.005 240.885 ;
        RECT 331.675 239.195 332.005 239.525 ;
        RECT 331.675 237.835 332.005 238.165 ;
        RECT 331.68 237.16 332 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 -1.525 332.005 -1.195 ;
        RECT 331.675 -2.885 332.005 -2.555 ;
        RECT 331.68 -3.56 332 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.035 246.76 333.365 247.89 ;
        RECT 333.035 241.915 333.365 242.245 ;
        RECT 333.035 240.555 333.365 240.885 ;
        RECT 333.035 239.195 333.365 239.525 ;
        RECT 333.035 237.835 333.365 238.165 ;
        RECT 333.04 237.16 333.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.035 -1.525 333.365 -1.195 ;
        RECT 333.035 -2.885 333.365 -2.555 ;
        RECT 333.04 -3.56 333.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 246.76 334.725 247.89 ;
        RECT 334.395 241.915 334.725 242.245 ;
        RECT 334.395 240.555 334.725 240.885 ;
        RECT 334.395 239.195 334.725 239.525 ;
        RECT 334.395 237.835 334.725 238.165 ;
        RECT 334.4 237.16 334.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 -1.525 334.725 -1.195 ;
        RECT 334.395 -2.885 334.725 -2.555 ;
        RECT 334.4 -3.56 334.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 -122.565 334.725 -122.235 ;
        RECT 334.395 -123.925 334.725 -123.595 ;
        RECT 334.395 -125.285 334.725 -124.955 ;
        RECT 334.395 -126.645 334.725 -126.315 ;
        RECT 334.395 -128.005 334.725 -127.675 ;
        RECT 334.395 -129.365 334.725 -129.035 ;
        RECT 334.395 -130.725 334.725 -130.395 ;
        RECT 334.395 -132.085 334.725 -131.755 ;
        RECT 334.395 -133.445 334.725 -133.115 ;
        RECT 334.395 -134.805 334.725 -134.475 ;
        RECT 334.395 -136.165 334.725 -135.835 ;
        RECT 334.395 -137.525 334.725 -137.195 ;
        RECT 334.395 -138.885 334.725 -138.555 ;
        RECT 334.395 -140.245 334.725 -139.915 ;
        RECT 334.395 -141.605 334.725 -141.275 ;
        RECT 334.395 -142.965 334.725 -142.635 ;
        RECT 334.395 -144.325 334.725 -143.995 ;
        RECT 334.395 -145.685 334.725 -145.355 ;
        RECT 334.395 -147.045 334.725 -146.715 ;
        RECT 334.395 -148.405 334.725 -148.075 ;
        RECT 334.395 -149.765 334.725 -149.435 ;
        RECT 334.395 -151.125 334.725 -150.795 ;
        RECT 334.395 -152.485 334.725 -152.155 ;
        RECT 334.395 -153.845 334.725 -153.515 ;
        RECT 334.395 -155.205 334.725 -154.875 ;
        RECT 334.395 -156.565 334.725 -156.235 ;
        RECT 334.395 -157.925 334.725 -157.595 ;
        RECT 334.395 -159.285 334.725 -158.955 ;
        RECT 334.395 -160.645 334.725 -160.315 ;
        RECT 334.395 -162.005 334.725 -161.675 ;
        RECT 334.395 -163.365 334.725 -163.035 ;
        RECT 334.395 -164.725 334.725 -164.395 ;
        RECT 334.395 -166.085 334.725 -165.755 ;
        RECT 334.395 -167.445 334.725 -167.115 ;
        RECT 334.395 -168.805 334.725 -168.475 ;
        RECT 334.395 -170.165 334.725 -169.835 ;
        RECT 334.395 -171.525 334.725 -171.195 ;
        RECT 334.395 -172.885 334.725 -172.555 ;
        RECT 334.395 -174.245 334.725 -173.915 ;
        RECT 334.395 -175.605 334.725 -175.275 ;
        RECT 334.395 -176.965 334.725 -176.635 ;
        RECT 334.395 -178.325 334.725 -177.995 ;
        RECT 334.395 -179.685 334.725 -179.355 ;
        RECT 334.395 -181.045 334.725 -180.715 ;
        RECT 334.395 -182.405 334.725 -182.075 ;
        RECT 334.395 -183.765 334.725 -183.435 ;
        RECT 334.395 -185.125 334.725 -184.795 ;
        RECT 334.395 -186.485 334.725 -186.155 ;
        RECT 334.395 -187.845 334.725 -187.515 ;
        RECT 334.395 -189.205 334.725 -188.875 ;
        RECT 334.395 -190.565 334.725 -190.235 ;
        RECT 334.395 -191.925 334.725 -191.595 ;
        RECT 334.395 -193.285 334.725 -192.955 ;
        RECT 334.395 -194.645 334.725 -194.315 ;
        RECT 334.395 -196.005 334.725 -195.675 ;
        RECT 334.395 -197.365 334.725 -197.035 ;
        RECT 334.395 -198.725 334.725 -198.395 ;
        RECT 334.395 -200.085 334.725 -199.755 ;
        RECT 334.395 -201.445 334.725 -201.115 ;
        RECT 334.395 -202.805 334.725 -202.475 ;
        RECT 334.395 -204.165 334.725 -203.835 ;
        RECT 334.395 -205.525 334.725 -205.195 ;
        RECT 334.395 -206.885 334.725 -206.555 ;
        RECT 334.395 -208.245 334.725 -207.915 ;
        RECT 334.395 -209.605 334.725 -209.275 ;
        RECT 334.395 -210.965 334.725 -210.635 ;
        RECT 334.395 -212.325 334.725 -211.995 ;
        RECT 334.395 -213.685 334.725 -213.355 ;
        RECT 334.395 -215.045 334.725 -214.715 ;
        RECT 334.395 -216.405 334.725 -216.075 ;
        RECT 334.395 -217.765 334.725 -217.435 ;
        RECT 334.395 -219.125 334.725 -218.795 ;
        RECT 334.395 -220.485 334.725 -220.155 ;
        RECT 334.395 -221.845 334.725 -221.515 ;
        RECT 334.395 -223.205 334.725 -222.875 ;
        RECT 334.395 -224.565 334.725 -224.235 ;
        RECT 334.395 -225.925 334.725 -225.595 ;
        RECT 334.395 -227.285 334.725 -226.955 ;
        RECT 334.395 -228.645 334.725 -228.315 ;
        RECT 334.395 -230.005 334.725 -229.675 ;
        RECT 334.395 -231.365 334.725 -231.035 ;
        RECT 334.395 -232.725 334.725 -232.395 ;
        RECT 334.395 -234.085 334.725 -233.755 ;
        RECT 334.395 -235.445 334.725 -235.115 ;
        RECT 334.395 -236.805 334.725 -236.475 ;
        RECT 334.395 -238.165 334.725 -237.835 ;
        RECT 334.395 -243.81 334.725 -242.68 ;
        RECT 334.4 -243.925 334.72 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 246.76 336.085 247.89 ;
        RECT 335.755 241.915 336.085 242.245 ;
        RECT 335.755 240.555 336.085 240.885 ;
        RECT 335.755 239.195 336.085 239.525 ;
        RECT 335.755 237.835 336.085 238.165 ;
        RECT 335.76 237.16 336.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 -1.525 336.085 -1.195 ;
        RECT 335.755 -2.885 336.085 -2.555 ;
        RECT 335.76 -3.56 336.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 -122.565 336.085 -122.235 ;
        RECT 335.755 -123.925 336.085 -123.595 ;
        RECT 335.755 -125.285 336.085 -124.955 ;
        RECT 335.755 -126.645 336.085 -126.315 ;
        RECT 335.755 -128.005 336.085 -127.675 ;
        RECT 335.755 -129.365 336.085 -129.035 ;
        RECT 335.755 -130.725 336.085 -130.395 ;
        RECT 335.755 -132.085 336.085 -131.755 ;
        RECT 335.755 -133.445 336.085 -133.115 ;
        RECT 335.755 -134.805 336.085 -134.475 ;
        RECT 335.755 -136.165 336.085 -135.835 ;
        RECT 335.755 -137.525 336.085 -137.195 ;
        RECT 335.755 -138.885 336.085 -138.555 ;
        RECT 335.755 -140.245 336.085 -139.915 ;
        RECT 335.755 -141.605 336.085 -141.275 ;
        RECT 335.755 -142.965 336.085 -142.635 ;
        RECT 335.755 -144.325 336.085 -143.995 ;
        RECT 335.755 -145.685 336.085 -145.355 ;
        RECT 335.755 -147.045 336.085 -146.715 ;
        RECT 335.755 -148.405 336.085 -148.075 ;
        RECT 335.755 -149.765 336.085 -149.435 ;
        RECT 335.755 -151.125 336.085 -150.795 ;
        RECT 335.755 -152.485 336.085 -152.155 ;
        RECT 335.755 -153.845 336.085 -153.515 ;
        RECT 335.755 -155.205 336.085 -154.875 ;
        RECT 335.755 -156.565 336.085 -156.235 ;
        RECT 335.755 -157.925 336.085 -157.595 ;
        RECT 335.755 -159.285 336.085 -158.955 ;
        RECT 335.755 -160.645 336.085 -160.315 ;
        RECT 335.755 -162.005 336.085 -161.675 ;
        RECT 335.755 -163.365 336.085 -163.035 ;
        RECT 335.755 -164.725 336.085 -164.395 ;
        RECT 335.755 -166.085 336.085 -165.755 ;
        RECT 335.755 -167.445 336.085 -167.115 ;
        RECT 335.755 -168.805 336.085 -168.475 ;
        RECT 335.755 -170.165 336.085 -169.835 ;
        RECT 335.755 -171.525 336.085 -171.195 ;
        RECT 335.755 -172.885 336.085 -172.555 ;
        RECT 335.755 -174.245 336.085 -173.915 ;
        RECT 335.755 -175.605 336.085 -175.275 ;
        RECT 335.755 -176.965 336.085 -176.635 ;
        RECT 335.755 -178.325 336.085 -177.995 ;
        RECT 335.755 -179.685 336.085 -179.355 ;
        RECT 335.755 -181.045 336.085 -180.715 ;
        RECT 335.755 -182.405 336.085 -182.075 ;
        RECT 335.755 -183.765 336.085 -183.435 ;
        RECT 335.755 -185.125 336.085 -184.795 ;
        RECT 335.755 -186.485 336.085 -186.155 ;
        RECT 335.755 -187.845 336.085 -187.515 ;
        RECT 335.755 -189.205 336.085 -188.875 ;
        RECT 335.755 -190.565 336.085 -190.235 ;
        RECT 335.755 -191.925 336.085 -191.595 ;
        RECT 335.755 -193.285 336.085 -192.955 ;
        RECT 335.755 -194.645 336.085 -194.315 ;
        RECT 335.755 -196.005 336.085 -195.675 ;
        RECT 335.755 -197.365 336.085 -197.035 ;
        RECT 335.755 -198.725 336.085 -198.395 ;
        RECT 335.755 -200.085 336.085 -199.755 ;
        RECT 335.755 -201.445 336.085 -201.115 ;
        RECT 335.755 -202.805 336.085 -202.475 ;
        RECT 335.755 -204.165 336.085 -203.835 ;
        RECT 335.755 -205.525 336.085 -205.195 ;
        RECT 335.755 -206.885 336.085 -206.555 ;
        RECT 335.755 -208.245 336.085 -207.915 ;
        RECT 335.755 -209.605 336.085 -209.275 ;
        RECT 335.755 -210.965 336.085 -210.635 ;
        RECT 335.755 -212.325 336.085 -211.995 ;
        RECT 335.755 -213.685 336.085 -213.355 ;
        RECT 335.755 -215.045 336.085 -214.715 ;
        RECT 335.755 -216.405 336.085 -216.075 ;
        RECT 335.755 -217.765 336.085 -217.435 ;
        RECT 335.755 -219.125 336.085 -218.795 ;
        RECT 335.755 -220.485 336.085 -220.155 ;
        RECT 335.755 -221.845 336.085 -221.515 ;
        RECT 335.755 -223.205 336.085 -222.875 ;
        RECT 335.755 -224.565 336.085 -224.235 ;
        RECT 335.755 -225.925 336.085 -225.595 ;
        RECT 335.755 -227.285 336.085 -226.955 ;
        RECT 335.755 -228.645 336.085 -228.315 ;
        RECT 335.755 -230.005 336.085 -229.675 ;
        RECT 335.755 -231.365 336.085 -231.035 ;
        RECT 335.755 -232.725 336.085 -232.395 ;
        RECT 335.755 -234.085 336.085 -233.755 ;
        RECT 335.755 -235.445 336.085 -235.115 ;
        RECT 335.755 -236.805 336.085 -236.475 ;
        RECT 335.755 -238.165 336.085 -237.835 ;
        RECT 335.755 -243.81 336.085 -242.68 ;
        RECT 335.76 -243.925 336.08 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 246.76 337.445 247.89 ;
        RECT 337.115 241.915 337.445 242.245 ;
        RECT 337.115 240.555 337.445 240.885 ;
        RECT 337.115 239.195 337.445 239.525 ;
        RECT 337.115 237.835 337.445 238.165 ;
        RECT 337.12 237.16 337.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 -1.525 337.445 -1.195 ;
        RECT 337.115 -2.885 337.445 -2.555 ;
        RECT 337.12 -3.56 337.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 -122.565 337.445 -122.235 ;
        RECT 337.115 -123.925 337.445 -123.595 ;
        RECT 337.115 -125.285 337.445 -124.955 ;
        RECT 337.115 -126.645 337.445 -126.315 ;
        RECT 337.115 -128.005 337.445 -127.675 ;
        RECT 337.115 -129.365 337.445 -129.035 ;
        RECT 337.115 -130.725 337.445 -130.395 ;
        RECT 337.115 -132.085 337.445 -131.755 ;
        RECT 337.115 -133.445 337.445 -133.115 ;
        RECT 337.115 -134.805 337.445 -134.475 ;
        RECT 337.115 -136.165 337.445 -135.835 ;
        RECT 337.115 -137.525 337.445 -137.195 ;
        RECT 337.115 -138.885 337.445 -138.555 ;
        RECT 337.115 -140.245 337.445 -139.915 ;
        RECT 337.115 -141.605 337.445 -141.275 ;
        RECT 337.115 -142.965 337.445 -142.635 ;
        RECT 337.115 -144.325 337.445 -143.995 ;
        RECT 337.115 -145.685 337.445 -145.355 ;
        RECT 337.115 -147.045 337.445 -146.715 ;
        RECT 337.115 -148.405 337.445 -148.075 ;
        RECT 337.115 -149.765 337.445 -149.435 ;
        RECT 337.115 -151.125 337.445 -150.795 ;
        RECT 337.115 -152.485 337.445 -152.155 ;
        RECT 337.115 -153.845 337.445 -153.515 ;
        RECT 337.115 -155.205 337.445 -154.875 ;
        RECT 337.115 -156.565 337.445 -156.235 ;
        RECT 337.115 -157.925 337.445 -157.595 ;
        RECT 337.115 -159.285 337.445 -158.955 ;
        RECT 337.115 -160.645 337.445 -160.315 ;
        RECT 337.115 -162.005 337.445 -161.675 ;
        RECT 337.115 -163.365 337.445 -163.035 ;
        RECT 337.115 -164.725 337.445 -164.395 ;
        RECT 337.115 -166.085 337.445 -165.755 ;
        RECT 337.115 -167.445 337.445 -167.115 ;
        RECT 337.115 -168.805 337.445 -168.475 ;
        RECT 337.115 -170.165 337.445 -169.835 ;
        RECT 337.115 -171.525 337.445 -171.195 ;
        RECT 337.115 -172.885 337.445 -172.555 ;
        RECT 337.115 -174.245 337.445 -173.915 ;
        RECT 337.115 -175.605 337.445 -175.275 ;
        RECT 337.115 -176.965 337.445 -176.635 ;
        RECT 337.115 -178.325 337.445 -177.995 ;
        RECT 337.115 -179.685 337.445 -179.355 ;
        RECT 337.115 -181.045 337.445 -180.715 ;
        RECT 337.115 -182.405 337.445 -182.075 ;
        RECT 337.115 -183.765 337.445 -183.435 ;
        RECT 337.115 -185.125 337.445 -184.795 ;
        RECT 337.115 -186.485 337.445 -186.155 ;
        RECT 337.115 -187.845 337.445 -187.515 ;
        RECT 337.115 -189.205 337.445 -188.875 ;
        RECT 337.115 -190.565 337.445 -190.235 ;
        RECT 337.115 -191.925 337.445 -191.595 ;
        RECT 337.115 -193.285 337.445 -192.955 ;
        RECT 337.115 -194.645 337.445 -194.315 ;
        RECT 337.115 -196.005 337.445 -195.675 ;
        RECT 337.115 -197.365 337.445 -197.035 ;
        RECT 337.115 -198.725 337.445 -198.395 ;
        RECT 337.115 -200.085 337.445 -199.755 ;
        RECT 337.115 -201.445 337.445 -201.115 ;
        RECT 337.115 -202.805 337.445 -202.475 ;
        RECT 337.115 -204.165 337.445 -203.835 ;
        RECT 337.115 -205.525 337.445 -205.195 ;
        RECT 337.115 -206.885 337.445 -206.555 ;
        RECT 337.115 -208.245 337.445 -207.915 ;
        RECT 337.115 -209.605 337.445 -209.275 ;
        RECT 337.115 -210.965 337.445 -210.635 ;
        RECT 337.115 -212.325 337.445 -211.995 ;
        RECT 337.115 -213.685 337.445 -213.355 ;
        RECT 337.115 -215.045 337.445 -214.715 ;
        RECT 337.115 -216.405 337.445 -216.075 ;
        RECT 337.115 -217.765 337.445 -217.435 ;
        RECT 337.115 -219.125 337.445 -218.795 ;
        RECT 337.115 -220.485 337.445 -220.155 ;
        RECT 337.115 -221.845 337.445 -221.515 ;
        RECT 337.115 -223.205 337.445 -222.875 ;
        RECT 337.115 -224.565 337.445 -224.235 ;
        RECT 337.115 -225.925 337.445 -225.595 ;
        RECT 337.115 -227.285 337.445 -226.955 ;
        RECT 337.115 -228.645 337.445 -228.315 ;
        RECT 337.115 -230.005 337.445 -229.675 ;
        RECT 337.115 -231.365 337.445 -231.035 ;
        RECT 337.115 -232.725 337.445 -232.395 ;
        RECT 337.115 -234.085 337.445 -233.755 ;
        RECT 337.115 -235.445 337.445 -235.115 ;
        RECT 337.115 -236.805 337.445 -236.475 ;
        RECT 337.115 -238.165 337.445 -237.835 ;
        RECT 337.115 -243.81 337.445 -242.68 ;
        RECT 337.12 -243.925 337.44 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 246.76 338.805 247.89 ;
        RECT 338.475 241.915 338.805 242.245 ;
        RECT 338.475 240.555 338.805 240.885 ;
        RECT 338.475 239.195 338.805 239.525 ;
        RECT 338.475 237.835 338.805 238.165 ;
        RECT 338.48 237.16 338.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 -1.525 338.805 -1.195 ;
        RECT 338.475 -2.885 338.805 -2.555 ;
        RECT 338.48 -3.56 338.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 -122.565 338.805 -122.235 ;
        RECT 338.475 -123.925 338.805 -123.595 ;
        RECT 338.475 -125.285 338.805 -124.955 ;
        RECT 338.475 -126.645 338.805 -126.315 ;
        RECT 338.475 -128.005 338.805 -127.675 ;
        RECT 338.475 -129.365 338.805 -129.035 ;
        RECT 338.475 -130.725 338.805 -130.395 ;
        RECT 338.475 -132.085 338.805 -131.755 ;
        RECT 338.475 -133.445 338.805 -133.115 ;
        RECT 338.475 -134.805 338.805 -134.475 ;
        RECT 338.475 -136.165 338.805 -135.835 ;
        RECT 338.475 -137.525 338.805 -137.195 ;
        RECT 338.475 -138.885 338.805 -138.555 ;
        RECT 338.475 -140.245 338.805 -139.915 ;
        RECT 338.475 -141.605 338.805 -141.275 ;
        RECT 338.475 -142.965 338.805 -142.635 ;
        RECT 338.475 -144.325 338.805 -143.995 ;
        RECT 338.475 -145.685 338.805 -145.355 ;
        RECT 338.475 -147.045 338.805 -146.715 ;
        RECT 338.475 -148.405 338.805 -148.075 ;
        RECT 338.475 -149.765 338.805 -149.435 ;
        RECT 338.475 -151.125 338.805 -150.795 ;
        RECT 338.475 -152.485 338.805 -152.155 ;
        RECT 338.475 -153.845 338.805 -153.515 ;
        RECT 338.475 -155.205 338.805 -154.875 ;
        RECT 338.475 -156.565 338.805 -156.235 ;
        RECT 338.475 -157.925 338.805 -157.595 ;
        RECT 338.475 -159.285 338.805 -158.955 ;
        RECT 338.475 -160.645 338.805 -160.315 ;
        RECT 338.475 -162.005 338.805 -161.675 ;
        RECT 338.475 -163.365 338.805 -163.035 ;
        RECT 338.475 -164.725 338.805 -164.395 ;
        RECT 338.475 -166.085 338.805 -165.755 ;
        RECT 338.475 -167.445 338.805 -167.115 ;
        RECT 338.475 -168.805 338.805 -168.475 ;
        RECT 338.475 -170.165 338.805 -169.835 ;
        RECT 338.475 -171.525 338.805 -171.195 ;
        RECT 338.475 -172.885 338.805 -172.555 ;
        RECT 338.475 -174.245 338.805 -173.915 ;
        RECT 338.475 -175.605 338.805 -175.275 ;
        RECT 338.475 -176.965 338.805 -176.635 ;
        RECT 338.475 -178.325 338.805 -177.995 ;
        RECT 338.475 -179.685 338.805 -179.355 ;
        RECT 338.475 -181.045 338.805 -180.715 ;
        RECT 338.475 -182.405 338.805 -182.075 ;
        RECT 338.475 -183.765 338.805 -183.435 ;
        RECT 338.475 -185.125 338.805 -184.795 ;
        RECT 338.475 -186.485 338.805 -186.155 ;
        RECT 338.475 -187.845 338.805 -187.515 ;
        RECT 338.475 -189.205 338.805 -188.875 ;
        RECT 338.475 -190.565 338.805 -190.235 ;
        RECT 338.475 -191.925 338.805 -191.595 ;
        RECT 338.475 -193.285 338.805 -192.955 ;
        RECT 338.475 -194.645 338.805 -194.315 ;
        RECT 338.475 -196.005 338.805 -195.675 ;
        RECT 338.475 -197.365 338.805 -197.035 ;
        RECT 338.475 -198.725 338.805 -198.395 ;
        RECT 338.475 -200.085 338.805 -199.755 ;
        RECT 338.475 -201.445 338.805 -201.115 ;
        RECT 338.475 -202.805 338.805 -202.475 ;
        RECT 338.475 -204.165 338.805 -203.835 ;
        RECT 338.475 -205.525 338.805 -205.195 ;
        RECT 338.475 -206.885 338.805 -206.555 ;
        RECT 338.475 -208.245 338.805 -207.915 ;
        RECT 338.475 -209.605 338.805 -209.275 ;
        RECT 338.475 -210.965 338.805 -210.635 ;
        RECT 338.475 -212.325 338.805 -211.995 ;
        RECT 338.475 -213.685 338.805 -213.355 ;
        RECT 338.475 -215.045 338.805 -214.715 ;
        RECT 338.475 -216.405 338.805 -216.075 ;
        RECT 338.475 -217.765 338.805 -217.435 ;
        RECT 338.475 -219.125 338.805 -218.795 ;
        RECT 338.475 -220.485 338.805 -220.155 ;
        RECT 338.475 -221.845 338.805 -221.515 ;
        RECT 338.475 -223.205 338.805 -222.875 ;
        RECT 338.475 -224.565 338.805 -224.235 ;
        RECT 338.475 -225.925 338.805 -225.595 ;
        RECT 338.475 -227.285 338.805 -226.955 ;
        RECT 338.475 -228.645 338.805 -228.315 ;
        RECT 338.475 -230.005 338.805 -229.675 ;
        RECT 338.475 -231.365 338.805 -231.035 ;
        RECT 338.475 -232.725 338.805 -232.395 ;
        RECT 338.475 -234.085 338.805 -233.755 ;
        RECT 338.475 -235.445 338.805 -235.115 ;
        RECT 338.475 -236.805 338.805 -236.475 ;
        RECT 338.475 -238.165 338.805 -237.835 ;
        RECT 338.475 -243.81 338.805 -242.68 ;
        RECT 338.48 -243.925 338.8 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 246.76 340.165 247.89 ;
        RECT 339.835 241.915 340.165 242.245 ;
        RECT 339.835 240.555 340.165 240.885 ;
        RECT 339.835 239.195 340.165 239.525 ;
        RECT 339.835 237.835 340.165 238.165 ;
        RECT 339.84 237.16 340.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 -1.525 340.165 -1.195 ;
        RECT 339.835 -2.885 340.165 -2.555 ;
        RECT 339.84 -3.56 340.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 -232.725 340.165 -232.395 ;
        RECT 339.835 -234.085 340.165 -233.755 ;
        RECT 339.835 -235.445 340.165 -235.115 ;
        RECT 339.835 -236.805 340.165 -236.475 ;
        RECT 339.835 -238.165 340.165 -237.835 ;
        RECT 339.835 -243.81 340.165 -242.68 ;
        RECT 339.84 -243.925 340.16 -122.235 ;
        RECT 339.835 -122.565 340.165 -122.235 ;
        RECT 339.835 -123.925 340.165 -123.595 ;
        RECT 339.835 -125.285 340.165 -124.955 ;
        RECT 339.835 -126.645 340.165 -126.315 ;
        RECT 339.835 -128.005 340.165 -127.675 ;
        RECT 339.835 -129.365 340.165 -129.035 ;
        RECT 339.835 -130.725 340.165 -130.395 ;
        RECT 339.835 -132.085 340.165 -131.755 ;
        RECT 339.835 -133.445 340.165 -133.115 ;
        RECT 339.835 -134.805 340.165 -134.475 ;
        RECT 339.835 -136.165 340.165 -135.835 ;
        RECT 339.835 -137.525 340.165 -137.195 ;
        RECT 339.835 -138.885 340.165 -138.555 ;
        RECT 339.835 -140.245 340.165 -139.915 ;
        RECT 339.835 -141.605 340.165 -141.275 ;
        RECT 339.835 -142.965 340.165 -142.635 ;
        RECT 339.835 -144.325 340.165 -143.995 ;
        RECT 339.835 -145.685 340.165 -145.355 ;
        RECT 339.835 -147.045 340.165 -146.715 ;
        RECT 339.835 -148.405 340.165 -148.075 ;
        RECT 339.835 -149.765 340.165 -149.435 ;
        RECT 339.835 -151.125 340.165 -150.795 ;
        RECT 339.835 -152.485 340.165 -152.155 ;
        RECT 339.835 -153.845 340.165 -153.515 ;
        RECT 339.835 -155.205 340.165 -154.875 ;
        RECT 339.835 -156.565 340.165 -156.235 ;
        RECT 339.835 -157.925 340.165 -157.595 ;
        RECT 339.835 -159.285 340.165 -158.955 ;
        RECT 339.835 -160.645 340.165 -160.315 ;
        RECT 339.835 -162.005 340.165 -161.675 ;
        RECT 339.835 -163.365 340.165 -163.035 ;
        RECT 339.835 -164.725 340.165 -164.395 ;
        RECT 339.835 -166.085 340.165 -165.755 ;
        RECT 339.835 -167.445 340.165 -167.115 ;
        RECT 339.835 -168.805 340.165 -168.475 ;
        RECT 339.835 -170.165 340.165 -169.835 ;
        RECT 339.835 -171.525 340.165 -171.195 ;
        RECT 339.835 -172.885 340.165 -172.555 ;
        RECT 339.835 -174.245 340.165 -173.915 ;
        RECT 339.835 -175.605 340.165 -175.275 ;
        RECT 339.835 -176.965 340.165 -176.635 ;
        RECT 339.835 -178.325 340.165 -177.995 ;
        RECT 339.835 -179.685 340.165 -179.355 ;
        RECT 339.835 -181.045 340.165 -180.715 ;
        RECT 339.835 -182.405 340.165 -182.075 ;
        RECT 339.835 -183.765 340.165 -183.435 ;
        RECT 339.835 -185.125 340.165 -184.795 ;
        RECT 339.835 -186.485 340.165 -186.155 ;
        RECT 339.835 -187.845 340.165 -187.515 ;
        RECT 339.835 -189.205 340.165 -188.875 ;
        RECT 339.835 -190.565 340.165 -190.235 ;
        RECT 339.835 -191.925 340.165 -191.595 ;
        RECT 339.835 -193.285 340.165 -192.955 ;
        RECT 339.835 -194.645 340.165 -194.315 ;
        RECT 339.835 -196.005 340.165 -195.675 ;
        RECT 339.835 -197.365 340.165 -197.035 ;
        RECT 339.835 -198.725 340.165 -198.395 ;
        RECT 339.835 -200.085 340.165 -199.755 ;
        RECT 339.835 -201.445 340.165 -201.115 ;
        RECT 339.835 -202.805 340.165 -202.475 ;
        RECT 339.835 -204.165 340.165 -203.835 ;
        RECT 339.835 -205.525 340.165 -205.195 ;
        RECT 339.835 -206.885 340.165 -206.555 ;
        RECT 339.835 -208.245 340.165 -207.915 ;
        RECT 339.835 -209.605 340.165 -209.275 ;
        RECT 339.835 -210.965 340.165 -210.635 ;
        RECT 339.835 -212.325 340.165 -211.995 ;
        RECT 339.835 -213.685 340.165 -213.355 ;
        RECT 339.835 -215.045 340.165 -214.715 ;
        RECT 339.835 -216.405 340.165 -216.075 ;
        RECT 339.835 -217.765 340.165 -217.435 ;
        RECT 339.835 -219.125 340.165 -218.795 ;
        RECT 339.835 -220.485 340.165 -220.155 ;
        RECT 339.835 -221.845 340.165 -221.515 ;
        RECT 339.835 -223.205 340.165 -222.875 ;
        RECT 339.835 -224.565 340.165 -224.235 ;
        RECT 339.835 -225.925 340.165 -225.595 ;
        RECT 339.835 -227.285 340.165 -226.955 ;
        RECT 339.835 -228.645 340.165 -228.315 ;
        RECT 339.835 -230.005 340.165 -229.675 ;
        RECT 339.835 -231.365 340.165 -231.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 246.76 303.445 247.89 ;
        RECT 303.115 241.915 303.445 242.245 ;
        RECT 303.115 240.555 303.445 240.885 ;
        RECT 303.115 239.195 303.445 239.525 ;
        RECT 303.115 237.835 303.445 238.165 ;
        RECT 303.12 237.16 303.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 -1.525 303.445 -1.195 ;
        RECT 303.115 -2.885 303.445 -2.555 ;
        RECT 303.12 -3.56 303.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 -122.565 303.445 -122.235 ;
        RECT 303.115 -123.925 303.445 -123.595 ;
        RECT 303.115 -125.285 303.445 -124.955 ;
        RECT 303.115 -126.645 303.445 -126.315 ;
        RECT 303.115 -128.005 303.445 -127.675 ;
        RECT 303.115 -129.365 303.445 -129.035 ;
        RECT 303.115 -130.725 303.445 -130.395 ;
        RECT 303.115 -132.085 303.445 -131.755 ;
        RECT 303.115 -133.445 303.445 -133.115 ;
        RECT 303.115 -134.805 303.445 -134.475 ;
        RECT 303.115 -136.165 303.445 -135.835 ;
        RECT 303.115 -137.525 303.445 -137.195 ;
        RECT 303.115 -138.885 303.445 -138.555 ;
        RECT 303.115 -140.245 303.445 -139.915 ;
        RECT 303.115 -141.605 303.445 -141.275 ;
        RECT 303.115 -142.965 303.445 -142.635 ;
        RECT 303.115 -144.325 303.445 -143.995 ;
        RECT 303.115 -145.685 303.445 -145.355 ;
        RECT 303.115 -147.045 303.445 -146.715 ;
        RECT 303.115 -148.405 303.445 -148.075 ;
        RECT 303.115 -149.765 303.445 -149.435 ;
        RECT 303.115 -151.125 303.445 -150.795 ;
        RECT 303.115 -152.485 303.445 -152.155 ;
        RECT 303.115 -153.845 303.445 -153.515 ;
        RECT 303.115 -155.205 303.445 -154.875 ;
        RECT 303.115 -156.565 303.445 -156.235 ;
        RECT 303.115 -157.925 303.445 -157.595 ;
        RECT 303.115 -159.285 303.445 -158.955 ;
        RECT 303.115 -160.645 303.445 -160.315 ;
        RECT 303.115 -162.005 303.445 -161.675 ;
        RECT 303.115 -163.365 303.445 -163.035 ;
        RECT 303.115 -164.725 303.445 -164.395 ;
        RECT 303.115 -166.085 303.445 -165.755 ;
        RECT 303.115 -167.445 303.445 -167.115 ;
        RECT 303.115 -168.805 303.445 -168.475 ;
        RECT 303.115 -170.165 303.445 -169.835 ;
        RECT 303.115 -171.525 303.445 -171.195 ;
        RECT 303.115 -172.885 303.445 -172.555 ;
        RECT 303.115 -174.245 303.445 -173.915 ;
        RECT 303.115 -175.605 303.445 -175.275 ;
        RECT 303.115 -176.965 303.445 -176.635 ;
        RECT 303.115 -178.325 303.445 -177.995 ;
        RECT 303.115 -179.685 303.445 -179.355 ;
        RECT 303.115 -181.045 303.445 -180.715 ;
        RECT 303.115 -182.405 303.445 -182.075 ;
        RECT 303.115 -183.765 303.445 -183.435 ;
        RECT 303.115 -185.125 303.445 -184.795 ;
        RECT 303.115 -186.485 303.445 -186.155 ;
        RECT 303.115 -187.845 303.445 -187.515 ;
        RECT 303.115 -189.205 303.445 -188.875 ;
        RECT 303.115 -190.565 303.445 -190.235 ;
        RECT 303.115 -191.925 303.445 -191.595 ;
        RECT 303.115 -193.285 303.445 -192.955 ;
        RECT 303.115 -194.645 303.445 -194.315 ;
        RECT 303.115 -196.005 303.445 -195.675 ;
        RECT 303.115 -197.365 303.445 -197.035 ;
        RECT 303.115 -198.725 303.445 -198.395 ;
        RECT 303.115 -200.085 303.445 -199.755 ;
        RECT 303.115 -201.445 303.445 -201.115 ;
        RECT 303.115 -202.805 303.445 -202.475 ;
        RECT 303.115 -204.165 303.445 -203.835 ;
        RECT 303.115 -205.525 303.445 -205.195 ;
        RECT 303.115 -206.885 303.445 -206.555 ;
        RECT 303.115 -208.245 303.445 -207.915 ;
        RECT 303.115 -209.605 303.445 -209.275 ;
        RECT 303.115 -210.965 303.445 -210.635 ;
        RECT 303.115 -212.325 303.445 -211.995 ;
        RECT 303.115 -213.685 303.445 -213.355 ;
        RECT 303.115 -215.045 303.445 -214.715 ;
        RECT 303.115 -216.405 303.445 -216.075 ;
        RECT 303.115 -217.765 303.445 -217.435 ;
        RECT 303.115 -219.125 303.445 -218.795 ;
        RECT 303.115 -220.485 303.445 -220.155 ;
        RECT 303.115 -221.845 303.445 -221.515 ;
        RECT 303.115 -223.205 303.445 -222.875 ;
        RECT 303.115 -224.565 303.445 -224.235 ;
        RECT 303.115 -225.925 303.445 -225.595 ;
        RECT 303.115 -227.285 303.445 -226.955 ;
        RECT 303.115 -228.645 303.445 -228.315 ;
        RECT 303.115 -230.005 303.445 -229.675 ;
        RECT 303.115 -231.365 303.445 -231.035 ;
        RECT 303.115 -232.725 303.445 -232.395 ;
        RECT 303.115 -234.085 303.445 -233.755 ;
        RECT 303.115 -235.445 303.445 -235.115 ;
        RECT 303.115 -236.805 303.445 -236.475 ;
        RECT 303.115 -238.165 303.445 -237.835 ;
        RECT 303.115 -243.81 303.445 -242.68 ;
        RECT 303.12 -243.925 303.44 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 246.76 304.805 247.89 ;
        RECT 304.475 241.915 304.805 242.245 ;
        RECT 304.475 240.555 304.805 240.885 ;
        RECT 304.475 239.195 304.805 239.525 ;
        RECT 304.475 237.835 304.805 238.165 ;
        RECT 304.48 237.16 304.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 -1.525 304.805 -1.195 ;
        RECT 304.475 -2.885 304.805 -2.555 ;
        RECT 304.48 -3.56 304.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 -122.565 304.805 -122.235 ;
        RECT 304.475 -123.925 304.805 -123.595 ;
        RECT 304.475 -125.285 304.805 -124.955 ;
        RECT 304.475 -126.645 304.805 -126.315 ;
        RECT 304.475 -128.005 304.805 -127.675 ;
        RECT 304.475 -129.365 304.805 -129.035 ;
        RECT 304.475 -130.725 304.805 -130.395 ;
        RECT 304.475 -132.085 304.805 -131.755 ;
        RECT 304.475 -133.445 304.805 -133.115 ;
        RECT 304.475 -134.805 304.805 -134.475 ;
        RECT 304.475 -136.165 304.805 -135.835 ;
        RECT 304.475 -137.525 304.805 -137.195 ;
        RECT 304.475 -138.885 304.805 -138.555 ;
        RECT 304.475 -140.245 304.805 -139.915 ;
        RECT 304.475 -141.605 304.805 -141.275 ;
        RECT 304.475 -142.965 304.805 -142.635 ;
        RECT 304.475 -144.325 304.805 -143.995 ;
        RECT 304.475 -145.685 304.805 -145.355 ;
        RECT 304.475 -147.045 304.805 -146.715 ;
        RECT 304.475 -148.405 304.805 -148.075 ;
        RECT 304.475 -149.765 304.805 -149.435 ;
        RECT 304.475 -151.125 304.805 -150.795 ;
        RECT 304.475 -152.485 304.805 -152.155 ;
        RECT 304.475 -153.845 304.805 -153.515 ;
        RECT 304.475 -155.205 304.805 -154.875 ;
        RECT 304.475 -156.565 304.805 -156.235 ;
        RECT 304.475 -157.925 304.805 -157.595 ;
        RECT 304.475 -159.285 304.805 -158.955 ;
        RECT 304.475 -160.645 304.805 -160.315 ;
        RECT 304.475 -162.005 304.805 -161.675 ;
        RECT 304.475 -163.365 304.805 -163.035 ;
        RECT 304.475 -164.725 304.805 -164.395 ;
        RECT 304.475 -166.085 304.805 -165.755 ;
        RECT 304.475 -167.445 304.805 -167.115 ;
        RECT 304.475 -168.805 304.805 -168.475 ;
        RECT 304.475 -170.165 304.805 -169.835 ;
        RECT 304.475 -171.525 304.805 -171.195 ;
        RECT 304.475 -172.885 304.805 -172.555 ;
        RECT 304.475 -174.245 304.805 -173.915 ;
        RECT 304.475 -175.605 304.805 -175.275 ;
        RECT 304.475 -176.965 304.805 -176.635 ;
        RECT 304.475 -178.325 304.805 -177.995 ;
        RECT 304.475 -179.685 304.805 -179.355 ;
        RECT 304.475 -181.045 304.805 -180.715 ;
        RECT 304.475 -182.405 304.805 -182.075 ;
        RECT 304.475 -183.765 304.805 -183.435 ;
        RECT 304.475 -185.125 304.805 -184.795 ;
        RECT 304.475 -186.485 304.805 -186.155 ;
        RECT 304.475 -187.845 304.805 -187.515 ;
        RECT 304.475 -189.205 304.805 -188.875 ;
        RECT 304.475 -190.565 304.805 -190.235 ;
        RECT 304.475 -191.925 304.805 -191.595 ;
        RECT 304.475 -193.285 304.805 -192.955 ;
        RECT 304.475 -194.645 304.805 -194.315 ;
        RECT 304.475 -196.005 304.805 -195.675 ;
        RECT 304.475 -197.365 304.805 -197.035 ;
        RECT 304.475 -198.725 304.805 -198.395 ;
        RECT 304.475 -200.085 304.805 -199.755 ;
        RECT 304.475 -201.445 304.805 -201.115 ;
        RECT 304.475 -202.805 304.805 -202.475 ;
        RECT 304.475 -204.165 304.805 -203.835 ;
        RECT 304.475 -205.525 304.805 -205.195 ;
        RECT 304.475 -206.885 304.805 -206.555 ;
        RECT 304.475 -208.245 304.805 -207.915 ;
        RECT 304.475 -209.605 304.805 -209.275 ;
        RECT 304.475 -210.965 304.805 -210.635 ;
        RECT 304.475 -212.325 304.805 -211.995 ;
        RECT 304.475 -213.685 304.805 -213.355 ;
        RECT 304.475 -215.045 304.805 -214.715 ;
        RECT 304.475 -216.405 304.805 -216.075 ;
        RECT 304.475 -217.765 304.805 -217.435 ;
        RECT 304.475 -219.125 304.805 -218.795 ;
        RECT 304.475 -220.485 304.805 -220.155 ;
        RECT 304.475 -221.845 304.805 -221.515 ;
        RECT 304.475 -223.205 304.805 -222.875 ;
        RECT 304.475 -224.565 304.805 -224.235 ;
        RECT 304.475 -225.925 304.805 -225.595 ;
        RECT 304.475 -227.285 304.805 -226.955 ;
        RECT 304.475 -228.645 304.805 -228.315 ;
        RECT 304.475 -230.005 304.805 -229.675 ;
        RECT 304.475 -231.365 304.805 -231.035 ;
        RECT 304.475 -232.725 304.805 -232.395 ;
        RECT 304.475 -234.085 304.805 -233.755 ;
        RECT 304.475 -235.445 304.805 -235.115 ;
        RECT 304.475 -236.805 304.805 -236.475 ;
        RECT 304.475 -238.165 304.805 -237.835 ;
        RECT 304.475 -243.81 304.805 -242.68 ;
        RECT 304.48 -243.925 304.8 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 246.76 306.165 247.89 ;
        RECT 305.835 241.915 306.165 242.245 ;
        RECT 305.835 240.555 306.165 240.885 ;
        RECT 305.835 239.195 306.165 239.525 ;
        RECT 305.835 237.835 306.165 238.165 ;
        RECT 305.84 237.16 306.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 -1.525 306.165 -1.195 ;
        RECT 305.835 -2.885 306.165 -2.555 ;
        RECT 305.84 -3.56 306.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 -122.565 306.165 -122.235 ;
        RECT 305.835 -123.925 306.165 -123.595 ;
        RECT 305.835 -125.285 306.165 -124.955 ;
        RECT 305.835 -126.645 306.165 -126.315 ;
        RECT 305.835 -128.005 306.165 -127.675 ;
        RECT 305.835 -129.365 306.165 -129.035 ;
        RECT 305.835 -130.725 306.165 -130.395 ;
        RECT 305.835 -132.085 306.165 -131.755 ;
        RECT 305.835 -133.445 306.165 -133.115 ;
        RECT 305.835 -134.805 306.165 -134.475 ;
        RECT 305.835 -136.165 306.165 -135.835 ;
        RECT 305.835 -137.525 306.165 -137.195 ;
        RECT 305.835 -138.885 306.165 -138.555 ;
        RECT 305.835 -140.245 306.165 -139.915 ;
        RECT 305.835 -141.605 306.165 -141.275 ;
        RECT 305.835 -142.965 306.165 -142.635 ;
        RECT 305.835 -144.325 306.165 -143.995 ;
        RECT 305.835 -145.685 306.165 -145.355 ;
        RECT 305.835 -147.045 306.165 -146.715 ;
        RECT 305.835 -148.405 306.165 -148.075 ;
        RECT 305.835 -149.765 306.165 -149.435 ;
        RECT 305.835 -151.125 306.165 -150.795 ;
        RECT 305.835 -152.485 306.165 -152.155 ;
        RECT 305.835 -153.845 306.165 -153.515 ;
        RECT 305.835 -155.205 306.165 -154.875 ;
        RECT 305.835 -156.565 306.165 -156.235 ;
        RECT 305.835 -157.925 306.165 -157.595 ;
        RECT 305.835 -159.285 306.165 -158.955 ;
        RECT 305.835 -160.645 306.165 -160.315 ;
        RECT 305.835 -162.005 306.165 -161.675 ;
        RECT 305.835 -163.365 306.165 -163.035 ;
        RECT 305.835 -164.725 306.165 -164.395 ;
        RECT 305.835 -166.085 306.165 -165.755 ;
        RECT 305.835 -167.445 306.165 -167.115 ;
        RECT 305.835 -168.805 306.165 -168.475 ;
        RECT 305.835 -170.165 306.165 -169.835 ;
        RECT 305.835 -171.525 306.165 -171.195 ;
        RECT 305.835 -172.885 306.165 -172.555 ;
        RECT 305.835 -174.245 306.165 -173.915 ;
        RECT 305.835 -175.605 306.165 -175.275 ;
        RECT 305.835 -176.965 306.165 -176.635 ;
        RECT 305.835 -178.325 306.165 -177.995 ;
        RECT 305.835 -179.685 306.165 -179.355 ;
        RECT 305.835 -181.045 306.165 -180.715 ;
        RECT 305.835 -182.405 306.165 -182.075 ;
        RECT 305.835 -183.765 306.165 -183.435 ;
        RECT 305.835 -185.125 306.165 -184.795 ;
        RECT 305.835 -186.485 306.165 -186.155 ;
        RECT 305.835 -187.845 306.165 -187.515 ;
        RECT 305.835 -189.205 306.165 -188.875 ;
        RECT 305.835 -190.565 306.165 -190.235 ;
        RECT 305.835 -191.925 306.165 -191.595 ;
        RECT 305.835 -193.285 306.165 -192.955 ;
        RECT 305.835 -194.645 306.165 -194.315 ;
        RECT 305.835 -196.005 306.165 -195.675 ;
        RECT 305.835 -197.365 306.165 -197.035 ;
        RECT 305.835 -198.725 306.165 -198.395 ;
        RECT 305.835 -200.085 306.165 -199.755 ;
        RECT 305.835 -201.445 306.165 -201.115 ;
        RECT 305.835 -202.805 306.165 -202.475 ;
        RECT 305.835 -204.165 306.165 -203.835 ;
        RECT 305.835 -205.525 306.165 -205.195 ;
        RECT 305.835 -206.885 306.165 -206.555 ;
        RECT 305.835 -208.245 306.165 -207.915 ;
        RECT 305.835 -209.605 306.165 -209.275 ;
        RECT 305.835 -210.965 306.165 -210.635 ;
        RECT 305.835 -212.325 306.165 -211.995 ;
        RECT 305.835 -213.685 306.165 -213.355 ;
        RECT 305.835 -215.045 306.165 -214.715 ;
        RECT 305.835 -216.405 306.165 -216.075 ;
        RECT 305.835 -217.765 306.165 -217.435 ;
        RECT 305.835 -219.125 306.165 -218.795 ;
        RECT 305.835 -220.485 306.165 -220.155 ;
        RECT 305.835 -221.845 306.165 -221.515 ;
        RECT 305.835 -223.205 306.165 -222.875 ;
        RECT 305.835 -224.565 306.165 -224.235 ;
        RECT 305.835 -225.925 306.165 -225.595 ;
        RECT 305.835 -227.285 306.165 -226.955 ;
        RECT 305.835 -228.645 306.165 -228.315 ;
        RECT 305.835 -230.005 306.165 -229.675 ;
        RECT 305.835 -231.365 306.165 -231.035 ;
        RECT 305.835 -232.725 306.165 -232.395 ;
        RECT 305.835 -234.085 306.165 -233.755 ;
        RECT 305.835 -235.445 306.165 -235.115 ;
        RECT 305.835 -236.805 306.165 -236.475 ;
        RECT 305.835 -238.165 306.165 -237.835 ;
        RECT 305.835 -243.81 306.165 -242.68 ;
        RECT 305.84 -243.925 306.16 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 246.76 307.525 247.89 ;
        RECT 307.195 241.915 307.525 242.245 ;
        RECT 307.195 240.555 307.525 240.885 ;
        RECT 307.195 239.195 307.525 239.525 ;
        RECT 307.195 237.835 307.525 238.165 ;
        RECT 307.2 237.16 307.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 -126.645 307.525 -126.315 ;
        RECT 307.195 -128.005 307.525 -127.675 ;
        RECT 307.195 -129.365 307.525 -129.035 ;
        RECT 307.195 -130.725 307.525 -130.395 ;
        RECT 307.195 -132.085 307.525 -131.755 ;
        RECT 307.195 -133.445 307.525 -133.115 ;
        RECT 307.195 -134.805 307.525 -134.475 ;
        RECT 307.195 -136.165 307.525 -135.835 ;
        RECT 307.195 -137.525 307.525 -137.195 ;
        RECT 307.195 -138.885 307.525 -138.555 ;
        RECT 307.195 -140.245 307.525 -139.915 ;
        RECT 307.195 -141.605 307.525 -141.275 ;
        RECT 307.195 -142.965 307.525 -142.635 ;
        RECT 307.195 -144.325 307.525 -143.995 ;
        RECT 307.195 -145.685 307.525 -145.355 ;
        RECT 307.195 -147.045 307.525 -146.715 ;
        RECT 307.195 -148.405 307.525 -148.075 ;
        RECT 307.195 -149.765 307.525 -149.435 ;
        RECT 307.195 -151.125 307.525 -150.795 ;
        RECT 307.195 -152.485 307.525 -152.155 ;
        RECT 307.195 -153.845 307.525 -153.515 ;
        RECT 307.195 -155.205 307.525 -154.875 ;
        RECT 307.195 -156.565 307.525 -156.235 ;
        RECT 307.195 -157.925 307.525 -157.595 ;
        RECT 307.195 -159.285 307.525 -158.955 ;
        RECT 307.195 -160.645 307.525 -160.315 ;
        RECT 307.195 -162.005 307.525 -161.675 ;
        RECT 307.195 -163.365 307.525 -163.035 ;
        RECT 307.195 -164.725 307.525 -164.395 ;
        RECT 307.195 -166.085 307.525 -165.755 ;
        RECT 307.195 -167.445 307.525 -167.115 ;
        RECT 307.195 -168.805 307.525 -168.475 ;
        RECT 307.195 -170.165 307.525 -169.835 ;
        RECT 307.195 -171.525 307.525 -171.195 ;
        RECT 307.195 -172.885 307.525 -172.555 ;
        RECT 307.195 -174.245 307.525 -173.915 ;
        RECT 307.195 -175.605 307.525 -175.275 ;
        RECT 307.195 -176.965 307.525 -176.635 ;
        RECT 307.195 -178.325 307.525 -177.995 ;
        RECT 307.195 -179.685 307.525 -179.355 ;
        RECT 307.195 -181.045 307.525 -180.715 ;
        RECT 307.195 -182.405 307.525 -182.075 ;
        RECT 307.195 -183.765 307.525 -183.435 ;
        RECT 307.195 -185.125 307.525 -184.795 ;
        RECT 307.195 -186.485 307.525 -186.155 ;
        RECT 307.195 -187.845 307.525 -187.515 ;
        RECT 307.195 -189.205 307.525 -188.875 ;
        RECT 307.195 -190.565 307.525 -190.235 ;
        RECT 307.195 -191.925 307.525 -191.595 ;
        RECT 307.195 -193.285 307.525 -192.955 ;
        RECT 307.195 -194.645 307.525 -194.315 ;
        RECT 307.195 -196.005 307.525 -195.675 ;
        RECT 307.195 -197.365 307.525 -197.035 ;
        RECT 307.195 -198.725 307.525 -198.395 ;
        RECT 307.195 -200.085 307.525 -199.755 ;
        RECT 307.195 -201.445 307.525 -201.115 ;
        RECT 307.195 -202.805 307.525 -202.475 ;
        RECT 307.195 -204.165 307.525 -203.835 ;
        RECT 307.195 -205.525 307.525 -205.195 ;
        RECT 307.195 -206.885 307.525 -206.555 ;
        RECT 307.195 -208.245 307.525 -207.915 ;
        RECT 307.195 -209.605 307.525 -209.275 ;
        RECT 307.195 -210.965 307.525 -210.635 ;
        RECT 307.195 -212.325 307.525 -211.995 ;
        RECT 307.195 -213.685 307.525 -213.355 ;
        RECT 307.195 -215.045 307.525 -214.715 ;
        RECT 307.195 -216.405 307.525 -216.075 ;
        RECT 307.195 -217.765 307.525 -217.435 ;
        RECT 307.195 -219.125 307.525 -218.795 ;
        RECT 307.195 -220.485 307.525 -220.155 ;
        RECT 307.195 -221.845 307.525 -221.515 ;
        RECT 307.195 -223.205 307.525 -222.875 ;
        RECT 307.195 -224.565 307.525 -224.235 ;
        RECT 307.195 -225.925 307.525 -225.595 ;
        RECT 307.195 -227.285 307.525 -226.955 ;
        RECT 307.195 -228.645 307.525 -228.315 ;
        RECT 307.195 -230.005 307.525 -229.675 ;
        RECT 307.195 -231.365 307.525 -231.035 ;
        RECT 307.195 -232.725 307.525 -232.395 ;
        RECT 307.195 -234.085 307.525 -233.755 ;
        RECT 307.195 -235.445 307.525 -235.115 ;
        RECT 307.195 -236.805 307.525 -236.475 ;
        RECT 307.195 -238.165 307.525 -237.835 ;
        RECT 307.195 -243.81 307.525 -242.68 ;
        RECT 307.2 -243.925 307.52 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.86 -125.535 308.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.555 246.76 308.885 247.89 ;
        RECT 308.555 241.915 308.885 242.245 ;
        RECT 308.555 240.555 308.885 240.885 ;
        RECT 308.555 239.195 308.885 239.525 ;
        RECT 308.555 237.835 308.885 238.165 ;
        RECT 308.56 237.16 308.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 246.76 310.245 247.89 ;
        RECT 309.915 241.915 310.245 242.245 ;
        RECT 309.915 240.555 310.245 240.885 ;
        RECT 309.915 239.195 310.245 239.525 ;
        RECT 309.915 237.835 310.245 238.165 ;
        RECT 309.92 237.16 310.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 -1.525 310.245 -1.195 ;
        RECT 309.915 -2.885 310.245 -2.555 ;
        RECT 309.92 -3.56 310.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 246.76 311.605 247.89 ;
        RECT 311.275 241.915 311.605 242.245 ;
        RECT 311.275 240.555 311.605 240.885 ;
        RECT 311.275 239.195 311.605 239.525 ;
        RECT 311.275 237.835 311.605 238.165 ;
        RECT 311.28 237.16 311.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 -1.525 311.605 -1.195 ;
        RECT 311.275 -2.885 311.605 -2.555 ;
        RECT 311.28 -3.56 311.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 246.76 312.965 247.89 ;
        RECT 312.635 241.915 312.965 242.245 ;
        RECT 312.635 240.555 312.965 240.885 ;
        RECT 312.635 239.195 312.965 239.525 ;
        RECT 312.635 237.835 312.965 238.165 ;
        RECT 312.64 237.16 312.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 -1.525 312.965 -1.195 ;
        RECT 312.635 -2.885 312.965 -2.555 ;
        RECT 312.64 -3.56 312.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 -122.565 312.965 -122.235 ;
        RECT 312.635 -123.925 312.965 -123.595 ;
        RECT 312.635 -125.285 312.965 -124.955 ;
        RECT 312.635 -126.645 312.965 -126.315 ;
        RECT 312.635 -128.005 312.965 -127.675 ;
        RECT 312.635 -129.365 312.965 -129.035 ;
        RECT 312.635 -130.725 312.965 -130.395 ;
        RECT 312.635 -132.085 312.965 -131.755 ;
        RECT 312.635 -133.445 312.965 -133.115 ;
        RECT 312.635 -134.805 312.965 -134.475 ;
        RECT 312.635 -136.165 312.965 -135.835 ;
        RECT 312.635 -137.525 312.965 -137.195 ;
        RECT 312.635 -138.885 312.965 -138.555 ;
        RECT 312.635 -140.245 312.965 -139.915 ;
        RECT 312.635 -141.605 312.965 -141.275 ;
        RECT 312.635 -142.965 312.965 -142.635 ;
        RECT 312.635 -144.325 312.965 -143.995 ;
        RECT 312.635 -145.685 312.965 -145.355 ;
        RECT 312.635 -147.045 312.965 -146.715 ;
        RECT 312.635 -148.405 312.965 -148.075 ;
        RECT 312.635 -149.765 312.965 -149.435 ;
        RECT 312.635 -151.125 312.965 -150.795 ;
        RECT 312.635 -152.485 312.965 -152.155 ;
        RECT 312.635 -153.845 312.965 -153.515 ;
        RECT 312.635 -155.205 312.965 -154.875 ;
        RECT 312.635 -156.565 312.965 -156.235 ;
        RECT 312.635 -157.925 312.965 -157.595 ;
        RECT 312.635 -159.285 312.965 -158.955 ;
        RECT 312.635 -160.645 312.965 -160.315 ;
        RECT 312.635 -162.005 312.965 -161.675 ;
        RECT 312.635 -163.365 312.965 -163.035 ;
        RECT 312.635 -164.725 312.965 -164.395 ;
        RECT 312.635 -166.085 312.965 -165.755 ;
        RECT 312.635 -167.445 312.965 -167.115 ;
        RECT 312.635 -168.805 312.965 -168.475 ;
        RECT 312.635 -170.165 312.965 -169.835 ;
        RECT 312.635 -171.525 312.965 -171.195 ;
        RECT 312.635 -172.885 312.965 -172.555 ;
        RECT 312.635 -174.245 312.965 -173.915 ;
        RECT 312.635 -175.605 312.965 -175.275 ;
        RECT 312.635 -176.965 312.965 -176.635 ;
        RECT 312.635 -178.325 312.965 -177.995 ;
        RECT 312.635 -179.685 312.965 -179.355 ;
        RECT 312.635 -181.045 312.965 -180.715 ;
        RECT 312.635 -182.405 312.965 -182.075 ;
        RECT 312.635 -183.765 312.965 -183.435 ;
        RECT 312.635 -185.125 312.965 -184.795 ;
        RECT 312.635 -186.485 312.965 -186.155 ;
        RECT 312.635 -187.845 312.965 -187.515 ;
        RECT 312.635 -189.205 312.965 -188.875 ;
        RECT 312.635 -190.565 312.965 -190.235 ;
        RECT 312.635 -191.925 312.965 -191.595 ;
        RECT 312.635 -193.285 312.965 -192.955 ;
        RECT 312.635 -194.645 312.965 -194.315 ;
        RECT 312.635 -196.005 312.965 -195.675 ;
        RECT 312.635 -197.365 312.965 -197.035 ;
        RECT 312.635 -198.725 312.965 -198.395 ;
        RECT 312.635 -200.085 312.965 -199.755 ;
        RECT 312.635 -201.445 312.965 -201.115 ;
        RECT 312.635 -202.805 312.965 -202.475 ;
        RECT 312.635 -204.165 312.965 -203.835 ;
        RECT 312.635 -205.525 312.965 -205.195 ;
        RECT 312.635 -206.885 312.965 -206.555 ;
        RECT 312.635 -208.245 312.965 -207.915 ;
        RECT 312.635 -209.605 312.965 -209.275 ;
        RECT 312.635 -210.965 312.965 -210.635 ;
        RECT 312.635 -212.325 312.965 -211.995 ;
        RECT 312.635 -213.685 312.965 -213.355 ;
        RECT 312.635 -215.045 312.965 -214.715 ;
        RECT 312.635 -216.405 312.965 -216.075 ;
        RECT 312.635 -217.765 312.965 -217.435 ;
        RECT 312.635 -219.125 312.965 -218.795 ;
        RECT 312.635 -220.485 312.965 -220.155 ;
        RECT 312.635 -221.845 312.965 -221.515 ;
        RECT 312.635 -223.205 312.965 -222.875 ;
        RECT 312.635 -224.565 312.965 -224.235 ;
        RECT 312.635 -225.925 312.965 -225.595 ;
        RECT 312.635 -227.285 312.965 -226.955 ;
        RECT 312.635 -228.645 312.965 -228.315 ;
        RECT 312.635 -230.005 312.965 -229.675 ;
        RECT 312.635 -231.365 312.965 -231.035 ;
        RECT 312.635 -232.725 312.965 -232.395 ;
        RECT 312.635 -234.085 312.965 -233.755 ;
        RECT 312.635 -235.445 312.965 -235.115 ;
        RECT 312.635 -236.805 312.965 -236.475 ;
        RECT 312.635 -238.165 312.965 -237.835 ;
        RECT 312.635 -243.81 312.965 -242.68 ;
        RECT 312.64 -243.925 312.96 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 246.76 314.325 247.89 ;
        RECT 313.995 241.915 314.325 242.245 ;
        RECT 313.995 240.555 314.325 240.885 ;
        RECT 313.995 239.195 314.325 239.525 ;
        RECT 313.995 237.835 314.325 238.165 ;
        RECT 314 237.16 314.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 -1.525 314.325 -1.195 ;
        RECT 313.995 -2.885 314.325 -2.555 ;
        RECT 314 -3.56 314.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 -122.565 314.325 -122.235 ;
        RECT 313.995 -123.925 314.325 -123.595 ;
        RECT 313.995 -125.285 314.325 -124.955 ;
        RECT 313.995 -126.645 314.325 -126.315 ;
        RECT 313.995 -128.005 314.325 -127.675 ;
        RECT 313.995 -129.365 314.325 -129.035 ;
        RECT 313.995 -130.725 314.325 -130.395 ;
        RECT 313.995 -132.085 314.325 -131.755 ;
        RECT 313.995 -133.445 314.325 -133.115 ;
        RECT 313.995 -134.805 314.325 -134.475 ;
        RECT 313.995 -136.165 314.325 -135.835 ;
        RECT 313.995 -137.525 314.325 -137.195 ;
        RECT 313.995 -138.885 314.325 -138.555 ;
        RECT 313.995 -140.245 314.325 -139.915 ;
        RECT 313.995 -141.605 314.325 -141.275 ;
        RECT 313.995 -142.965 314.325 -142.635 ;
        RECT 313.995 -144.325 314.325 -143.995 ;
        RECT 313.995 -145.685 314.325 -145.355 ;
        RECT 313.995 -147.045 314.325 -146.715 ;
        RECT 313.995 -148.405 314.325 -148.075 ;
        RECT 313.995 -149.765 314.325 -149.435 ;
        RECT 313.995 -151.125 314.325 -150.795 ;
        RECT 313.995 -152.485 314.325 -152.155 ;
        RECT 313.995 -153.845 314.325 -153.515 ;
        RECT 313.995 -155.205 314.325 -154.875 ;
        RECT 313.995 -156.565 314.325 -156.235 ;
        RECT 313.995 -157.925 314.325 -157.595 ;
        RECT 313.995 -159.285 314.325 -158.955 ;
        RECT 313.995 -160.645 314.325 -160.315 ;
        RECT 313.995 -162.005 314.325 -161.675 ;
        RECT 313.995 -163.365 314.325 -163.035 ;
        RECT 313.995 -164.725 314.325 -164.395 ;
        RECT 313.995 -166.085 314.325 -165.755 ;
        RECT 313.995 -167.445 314.325 -167.115 ;
        RECT 313.995 -168.805 314.325 -168.475 ;
        RECT 313.995 -170.165 314.325 -169.835 ;
        RECT 313.995 -171.525 314.325 -171.195 ;
        RECT 313.995 -172.885 314.325 -172.555 ;
        RECT 313.995 -174.245 314.325 -173.915 ;
        RECT 313.995 -175.605 314.325 -175.275 ;
        RECT 313.995 -176.965 314.325 -176.635 ;
        RECT 313.995 -178.325 314.325 -177.995 ;
        RECT 313.995 -179.685 314.325 -179.355 ;
        RECT 313.995 -181.045 314.325 -180.715 ;
        RECT 313.995 -182.405 314.325 -182.075 ;
        RECT 313.995 -183.765 314.325 -183.435 ;
        RECT 313.995 -185.125 314.325 -184.795 ;
        RECT 313.995 -186.485 314.325 -186.155 ;
        RECT 313.995 -187.845 314.325 -187.515 ;
        RECT 313.995 -189.205 314.325 -188.875 ;
        RECT 313.995 -190.565 314.325 -190.235 ;
        RECT 313.995 -191.925 314.325 -191.595 ;
        RECT 313.995 -193.285 314.325 -192.955 ;
        RECT 313.995 -194.645 314.325 -194.315 ;
        RECT 313.995 -196.005 314.325 -195.675 ;
        RECT 313.995 -197.365 314.325 -197.035 ;
        RECT 313.995 -198.725 314.325 -198.395 ;
        RECT 313.995 -200.085 314.325 -199.755 ;
        RECT 313.995 -201.445 314.325 -201.115 ;
        RECT 313.995 -202.805 314.325 -202.475 ;
        RECT 313.995 -204.165 314.325 -203.835 ;
        RECT 313.995 -205.525 314.325 -205.195 ;
        RECT 313.995 -206.885 314.325 -206.555 ;
        RECT 313.995 -208.245 314.325 -207.915 ;
        RECT 313.995 -209.605 314.325 -209.275 ;
        RECT 313.995 -210.965 314.325 -210.635 ;
        RECT 313.995 -212.325 314.325 -211.995 ;
        RECT 313.995 -213.685 314.325 -213.355 ;
        RECT 313.995 -215.045 314.325 -214.715 ;
        RECT 313.995 -216.405 314.325 -216.075 ;
        RECT 313.995 -217.765 314.325 -217.435 ;
        RECT 313.995 -219.125 314.325 -218.795 ;
        RECT 313.995 -220.485 314.325 -220.155 ;
        RECT 313.995 -221.845 314.325 -221.515 ;
        RECT 313.995 -223.205 314.325 -222.875 ;
        RECT 313.995 -224.565 314.325 -224.235 ;
        RECT 313.995 -225.925 314.325 -225.595 ;
        RECT 313.995 -227.285 314.325 -226.955 ;
        RECT 313.995 -228.645 314.325 -228.315 ;
        RECT 313.995 -230.005 314.325 -229.675 ;
        RECT 313.995 -231.365 314.325 -231.035 ;
        RECT 313.995 -232.725 314.325 -232.395 ;
        RECT 313.995 -234.085 314.325 -233.755 ;
        RECT 313.995 -235.445 314.325 -235.115 ;
        RECT 313.995 -236.805 314.325 -236.475 ;
        RECT 313.995 -238.165 314.325 -237.835 ;
        RECT 313.995 -243.81 314.325 -242.68 ;
        RECT 314 -243.925 314.32 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 246.76 315.685 247.89 ;
        RECT 315.355 241.915 315.685 242.245 ;
        RECT 315.355 240.555 315.685 240.885 ;
        RECT 315.355 239.195 315.685 239.525 ;
        RECT 315.355 237.835 315.685 238.165 ;
        RECT 315.36 237.16 315.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 -1.525 315.685 -1.195 ;
        RECT 315.355 -2.885 315.685 -2.555 ;
        RECT 315.36 -3.56 315.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 -122.565 315.685 -122.235 ;
        RECT 315.355 -123.925 315.685 -123.595 ;
        RECT 315.355 -125.285 315.685 -124.955 ;
        RECT 315.355 -126.645 315.685 -126.315 ;
        RECT 315.355 -128.005 315.685 -127.675 ;
        RECT 315.355 -129.365 315.685 -129.035 ;
        RECT 315.355 -130.725 315.685 -130.395 ;
        RECT 315.355 -132.085 315.685 -131.755 ;
        RECT 315.355 -133.445 315.685 -133.115 ;
        RECT 315.355 -134.805 315.685 -134.475 ;
        RECT 315.355 -136.165 315.685 -135.835 ;
        RECT 315.355 -137.525 315.685 -137.195 ;
        RECT 315.355 -138.885 315.685 -138.555 ;
        RECT 315.355 -140.245 315.685 -139.915 ;
        RECT 315.355 -141.605 315.685 -141.275 ;
        RECT 315.355 -142.965 315.685 -142.635 ;
        RECT 315.355 -144.325 315.685 -143.995 ;
        RECT 315.355 -145.685 315.685 -145.355 ;
        RECT 315.355 -147.045 315.685 -146.715 ;
        RECT 315.355 -148.405 315.685 -148.075 ;
        RECT 315.355 -149.765 315.685 -149.435 ;
        RECT 315.355 -151.125 315.685 -150.795 ;
        RECT 315.355 -152.485 315.685 -152.155 ;
        RECT 315.355 -153.845 315.685 -153.515 ;
        RECT 315.355 -155.205 315.685 -154.875 ;
        RECT 315.355 -156.565 315.685 -156.235 ;
        RECT 315.355 -157.925 315.685 -157.595 ;
        RECT 315.355 -159.285 315.685 -158.955 ;
        RECT 315.355 -160.645 315.685 -160.315 ;
        RECT 315.355 -162.005 315.685 -161.675 ;
        RECT 315.355 -163.365 315.685 -163.035 ;
        RECT 315.355 -164.725 315.685 -164.395 ;
        RECT 315.355 -166.085 315.685 -165.755 ;
        RECT 315.355 -167.445 315.685 -167.115 ;
        RECT 315.355 -168.805 315.685 -168.475 ;
        RECT 315.355 -170.165 315.685 -169.835 ;
        RECT 315.355 -171.525 315.685 -171.195 ;
        RECT 315.355 -172.885 315.685 -172.555 ;
        RECT 315.355 -174.245 315.685 -173.915 ;
        RECT 315.355 -175.605 315.685 -175.275 ;
        RECT 315.355 -176.965 315.685 -176.635 ;
        RECT 315.355 -178.325 315.685 -177.995 ;
        RECT 315.355 -179.685 315.685 -179.355 ;
        RECT 315.355 -181.045 315.685 -180.715 ;
        RECT 315.355 -182.405 315.685 -182.075 ;
        RECT 315.355 -183.765 315.685 -183.435 ;
        RECT 315.355 -185.125 315.685 -184.795 ;
        RECT 315.355 -186.485 315.685 -186.155 ;
        RECT 315.355 -187.845 315.685 -187.515 ;
        RECT 315.355 -189.205 315.685 -188.875 ;
        RECT 315.355 -190.565 315.685 -190.235 ;
        RECT 315.355 -191.925 315.685 -191.595 ;
        RECT 315.355 -193.285 315.685 -192.955 ;
        RECT 315.355 -194.645 315.685 -194.315 ;
        RECT 315.355 -196.005 315.685 -195.675 ;
        RECT 315.355 -197.365 315.685 -197.035 ;
        RECT 315.355 -198.725 315.685 -198.395 ;
        RECT 315.355 -200.085 315.685 -199.755 ;
        RECT 315.355 -201.445 315.685 -201.115 ;
        RECT 315.355 -202.805 315.685 -202.475 ;
        RECT 315.355 -204.165 315.685 -203.835 ;
        RECT 315.355 -205.525 315.685 -205.195 ;
        RECT 315.355 -206.885 315.685 -206.555 ;
        RECT 315.355 -208.245 315.685 -207.915 ;
        RECT 315.355 -209.605 315.685 -209.275 ;
        RECT 315.355 -210.965 315.685 -210.635 ;
        RECT 315.355 -212.325 315.685 -211.995 ;
        RECT 315.355 -213.685 315.685 -213.355 ;
        RECT 315.355 -215.045 315.685 -214.715 ;
        RECT 315.355 -216.405 315.685 -216.075 ;
        RECT 315.355 -217.765 315.685 -217.435 ;
        RECT 315.355 -219.125 315.685 -218.795 ;
        RECT 315.355 -220.485 315.685 -220.155 ;
        RECT 315.355 -221.845 315.685 -221.515 ;
        RECT 315.355 -223.205 315.685 -222.875 ;
        RECT 315.355 -224.565 315.685 -224.235 ;
        RECT 315.355 -225.925 315.685 -225.595 ;
        RECT 315.355 -227.285 315.685 -226.955 ;
        RECT 315.355 -228.645 315.685 -228.315 ;
        RECT 315.355 -230.005 315.685 -229.675 ;
        RECT 315.355 -231.365 315.685 -231.035 ;
        RECT 315.355 -232.725 315.685 -232.395 ;
        RECT 315.355 -234.085 315.685 -233.755 ;
        RECT 315.355 -235.445 315.685 -235.115 ;
        RECT 315.355 -236.805 315.685 -236.475 ;
        RECT 315.355 -238.165 315.685 -237.835 ;
        RECT 315.355 -243.81 315.685 -242.68 ;
        RECT 315.36 -243.925 315.68 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 246.76 317.045 247.89 ;
        RECT 316.715 241.915 317.045 242.245 ;
        RECT 316.715 240.555 317.045 240.885 ;
        RECT 316.715 239.195 317.045 239.525 ;
        RECT 316.715 237.835 317.045 238.165 ;
        RECT 316.72 237.16 317.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 -1.525 317.045 -1.195 ;
        RECT 316.715 -2.885 317.045 -2.555 ;
        RECT 316.72 -3.56 317.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 -122.565 317.045 -122.235 ;
        RECT 316.715 -123.925 317.045 -123.595 ;
        RECT 316.715 -125.285 317.045 -124.955 ;
        RECT 316.715 -126.645 317.045 -126.315 ;
        RECT 316.715 -128.005 317.045 -127.675 ;
        RECT 316.715 -129.365 317.045 -129.035 ;
        RECT 316.715 -130.725 317.045 -130.395 ;
        RECT 316.715 -132.085 317.045 -131.755 ;
        RECT 316.715 -133.445 317.045 -133.115 ;
        RECT 316.715 -134.805 317.045 -134.475 ;
        RECT 316.715 -136.165 317.045 -135.835 ;
        RECT 316.715 -137.525 317.045 -137.195 ;
        RECT 316.715 -138.885 317.045 -138.555 ;
        RECT 316.715 -140.245 317.045 -139.915 ;
        RECT 316.715 -141.605 317.045 -141.275 ;
        RECT 316.715 -142.965 317.045 -142.635 ;
        RECT 316.715 -144.325 317.045 -143.995 ;
        RECT 316.715 -145.685 317.045 -145.355 ;
        RECT 316.715 -147.045 317.045 -146.715 ;
        RECT 316.715 -148.405 317.045 -148.075 ;
        RECT 316.715 -149.765 317.045 -149.435 ;
        RECT 316.715 -151.125 317.045 -150.795 ;
        RECT 316.715 -152.485 317.045 -152.155 ;
        RECT 316.715 -153.845 317.045 -153.515 ;
        RECT 316.715 -155.205 317.045 -154.875 ;
        RECT 316.715 -156.565 317.045 -156.235 ;
        RECT 316.715 -157.925 317.045 -157.595 ;
        RECT 316.715 -159.285 317.045 -158.955 ;
        RECT 316.715 -160.645 317.045 -160.315 ;
        RECT 316.715 -162.005 317.045 -161.675 ;
        RECT 316.715 -163.365 317.045 -163.035 ;
        RECT 316.715 -164.725 317.045 -164.395 ;
        RECT 316.715 -166.085 317.045 -165.755 ;
        RECT 316.715 -167.445 317.045 -167.115 ;
        RECT 316.715 -168.805 317.045 -168.475 ;
        RECT 316.715 -170.165 317.045 -169.835 ;
        RECT 316.715 -171.525 317.045 -171.195 ;
        RECT 316.715 -172.885 317.045 -172.555 ;
        RECT 316.715 -174.245 317.045 -173.915 ;
        RECT 316.715 -175.605 317.045 -175.275 ;
        RECT 316.715 -176.965 317.045 -176.635 ;
        RECT 316.715 -178.325 317.045 -177.995 ;
        RECT 316.715 -179.685 317.045 -179.355 ;
        RECT 316.715 -181.045 317.045 -180.715 ;
        RECT 316.715 -182.405 317.045 -182.075 ;
        RECT 316.715 -183.765 317.045 -183.435 ;
        RECT 316.715 -185.125 317.045 -184.795 ;
        RECT 316.715 -186.485 317.045 -186.155 ;
        RECT 316.715 -187.845 317.045 -187.515 ;
        RECT 316.715 -189.205 317.045 -188.875 ;
        RECT 316.715 -190.565 317.045 -190.235 ;
        RECT 316.715 -191.925 317.045 -191.595 ;
        RECT 316.715 -193.285 317.045 -192.955 ;
        RECT 316.715 -194.645 317.045 -194.315 ;
        RECT 316.715 -196.005 317.045 -195.675 ;
        RECT 316.715 -197.365 317.045 -197.035 ;
        RECT 316.715 -198.725 317.045 -198.395 ;
        RECT 316.715 -200.085 317.045 -199.755 ;
        RECT 316.715 -201.445 317.045 -201.115 ;
        RECT 316.715 -202.805 317.045 -202.475 ;
        RECT 316.715 -204.165 317.045 -203.835 ;
        RECT 316.715 -205.525 317.045 -205.195 ;
        RECT 316.715 -206.885 317.045 -206.555 ;
        RECT 316.715 -208.245 317.045 -207.915 ;
        RECT 316.715 -209.605 317.045 -209.275 ;
        RECT 316.715 -210.965 317.045 -210.635 ;
        RECT 316.715 -212.325 317.045 -211.995 ;
        RECT 316.715 -213.685 317.045 -213.355 ;
        RECT 316.715 -215.045 317.045 -214.715 ;
        RECT 316.715 -216.405 317.045 -216.075 ;
        RECT 316.715 -217.765 317.045 -217.435 ;
        RECT 316.715 -219.125 317.045 -218.795 ;
        RECT 316.715 -220.485 317.045 -220.155 ;
        RECT 316.715 -221.845 317.045 -221.515 ;
        RECT 316.715 -223.205 317.045 -222.875 ;
        RECT 316.715 -224.565 317.045 -224.235 ;
        RECT 316.715 -225.925 317.045 -225.595 ;
        RECT 316.715 -227.285 317.045 -226.955 ;
        RECT 316.715 -228.645 317.045 -228.315 ;
        RECT 316.715 -230.005 317.045 -229.675 ;
        RECT 316.715 -231.365 317.045 -231.035 ;
        RECT 316.715 -232.725 317.045 -232.395 ;
        RECT 316.715 -234.085 317.045 -233.755 ;
        RECT 316.715 -235.445 317.045 -235.115 ;
        RECT 316.715 -236.805 317.045 -236.475 ;
        RECT 316.715 -238.165 317.045 -237.835 ;
        RECT 316.715 -243.81 317.045 -242.68 ;
        RECT 316.72 -243.925 317.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 246.76 318.405 247.89 ;
        RECT 318.075 241.915 318.405 242.245 ;
        RECT 318.075 240.555 318.405 240.885 ;
        RECT 318.075 239.195 318.405 239.525 ;
        RECT 318.075 237.835 318.405 238.165 ;
        RECT 318.08 237.16 318.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 -1.525 318.405 -1.195 ;
        RECT 318.075 -2.885 318.405 -2.555 ;
        RECT 318.08 -3.56 318.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 -122.565 318.405 -122.235 ;
        RECT 318.075 -123.925 318.405 -123.595 ;
        RECT 318.075 -125.285 318.405 -124.955 ;
        RECT 318.075 -126.645 318.405 -126.315 ;
        RECT 318.075 -128.005 318.405 -127.675 ;
        RECT 318.075 -129.365 318.405 -129.035 ;
        RECT 318.075 -130.725 318.405 -130.395 ;
        RECT 318.075 -132.085 318.405 -131.755 ;
        RECT 318.075 -133.445 318.405 -133.115 ;
        RECT 318.075 -134.805 318.405 -134.475 ;
        RECT 318.075 -136.165 318.405 -135.835 ;
        RECT 318.075 -137.525 318.405 -137.195 ;
        RECT 318.075 -138.885 318.405 -138.555 ;
        RECT 318.075 -140.245 318.405 -139.915 ;
        RECT 318.075 -141.605 318.405 -141.275 ;
        RECT 318.075 -142.965 318.405 -142.635 ;
        RECT 318.075 -144.325 318.405 -143.995 ;
        RECT 318.075 -145.685 318.405 -145.355 ;
        RECT 318.075 -147.045 318.405 -146.715 ;
        RECT 318.075 -148.405 318.405 -148.075 ;
        RECT 318.075 -149.765 318.405 -149.435 ;
        RECT 318.075 -151.125 318.405 -150.795 ;
        RECT 318.075 -152.485 318.405 -152.155 ;
        RECT 318.075 -153.845 318.405 -153.515 ;
        RECT 318.075 -155.205 318.405 -154.875 ;
        RECT 318.075 -156.565 318.405 -156.235 ;
        RECT 318.075 -157.925 318.405 -157.595 ;
        RECT 318.075 -159.285 318.405 -158.955 ;
        RECT 318.075 -160.645 318.405 -160.315 ;
        RECT 318.075 -162.005 318.405 -161.675 ;
        RECT 318.075 -163.365 318.405 -163.035 ;
        RECT 318.075 -164.725 318.405 -164.395 ;
        RECT 318.075 -166.085 318.405 -165.755 ;
        RECT 318.075 -167.445 318.405 -167.115 ;
        RECT 318.075 -168.805 318.405 -168.475 ;
        RECT 318.075 -170.165 318.405 -169.835 ;
        RECT 318.075 -171.525 318.405 -171.195 ;
        RECT 318.075 -172.885 318.405 -172.555 ;
        RECT 318.075 -174.245 318.405 -173.915 ;
        RECT 318.075 -175.605 318.405 -175.275 ;
        RECT 318.075 -176.965 318.405 -176.635 ;
        RECT 318.075 -178.325 318.405 -177.995 ;
        RECT 318.075 -179.685 318.405 -179.355 ;
        RECT 318.075 -181.045 318.405 -180.715 ;
        RECT 318.075 -182.405 318.405 -182.075 ;
        RECT 318.075 -183.765 318.405 -183.435 ;
        RECT 318.075 -185.125 318.405 -184.795 ;
        RECT 318.075 -186.485 318.405 -186.155 ;
        RECT 318.075 -187.845 318.405 -187.515 ;
        RECT 318.075 -189.205 318.405 -188.875 ;
        RECT 318.075 -190.565 318.405 -190.235 ;
        RECT 318.075 -191.925 318.405 -191.595 ;
        RECT 318.075 -193.285 318.405 -192.955 ;
        RECT 318.075 -194.645 318.405 -194.315 ;
        RECT 318.075 -196.005 318.405 -195.675 ;
        RECT 318.075 -197.365 318.405 -197.035 ;
        RECT 318.075 -198.725 318.405 -198.395 ;
        RECT 318.075 -200.085 318.405 -199.755 ;
        RECT 318.075 -201.445 318.405 -201.115 ;
        RECT 318.075 -202.805 318.405 -202.475 ;
        RECT 318.075 -204.165 318.405 -203.835 ;
        RECT 318.075 -205.525 318.405 -205.195 ;
        RECT 318.075 -206.885 318.405 -206.555 ;
        RECT 318.075 -208.245 318.405 -207.915 ;
        RECT 318.075 -209.605 318.405 -209.275 ;
        RECT 318.075 -210.965 318.405 -210.635 ;
        RECT 318.075 -212.325 318.405 -211.995 ;
        RECT 318.075 -213.685 318.405 -213.355 ;
        RECT 318.075 -215.045 318.405 -214.715 ;
        RECT 318.075 -216.405 318.405 -216.075 ;
        RECT 318.075 -217.765 318.405 -217.435 ;
        RECT 318.075 -219.125 318.405 -218.795 ;
        RECT 318.075 -220.485 318.405 -220.155 ;
        RECT 318.075 -221.845 318.405 -221.515 ;
        RECT 318.075 -223.205 318.405 -222.875 ;
        RECT 318.075 -224.565 318.405 -224.235 ;
        RECT 318.075 -225.925 318.405 -225.595 ;
        RECT 318.075 -227.285 318.405 -226.955 ;
        RECT 318.075 -228.645 318.405 -228.315 ;
        RECT 318.075 -230.005 318.405 -229.675 ;
        RECT 318.075 -231.365 318.405 -231.035 ;
        RECT 318.075 -232.725 318.405 -232.395 ;
        RECT 318.075 -234.085 318.405 -233.755 ;
        RECT 318.075 -235.445 318.405 -235.115 ;
        RECT 318.075 -236.805 318.405 -236.475 ;
        RECT 318.075 -238.165 318.405 -237.835 ;
        RECT 318.075 -243.81 318.405 -242.68 ;
        RECT 318.08 -243.925 318.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.76 -125.535 319.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.435 246.76 319.765 247.89 ;
        RECT 319.435 241.915 319.765 242.245 ;
        RECT 319.435 240.555 319.765 240.885 ;
        RECT 319.435 239.195 319.765 239.525 ;
        RECT 319.435 237.835 319.765 238.165 ;
        RECT 319.44 237.16 319.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.795 246.76 321.125 247.89 ;
        RECT 320.795 241.915 321.125 242.245 ;
        RECT 320.795 240.555 321.125 240.885 ;
        RECT 320.795 239.195 321.125 239.525 ;
        RECT 320.795 237.835 321.125 238.165 ;
        RECT 320.8 237.16 321.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.795 -1.525 321.125 -1.195 ;
        RECT 320.795 -2.885 321.125 -2.555 ;
        RECT 320.8 -3.56 321.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 246.76 322.485 247.89 ;
        RECT 322.155 241.915 322.485 242.245 ;
        RECT 322.155 240.555 322.485 240.885 ;
        RECT 322.155 239.195 322.485 239.525 ;
        RECT 322.155 237.835 322.485 238.165 ;
        RECT 322.16 237.16 322.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 -2.885 322.485 -2.555 ;
        RECT 322.16 -3.56 322.48 -0.52 ;
        RECT 322.155 -1.525 322.485 -1.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 246.76 283.045 247.89 ;
        RECT 282.715 241.915 283.045 242.245 ;
        RECT 282.715 240.555 283.045 240.885 ;
        RECT 282.715 239.195 283.045 239.525 ;
        RECT 282.715 237.835 283.045 238.165 ;
        RECT 282.72 237.16 283.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 -1.525 283.045 -1.195 ;
        RECT 282.715 -2.885 283.045 -2.555 ;
        RECT 282.72 -3.56 283.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 -122.565 283.045 -122.235 ;
        RECT 282.715 -123.925 283.045 -123.595 ;
        RECT 282.715 -125.285 283.045 -124.955 ;
        RECT 282.715 -126.645 283.045 -126.315 ;
        RECT 282.715 -128.005 283.045 -127.675 ;
        RECT 282.715 -129.365 283.045 -129.035 ;
        RECT 282.715 -130.725 283.045 -130.395 ;
        RECT 282.715 -132.085 283.045 -131.755 ;
        RECT 282.715 -133.445 283.045 -133.115 ;
        RECT 282.715 -134.805 283.045 -134.475 ;
        RECT 282.715 -136.165 283.045 -135.835 ;
        RECT 282.715 -137.525 283.045 -137.195 ;
        RECT 282.715 -138.885 283.045 -138.555 ;
        RECT 282.715 -140.245 283.045 -139.915 ;
        RECT 282.715 -141.605 283.045 -141.275 ;
        RECT 282.715 -142.965 283.045 -142.635 ;
        RECT 282.715 -144.325 283.045 -143.995 ;
        RECT 282.715 -145.685 283.045 -145.355 ;
        RECT 282.715 -147.045 283.045 -146.715 ;
        RECT 282.715 -148.405 283.045 -148.075 ;
        RECT 282.715 -149.765 283.045 -149.435 ;
        RECT 282.715 -151.125 283.045 -150.795 ;
        RECT 282.715 -152.485 283.045 -152.155 ;
        RECT 282.715 -153.845 283.045 -153.515 ;
        RECT 282.715 -155.205 283.045 -154.875 ;
        RECT 282.715 -156.565 283.045 -156.235 ;
        RECT 282.715 -157.925 283.045 -157.595 ;
        RECT 282.715 -159.285 283.045 -158.955 ;
        RECT 282.715 -160.645 283.045 -160.315 ;
        RECT 282.715 -162.005 283.045 -161.675 ;
        RECT 282.715 -163.365 283.045 -163.035 ;
        RECT 282.715 -164.725 283.045 -164.395 ;
        RECT 282.715 -166.085 283.045 -165.755 ;
        RECT 282.715 -167.445 283.045 -167.115 ;
        RECT 282.715 -168.805 283.045 -168.475 ;
        RECT 282.715 -170.165 283.045 -169.835 ;
        RECT 282.715 -171.525 283.045 -171.195 ;
        RECT 282.715 -172.885 283.045 -172.555 ;
        RECT 282.715 -174.245 283.045 -173.915 ;
        RECT 282.715 -175.605 283.045 -175.275 ;
        RECT 282.715 -176.965 283.045 -176.635 ;
        RECT 282.715 -178.325 283.045 -177.995 ;
        RECT 282.715 -179.685 283.045 -179.355 ;
        RECT 282.715 -181.045 283.045 -180.715 ;
        RECT 282.715 -182.405 283.045 -182.075 ;
        RECT 282.715 -183.765 283.045 -183.435 ;
        RECT 282.715 -185.125 283.045 -184.795 ;
        RECT 282.715 -186.485 283.045 -186.155 ;
        RECT 282.715 -187.845 283.045 -187.515 ;
        RECT 282.715 -189.205 283.045 -188.875 ;
        RECT 282.715 -190.565 283.045 -190.235 ;
        RECT 282.715 -191.925 283.045 -191.595 ;
        RECT 282.715 -193.285 283.045 -192.955 ;
        RECT 282.715 -194.645 283.045 -194.315 ;
        RECT 282.715 -196.005 283.045 -195.675 ;
        RECT 282.715 -197.365 283.045 -197.035 ;
        RECT 282.715 -198.725 283.045 -198.395 ;
        RECT 282.715 -200.085 283.045 -199.755 ;
        RECT 282.715 -201.445 283.045 -201.115 ;
        RECT 282.715 -202.805 283.045 -202.475 ;
        RECT 282.715 -204.165 283.045 -203.835 ;
        RECT 282.715 -205.525 283.045 -205.195 ;
        RECT 282.715 -206.885 283.045 -206.555 ;
        RECT 282.715 -208.245 283.045 -207.915 ;
        RECT 282.715 -209.605 283.045 -209.275 ;
        RECT 282.715 -210.965 283.045 -210.635 ;
        RECT 282.715 -212.325 283.045 -211.995 ;
        RECT 282.715 -213.685 283.045 -213.355 ;
        RECT 282.715 -215.045 283.045 -214.715 ;
        RECT 282.715 -216.405 283.045 -216.075 ;
        RECT 282.715 -217.765 283.045 -217.435 ;
        RECT 282.715 -219.125 283.045 -218.795 ;
        RECT 282.715 -220.485 283.045 -220.155 ;
        RECT 282.715 -221.845 283.045 -221.515 ;
        RECT 282.715 -223.205 283.045 -222.875 ;
        RECT 282.715 -224.565 283.045 -224.235 ;
        RECT 282.715 -225.925 283.045 -225.595 ;
        RECT 282.715 -227.285 283.045 -226.955 ;
        RECT 282.715 -228.645 283.045 -228.315 ;
        RECT 282.715 -230.005 283.045 -229.675 ;
        RECT 282.715 -231.365 283.045 -231.035 ;
        RECT 282.715 -232.725 283.045 -232.395 ;
        RECT 282.715 -234.085 283.045 -233.755 ;
        RECT 282.715 -235.445 283.045 -235.115 ;
        RECT 282.715 -236.805 283.045 -236.475 ;
        RECT 282.715 -238.165 283.045 -237.835 ;
        RECT 282.715 -243.81 283.045 -242.68 ;
        RECT 282.72 -243.925 283.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 246.76 284.405 247.89 ;
        RECT 284.075 241.915 284.405 242.245 ;
        RECT 284.075 240.555 284.405 240.885 ;
        RECT 284.075 239.195 284.405 239.525 ;
        RECT 284.075 237.835 284.405 238.165 ;
        RECT 284.08 237.16 284.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 -1.525 284.405 -1.195 ;
        RECT 284.075 -2.885 284.405 -2.555 ;
        RECT 284.08 -3.56 284.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 -122.565 284.405 -122.235 ;
        RECT 284.075 -123.925 284.405 -123.595 ;
        RECT 284.075 -125.285 284.405 -124.955 ;
        RECT 284.075 -126.645 284.405 -126.315 ;
        RECT 284.075 -128.005 284.405 -127.675 ;
        RECT 284.075 -129.365 284.405 -129.035 ;
        RECT 284.075 -130.725 284.405 -130.395 ;
        RECT 284.075 -132.085 284.405 -131.755 ;
        RECT 284.075 -133.445 284.405 -133.115 ;
        RECT 284.075 -134.805 284.405 -134.475 ;
        RECT 284.075 -136.165 284.405 -135.835 ;
        RECT 284.075 -137.525 284.405 -137.195 ;
        RECT 284.075 -138.885 284.405 -138.555 ;
        RECT 284.075 -140.245 284.405 -139.915 ;
        RECT 284.075 -141.605 284.405 -141.275 ;
        RECT 284.075 -142.965 284.405 -142.635 ;
        RECT 284.075 -144.325 284.405 -143.995 ;
        RECT 284.075 -145.685 284.405 -145.355 ;
        RECT 284.075 -147.045 284.405 -146.715 ;
        RECT 284.075 -148.405 284.405 -148.075 ;
        RECT 284.075 -149.765 284.405 -149.435 ;
        RECT 284.075 -151.125 284.405 -150.795 ;
        RECT 284.075 -152.485 284.405 -152.155 ;
        RECT 284.075 -153.845 284.405 -153.515 ;
        RECT 284.075 -155.205 284.405 -154.875 ;
        RECT 284.075 -156.565 284.405 -156.235 ;
        RECT 284.075 -157.925 284.405 -157.595 ;
        RECT 284.075 -159.285 284.405 -158.955 ;
        RECT 284.075 -160.645 284.405 -160.315 ;
        RECT 284.075 -162.005 284.405 -161.675 ;
        RECT 284.075 -163.365 284.405 -163.035 ;
        RECT 284.075 -164.725 284.405 -164.395 ;
        RECT 284.075 -166.085 284.405 -165.755 ;
        RECT 284.075 -167.445 284.405 -167.115 ;
        RECT 284.075 -168.805 284.405 -168.475 ;
        RECT 284.075 -170.165 284.405 -169.835 ;
        RECT 284.075 -171.525 284.405 -171.195 ;
        RECT 284.075 -172.885 284.405 -172.555 ;
        RECT 284.075 -174.245 284.405 -173.915 ;
        RECT 284.075 -175.605 284.405 -175.275 ;
        RECT 284.075 -176.965 284.405 -176.635 ;
        RECT 284.075 -178.325 284.405 -177.995 ;
        RECT 284.075 -179.685 284.405 -179.355 ;
        RECT 284.075 -181.045 284.405 -180.715 ;
        RECT 284.075 -182.405 284.405 -182.075 ;
        RECT 284.075 -183.765 284.405 -183.435 ;
        RECT 284.075 -185.125 284.405 -184.795 ;
        RECT 284.075 -186.485 284.405 -186.155 ;
        RECT 284.075 -187.845 284.405 -187.515 ;
        RECT 284.075 -189.205 284.405 -188.875 ;
        RECT 284.075 -190.565 284.405 -190.235 ;
        RECT 284.075 -191.925 284.405 -191.595 ;
        RECT 284.075 -193.285 284.405 -192.955 ;
        RECT 284.075 -194.645 284.405 -194.315 ;
        RECT 284.075 -196.005 284.405 -195.675 ;
        RECT 284.075 -197.365 284.405 -197.035 ;
        RECT 284.075 -198.725 284.405 -198.395 ;
        RECT 284.075 -200.085 284.405 -199.755 ;
        RECT 284.075 -201.445 284.405 -201.115 ;
        RECT 284.075 -202.805 284.405 -202.475 ;
        RECT 284.075 -204.165 284.405 -203.835 ;
        RECT 284.075 -205.525 284.405 -205.195 ;
        RECT 284.075 -206.885 284.405 -206.555 ;
        RECT 284.075 -208.245 284.405 -207.915 ;
        RECT 284.075 -209.605 284.405 -209.275 ;
        RECT 284.075 -210.965 284.405 -210.635 ;
        RECT 284.075 -212.325 284.405 -211.995 ;
        RECT 284.075 -213.685 284.405 -213.355 ;
        RECT 284.075 -215.045 284.405 -214.715 ;
        RECT 284.075 -216.405 284.405 -216.075 ;
        RECT 284.075 -217.765 284.405 -217.435 ;
        RECT 284.075 -219.125 284.405 -218.795 ;
        RECT 284.075 -220.485 284.405 -220.155 ;
        RECT 284.075 -221.845 284.405 -221.515 ;
        RECT 284.075 -223.205 284.405 -222.875 ;
        RECT 284.075 -224.565 284.405 -224.235 ;
        RECT 284.075 -225.925 284.405 -225.595 ;
        RECT 284.075 -227.285 284.405 -226.955 ;
        RECT 284.075 -228.645 284.405 -228.315 ;
        RECT 284.075 -230.005 284.405 -229.675 ;
        RECT 284.075 -231.365 284.405 -231.035 ;
        RECT 284.075 -232.725 284.405 -232.395 ;
        RECT 284.075 -234.085 284.405 -233.755 ;
        RECT 284.075 -235.445 284.405 -235.115 ;
        RECT 284.075 -236.805 284.405 -236.475 ;
        RECT 284.075 -238.165 284.405 -237.835 ;
        RECT 284.075 -243.81 284.405 -242.68 ;
        RECT 284.08 -243.925 284.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 246.76 285.765 247.89 ;
        RECT 285.435 241.915 285.765 242.245 ;
        RECT 285.435 240.555 285.765 240.885 ;
        RECT 285.435 239.195 285.765 239.525 ;
        RECT 285.435 237.835 285.765 238.165 ;
        RECT 285.44 237.16 285.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 -126.645 285.765 -126.315 ;
        RECT 285.435 -128.005 285.765 -127.675 ;
        RECT 285.435 -129.365 285.765 -129.035 ;
        RECT 285.435 -130.725 285.765 -130.395 ;
        RECT 285.435 -132.085 285.765 -131.755 ;
        RECT 285.435 -133.445 285.765 -133.115 ;
        RECT 285.435 -134.805 285.765 -134.475 ;
        RECT 285.435 -136.165 285.765 -135.835 ;
        RECT 285.435 -137.525 285.765 -137.195 ;
        RECT 285.435 -138.885 285.765 -138.555 ;
        RECT 285.435 -140.245 285.765 -139.915 ;
        RECT 285.435 -141.605 285.765 -141.275 ;
        RECT 285.435 -142.965 285.765 -142.635 ;
        RECT 285.435 -144.325 285.765 -143.995 ;
        RECT 285.435 -145.685 285.765 -145.355 ;
        RECT 285.435 -147.045 285.765 -146.715 ;
        RECT 285.435 -148.405 285.765 -148.075 ;
        RECT 285.435 -149.765 285.765 -149.435 ;
        RECT 285.435 -151.125 285.765 -150.795 ;
        RECT 285.435 -152.485 285.765 -152.155 ;
        RECT 285.435 -153.845 285.765 -153.515 ;
        RECT 285.435 -155.205 285.765 -154.875 ;
        RECT 285.435 -156.565 285.765 -156.235 ;
        RECT 285.435 -157.925 285.765 -157.595 ;
        RECT 285.435 -159.285 285.765 -158.955 ;
        RECT 285.435 -160.645 285.765 -160.315 ;
        RECT 285.435 -162.005 285.765 -161.675 ;
        RECT 285.435 -163.365 285.765 -163.035 ;
        RECT 285.435 -164.725 285.765 -164.395 ;
        RECT 285.435 -166.085 285.765 -165.755 ;
        RECT 285.435 -167.445 285.765 -167.115 ;
        RECT 285.435 -168.805 285.765 -168.475 ;
        RECT 285.435 -170.165 285.765 -169.835 ;
        RECT 285.435 -171.525 285.765 -171.195 ;
        RECT 285.435 -172.885 285.765 -172.555 ;
        RECT 285.435 -174.245 285.765 -173.915 ;
        RECT 285.435 -175.605 285.765 -175.275 ;
        RECT 285.435 -176.965 285.765 -176.635 ;
        RECT 285.435 -178.325 285.765 -177.995 ;
        RECT 285.435 -179.685 285.765 -179.355 ;
        RECT 285.435 -181.045 285.765 -180.715 ;
        RECT 285.435 -182.405 285.765 -182.075 ;
        RECT 285.435 -183.765 285.765 -183.435 ;
        RECT 285.435 -185.125 285.765 -184.795 ;
        RECT 285.435 -186.485 285.765 -186.155 ;
        RECT 285.435 -187.845 285.765 -187.515 ;
        RECT 285.435 -189.205 285.765 -188.875 ;
        RECT 285.435 -190.565 285.765 -190.235 ;
        RECT 285.435 -191.925 285.765 -191.595 ;
        RECT 285.435 -193.285 285.765 -192.955 ;
        RECT 285.435 -194.645 285.765 -194.315 ;
        RECT 285.435 -196.005 285.765 -195.675 ;
        RECT 285.435 -197.365 285.765 -197.035 ;
        RECT 285.435 -198.725 285.765 -198.395 ;
        RECT 285.435 -200.085 285.765 -199.755 ;
        RECT 285.435 -201.445 285.765 -201.115 ;
        RECT 285.435 -202.805 285.765 -202.475 ;
        RECT 285.435 -204.165 285.765 -203.835 ;
        RECT 285.435 -205.525 285.765 -205.195 ;
        RECT 285.435 -206.885 285.765 -206.555 ;
        RECT 285.435 -208.245 285.765 -207.915 ;
        RECT 285.435 -209.605 285.765 -209.275 ;
        RECT 285.435 -210.965 285.765 -210.635 ;
        RECT 285.435 -212.325 285.765 -211.995 ;
        RECT 285.435 -213.685 285.765 -213.355 ;
        RECT 285.435 -215.045 285.765 -214.715 ;
        RECT 285.435 -216.405 285.765 -216.075 ;
        RECT 285.435 -217.765 285.765 -217.435 ;
        RECT 285.435 -219.125 285.765 -218.795 ;
        RECT 285.435 -220.485 285.765 -220.155 ;
        RECT 285.435 -221.845 285.765 -221.515 ;
        RECT 285.435 -223.205 285.765 -222.875 ;
        RECT 285.435 -224.565 285.765 -224.235 ;
        RECT 285.435 -225.925 285.765 -225.595 ;
        RECT 285.435 -227.285 285.765 -226.955 ;
        RECT 285.435 -228.645 285.765 -228.315 ;
        RECT 285.435 -230.005 285.765 -229.675 ;
        RECT 285.435 -231.365 285.765 -231.035 ;
        RECT 285.435 -232.725 285.765 -232.395 ;
        RECT 285.435 -234.085 285.765 -233.755 ;
        RECT 285.435 -235.445 285.765 -235.115 ;
        RECT 285.435 -236.805 285.765 -236.475 ;
        RECT 285.435 -238.165 285.765 -237.835 ;
        RECT 285.435 -243.81 285.765 -242.68 ;
        RECT 285.44 -243.925 285.76 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.06 -125.535 286.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.795 246.76 287.125 247.89 ;
        RECT 286.795 241.915 287.125 242.245 ;
        RECT 286.795 240.555 287.125 240.885 ;
        RECT 286.795 239.195 287.125 239.525 ;
        RECT 286.795 237.835 287.125 238.165 ;
        RECT 286.8 237.16 287.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 246.76 288.485 247.89 ;
        RECT 288.155 241.915 288.485 242.245 ;
        RECT 288.155 240.555 288.485 240.885 ;
        RECT 288.155 239.195 288.485 239.525 ;
        RECT 288.155 237.835 288.485 238.165 ;
        RECT 288.16 237.16 288.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 -1.525 288.485 -1.195 ;
        RECT 288.155 -2.885 288.485 -2.555 ;
        RECT 288.16 -3.56 288.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 -122.565 288.485 -122.235 ;
        RECT 288.155 -123.925 288.485 -123.595 ;
        RECT 288.155 -125.285 288.485 -124.955 ;
        RECT 288.155 -126.645 288.485 -126.315 ;
        RECT 288.155 -128.005 288.485 -127.675 ;
        RECT 288.155 -129.365 288.485 -129.035 ;
        RECT 288.155 -130.725 288.485 -130.395 ;
        RECT 288.155 -132.085 288.485 -131.755 ;
        RECT 288.155 -133.445 288.485 -133.115 ;
        RECT 288.155 -134.805 288.485 -134.475 ;
        RECT 288.155 -136.165 288.485 -135.835 ;
        RECT 288.155 -137.525 288.485 -137.195 ;
        RECT 288.155 -138.885 288.485 -138.555 ;
        RECT 288.155 -140.245 288.485 -139.915 ;
        RECT 288.155 -141.605 288.485 -141.275 ;
        RECT 288.155 -142.965 288.485 -142.635 ;
        RECT 288.155 -144.325 288.485 -143.995 ;
        RECT 288.155 -145.685 288.485 -145.355 ;
        RECT 288.155 -147.045 288.485 -146.715 ;
        RECT 288.155 -148.405 288.485 -148.075 ;
        RECT 288.155 -149.765 288.485 -149.435 ;
        RECT 288.155 -151.125 288.485 -150.795 ;
        RECT 288.155 -152.485 288.485 -152.155 ;
        RECT 288.155 -153.845 288.485 -153.515 ;
        RECT 288.155 -155.205 288.485 -154.875 ;
        RECT 288.155 -156.565 288.485 -156.235 ;
        RECT 288.155 -157.925 288.485 -157.595 ;
        RECT 288.155 -159.285 288.485 -158.955 ;
        RECT 288.155 -160.645 288.485 -160.315 ;
        RECT 288.155 -162.005 288.485 -161.675 ;
        RECT 288.155 -163.365 288.485 -163.035 ;
        RECT 288.155 -164.725 288.485 -164.395 ;
        RECT 288.155 -166.085 288.485 -165.755 ;
        RECT 288.155 -167.445 288.485 -167.115 ;
        RECT 288.155 -168.805 288.485 -168.475 ;
        RECT 288.155 -170.165 288.485 -169.835 ;
        RECT 288.155 -171.525 288.485 -171.195 ;
        RECT 288.155 -172.885 288.485 -172.555 ;
        RECT 288.155 -174.245 288.485 -173.915 ;
        RECT 288.155 -175.605 288.485 -175.275 ;
        RECT 288.155 -176.965 288.485 -176.635 ;
        RECT 288.155 -178.325 288.485 -177.995 ;
        RECT 288.155 -179.685 288.485 -179.355 ;
        RECT 288.155 -181.045 288.485 -180.715 ;
        RECT 288.155 -182.405 288.485 -182.075 ;
        RECT 288.155 -183.765 288.485 -183.435 ;
        RECT 288.155 -185.125 288.485 -184.795 ;
        RECT 288.155 -186.485 288.485 -186.155 ;
        RECT 288.155 -187.845 288.485 -187.515 ;
        RECT 288.155 -189.205 288.485 -188.875 ;
        RECT 288.155 -190.565 288.485 -190.235 ;
        RECT 288.155 -191.925 288.485 -191.595 ;
        RECT 288.155 -193.285 288.485 -192.955 ;
        RECT 288.155 -194.645 288.485 -194.315 ;
        RECT 288.155 -196.005 288.485 -195.675 ;
        RECT 288.155 -197.365 288.485 -197.035 ;
        RECT 288.155 -198.725 288.485 -198.395 ;
        RECT 288.155 -200.085 288.485 -199.755 ;
        RECT 288.155 -201.445 288.485 -201.115 ;
        RECT 288.155 -202.805 288.485 -202.475 ;
        RECT 288.155 -204.165 288.485 -203.835 ;
        RECT 288.155 -205.525 288.485 -205.195 ;
        RECT 288.155 -206.885 288.485 -206.555 ;
        RECT 288.155 -208.245 288.485 -207.915 ;
        RECT 288.155 -209.605 288.485 -209.275 ;
        RECT 288.155 -210.965 288.485 -210.635 ;
        RECT 288.155 -212.325 288.485 -211.995 ;
        RECT 288.155 -213.685 288.485 -213.355 ;
        RECT 288.155 -215.045 288.485 -214.715 ;
        RECT 288.155 -216.405 288.485 -216.075 ;
        RECT 288.155 -217.765 288.485 -217.435 ;
        RECT 288.155 -219.125 288.485 -218.795 ;
        RECT 288.155 -220.485 288.485 -220.155 ;
        RECT 288.155 -221.845 288.485 -221.515 ;
        RECT 288.155 -223.205 288.485 -222.875 ;
        RECT 288.155 -224.565 288.485 -224.235 ;
        RECT 288.155 -225.925 288.485 -225.595 ;
        RECT 288.155 -227.285 288.485 -226.955 ;
        RECT 288.155 -228.645 288.485 -228.315 ;
        RECT 288.155 -230.005 288.485 -229.675 ;
        RECT 288.155 -231.365 288.485 -231.035 ;
        RECT 288.155 -232.725 288.485 -232.395 ;
        RECT 288.155 -234.085 288.485 -233.755 ;
        RECT 288.155 -235.445 288.485 -235.115 ;
        RECT 288.155 -236.805 288.485 -236.475 ;
        RECT 288.155 -238.165 288.485 -237.835 ;
        RECT 288.155 -243.81 288.485 -242.68 ;
        RECT 288.16 -243.925 288.48 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 246.76 289.845 247.89 ;
        RECT 289.515 241.915 289.845 242.245 ;
        RECT 289.515 240.555 289.845 240.885 ;
        RECT 289.515 239.195 289.845 239.525 ;
        RECT 289.515 237.835 289.845 238.165 ;
        RECT 289.52 237.16 289.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 -1.525 289.845 -1.195 ;
        RECT 289.515 -2.885 289.845 -2.555 ;
        RECT 289.52 -3.56 289.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 246.76 291.205 247.89 ;
        RECT 290.875 241.915 291.205 242.245 ;
        RECT 290.875 240.555 291.205 240.885 ;
        RECT 290.875 239.195 291.205 239.525 ;
        RECT 290.875 237.835 291.205 238.165 ;
        RECT 290.88 237.16 291.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 -1.525 291.205 -1.195 ;
        RECT 290.875 -2.885 291.205 -2.555 ;
        RECT 290.88 -3.56 291.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 -122.565 291.205 -122.235 ;
        RECT 290.875 -123.925 291.205 -123.595 ;
        RECT 290.875 -125.285 291.205 -124.955 ;
        RECT 290.875 -126.645 291.205 -126.315 ;
        RECT 290.875 -128.005 291.205 -127.675 ;
        RECT 290.875 -129.365 291.205 -129.035 ;
        RECT 290.875 -130.725 291.205 -130.395 ;
        RECT 290.875 -132.085 291.205 -131.755 ;
        RECT 290.875 -133.445 291.205 -133.115 ;
        RECT 290.875 -134.805 291.205 -134.475 ;
        RECT 290.875 -136.165 291.205 -135.835 ;
        RECT 290.875 -137.525 291.205 -137.195 ;
        RECT 290.875 -138.885 291.205 -138.555 ;
        RECT 290.875 -140.245 291.205 -139.915 ;
        RECT 290.875 -141.605 291.205 -141.275 ;
        RECT 290.875 -142.965 291.205 -142.635 ;
        RECT 290.875 -144.325 291.205 -143.995 ;
        RECT 290.875 -145.685 291.205 -145.355 ;
        RECT 290.875 -147.045 291.205 -146.715 ;
        RECT 290.875 -148.405 291.205 -148.075 ;
        RECT 290.875 -149.765 291.205 -149.435 ;
        RECT 290.875 -151.125 291.205 -150.795 ;
        RECT 290.875 -152.485 291.205 -152.155 ;
        RECT 290.875 -153.845 291.205 -153.515 ;
        RECT 290.875 -155.205 291.205 -154.875 ;
        RECT 290.875 -156.565 291.205 -156.235 ;
        RECT 290.875 -157.925 291.205 -157.595 ;
        RECT 290.875 -159.285 291.205 -158.955 ;
        RECT 290.875 -160.645 291.205 -160.315 ;
        RECT 290.875 -162.005 291.205 -161.675 ;
        RECT 290.875 -163.365 291.205 -163.035 ;
        RECT 290.875 -164.725 291.205 -164.395 ;
        RECT 290.875 -166.085 291.205 -165.755 ;
        RECT 290.875 -167.445 291.205 -167.115 ;
        RECT 290.875 -168.805 291.205 -168.475 ;
        RECT 290.875 -170.165 291.205 -169.835 ;
        RECT 290.875 -171.525 291.205 -171.195 ;
        RECT 290.875 -172.885 291.205 -172.555 ;
        RECT 290.875 -174.245 291.205 -173.915 ;
        RECT 290.875 -175.605 291.205 -175.275 ;
        RECT 290.875 -176.965 291.205 -176.635 ;
        RECT 290.875 -178.325 291.205 -177.995 ;
        RECT 290.875 -179.685 291.205 -179.355 ;
        RECT 290.875 -181.045 291.205 -180.715 ;
        RECT 290.875 -182.405 291.205 -182.075 ;
        RECT 290.875 -183.765 291.205 -183.435 ;
        RECT 290.875 -185.125 291.205 -184.795 ;
        RECT 290.875 -186.485 291.205 -186.155 ;
        RECT 290.875 -187.845 291.205 -187.515 ;
        RECT 290.875 -189.205 291.205 -188.875 ;
        RECT 290.875 -190.565 291.205 -190.235 ;
        RECT 290.875 -191.925 291.205 -191.595 ;
        RECT 290.875 -193.285 291.205 -192.955 ;
        RECT 290.875 -194.645 291.205 -194.315 ;
        RECT 290.875 -196.005 291.205 -195.675 ;
        RECT 290.875 -197.365 291.205 -197.035 ;
        RECT 290.875 -198.725 291.205 -198.395 ;
        RECT 290.875 -200.085 291.205 -199.755 ;
        RECT 290.875 -201.445 291.205 -201.115 ;
        RECT 290.875 -202.805 291.205 -202.475 ;
        RECT 290.875 -204.165 291.205 -203.835 ;
        RECT 290.875 -205.525 291.205 -205.195 ;
        RECT 290.875 -206.885 291.205 -206.555 ;
        RECT 290.875 -208.245 291.205 -207.915 ;
        RECT 290.875 -209.605 291.205 -209.275 ;
        RECT 290.875 -210.965 291.205 -210.635 ;
        RECT 290.875 -212.325 291.205 -211.995 ;
        RECT 290.875 -213.685 291.205 -213.355 ;
        RECT 290.875 -215.045 291.205 -214.715 ;
        RECT 290.875 -216.405 291.205 -216.075 ;
        RECT 290.875 -217.765 291.205 -217.435 ;
        RECT 290.875 -219.125 291.205 -218.795 ;
        RECT 290.875 -220.485 291.205 -220.155 ;
        RECT 290.875 -221.845 291.205 -221.515 ;
        RECT 290.875 -223.205 291.205 -222.875 ;
        RECT 290.875 -224.565 291.205 -224.235 ;
        RECT 290.875 -225.925 291.205 -225.595 ;
        RECT 290.875 -227.285 291.205 -226.955 ;
        RECT 290.875 -228.645 291.205 -228.315 ;
        RECT 290.875 -230.005 291.205 -229.675 ;
        RECT 290.875 -231.365 291.205 -231.035 ;
        RECT 290.875 -232.725 291.205 -232.395 ;
        RECT 290.875 -234.085 291.205 -233.755 ;
        RECT 290.875 -235.445 291.205 -235.115 ;
        RECT 290.875 -236.805 291.205 -236.475 ;
        RECT 290.875 -238.165 291.205 -237.835 ;
        RECT 290.875 -243.81 291.205 -242.68 ;
        RECT 290.88 -243.925 291.2 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 246.76 292.565 247.89 ;
        RECT 292.235 241.915 292.565 242.245 ;
        RECT 292.235 240.555 292.565 240.885 ;
        RECT 292.235 239.195 292.565 239.525 ;
        RECT 292.235 237.835 292.565 238.165 ;
        RECT 292.24 237.16 292.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 -1.525 292.565 -1.195 ;
        RECT 292.235 -2.885 292.565 -2.555 ;
        RECT 292.24 -3.56 292.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 -122.565 292.565 -122.235 ;
        RECT 292.235 -123.925 292.565 -123.595 ;
        RECT 292.235 -125.285 292.565 -124.955 ;
        RECT 292.235 -126.645 292.565 -126.315 ;
        RECT 292.235 -128.005 292.565 -127.675 ;
        RECT 292.235 -129.365 292.565 -129.035 ;
        RECT 292.235 -130.725 292.565 -130.395 ;
        RECT 292.235 -132.085 292.565 -131.755 ;
        RECT 292.235 -133.445 292.565 -133.115 ;
        RECT 292.235 -134.805 292.565 -134.475 ;
        RECT 292.235 -136.165 292.565 -135.835 ;
        RECT 292.235 -137.525 292.565 -137.195 ;
        RECT 292.235 -138.885 292.565 -138.555 ;
        RECT 292.235 -140.245 292.565 -139.915 ;
        RECT 292.235 -141.605 292.565 -141.275 ;
        RECT 292.235 -142.965 292.565 -142.635 ;
        RECT 292.235 -144.325 292.565 -143.995 ;
        RECT 292.235 -145.685 292.565 -145.355 ;
        RECT 292.235 -147.045 292.565 -146.715 ;
        RECT 292.235 -148.405 292.565 -148.075 ;
        RECT 292.235 -149.765 292.565 -149.435 ;
        RECT 292.235 -151.125 292.565 -150.795 ;
        RECT 292.235 -152.485 292.565 -152.155 ;
        RECT 292.235 -153.845 292.565 -153.515 ;
        RECT 292.235 -155.205 292.565 -154.875 ;
        RECT 292.235 -156.565 292.565 -156.235 ;
        RECT 292.235 -157.925 292.565 -157.595 ;
        RECT 292.235 -159.285 292.565 -158.955 ;
        RECT 292.235 -160.645 292.565 -160.315 ;
        RECT 292.235 -162.005 292.565 -161.675 ;
        RECT 292.235 -163.365 292.565 -163.035 ;
        RECT 292.235 -164.725 292.565 -164.395 ;
        RECT 292.235 -166.085 292.565 -165.755 ;
        RECT 292.235 -167.445 292.565 -167.115 ;
        RECT 292.235 -168.805 292.565 -168.475 ;
        RECT 292.235 -170.165 292.565 -169.835 ;
        RECT 292.235 -171.525 292.565 -171.195 ;
        RECT 292.235 -172.885 292.565 -172.555 ;
        RECT 292.235 -174.245 292.565 -173.915 ;
        RECT 292.235 -175.605 292.565 -175.275 ;
        RECT 292.235 -176.965 292.565 -176.635 ;
        RECT 292.235 -178.325 292.565 -177.995 ;
        RECT 292.235 -179.685 292.565 -179.355 ;
        RECT 292.235 -181.045 292.565 -180.715 ;
        RECT 292.235 -182.405 292.565 -182.075 ;
        RECT 292.235 -183.765 292.565 -183.435 ;
        RECT 292.235 -185.125 292.565 -184.795 ;
        RECT 292.235 -186.485 292.565 -186.155 ;
        RECT 292.235 -187.845 292.565 -187.515 ;
        RECT 292.235 -189.205 292.565 -188.875 ;
        RECT 292.235 -190.565 292.565 -190.235 ;
        RECT 292.235 -191.925 292.565 -191.595 ;
        RECT 292.235 -193.285 292.565 -192.955 ;
        RECT 292.235 -194.645 292.565 -194.315 ;
        RECT 292.235 -196.005 292.565 -195.675 ;
        RECT 292.235 -197.365 292.565 -197.035 ;
        RECT 292.235 -198.725 292.565 -198.395 ;
        RECT 292.235 -200.085 292.565 -199.755 ;
        RECT 292.235 -201.445 292.565 -201.115 ;
        RECT 292.235 -202.805 292.565 -202.475 ;
        RECT 292.235 -204.165 292.565 -203.835 ;
        RECT 292.235 -205.525 292.565 -205.195 ;
        RECT 292.235 -206.885 292.565 -206.555 ;
        RECT 292.235 -208.245 292.565 -207.915 ;
        RECT 292.235 -209.605 292.565 -209.275 ;
        RECT 292.235 -210.965 292.565 -210.635 ;
        RECT 292.235 -212.325 292.565 -211.995 ;
        RECT 292.235 -213.685 292.565 -213.355 ;
        RECT 292.235 -215.045 292.565 -214.715 ;
        RECT 292.235 -216.405 292.565 -216.075 ;
        RECT 292.235 -217.765 292.565 -217.435 ;
        RECT 292.235 -219.125 292.565 -218.795 ;
        RECT 292.235 -220.485 292.565 -220.155 ;
        RECT 292.235 -221.845 292.565 -221.515 ;
        RECT 292.235 -223.205 292.565 -222.875 ;
        RECT 292.235 -224.565 292.565 -224.235 ;
        RECT 292.235 -225.925 292.565 -225.595 ;
        RECT 292.235 -227.285 292.565 -226.955 ;
        RECT 292.235 -228.645 292.565 -228.315 ;
        RECT 292.235 -230.005 292.565 -229.675 ;
        RECT 292.235 -231.365 292.565 -231.035 ;
        RECT 292.235 -232.725 292.565 -232.395 ;
        RECT 292.235 -234.085 292.565 -233.755 ;
        RECT 292.235 -235.445 292.565 -235.115 ;
        RECT 292.235 -236.805 292.565 -236.475 ;
        RECT 292.235 -238.165 292.565 -237.835 ;
        RECT 292.235 -243.81 292.565 -242.68 ;
        RECT 292.24 -243.925 292.56 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 246.76 293.925 247.89 ;
        RECT 293.595 241.915 293.925 242.245 ;
        RECT 293.595 240.555 293.925 240.885 ;
        RECT 293.595 239.195 293.925 239.525 ;
        RECT 293.595 237.835 293.925 238.165 ;
        RECT 293.6 237.16 293.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 -1.525 293.925 -1.195 ;
        RECT 293.595 -2.885 293.925 -2.555 ;
        RECT 293.6 -3.56 293.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 -122.565 293.925 -122.235 ;
        RECT 293.595 -123.925 293.925 -123.595 ;
        RECT 293.595 -125.285 293.925 -124.955 ;
        RECT 293.595 -126.645 293.925 -126.315 ;
        RECT 293.595 -128.005 293.925 -127.675 ;
        RECT 293.595 -129.365 293.925 -129.035 ;
        RECT 293.595 -130.725 293.925 -130.395 ;
        RECT 293.595 -132.085 293.925 -131.755 ;
        RECT 293.595 -133.445 293.925 -133.115 ;
        RECT 293.595 -134.805 293.925 -134.475 ;
        RECT 293.595 -136.165 293.925 -135.835 ;
        RECT 293.595 -137.525 293.925 -137.195 ;
        RECT 293.595 -138.885 293.925 -138.555 ;
        RECT 293.595 -140.245 293.925 -139.915 ;
        RECT 293.595 -141.605 293.925 -141.275 ;
        RECT 293.595 -142.965 293.925 -142.635 ;
        RECT 293.595 -144.325 293.925 -143.995 ;
        RECT 293.595 -145.685 293.925 -145.355 ;
        RECT 293.595 -147.045 293.925 -146.715 ;
        RECT 293.595 -148.405 293.925 -148.075 ;
        RECT 293.595 -149.765 293.925 -149.435 ;
        RECT 293.595 -151.125 293.925 -150.795 ;
        RECT 293.595 -152.485 293.925 -152.155 ;
        RECT 293.595 -153.845 293.925 -153.515 ;
        RECT 293.595 -155.205 293.925 -154.875 ;
        RECT 293.595 -156.565 293.925 -156.235 ;
        RECT 293.595 -157.925 293.925 -157.595 ;
        RECT 293.595 -159.285 293.925 -158.955 ;
        RECT 293.595 -160.645 293.925 -160.315 ;
        RECT 293.595 -162.005 293.925 -161.675 ;
        RECT 293.595 -163.365 293.925 -163.035 ;
        RECT 293.595 -164.725 293.925 -164.395 ;
        RECT 293.595 -166.085 293.925 -165.755 ;
        RECT 293.595 -167.445 293.925 -167.115 ;
        RECT 293.595 -168.805 293.925 -168.475 ;
        RECT 293.595 -170.165 293.925 -169.835 ;
        RECT 293.595 -171.525 293.925 -171.195 ;
        RECT 293.595 -172.885 293.925 -172.555 ;
        RECT 293.595 -174.245 293.925 -173.915 ;
        RECT 293.595 -175.605 293.925 -175.275 ;
        RECT 293.595 -176.965 293.925 -176.635 ;
        RECT 293.595 -178.325 293.925 -177.995 ;
        RECT 293.595 -179.685 293.925 -179.355 ;
        RECT 293.595 -181.045 293.925 -180.715 ;
        RECT 293.595 -182.405 293.925 -182.075 ;
        RECT 293.595 -183.765 293.925 -183.435 ;
        RECT 293.595 -185.125 293.925 -184.795 ;
        RECT 293.595 -186.485 293.925 -186.155 ;
        RECT 293.595 -187.845 293.925 -187.515 ;
        RECT 293.595 -189.205 293.925 -188.875 ;
        RECT 293.595 -190.565 293.925 -190.235 ;
        RECT 293.595 -191.925 293.925 -191.595 ;
        RECT 293.595 -193.285 293.925 -192.955 ;
        RECT 293.595 -194.645 293.925 -194.315 ;
        RECT 293.595 -196.005 293.925 -195.675 ;
        RECT 293.595 -197.365 293.925 -197.035 ;
        RECT 293.595 -198.725 293.925 -198.395 ;
        RECT 293.595 -200.085 293.925 -199.755 ;
        RECT 293.595 -201.445 293.925 -201.115 ;
        RECT 293.595 -202.805 293.925 -202.475 ;
        RECT 293.595 -204.165 293.925 -203.835 ;
        RECT 293.595 -205.525 293.925 -205.195 ;
        RECT 293.595 -206.885 293.925 -206.555 ;
        RECT 293.595 -208.245 293.925 -207.915 ;
        RECT 293.595 -209.605 293.925 -209.275 ;
        RECT 293.595 -210.965 293.925 -210.635 ;
        RECT 293.595 -212.325 293.925 -211.995 ;
        RECT 293.595 -213.685 293.925 -213.355 ;
        RECT 293.595 -215.045 293.925 -214.715 ;
        RECT 293.595 -216.405 293.925 -216.075 ;
        RECT 293.595 -217.765 293.925 -217.435 ;
        RECT 293.595 -219.125 293.925 -218.795 ;
        RECT 293.595 -220.485 293.925 -220.155 ;
        RECT 293.595 -221.845 293.925 -221.515 ;
        RECT 293.595 -223.205 293.925 -222.875 ;
        RECT 293.595 -224.565 293.925 -224.235 ;
        RECT 293.595 -225.925 293.925 -225.595 ;
        RECT 293.595 -227.285 293.925 -226.955 ;
        RECT 293.595 -228.645 293.925 -228.315 ;
        RECT 293.595 -230.005 293.925 -229.675 ;
        RECT 293.595 -231.365 293.925 -231.035 ;
        RECT 293.595 -232.725 293.925 -232.395 ;
        RECT 293.595 -234.085 293.925 -233.755 ;
        RECT 293.595 -235.445 293.925 -235.115 ;
        RECT 293.595 -236.805 293.925 -236.475 ;
        RECT 293.595 -238.165 293.925 -237.835 ;
        RECT 293.595 -243.81 293.925 -242.68 ;
        RECT 293.6 -243.925 293.92 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 246.76 295.285 247.89 ;
        RECT 294.955 241.915 295.285 242.245 ;
        RECT 294.955 240.555 295.285 240.885 ;
        RECT 294.955 239.195 295.285 239.525 ;
        RECT 294.955 237.835 295.285 238.165 ;
        RECT 294.96 237.16 295.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 -1.525 295.285 -1.195 ;
        RECT 294.955 -2.885 295.285 -2.555 ;
        RECT 294.96 -3.56 295.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 -122.565 295.285 -122.235 ;
        RECT 294.955 -123.925 295.285 -123.595 ;
        RECT 294.955 -125.285 295.285 -124.955 ;
        RECT 294.955 -126.645 295.285 -126.315 ;
        RECT 294.955 -128.005 295.285 -127.675 ;
        RECT 294.955 -129.365 295.285 -129.035 ;
        RECT 294.955 -130.725 295.285 -130.395 ;
        RECT 294.955 -132.085 295.285 -131.755 ;
        RECT 294.955 -133.445 295.285 -133.115 ;
        RECT 294.955 -134.805 295.285 -134.475 ;
        RECT 294.955 -136.165 295.285 -135.835 ;
        RECT 294.955 -137.525 295.285 -137.195 ;
        RECT 294.955 -138.885 295.285 -138.555 ;
        RECT 294.955 -140.245 295.285 -139.915 ;
        RECT 294.955 -141.605 295.285 -141.275 ;
        RECT 294.955 -142.965 295.285 -142.635 ;
        RECT 294.955 -144.325 295.285 -143.995 ;
        RECT 294.955 -145.685 295.285 -145.355 ;
        RECT 294.955 -147.045 295.285 -146.715 ;
        RECT 294.955 -148.405 295.285 -148.075 ;
        RECT 294.955 -149.765 295.285 -149.435 ;
        RECT 294.955 -151.125 295.285 -150.795 ;
        RECT 294.955 -152.485 295.285 -152.155 ;
        RECT 294.955 -153.845 295.285 -153.515 ;
        RECT 294.955 -155.205 295.285 -154.875 ;
        RECT 294.955 -156.565 295.285 -156.235 ;
        RECT 294.955 -157.925 295.285 -157.595 ;
        RECT 294.955 -159.285 295.285 -158.955 ;
        RECT 294.955 -160.645 295.285 -160.315 ;
        RECT 294.955 -162.005 295.285 -161.675 ;
        RECT 294.955 -163.365 295.285 -163.035 ;
        RECT 294.955 -164.725 295.285 -164.395 ;
        RECT 294.955 -166.085 295.285 -165.755 ;
        RECT 294.955 -167.445 295.285 -167.115 ;
        RECT 294.955 -168.805 295.285 -168.475 ;
        RECT 294.955 -170.165 295.285 -169.835 ;
        RECT 294.955 -171.525 295.285 -171.195 ;
        RECT 294.955 -172.885 295.285 -172.555 ;
        RECT 294.955 -174.245 295.285 -173.915 ;
        RECT 294.955 -175.605 295.285 -175.275 ;
        RECT 294.955 -176.965 295.285 -176.635 ;
        RECT 294.955 -178.325 295.285 -177.995 ;
        RECT 294.955 -179.685 295.285 -179.355 ;
        RECT 294.955 -181.045 295.285 -180.715 ;
        RECT 294.955 -182.405 295.285 -182.075 ;
        RECT 294.955 -183.765 295.285 -183.435 ;
        RECT 294.955 -185.125 295.285 -184.795 ;
        RECT 294.955 -186.485 295.285 -186.155 ;
        RECT 294.955 -187.845 295.285 -187.515 ;
        RECT 294.955 -189.205 295.285 -188.875 ;
        RECT 294.955 -190.565 295.285 -190.235 ;
        RECT 294.955 -191.925 295.285 -191.595 ;
        RECT 294.955 -193.285 295.285 -192.955 ;
        RECT 294.955 -194.645 295.285 -194.315 ;
        RECT 294.955 -196.005 295.285 -195.675 ;
        RECT 294.955 -197.365 295.285 -197.035 ;
        RECT 294.955 -198.725 295.285 -198.395 ;
        RECT 294.955 -200.085 295.285 -199.755 ;
        RECT 294.955 -201.445 295.285 -201.115 ;
        RECT 294.955 -202.805 295.285 -202.475 ;
        RECT 294.955 -204.165 295.285 -203.835 ;
        RECT 294.955 -205.525 295.285 -205.195 ;
        RECT 294.955 -206.885 295.285 -206.555 ;
        RECT 294.955 -208.245 295.285 -207.915 ;
        RECT 294.955 -209.605 295.285 -209.275 ;
        RECT 294.955 -210.965 295.285 -210.635 ;
        RECT 294.955 -212.325 295.285 -211.995 ;
        RECT 294.955 -213.685 295.285 -213.355 ;
        RECT 294.955 -215.045 295.285 -214.715 ;
        RECT 294.955 -216.405 295.285 -216.075 ;
        RECT 294.955 -217.765 295.285 -217.435 ;
        RECT 294.955 -219.125 295.285 -218.795 ;
        RECT 294.955 -220.485 295.285 -220.155 ;
        RECT 294.955 -221.845 295.285 -221.515 ;
        RECT 294.955 -223.205 295.285 -222.875 ;
        RECT 294.955 -224.565 295.285 -224.235 ;
        RECT 294.955 -225.925 295.285 -225.595 ;
        RECT 294.955 -227.285 295.285 -226.955 ;
        RECT 294.955 -228.645 295.285 -228.315 ;
        RECT 294.955 -230.005 295.285 -229.675 ;
        RECT 294.955 -231.365 295.285 -231.035 ;
        RECT 294.955 -232.725 295.285 -232.395 ;
        RECT 294.955 -234.085 295.285 -233.755 ;
        RECT 294.955 -235.445 295.285 -235.115 ;
        RECT 294.955 -236.805 295.285 -236.475 ;
        RECT 294.955 -238.165 295.285 -237.835 ;
        RECT 294.955 -243.81 295.285 -242.68 ;
        RECT 294.96 -243.925 295.28 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.315 246.76 296.645 247.89 ;
        RECT 296.315 241.915 296.645 242.245 ;
        RECT 296.315 240.555 296.645 240.885 ;
        RECT 296.315 239.195 296.645 239.525 ;
        RECT 296.315 237.835 296.645 238.165 ;
        RECT 296.32 237.16 296.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.315 -126.645 296.645 -126.315 ;
        RECT 296.315 -128.005 296.645 -127.675 ;
        RECT 296.315 -129.365 296.645 -129.035 ;
        RECT 296.315 -130.725 296.645 -130.395 ;
        RECT 296.315 -132.085 296.645 -131.755 ;
        RECT 296.315 -133.445 296.645 -133.115 ;
        RECT 296.315 -134.805 296.645 -134.475 ;
        RECT 296.315 -136.165 296.645 -135.835 ;
        RECT 296.315 -137.525 296.645 -137.195 ;
        RECT 296.315 -138.885 296.645 -138.555 ;
        RECT 296.315 -140.245 296.645 -139.915 ;
        RECT 296.315 -141.605 296.645 -141.275 ;
        RECT 296.315 -142.965 296.645 -142.635 ;
        RECT 296.315 -144.325 296.645 -143.995 ;
        RECT 296.315 -145.685 296.645 -145.355 ;
        RECT 296.315 -147.045 296.645 -146.715 ;
        RECT 296.315 -148.405 296.645 -148.075 ;
        RECT 296.315 -149.765 296.645 -149.435 ;
        RECT 296.315 -151.125 296.645 -150.795 ;
        RECT 296.315 -152.485 296.645 -152.155 ;
        RECT 296.315 -153.845 296.645 -153.515 ;
        RECT 296.315 -155.205 296.645 -154.875 ;
        RECT 296.315 -156.565 296.645 -156.235 ;
        RECT 296.315 -157.925 296.645 -157.595 ;
        RECT 296.315 -159.285 296.645 -158.955 ;
        RECT 296.315 -160.645 296.645 -160.315 ;
        RECT 296.315 -162.005 296.645 -161.675 ;
        RECT 296.315 -163.365 296.645 -163.035 ;
        RECT 296.315 -164.725 296.645 -164.395 ;
        RECT 296.315 -166.085 296.645 -165.755 ;
        RECT 296.315 -167.445 296.645 -167.115 ;
        RECT 296.315 -168.805 296.645 -168.475 ;
        RECT 296.315 -170.165 296.645 -169.835 ;
        RECT 296.315 -171.525 296.645 -171.195 ;
        RECT 296.315 -172.885 296.645 -172.555 ;
        RECT 296.315 -174.245 296.645 -173.915 ;
        RECT 296.315 -175.605 296.645 -175.275 ;
        RECT 296.315 -176.965 296.645 -176.635 ;
        RECT 296.315 -178.325 296.645 -177.995 ;
        RECT 296.315 -179.685 296.645 -179.355 ;
        RECT 296.315 -181.045 296.645 -180.715 ;
        RECT 296.315 -182.405 296.645 -182.075 ;
        RECT 296.315 -183.765 296.645 -183.435 ;
        RECT 296.315 -185.125 296.645 -184.795 ;
        RECT 296.315 -186.485 296.645 -186.155 ;
        RECT 296.315 -187.845 296.645 -187.515 ;
        RECT 296.315 -189.205 296.645 -188.875 ;
        RECT 296.315 -190.565 296.645 -190.235 ;
        RECT 296.315 -191.925 296.645 -191.595 ;
        RECT 296.315 -193.285 296.645 -192.955 ;
        RECT 296.315 -194.645 296.645 -194.315 ;
        RECT 296.315 -196.005 296.645 -195.675 ;
        RECT 296.315 -197.365 296.645 -197.035 ;
        RECT 296.315 -198.725 296.645 -198.395 ;
        RECT 296.315 -200.085 296.645 -199.755 ;
        RECT 296.315 -201.445 296.645 -201.115 ;
        RECT 296.315 -202.805 296.645 -202.475 ;
        RECT 296.315 -204.165 296.645 -203.835 ;
        RECT 296.315 -205.525 296.645 -205.195 ;
        RECT 296.315 -206.885 296.645 -206.555 ;
        RECT 296.315 -208.245 296.645 -207.915 ;
        RECT 296.315 -209.605 296.645 -209.275 ;
        RECT 296.315 -210.965 296.645 -210.635 ;
        RECT 296.315 -212.325 296.645 -211.995 ;
        RECT 296.315 -213.685 296.645 -213.355 ;
        RECT 296.315 -215.045 296.645 -214.715 ;
        RECT 296.315 -216.405 296.645 -216.075 ;
        RECT 296.315 -217.765 296.645 -217.435 ;
        RECT 296.315 -219.125 296.645 -218.795 ;
        RECT 296.315 -220.485 296.645 -220.155 ;
        RECT 296.315 -221.845 296.645 -221.515 ;
        RECT 296.315 -223.205 296.645 -222.875 ;
        RECT 296.315 -224.565 296.645 -224.235 ;
        RECT 296.315 -225.925 296.645 -225.595 ;
        RECT 296.315 -227.285 296.645 -226.955 ;
        RECT 296.315 -228.645 296.645 -228.315 ;
        RECT 296.315 -230.005 296.645 -229.675 ;
        RECT 296.315 -231.365 296.645 -231.035 ;
        RECT 296.315 -232.725 296.645 -232.395 ;
        RECT 296.315 -234.085 296.645 -233.755 ;
        RECT 296.315 -235.445 296.645 -235.115 ;
        RECT 296.315 -236.805 296.645 -236.475 ;
        RECT 296.315 -238.165 296.645 -237.835 ;
        RECT 296.315 -243.81 296.645 -242.68 ;
        RECT 296.32 -243.925 296.64 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.96 -125.535 297.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.675 246.76 298.005 247.89 ;
        RECT 297.675 241.915 298.005 242.245 ;
        RECT 297.675 240.555 298.005 240.885 ;
        RECT 297.675 239.195 298.005 239.525 ;
        RECT 297.675 237.835 298.005 238.165 ;
        RECT 297.68 237.16 298 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 246.76 299.365 247.89 ;
        RECT 299.035 241.915 299.365 242.245 ;
        RECT 299.035 240.555 299.365 240.885 ;
        RECT 299.035 239.195 299.365 239.525 ;
        RECT 299.035 237.835 299.365 238.165 ;
        RECT 299.04 237.16 299.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 -1.525 299.365 -1.195 ;
        RECT 299.035 -2.885 299.365 -2.555 ;
        RECT 299.04 -3.56 299.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 246.76 300.725 247.89 ;
        RECT 300.395 241.915 300.725 242.245 ;
        RECT 300.395 240.555 300.725 240.885 ;
        RECT 300.395 239.195 300.725 239.525 ;
        RECT 300.395 237.835 300.725 238.165 ;
        RECT 300.4 237.16 300.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 -1.525 300.725 -1.195 ;
        RECT 300.395 -2.885 300.725 -2.555 ;
        RECT 300.4 -3.56 300.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 246.76 302.085 247.89 ;
        RECT 301.755 241.915 302.085 242.245 ;
        RECT 301.755 240.555 302.085 240.885 ;
        RECT 301.755 239.195 302.085 239.525 ;
        RECT 301.755 237.835 302.085 238.165 ;
        RECT 301.76 237.16 302.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 -1.525 302.085 -1.195 ;
        RECT 301.755 -2.885 302.085 -2.555 ;
        RECT 301.76 -3.56 302.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 -236.805 302.085 -236.475 ;
        RECT 301.755 -238.165 302.085 -237.835 ;
        RECT 301.755 -243.81 302.085 -242.68 ;
        RECT 301.76 -243.925 302.08 -122.235 ;
        RECT 301.755 -122.565 302.085 -122.235 ;
        RECT 301.755 -123.925 302.085 -123.595 ;
        RECT 301.755 -125.285 302.085 -124.955 ;
        RECT 301.755 -126.645 302.085 -126.315 ;
        RECT 301.755 -128.005 302.085 -127.675 ;
        RECT 301.755 -129.365 302.085 -129.035 ;
        RECT 301.755 -130.725 302.085 -130.395 ;
        RECT 301.755 -132.085 302.085 -131.755 ;
        RECT 301.755 -133.445 302.085 -133.115 ;
        RECT 301.755 -134.805 302.085 -134.475 ;
        RECT 301.755 -136.165 302.085 -135.835 ;
        RECT 301.755 -137.525 302.085 -137.195 ;
        RECT 301.755 -138.885 302.085 -138.555 ;
        RECT 301.755 -140.245 302.085 -139.915 ;
        RECT 301.755 -141.605 302.085 -141.275 ;
        RECT 301.755 -142.965 302.085 -142.635 ;
        RECT 301.755 -144.325 302.085 -143.995 ;
        RECT 301.755 -145.685 302.085 -145.355 ;
        RECT 301.755 -147.045 302.085 -146.715 ;
        RECT 301.755 -148.405 302.085 -148.075 ;
        RECT 301.755 -149.765 302.085 -149.435 ;
        RECT 301.755 -151.125 302.085 -150.795 ;
        RECT 301.755 -152.485 302.085 -152.155 ;
        RECT 301.755 -153.845 302.085 -153.515 ;
        RECT 301.755 -155.205 302.085 -154.875 ;
        RECT 301.755 -156.565 302.085 -156.235 ;
        RECT 301.755 -157.925 302.085 -157.595 ;
        RECT 301.755 -159.285 302.085 -158.955 ;
        RECT 301.755 -160.645 302.085 -160.315 ;
        RECT 301.755 -162.005 302.085 -161.675 ;
        RECT 301.755 -163.365 302.085 -163.035 ;
        RECT 301.755 -164.725 302.085 -164.395 ;
        RECT 301.755 -166.085 302.085 -165.755 ;
        RECT 301.755 -167.445 302.085 -167.115 ;
        RECT 301.755 -168.805 302.085 -168.475 ;
        RECT 301.755 -170.165 302.085 -169.835 ;
        RECT 301.755 -171.525 302.085 -171.195 ;
        RECT 301.755 -172.885 302.085 -172.555 ;
        RECT 301.755 -174.245 302.085 -173.915 ;
        RECT 301.755 -175.605 302.085 -175.275 ;
        RECT 301.755 -176.965 302.085 -176.635 ;
        RECT 301.755 -178.325 302.085 -177.995 ;
        RECT 301.755 -179.685 302.085 -179.355 ;
        RECT 301.755 -181.045 302.085 -180.715 ;
        RECT 301.755 -182.405 302.085 -182.075 ;
        RECT 301.755 -183.765 302.085 -183.435 ;
        RECT 301.755 -185.125 302.085 -184.795 ;
        RECT 301.755 -186.485 302.085 -186.155 ;
        RECT 301.755 -187.845 302.085 -187.515 ;
        RECT 301.755 -189.205 302.085 -188.875 ;
        RECT 301.755 -190.565 302.085 -190.235 ;
        RECT 301.755 -191.925 302.085 -191.595 ;
        RECT 301.755 -193.285 302.085 -192.955 ;
        RECT 301.755 -194.645 302.085 -194.315 ;
        RECT 301.755 -196.005 302.085 -195.675 ;
        RECT 301.755 -197.365 302.085 -197.035 ;
        RECT 301.755 -198.725 302.085 -198.395 ;
        RECT 301.755 -200.085 302.085 -199.755 ;
        RECT 301.755 -201.445 302.085 -201.115 ;
        RECT 301.755 -202.805 302.085 -202.475 ;
        RECT 301.755 -204.165 302.085 -203.835 ;
        RECT 301.755 -205.525 302.085 -205.195 ;
        RECT 301.755 -206.885 302.085 -206.555 ;
        RECT 301.755 -208.245 302.085 -207.915 ;
        RECT 301.755 -209.605 302.085 -209.275 ;
        RECT 301.755 -210.965 302.085 -210.635 ;
        RECT 301.755 -212.325 302.085 -211.995 ;
        RECT 301.755 -213.685 302.085 -213.355 ;
        RECT 301.755 -215.045 302.085 -214.715 ;
        RECT 301.755 -216.405 302.085 -216.075 ;
        RECT 301.755 -217.765 302.085 -217.435 ;
        RECT 301.755 -219.125 302.085 -218.795 ;
        RECT 301.755 -220.485 302.085 -220.155 ;
        RECT 301.755 -221.845 302.085 -221.515 ;
        RECT 301.755 -223.205 302.085 -222.875 ;
        RECT 301.755 -224.565 302.085 -224.235 ;
        RECT 301.755 -225.925 302.085 -225.595 ;
        RECT 301.755 -227.285 302.085 -226.955 ;
        RECT 301.755 -228.645 302.085 -228.315 ;
        RECT 301.755 -230.005 302.085 -229.675 ;
        RECT 301.755 -231.365 302.085 -231.035 ;
        RECT 301.755 -232.725 302.085 -232.395 ;
        RECT 301.755 -234.085 302.085 -233.755 ;
        RECT 301.755 -235.445 302.085 -235.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 -1.525 262.645 -1.195 ;
        RECT 262.315 -2.885 262.645 -2.555 ;
        RECT 262.32 -3.56 262.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 -122.565 262.645 -122.235 ;
        RECT 262.315 -123.925 262.645 -123.595 ;
        RECT 262.315 -125.285 262.645 -124.955 ;
        RECT 262.315 -126.645 262.645 -126.315 ;
        RECT 262.315 -128.005 262.645 -127.675 ;
        RECT 262.315 -129.365 262.645 -129.035 ;
        RECT 262.315 -130.725 262.645 -130.395 ;
        RECT 262.315 -132.085 262.645 -131.755 ;
        RECT 262.315 -133.445 262.645 -133.115 ;
        RECT 262.315 -134.805 262.645 -134.475 ;
        RECT 262.315 -136.165 262.645 -135.835 ;
        RECT 262.315 -137.525 262.645 -137.195 ;
        RECT 262.315 -138.885 262.645 -138.555 ;
        RECT 262.315 -140.245 262.645 -139.915 ;
        RECT 262.315 -141.605 262.645 -141.275 ;
        RECT 262.315 -142.965 262.645 -142.635 ;
        RECT 262.315 -144.325 262.645 -143.995 ;
        RECT 262.315 -145.685 262.645 -145.355 ;
        RECT 262.315 -147.045 262.645 -146.715 ;
        RECT 262.315 -148.405 262.645 -148.075 ;
        RECT 262.315 -149.765 262.645 -149.435 ;
        RECT 262.315 -151.125 262.645 -150.795 ;
        RECT 262.315 -152.485 262.645 -152.155 ;
        RECT 262.315 -153.845 262.645 -153.515 ;
        RECT 262.315 -155.205 262.645 -154.875 ;
        RECT 262.315 -156.565 262.645 -156.235 ;
        RECT 262.315 -157.925 262.645 -157.595 ;
        RECT 262.315 -159.285 262.645 -158.955 ;
        RECT 262.315 -160.645 262.645 -160.315 ;
        RECT 262.315 -162.005 262.645 -161.675 ;
        RECT 262.315 -163.365 262.645 -163.035 ;
        RECT 262.315 -164.725 262.645 -164.395 ;
        RECT 262.315 -166.085 262.645 -165.755 ;
        RECT 262.315 -167.445 262.645 -167.115 ;
        RECT 262.315 -168.805 262.645 -168.475 ;
        RECT 262.315 -170.165 262.645 -169.835 ;
        RECT 262.315 -171.525 262.645 -171.195 ;
        RECT 262.315 -172.885 262.645 -172.555 ;
        RECT 262.315 -174.245 262.645 -173.915 ;
        RECT 262.315 -175.605 262.645 -175.275 ;
        RECT 262.315 -176.965 262.645 -176.635 ;
        RECT 262.315 -178.325 262.645 -177.995 ;
        RECT 262.315 -179.685 262.645 -179.355 ;
        RECT 262.315 -181.045 262.645 -180.715 ;
        RECT 262.315 -182.405 262.645 -182.075 ;
        RECT 262.315 -183.765 262.645 -183.435 ;
        RECT 262.315 -185.125 262.645 -184.795 ;
        RECT 262.315 -186.485 262.645 -186.155 ;
        RECT 262.315 -187.845 262.645 -187.515 ;
        RECT 262.315 -189.205 262.645 -188.875 ;
        RECT 262.315 -190.565 262.645 -190.235 ;
        RECT 262.315 -191.925 262.645 -191.595 ;
        RECT 262.315 -193.285 262.645 -192.955 ;
        RECT 262.315 -194.645 262.645 -194.315 ;
        RECT 262.315 -196.005 262.645 -195.675 ;
        RECT 262.315 -197.365 262.645 -197.035 ;
        RECT 262.315 -198.725 262.645 -198.395 ;
        RECT 262.315 -200.085 262.645 -199.755 ;
        RECT 262.315 -201.445 262.645 -201.115 ;
        RECT 262.315 -202.805 262.645 -202.475 ;
        RECT 262.315 -204.165 262.645 -203.835 ;
        RECT 262.315 -205.525 262.645 -205.195 ;
        RECT 262.315 -206.885 262.645 -206.555 ;
        RECT 262.315 -208.245 262.645 -207.915 ;
        RECT 262.315 -209.605 262.645 -209.275 ;
        RECT 262.315 -210.965 262.645 -210.635 ;
        RECT 262.315 -212.325 262.645 -211.995 ;
        RECT 262.315 -213.685 262.645 -213.355 ;
        RECT 262.315 -215.045 262.645 -214.715 ;
        RECT 262.315 -216.405 262.645 -216.075 ;
        RECT 262.315 -217.765 262.645 -217.435 ;
        RECT 262.315 -219.125 262.645 -218.795 ;
        RECT 262.315 -220.485 262.645 -220.155 ;
        RECT 262.315 -221.845 262.645 -221.515 ;
        RECT 262.315 -223.205 262.645 -222.875 ;
        RECT 262.315 -224.565 262.645 -224.235 ;
        RECT 262.315 -225.925 262.645 -225.595 ;
        RECT 262.315 -227.285 262.645 -226.955 ;
        RECT 262.315 -228.645 262.645 -228.315 ;
        RECT 262.315 -230.005 262.645 -229.675 ;
        RECT 262.315 -231.365 262.645 -231.035 ;
        RECT 262.315 -232.725 262.645 -232.395 ;
        RECT 262.315 -234.085 262.645 -233.755 ;
        RECT 262.315 -235.445 262.645 -235.115 ;
        RECT 262.315 -236.805 262.645 -236.475 ;
        RECT 262.315 -238.165 262.645 -237.835 ;
        RECT 262.315 -243.81 262.645 -242.68 ;
        RECT 262.32 -243.925 262.64 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 246.76 264.005 247.89 ;
        RECT 263.675 241.915 264.005 242.245 ;
        RECT 263.675 240.555 264.005 240.885 ;
        RECT 263.675 239.195 264.005 239.525 ;
        RECT 263.675 237.835 264.005 238.165 ;
        RECT 263.68 237.16 264 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 -126.645 264.005 -126.315 ;
        RECT 263.675 -128.005 264.005 -127.675 ;
        RECT 263.675 -129.365 264.005 -129.035 ;
        RECT 263.675 -130.725 264.005 -130.395 ;
        RECT 263.675 -132.085 264.005 -131.755 ;
        RECT 263.675 -133.445 264.005 -133.115 ;
        RECT 263.675 -134.805 264.005 -134.475 ;
        RECT 263.675 -136.165 264.005 -135.835 ;
        RECT 263.675 -137.525 264.005 -137.195 ;
        RECT 263.675 -138.885 264.005 -138.555 ;
        RECT 263.675 -140.245 264.005 -139.915 ;
        RECT 263.675 -141.605 264.005 -141.275 ;
        RECT 263.675 -142.965 264.005 -142.635 ;
        RECT 263.675 -144.325 264.005 -143.995 ;
        RECT 263.675 -145.685 264.005 -145.355 ;
        RECT 263.675 -147.045 264.005 -146.715 ;
        RECT 263.675 -148.405 264.005 -148.075 ;
        RECT 263.675 -149.765 264.005 -149.435 ;
        RECT 263.675 -151.125 264.005 -150.795 ;
        RECT 263.675 -152.485 264.005 -152.155 ;
        RECT 263.675 -153.845 264.005 -153.515 ;
        RECT 263.675 -155.205 264.005 -154.875 ;
        RECT 263.675 -156.565 264.005 -156.235 ;
        RECT 263.675 -157.925 264.005 -157.595 ;
        RECT 263.675 -159.285 264.005 -158.955 ;
        RECT 263.675 -160.645 264.005 -160.315 ;
        RECT 263.675 -162.005 264.005 -161.675 ;
        RECT 263.675 -163.365 264.005 -163.035 ;
        RECT 263.675 -164.725 264.005 -164.395 ;
        RECT 263.675 -166.085 264.005 -165.755 ;
        RECT 263.675 -167.445 264.005 -167.115 ;
        RECT 263.675 -168.805 264.005 -168.475 ;
        RECT 263.675 -170.165 264.005 -169.835 ;
        RECT 263.675 -171.525 264.005 -171.195 ;
        RECT 263.675 -172.885 264.005 -172.555 ;
        RECT 263.675 -174.245 264.005 -173.915 ;
        RECT 263.675 -175.605 264.005 -175.275 ;
        RECT 263.675 -176.965 264.005 -176.635 ;
        RECT 263.675 -178.325 264.005 -177.995 ;
        RECT 263.675 -179.685 264.005 -179.355 ;
        RECT 263.675 -181.045 264.005 -180.715 ;
        RECT 263.675 -182.405 264.005 -182.075 ;
        RECT 263.675 -183.765 264.005 -183.435 ;
        RECT 263.675 -185.125 264.005 -184.795 ;
        RECT 263.675 -186.485 264.005 -186.155 ;
        RECT 263.675 -187.845 264.005 -187.515 ;
        RECT 263.675 -189.205 264.005 -188.875 ;
        RECT 263.675 -190.565 264.005 -190.235 ;
        RECT 263.675 -191.925 264.005 -191.595 ;
        RECT 263.675 -193.285 264.005 -192.955 ;
        RECT 263.675 -194.645 264.005 -194.315 ;
        RECT 263.675 -196.005 264.005 -195.675 ;
        RECT 263.675 -197.365 264.005 -197.035 ;
        RECT 263.675 -198.725 264.005 -198.395 ;
        RECT 263.675 -200.085 264.005 -199.755 ;
        RECT 263.675 -201.445 264.005 -201.115 ;
        RECT 263.675 -202.805 264.005 -202.475 ;
        RECT 263.675 -204.165 264.005 -203.835 ;
        RECT 263.675 -205.525 264.005 -205.195 ;
        RECT 263.675 -206.885 264.005 -206.555 ;
        RECT 263.675 -208.245 264.005 -207.915 ;
        RECT 263.675 -209.605 264.005 -209.275 ;
        RECT 263.675 -210.965 264.005 -210.635 ;
        RECT 263.675 -212.325 264.005 -211.995 ;
        RECT 263.675 -213.685 264.005 -213.355 ;
        RECT 263.675 -215.045 264.005 -214.715 ;
        RECT 263.675 -216.405 264.005 -216.075 ;
        RECT 263.675 -217.765 264.005 -217.435 ;
        RECT 263.675 -219.125 264.005 -218.795 ;
        RECT 263.675 -220.485 264.005 -220.155 ;
        RECT 263.675 -221.845 264.005 -221.515 ;
        RECT 263.675 -223.205 264.005 -222.875 ;
        RECT 263.675 -224.565 264.005 -224.235 ;
        RECT 263.675 -225.925 264.005 -225.595 ;
        RECT 263.675 -227.285 264.005 -226.955 ;
        RECT 263.675 -228.645 264.005 -228.315 ;
        RECT 263.675 -230.005 264.005 -229.675 ;
        RECT 263.675 -231.365 264.005 -231.035 ;
        RECT 263.675 -232.725 264.005 -232.395 ;
        RECT 263.675 -234.085 264.005 -233.755 ;
        RECT 263.675 -235.445 264.005 -235.115 ;
        RECT 263.675 -236.805 264.005 -236.475 ;
        RECT 263.675 -238.165 264.005 -237.835 ;
        RECT 263.675 -243.81 264.005 -242.68 ;
        RECT 263.68 -243.925 264 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.26 -125.535 264.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.035 246.76 265.365 247.89 ;
        RECT 265.035 241.915 265.365 242.245 ;
        RECT 265.035 240.555 265.365 240.885 ;
        RECT 265.035 239.195 265.365 239.525 ;
        RECT 265.035 237.835 265.365 238.165 ;
        RECT 265.04 237.16 265.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 246.76 266.725 247.89 ;
        RECT 266.395 241.915 266.725 242.245 ;
        RECT 266.395 240.555 266.725 240.885 ;
        RECT 266.395 239.195 266.725 239.525 ;
        RECT 266.395 237.835 266.725 238.165 ;
        RECT 266.4 237.16 266.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 -1.525 266.725 -1.195 ;
        RECT 266.395 -2.885 266.725 -2.555 ;
        RECT 266.4 -3.56 266.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 -122.565 266.725 -122.235 ;
        RECT 266.395 -123.925 266.725 -123.595 ;
        RECT 266.395 -125.285 266.725 -124.955 ;
        RECT 266.395 -126.645 266.725 -126.315 ;
        RECT 266.395 -128.005 266.725 -127.675 ;
        RECT 266.395 -129.365 266.725 -129.035 ;
        RECT 266.395 -130.725 266.725 -130.395 ;
        RECT 266.395 -132.085 266.725 -131.755 ;
        RECT 266.395 -133.445 266.725 -133.115 ;
        RECT 266.395 -134.805 266.725 -134.475 ;
        RECT 266.395 -136.165 266.725 -135.835 ;
        RECT 266.395 -137.525 266.725 -137.195 ;
        RECT 266.395 -138.885 266.725 -138.555 ;
        RECT 266.395 -140.245 266.725 -139.915 ;
        RECT 266.395 -141.605 266.725 -141.275 ;
        RECT 266.395 -142.965 266.725 -142.635 ;
        RECT 266.395 -144.325 266.725 -143.995 ;
        RECT 266.395 -145.685 266.725 -145.355 ;
        RECT 266.395 -147.045 266.725 -146.715 ;
        RECT 266.395 -148.405 266.725 -148.075 ;
        RECT 266.395 -149.765 266.725 -149.435 ;
        RECT 266.395 -151.125 266.725 -150.795 ;
        RECT 266.395 -152.485 266.725 -152.155 ;
        RECT 266.395 -153.845 266.725 -153.515 ;
        RECT 266.395 -155.205 266.725 -154.875 ;
        RECT 266.395 -156.565 266.725 -156.235 ;
        RECT 266.395 -157.925 266.725 -157.595 ;
        RECT 266.395 -159.285 266.725 -158.955 ;
        RECT 266.395 -160.645 266.725 -160.315 ;
        RECT 266.395 -162.005 266.725 -161.675 ;
        RECT 266.395 -163.365 266.725 -163.035 ;
        RECT 266.395 -164.725 266.725 -164.395 ;
        RECT 266.395 -166.085 266.725 -165.755 ;
        RECT 266.395 -167.445 266.725 -167.115 ;
        RECT 266.395 -168.805 266.725 -168.475 ;
        RECT 266.395 -170.165 266.725 -169.835 ;
        RECT 266.395 -171.525 266.725 -171.195 ;
        RECT 266.395 -172.885 266.725 -172.555 ;
        RECT 266.395 -174.245 266.725 -173.915 ;
        RECT 266.395 -175.605 266.725 -175.275 ;
        RECT 266.395 -176.965 266.725 -176.635 ;
        RECT 266.395 -178.325 266.725 -177.995 ;
        RECT 266.395 -179.685 266.725 -179.355 ;
        RECT 266.395 -181.045 266.725 -180.715 ;
        RECT 266.395 -182.405 266.725 -182.075 ;
        RECT 266.395 -183.765 266.725 -183.435 ;
        RECT 266.395 -185.125 266.725 -184.795 ;
        RECT 266.395 -186.485 266.725 -186.155 ;
        RECT 266.395 -187.845 266.725 -187.515 ;
        RECT 266.395 -189.205 266.725 -188.875 ;
        RECT 266.395 -190.565 266.725 -190.235 ;
        RECT 266.395 -191.925 266.725 -191.595 ;
        RECT 266.395 -193.285 266.725 -192.955 ;
        RECT 266.395 -194.645 266.725 -194.315 ;
        RECT 266.395 -196.005 266.725 -195.675 ;
        RECT 266.395 -197.365 266.725 -197.035 ;
        RECT 266.395 -198.725 266.725 -198.395 ;
        RECT 266.395 -200.085 266.725 -199.755 ;
        RECT 266.395 -201.445 266.725 -201.115 ;
        RECT 266.395 -202.805 266.725 -202.475 ;
        RECT 266.395 -204.165 266.725 -203.835 ;
        RECT 266.395 -205.525 266.725 -205.195 ;
        RECT 266.395 -206.885 266.725 -206.555 ;
        RECT 266.395 -208.245 266.725 -207.915 ;
        RECT 266.395 -209.605 266.725 -209.275 ;
        RECT 266.395 -210.965 266.725 -210.635 ;
        RECT 266.395 -212.325 266.725 -211.995 ;
        RECT 266.395 -213.685 266.725 -213.355 ;
        RECT 266.395 -215.045 266.725 -214.715 ;
        RECT 266.395 -216.405 266.725 -216.075 ;
        RECT 266.395 -217.765 266.725 -217.435 ;
        RECT 266.395 -219.125 266.725 -218.795 ;
        RECT 266.395 -220.485 266.725 -220.155 ;
        RECT 266.395 -221.845 266.725 -221.515 ;
        RECT 266.395 -223.205 266.725 -222.875 ;
        RECT 266.395 -224.565 266.725 -224.235 ;
        RECT 266.395 -225.925 266.725 -225.595 ;
        RECT 266.395 -227.285 266.725 -226.955 ;
        RECT 266.395 -228.645 266.725 -228.315 ;
        RECT 266.395 -230.005 266.725 -229.675 ;
        RECT 266.395 -231.365 266.725 -231.035 ;
        RECT 266.395 -232.725 266.725 -232.395 ;
        RECT 266.395 -234.085 266.725 -233.755 ;
        RECT 266.395 -235.445 266.725 -235.115 ;
        RECT 266.395 -236.805 266.725 -236.475 ;
        RECT 266.395 -238.165 266.725 -237.835 ;
        RECT 266.395 -243.81 266.725 -242.68 ;
        RECT 266.4 -243.925 266.72 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 246.76 268.085 247.89 ;
        RECT 267.755 241.915 268.085 242.245 ;
        RECT 267.755 240.555 268.085 240.885 ;
        RECT 267.755 239.195 268.085 239.525 ;
        RECT 267.755 237.835 268.085 238.165 ;
        RECT 267.76 237.16 268.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 -1.525 268.085 -1.195 ;
        RECT 267.755 -2.885 268.085 -2.555 ;
        RECT 267.76 -3.56 268.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 246.76 269.445 247.89 ;
        RECT 269.115 241.915 269.445 242.245 ;
        RECT 269.115 240.555 269.445 240.885 ;
        RECT 269.115 239.195 269.445 239.525 ;
        RECT 269.115 237.835 269.445 238.165 ;
        RECT 269.12 237.16 269.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 -1.525 269.445 -1.195 ;
        RECT 269.115 -2.885 269.445 -2.555 ;
        RECT 269.12 -3.56 269.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 -122.565 269.445 -122.235 ;
        RECT 269.115 -123.925 269.445 -123.595 ;
        RECT 269.115 -125.285 269.445 -124.955 ;
        RECT 269.115 -126.645 269.445 -126.315 ;
        RECT 269.115 -128.005 269.445 -127.675 ;
        RECT 269.115 -129.365 269.445 -129.035 ;
        RECT 269.115 -130.725 269.445 -130.395 ;
        RECT 269.115 -132.085 269.445 -131.755 ;
        RECT 269.115 -133.445 269.445 -133.115 ;
        RECT 269.115 -134.805 269.445 -134.475 ;
        RECT 269.115 -136.165 269.445 -135.835 ;
        RECT 269.115 -137.525 269.445 -137.195 ;
        RECT 269.115 -138.885 269.445 -138.555 ;
        RECT 269.115 -140.245 269.445 -139.915 ;
        RECT 269.115 -141.605 269.445 -141.275 ;
        RECT 269.115 -142.965 269.445 -142.635 ;
        RECT 269.115 -144.325 269.445 -143.995 ;
        RECT 269.115 -145.685 269.445 -145.355 ;
        RECT 269.115 -147.045 269.445 -146.715 ;
        RECT 269.115 -148.405 269.445 -148.075 ;
        RECT 269.115 -149.765 269.445 -149.435 ;
        RECT 269.115 -151.125 269.445 -150.795 ;
        RECT 269.115 -152.485 269.445 -152.155 ;
        RECT 269.115 -153.845 269.445 -153.515 ;
        RECT 269.115 -155.205 269.445 -154.875 ;
        RECT 269.115 -156.565 269.445 -156.235 ;
        RECT 269.115 -157.925 269.445 -157.595 ;
        RECT 269.115 -159.285 269.445 -158.955 ;
        RECT 269.115 -160.645 269.445 -160.315 ;
        RECT 269.115 -162.005 269.445 -161.675 ;
        RECT 269.115 -163.365 269.445 -163.035 ;
        RECT 269.115 -164.725 269.445 -164.395 ;
        RECT 269.115 -166.085 269.445 -165.755 ;
        RECT 269.115 -167.445 269.445 -167.115 ;
        RECT 269.115 -168.805 269.445 -168.475 ;
        RECT 269.115 -170.165 269.445 -169.835 ;
        RECT 269.115 -171.525 269.445 -171.195 ;
        RECT 269.115 -172.885 269.445 -172.555 ;
        RECT 269.115 -174.245 269.445 -173.915 ;
        RECT 269.115 -175.605 269.445 -175.275 ;
        RECT 269.115 -176.965 269.445 -176.635 ;
        RECT 269.115 -178.325 269.445 -177.995 ;
        RECT 269.115 -179.685 269.445 -179.355 ;
        RECT 269.115 -181.045 269.445 -180.715 ;
        RECT 269.115 -182.405 269.445 -182.075 ;
        RECT 269.115 -183.765 269.445 -183.435 ;
        RECT 269.115 -185.125 269.445 -184.795 ;
        RECT 269.115 -186.485 269.445 -186.155 ;
        RECT 269.115 -187.845 269.445 -187.515 ;
        RECT 269.115 -189.205 269.445 -188.875 ;
        RECT 269.115 -190.565 269.445 -190.235 ;
        RECT 269.115 -191.925 269.445 -191.595 ;
        RECT 269.115 -193.285 269.445 -192.955 ;
        RECT 269.115 -194.645 269.445 -194.315 ;
        RECT 269.115 -196.005 269.445 -195.675 ;
        RECT 269.115 -197.365 269.445 -197.035 ;
        RECT 269.115 -198.725 269.445 -198.395 ;
        RECT 269.115 -200.085 269.445 -199.755 ;
        RECT 269.115 -201.445 269.445 -201.115 ;
        RECT 269.115 -202.805 269.445 -202.475 ;
        RECT 269.115 -204.165 269.445 -203.835 ;
        RECT 269.115 -205.525 269.445 -205.195 ;
        RECT 269.115 -206.885 269.445 -206.555 ;
        RECT 269.115 -208.245 269.445 -207.915 ;
        RECT 269.115 -209.605 269.445 -209.275 ;
        RECT 269.115 -210.965 269.445 -210.635 ;
        RECT 269.115 -212.325 269.445 -211.995 ;
        RECT 269.115 -213.685 269.445 -213.355 ;
        RECT 269.115 -215.045 269.445 -214.715 ;
        RECT 269.115 -216.405 269.445 -216.075 ;
        RECT 269.115 -217.765 269.445 -217.435 ;
        RECT 269.115 -219.125 269.445 -218.795 ;
        RECT 269.115 -220.485 269.445 -220.155 ;
        RECT 269.115 -221.845 269.445 -221.515 ;
        RECT 269.115 -223.205 269.445 -222.875 ;
        RECT 269.115 -224.565 269.445 -224.235 ;
        RECT 269.115 -225.925 269.445 -225.595 ;
        RECT 269.115 -227.285 269.445 -226.955 ;
        RECT 269.115 -228.645 269.445 -228.315 ;
        RECT 269.115 -230.005 269.445 -229.675 ;
        RECT 269.115 -231.365 269.445 -231.035 ;
        RECT 269.115 -232.725 269.445 -232.395 ;
        RECT 269.115 -234.085 269.445 -233.755 ;
        RECT 269.115 -235.445 269.445 -235.115 ;
        RECT 269.115 -236.805 269.445 -236.475 ;
        RECT 269.115 -238.165 269.445 -237.835 ;
        RECT 269.115 -243.81 269.445 -242.68 ;
        RECT 269.12 -243.925 269.44 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 246.76 270.805 247.89 ;
        RECT 270.475 241.915 270.805 242.245 ;
        RECT 270.475 240.555 270.805 240.885 ;
        RECT 270.475 239.195 270.805 239.525 ;
        RECT 270.475 237.835 270.805 238.165 ;
        RECT 270.48 237.16 270.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 -1.525 270.805 -1.195 ;
        RECT 270.475 -2.885 270.805 -2.555 ;
        RECT 270.48 -3.56 270.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 -122.565 270.805 -122.235 ;
        RECT 270.475 -123.925 270.805 -123.595 ;
        RECT 270.475 -125.285 270.805 -124.955 ;
        RECT 270.475 -126.645 270.805 -126.315 ;
        RECT 270.475 -128.005 270.805 -127.675 ;
        RECT 270.475 -129.365 270.805 -129.035 ;
        RECT 270.475 -130.725 270.805 -130.395 ;
        RECT 270.475 -132.085 270.805 -131.755 ;
        RECT 270.475 -133.445 270.805 -133.115 ;
        RECT 270.475 -134.805 270.805 -134.475 ;
        RECT 270.475 -136.165 270.805 -135.835 ;
        RECT 270.475 -137.525 270.805 -137.195 ;
        RECT 270.475 -138.885 270.805 -138.555 ;
        RECT 270.475 -140.245 270.805 -139.915 ;
        RECT 270.475 -141.605 270.805 -141.275 ;
        RECT 270.475 -142.965 270.805 -142.635 ;
        RECT 270.475 -144.325 270.805 -143.995 ;
        RECT 270.475 -145.685 270.805 -145.355 ;
        RECT 270.475 -147.045 270.805 -146.715 ;
        RECT 270.475 -148.405 270.805 -148.075 ;
        RECT 270.475 -149.765 270.805 -149.435 ;
        RECT 270.475 -151.125 270.805 -150.795 ;
        RECT 270.475 -152.485 270.805 -152.155 ;
        RECT 270.475 -153.845 270.805 -153.515 ;
        RECT 270.475 -155.205 270.805 -154.875 ;
        RECT 270.475 -156.565 270.805 -156.235 ;
        RECT 270.475 -157.925 270.805 -157.595 ;
        RECT 270.475 -159.285 270.805 -158.955 ;
        RECT 270.475 -160.645 270.805 -160.315 ;
        RECT 270.475 -162.005 270.805 -161.675 ;
        RECT 270.475 -163.365 270.805 -163.035 ;
        RECT 270.475 -164.725 270.805 -164.395 ;
        RECT 270.475 -166.085 270.805 -165.755 ;
        RECT 270.475 -167.445 270.805 -167.115 ;
        RECT 270.475 -168.805 270.805 -168.475 ;
        RECT 270.475 -170.165 270.805 -169.835 ;
        RECT 270.475 -171.525 270.805 -171.195 ;
        RECT 270.475 -172.885 270.805 -172.555 ;
        RECT 270.475 -174.245 270.805 -173.915 ;
        RECT 270.475 -175.605 270.805 -175.275 ;
        RECT 270.475 -176.965 270.805 -176.635 ;
        RECT 270.475 -178.325 270.805 -177.995 ;
        RECT 270.475 -179.685 270.805 -179.355 ;
        RECT 270.475 -181.045 270.805 -180.715 ;
        RECT 270.475 -182.405 270.805 -182.075 ;
        RECT 270.475 -183.765 270.805 -183.435 ;
        RECT 270.475 -185.125 270.805 -184.795 ;
        RECT 270.475 -186.485 270.805 -186.155 ;
        RECT 270.475 -187.845 270.805 -187.515 ;
        RECT 270.475 -189.205 270.805 -188.875 ;
        RECT 270.475 -190.565 270.805 -190.235 ;
        RECT 270.475 -191.925 270.805 -191.595 ;
        RECT 270.475 -193.285 270.805 -192.955 ;
        RECT 270.475 -194.645 270.805 -194.315 ;
        RECT 270.475 -196.005 270.805 -195.675 ;
        RECT 270.475 -197.365 270.805 -197.035 ;
        RECT 270.475 -198.725 270.805 -198.395 ;
        RECT 270.475 -200.085 270.805 -199.755 ;
        RECT 270.475 -201.445 270.805 -201.115 ;
        RECT 270.475 -202.805 270.805 -202.475 ;
        RECT 270.475 -204.165 270.805 -203.835 ;
        RECT 270.475 -205.525 270.805 -205.195 ;
        RECT 270.475 -206.885 270.805 -206.555 ;
        RECT 270.475 -208.245 270.805 -207.915 ;
        RECT 270.475 -209.605 270.805 -209.275 ;
        RECT 270.475 -210.965 270.805 -210.635 ;
        RECT 270.475 -212.325 270.805 -211.995 ;
        RECT 270.475 -213.685 270.805 -213.355 ;
        RECT 270.475 -215.045 270.805 -214.715 ;
        RECT 270.475 -216.405 270.805 -216.075 ;
        RECT 270.475 -217.765 270.805 -217.435 ;
        RECT 270.475 -219.125 270.805 -218.795 ;
        RECT 270.475 -220.485 270.805 -220.155 ;
        RECT 270.475 -221.845 270.805 -221.515 ;
        RECT 270.475 -223.205 270.805 -222.875 ;
        RECT 270.475 -224.565 270.805 -224.235 ;
        RECT 270.475 -225.925 270.805 -225.595 ;
        RECT 270.475 -227.285 270.805 -226.955 ;
        RECT 270.475 -228.645 270.805 -228.315 ;
        RECT 270.475 -230.005 270.805 -229.675 ;
        RECT 270.475 -231.365 270.805 -231.035 ;
        RECT 270.475 -232.725 270.805 -232.395 ;
        RECT 270.475 -234.085 270.805 -233.755 ;
        RECT 270.475 -235.445 270.805 -235.115 ;
        RECT 270.475 -236.805 270.805 -236.475 ;
        RECT 270.475 -238.165 270.805 -237.835 ;
        RECT 270.475 -243.81 270.805 -242.68 ;
        RECT 270.48 -243.925 270.8 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 246.76 272.165 247.89 ;
        RECT 271.835 241.915 272.165 242.245 ;
        RECT 271.835 240.555 272.165 240.885 ;
        RECT 271.835 239.195 272.165 239.525 ;
        RECT 271.835 237.835 272.165 238.165 ;
        RECT 271.84 237.16 272.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 -1.525 272.165 -1.195 ;
        RECT 271.835 -2.885 272.165 -2.555 ;
        RECT 271.84 -3.56 272.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 -122.565 272.165 -122.235 ;
        RECT 271.835 -123.925 272.165 -123.595 ;
        RECT 271.835 -125.285 272.165 -124.955 ;
        RECT 271.835 -126.645 272.165 -126.315 ;
        RECT 271.835 -128.005 272.165 -127.675 ;
        RECT 271.835 -129.365 272.165 -129.035 ;
        RECT 271.835 -130.725 272.165 -130.395 ;
        RECT 271.835 -132.085 272.165 -131.755 ;
        RECT 271.835 -133.445 272.165 -133.115 ;
        RECT 271.835 -134.805 272.165 -134.475 ;
        RECT 271.835 -136.165 272.165 -135.835 ;
        RECT 271.835 -137.525 272.165 -137.195 ;
        RECT 271.835 -138.885 272.165 -138.555 ;
        RECT 271.835 -140.245 272.165 -139.915 ;
        RECT 271.835 -141.605 272.165 -141.275 ;
        RECT 271.835 -142.965 272.165 -142.635 ;
        RECT 271.835 -144.325 272.165 -143.995 ;
        RECT 271.835 -145.685 272.165 -145.355 ;
        RECT 271.835 -147.045 272.165 -146.715 ;
        RECT 271.835 -148.405 272.165 -148.075 ;
        RECT 271.835 -149.765 272.165 -149.435 ;
        RECT 271.835 -151.125 272.165 -150.795 ;
        RECT 271.835 -152.485 272.165 -152.155 ;
        RECT 271.835 -153.845 272.165 -153.515 ;
        RECT 271.835 -155.205 272.165 -154.875 ;
        RECT 271.835 -156.565 272.165 -156.235 ;
        RECT 271.835 -157.925 272.165 -157.595 ;
        RECT 271.835 -159.285 272.165 -158.955 ;
        RECT 271.835 -160.645 272.165 -160.315 ;
        RECT 271.835 -162.005 272.165 -161.675 ;
        RECT 271.835 -163.365 272.165 -163.035 ;
        RECT 271.835 -164.725 272.165 -164.395 ;
        RECT 271.835 -166.085 272.165 -165.755 ;
        RECT 271.835 -167.445 272.165 -167.115 ;
        RECT 271.835 -168.805 272.165 -168.475 ;
        RECT 271.835 -170.165 272.165 -169.835 ;
        RECT 271.835 -171.525 272.165 -171.195 ;
        RECT 271.835 -172.885 272.165 -172.555 ;
        RECT 271.835 -174.245 272.165 -173.915 ;
        RECT 271.835 -175.605 272.165 -175.275 ;
        RECT 271.835 -176.965 272.165 -176.635 ;
        RECT 271.835 -178.325 272.165 -177.995 ;
        RECT 271.835 -179.685 272.165 -179.355 ;
        RECT 271.835 -181.045 272.165 -180.715 ;
        RECT 271.835 -182.405 272.165 -182.075 ;
        RECT 271.835 -183.765 272.165 -183.435 ;
        RECT 271.835 -185.125 272.165 -184.795 ;
        RECT 271.835 -186.485 272.165 -186.155 ;
        RECT 271.835 -187.845 272.165 -187.515 ;
        RECT 271.835 -189.205 272.165 -188.875 ;
        RECT 271.835 -190.565 272.165 -190.235 ;
        RECT 271.835 -191.925 272.165 -191.595 ;
        RECT 271.835 -193.285 272.165 -192.955 ;
        RECT 271.835 -194.645 272.165 -194.315 ;
        RECT 271.835 -196.005 272.165 -195.675 ;
        RECT 271.835 -197.365 272.165 -197.035 ;
        RECT 271.835 -198.725 272.165 -198.395 ;
        RECT 271.835 -200.085 272.165 -199.755 ;
        RECT 271.835 -201.445 272.165 -201.115 ;
        RECT 271.835 -202.805 272.165 -202.475 ;
        RECT 271.835 -204.165 272.165 -203.835 ;
        RECT 271.835 -205.525 272.165 -205.195 ;
        RECT 271.835 -206.885 272.165 -206.555 ;
        RECT 271.835 -208.245 272.165 -207.915 ;
        RECT 271.835 -209.605 272.165 -209.275 ;
        RECT 271.835 -210.965 272.165 -210.635 ;
        RECT 271.835 -212.325 272.165 -211.995 ;
        RECT 271.835 -213.685 272.165 -213.355 ;
        RECT 271.835 -215.045 272.165 -214.715 ;
        RECT 271.835 -216.405 272.165 -216.075 ;
        RECT 271.835 -217.765 272.165 -217.435 ;
        RECT 271.835 -219.125 272.165 -218.795 ;
        RECT 271.835 -220.485 272.165 -220.155 ;
        RECT 271.835 -221.845 272.165 -221.515 ;
        RECT 271.835 -223.205 272.165 -222.875 ;
        RECT 271.835 -224.565 272.165 -224.235 ;
        RECT 271.835 -225.925 272.165 -225.595 ;
        RECT 271.835 -227.285 272.165 -226.955 ;
        RECT 271.835 -228.645 272.165 -228.315 ;
        RECT 271.835 -230.005 272.165 -229.675 ;
        RECT 271.835 -231.365 272.165 -231.035 ;
        RECT 271.835 -232.725 272.165 -232.395 ;
        RECT 271.835 -234.085 272.165 -233.755 ;
        RECT 271.835 -235.445 272.165 -235.115 ;
        RECT 271.835 -236.805 272.165 -236.475 ;
        RECT 271.835 -238.165 272.165 -237.835 ;
        RECT 271.835 -243.81 272.165 -242.68 ;
        RECT 271.84 -243.925 272.16 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 246.76 273.525 247.89 ;
        RECT 273.195 241.915 273.525 242.245 ;
        RECT 273.195 240.555 273.525 240.885 ;
        RECT 273.195 239.195 273.525 239.525 ;
        RECT 273.195 237.835 273.525 238.165 ;
        RECT 273.2 237.16 273.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 -1.525 273.525 -1.195 ;
        RECT 273.195 -2.885 273.525 -2.555 ;
        RECT 273.2 -3.56 273.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 -122.565 273.525 -122.235 ;
        RECT 273.195 -123.925 273.525 -123.595 ;
        RECT 273.195 -125.285 273.525 -124.955 ;
        RECT 273.195 -126.645 273.525 -126.315 ;
        RECT 273.195 -128.005 273.525 -127.675 ;
        RECT 273.195 -129.365 273.525 -129.035 ;
        RECT 273.195 -130.725 273.525 -130.395 ;
        RECT 273.195 -132.085 273.525 -131.755 ;
        RECT 273.195 -133.445 273.525 -133.115 ;
        RECT 273.195 -134.805 273.525 -134.475 ;
        RECT 273.195 -136.165 273.525 -135.835 ;
        RECT 273.195 -137.525 273.525 -137.195 ;
        RECT 273.195 -138.885 273.525 -138.555 ;
        RECT 273.195 -140.245 273.525 -139.915 ;
        RECT 273.195 -141.605 273.525 -141.275 ;
        RECT 273.195 -142.965 273.525 -142.635 ;
        RECT 273.195 -144.325 273.525 -143.995 ;
        RECT 273.195 -145.685 273.525 -145.355 ;
        RECT 273.195 -147.045 273.525 -146.715 ;
        RECT 273.195 -148.405 273.525 -148.075 ;
        RECT 273.195 -149.765 273.525 -149.435 ;
        RECT 273.195 -151.125 273.525 -150.795 ;
        RECT 273.195 -152.485 273.525 -152.155 ;
        RECT 273.195 -153.845 273.525 -153.515 ;
        RECT 273.195 -155.205 273.525 -154.875 ;
        RECT 273.195 -156.565 273.525 -156.235 ;
        RECT 273.195 -157.925 273.525 -157.595 ;
        RECT 273.195 -159.285 273.525 -158.955 ;
        RECT 273.195 -160.645 273.525 -160.315 ;
        RECT 273.195 -162.005 273.525 -161.675 ;
        RECT 273.195 -163.365 273.525 -163.035 ;
        RECT 273.195 -164.725 273.525 -164.395 ;
        RECT 273.195 -166.085 273.525 -165.755 ;
        RECT 273.195 -167.445 273.525 -167.115 ;
        RECT 273.195 -168.805 273.525 -168.475 ;
        RECT 273.195 -170.165 273.525 -169.835 ;
        RECT 273.195 -171.525 273.525 -171.195 ;
        RECT 273.195 -172.885 273.525 -172.555 ;
        RECT 273.195 -174.245 273.525 -173.915 ;
        RECT 273.195 -175.605 273.525 -175.275 ;
        RECT 273.195 -176.965 273.525 -176.635 ;
        RECT 273.195 -178.325 273.525 -177.995 ;
        RECT 273.195 -179.685 273.525 -179.355 ;
        RECT 273.195 -181.045 273.525 -180.715 ;
        RECT 273.195 -182.405 273.525 -182.075 ;
        RECT 273.195 -183.765 273.525 -183.435 ;
        RECT 273.195 -185.125 273.525 -184.795 ;
        RECT 273.195 -186.485 273.525 -186.155 ;
        RECT 273.195 -187.845 273.525 -187.515 ;
        RECT 273.195 -189.205 273.525 -188.875 ;
        RECT 273.195 -190.565 273.525 -190.235 ;
        RECT 273.195 -191.925 273.525 -191.595 ;
        RECT 273.195 -193.285 273.525 -192.955 ;
        RECT 273.195 -194.645 273.525 -194.315 ;
        RECT 273.195 -196.005 273.525 -195.675 ;
        RECT 273.195 -197.365 273.525 -197.035 ;
        RECT 273.195 -198.725 273.525 -198.395 ;
        RECT 273.195 -200.085 273.525 -199.755 ;
        RECT 273.195 -201.445 273.525 -201.115 ;
        RECT 273.195 -202.805 273.525 -202.475 ;
        RECT 273.195 -204.165 273.525 -203.835 ;
        RECT 273.195 -205.525 273.525 -205.195 ;
        RECT 273.195 -206.885 273.525 -206.555 ;
        RECT 273.195 -208.245 273.525 -207.915 ;
        RECT 273.195 -209.605 273.525 -209.275 ;
        RECT 273.195 -210.965 273.525 -210.635 ;
        RECT 273.195 -212.325 273.525 -211.995 ;
        RECT 273.195 -213.685 273.525 -213.355 ;
        RECT 273.195 -215.045 273.525 -214.715 ;
        RECT 273.195 -216.405 273.525 -216.075 ;
        RECT 273.195 -217.765 273.525 -217.435 ;
        RECT 273.195 -219.125 273.525 -218.795 ;
        RECT 273.195 -220.485 273.525 -220.155 ;
        RECT 273.195 -221.845 273.525 -221.515 ;
        RECT 273.195 -223.205 273.525 -222.875 ;
        RECT 273.195 -224.565 273.525 -224.235 ;
        RECT 273.195 -225.925 273.525 -225.595 ;
        RECT 273.195 -227.285 273.525 -226.955 ;
        RECT 273.195 -228.645 273.525 -228.315 ;
        RECT 273.195 -230.005 273.525 -229.675 ;
        RECT 273.195 -231.365 273.525 -231.035 ;
        RECT 273.195 -232.725 273.525 -232.395 ;
        RECT 273.195 -234.085 273.525 -233.755 ;
        RECT 273.195 -235.445 273.525 -235.115 ;
        RECT 273.195 -236.805 273.525 -236.475 ;
        RECT 273.195 -238.165 273.525 -237.835 ;
        RECT 273.195 -243.81 273.525 -242.68 ;
        RECT 273.2 -243.925 273.52 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 246.76 274.885 247.89 ;
        RECT 274.555 241.915 274.885 242.245 ;
        RECT 274.555 240.555 274.885 240.885 ;
        RECT 274.555 239.195 274.885 239.525 ;
        RECT 274.555 237.835 274.885 238.165 ;
        RECT 274.56 237.16 274.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 -126.645 274.885 -126.315 ;
        RECT 274.555 -128.005 274.885 -127.675 ;
        RECT 274.555 -129.365 274.885 -129.035 ;
        RECT 274.555 -130.725 274.885 -130.395 ;
        RECT 274.555 -132.085 274.885 -131.755 ;
        RECT 274.555 -133.445 274.885 -133.115 ;
        RECT 274.555 -134.805 274.885 -134.475 ;
        RECT 274.555 -136.165 274.885 -135.835 ;
        RECT 274.555 -137.525 274.885 -137.195 ;
        RECT 274.555 -138.885 274.885 -138.555 ;
        RECT 274.555 -140.245 274.885 -139.915 ;
        RECT 274.555 -141.605 274.885 -141.275 ;
        RECT 274.555 -142.965 274.885 -142.635 ;
        RECT 274.555 -144.325 274.885 -143.995 ;
        RECT 274.555 -145.685 274.885 -145.355 ;
        RECT 274.555 -147.045 274.885 -146.715 ;
        RECT 274.555 -148.405 274.885 -148.075 ;
        RECT 274.555 -149.765 274.885 -149.435 ;
        RECT 274.555 -151.125 274.885 -150.795 ;
        RECT 274.555 -152.485 274.885 -152.155 ;
        RECT 274.555 -153.845 274.885 -153.515 ;
        RECT 274.555 -155.205 274.885 -154.875 ;
        RECT 274.555 -156.565 274.885 -156.235 ;
        RECT 274.555 -157.925 274.885 -157.595 ;
        RECT 274.555 -159.285 274.885 -158.955 ;
        RECT 274.555 -160.645 274.885 -160.315 ;
        RECT 274.555 -162.005 274.885 -161.675 ;
        RECT 274.555 -163.365 274.885 -163.035 ;
        RECT 274.555 -164.725 274.885 -164.395 ;
        RECT 274.555 -166.085 274.885 -165.755 ;
        RECT 274.555 -167.445 274.885 -167.115 ;
        RECT 274.555 -168.805 274.885 -168.475 ;
        RECT 274.555 -170.165 274.885 -169.835 ;
        RECT 274.555 -171.525 274.885 -171.195 ;
        RECT 274.555 -172.885 274.885 -172.555 ;
        RECT 274.555 -174.245 274.885 -173.915 ;
        RECT 274.555 -175.605 274.885 -175.275 ;
        RECT 274.555 -176.965 274.885 -176.635 ;
        RECT 274.555 -178.325 274.885 -177.995 ;
        RECT 274.555 -179.685 274.885 -179.355 ;
        RECT 274.555 -181.045 274.885 -180.715 ;
        RECT 274.555 -182.405 274.885 -182.075 ;
        RECT 274.555 -183.765 274.885 -183.435 ;
        RECT 274.555 -185.125 274.885 -184.795 ;
        RECT 274.555 -186.485 274.885 -186.155 ;
        RECT 274.555 -187.845 274.885 -187.515 ;
        RECT 274.555 -189.205 274.885 -188.875 ;
        RECT 274.555 -190.565 274.885 -190.235 ;
        RECT 274.555 -191.925 274.885 -191.595 ;
        RECT 274.555 -193.285 274.885 -192.955 ;
        RECT 274.555 -194.645 274.885 -194.315 ;
        RECT 274.555 -196.005 274.885 -195.675 ;
        RECT 274.555 -197.365 274.885 -197.035 ;
        RECT 274.555 -198.725 274.885 -198.395 ;
        RECT 274.555 -200.085 274.885 -199.755 ;
        RECT 274.555 -201.445 274.885 -201.115 ;
        RECT 274.555 -202.805 274.885 -202.475 ;
        RECT 274.555 -204.165 274.885 -203.835 ;
        RECT 274.555 -205.525 274.885 -205.195 ;
        RECT 274.555 -206.885 274.885 -206.555 ;
        RECT 274.555 -208.245 274.885 -207.915 ;
        RECT 274.555 -209.605 274.885 -209.275 ;
        RECT 274.555 -210.965 274.885 -210.635 ;
        RECT 274.555 -212.325 274.885 -211.995 ;
        RECT 274.555 -213.685 274.885 -213.355 ;
        RECT 274.555 -215.045 274.885 -214.715 ;
        RECT 274.555 -216.405 274.885 -216.075 ;
        RECT 274.555 -217.765 274.885 -217.435 ;
        RECT 274.555 -219.125 274.885 -218.795 ;
        RECT 274.555 -220.485 274.885 -220.155 ;
        RECT 274.555 -221.845 274.885 -221.515 ;
        RECT 274.555 -223.205 274.885 -222.875 ;
        RECT 274.555 -224.565 274.885 -224.235 ;
        RECT 274.555 -225.925 274.885 -225.595 ;
        RECT 274.555 -227.285 274.885 -226.955 ;
        RECT 274.555 -228.645 274.885 -228.315 ;
        RECT 274.555 -230.005 274.885 -229.675 ;
        RECT 274.555 -231.365 274.885 -231.035 ;
        RECT 274.555 -232.725 274.885 -232.395 ;
        RECT 274.555 -234.085 274.885 -233.755 ;
        RECT 274.555 -235.445 274.885 -235.115 ;
        RECT 274.555 -236.805 274.885 -236.475 ;
        RECT 274.555 -238.165 274.885 -237.835 ;
        RECT 274.555 -243.81 274.885 -242.68 ;
        RECT 274.56 -243.925 274.88 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.16 -125.535 275.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.915 246.76 276.245 247.89 ;
        RECT 275.915 241.915 276.245 242.245 ;
        RECT 275.915 240.555 276.245 240.885 ;
        RECT 275.915 239.195 276.245 239.525 ;
        RECT 275.915 237.835 276.245 238.165 ;
        RECT 275.92 237.16 276.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 246.76 277.605 247.89 ;
        RECT 277.275 241.915 277.605 242.245 ;
        RECT 277.275 240.555 277.605 240.885 ;
        RECT 277.275 239.195 277.605 239.525 ;
        RECT 277.275 237.835 277.605 238.165 ;
        RECT 277.28 237.16 277.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 -1.525 277.605 -1.195 ;
        RECT 277.275 -2.885 277.605 -2.555 ;
        RECT 277.28 -3.56 277.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 -122.565 277.605 -122.235 ;
        RECT 277.275 -123.925 277.605 -123.595 ;
        RECT 277.275 -125.285 277.605 -124.955 ;
        RECT 277.275 -126.645 277.605 -126.315 ;
        RECT 277.275 -128.005 277.605 -127.675 ;
        RECT 277.275 -129.365 277.605 -129.035 ;
        RECT 277.275 -130.725 277.605 -130.395 ;
        RECT 277.275 -132.085 277.605 -131.755 ;
        RECT 277.275 -133.445 277.605 -133.115 ;
        RECT 277.275 -134.805 277.605 -134.475 ;
        RECT 277.275 -136.165 277.605 -135.835 ;
        RECT 277.275 -137.525 277.605 -137.195 ;
        RECT 277.275 -138.885 277.605 -138.555 ;
        RECT 277.275 -140.245 277.605 -139.915 ;
        RECT 277.275 -141.605 277.605 -141.275 ;
        RECT 277.275 -142.965 277.605 -142.635 ;
        RECT 277.275 -144.325 277.605 -143.995 ;
        RECT 277.275 -145.685 277.605 -145.355 ;
        RECT 277.275 -147.045 277.605 -146.715 ;
        RECT 277.275 -148.405 277.605 -148.075 ;
        RECT 277.275 -149.765 277.605 -149.435 ;
        RECT 277.275 -151.125 277.605 -150.795 ;
        RECT 277.275 -152.485 277.605 -152.155 ;
        RECT 277.275 -153.845 277.605 -153.515 ;
        RECT 277.275 -155.205 277.605 -154.875 ;
        RECT 277.275 -156.565 277.605 -156.235 ;
        RECT 277.275 -157.925 277.605 -157.595 ;
        RECT 277.275 -159.285 277.605 -158.955 ;
        RECT 277.275 -160.645 277.605 -160.315 ;
        RECT 277.275 -162.005 277.605 -161.675 ;
        RECT 277.275 -163.365 277.605 -163.035 ;
        RECT 277.275 -164.725 277.605 -164.395 ;
        RECT 277.275 -166.085 277.605 -165.755 ;
        RECT 277.275 -167.445 277.605 -167.115 ;
        RECT 277.275 -168.805 277.605 -168.475 ;
        RECT 277.275 -170.165 277.605 -169.835 ;
        RECT 277.275 -171.525 277.605 -171.195 ;
        RECT 277.275 -172.885 277.605 -172.555 ;
        RECT 277.275 -174.245 277.605 -173.915 ;
        RECT 277.275 -175.605 277.605 -175.275 ;
        RECT 277.275 -176.965 277.605 -176.635 ;
        RECT 277.275 -178.325 277.605 -177.995 ;
        RECT 277.275 -179.685 277.605 -179.355 ;
        RECT 277.275 -181.045 277.605 -180.715 ;
        RECT 277.275 -182.405 277.605 -182.075 ;
        RECT 277.275 -183.765 277.605 -183.435 ;
        RECT 277.275 -185.125 277.605 -184.795 ;
        RECT 277.275 -186.485 277.605 -186.155 ;
        RECT 277.275 -187.845 277.605 -187.515 ;
        RECT 277.275 -189.205 277.605 -188.875 ;
        RECT 277.275 -190.565 277.605 -190.235 ;
        RECT 277.275 -191.925 277.605 -191.595 ;
        RECT 277.275 -193.285 277.605 -192.955 ;
        RECT 277.275 -194.645 277.605 -194.315 ;
        RECT 277.275 -196.005 277.605 -195.675 ;
        RECT 277.275 -197.365 277.605 -197.035 ;
        RECT 277.275 -198.725 277.605 -198.395 ;
        RECT 277.275 -200.085 277.605 -199.755 ;
        RECT 277.275 -201.445 277.605 -201.115 ;
        RECT 277.275 -202.805 277.605 -202.475 ;
        RECT 277.275 -204.165 277.605 -203.835 ;
        RECT 277.275 -205.525 277.605 -205.195 ;
        RECT 277.275 -206.885 277.605 -206.555 ;
        RECT 277.275 -208.245 277.605 -207.915 ;
        RECT 277.275 -209.605 277.605 -209.275 ;
        RECT 277.275 -210.965 277.605 -210.635 ;
        RECT 277.275 -212.325 277.605 -211.995 ;
        RECT 277.275 -213.685 277.605 -213.355 ;
        RECT 277.275 -215.045 277.605 -214.715 ;
        RECT 277.275 -216.405 277.605 -216.075 ;
        RECT 277.275 -217.765 277.605 -217.435 ;
        RECT 277.275 -219.125 277.605 -218.795 ;
        RECT 277.275 -220.485 277.605 -220.155 ;
        RECT 277.275 -221.845 277.605 -221.515 ;
        RECT 277.275 -223.205 277.605 -222.875 ;
        RECT 277.275 -224.565 277.605 -224.235 ;
        RECT 277.275 -225.925 277.605 -225.595 ;
        RECT 277.275 -227.285 277.605 -226.955 ;
        RECT 277.275 -228.645 277.605 -228.315 ;
        RECT 277.275 -230.005 277.605 -229.675 ;
        RECT 277.275 -231.365 277.605 -231.035 ;
        RECT 277.275 -232.725 277.605 -232.395 ;
        RECT 277.275 -234.085 277.605 -233.755 ;
        RECT 277.275 -235.445 277.605 -235.115 ;
        RECT 277.275 -236.805 277.605 -236.475 ;
        RECT 277.275 -238.165 277.605 -237.835 ;
        RECT 277.275 -243.81 277.605 -242.68 ;
        RECT 277.28 -243.925 277.6 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 246.76 278.965 247.89 ;
        RECT 278.635 241.915 278.965 242.245 ;
        RECT 278.635 240.555 278.965 240.885 ;
        RECT 278.635 239.195 278.965 239.525 ;
        RECT 278.635 237.835 278.965 238.165 ;
        RECT 278.64 237.16 278.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 -1.525 278.965 -1.195 ;
        RECT 278.635 -2.885 278.965 -2.555 ;
        RECT 278.64 -3.56 278.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 246.76 280.325 247.89 ;
        RECT 279.995 241.915 280.325 242.245 ;
        RECT 279.995 240.555 280.325 240.885 ;
        RECT 279.995 239.195 280.325 239.525 ;
        RECT 279.995 237.835 280.325 238.165 ;
        RECT 280 237.16 280.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 -1.525 280.325 -1.195 ;
        RECT 279.995 -2.885 280.325 -2.555 ;
        RECT 280 -3.56 280.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 -122.565 280.325 -122.235 ;
        RECT 279.995 -123.925 280.325 -123.595 ;
        RECT 279.995 -125.285 280.325 -124.955 ;
        RECT 279.995 -126.645 280.325 -126.315 ;
        RECT 279.995 -128.005 280.325 -127.675 ;
        RECT 279.995 -129.365 280.325 -129.035 ;
        RECT 279.995 -130.725 280.325 -130.395 ;
        RECT 279.995 -132.085 280.325 -131.755 ;
        RECT 279.995 -133.445 280.325 -133.115 ;
        RECT 279.995 -134.805 280.325 -134.475 ;
        RECT 279.995 -136.165 280.325 -135.835 ;
        RECT 279.995 -137.525 280.325 -137.195 ;
        RECT 279.995 -138.885 280.325 -138.555 ;
        RECT 279.995 -140.245 280.325 -139.915 ;
        RECT 279.995 -141.605 280.325 -141.275 ;
        RECT 279.995 -142.965 280.325 -142.635 ;
        RECT 279.995 -144.325 280.325 -143.995 ;
        RECT 279.995 -145.685 280.325 -145.355 ;
        RECT 279.995 -147.045 280.325 -146.715 ;
        RECT 279.995 -148.405 280.325 -148.075 ;
        RECT 279.995 -149.765 280.325 -149.435 ;
        RECT 279.995 -151.125 280.325 -150.795 ;
        RECT 279.995 -152.485 280.325 -152.155 ;
        RECT 279.995 -153.845 280.325 -153.515 ;
        RECT 279.995 -155.205 280.325 -154.875 ;
        RECT 279.995 -156.565 280.325 -156.235 ;
        RECT 279.995 -157.925 280.325 -157.595 ;
        RECT 279.995 -159.285 280.325 -158.955 ;
        RECT 279.995 -160.645 280.325 -160.315 ;
        RECT 279.995 -162.005 280.325 -161.675 ;
        RECT 279.995 -163.365 280.325 -163.035 ;
        RECT 279.995 -164.725 280.325 -164.395 ;
        RECT 279.995 -166.085 280.325 -165.755 ;
        RECT 279.995 -167.445 280.325 -167.115 ;
        RECT 279.995 -168.805 280.325 -168.475 ;
        RECT 279.995 -170.165 280.325 -169.835 ;
        RECT 279.995 -171.525 280.325 -171.195 ;
        RECT 279.995 -172.885 280.325 -172.555 ;
        RECT 279.995 -174.245 280.325 -173.915 ;
        RECT 279.995 -175.605 280.325 -175.275 ;
        RECT 279.995 -176.965 280.325 -176.635 ;
        RECT 279.995 -178.325 280.325 -177.995 ;
        RECT 279.995 -179.685 280.325 -179.355 ;
        RECT 279.995 -181.045 280.325 -180.715 ;
        RECT 279.995 -182.405 280.325 -182.075 ;
        RECT 279.995 -183.765 280.325 -183.435 ;
        RECT 279.995 -185.125 280.325 -184.795 ;
        RECT 279.995 -186.485 280.325 -186.155 ;
        RECT 279.995 -187.845 280.325 -187.515 ;
        RECT 279.995 -189.205 280.325 -188.875 ;
        RECT 279.995 -190.565 280.325 -190.235 ;
        RECT 279.995 -191.925 280.325 -191.595 ;
        RECT 279.995 -193.285 280.325 -192.955 ;
        RECT 279.995 -194.645 280.325 -194.315 ;
        RECT 279.995 -196.005 280.325 -195.675 ;
        RECT 279.995 -197.365 280.325 -197.035 ;
        RECT 279.995 -198.725 280.325 -198.395 ;
        RECT 279.995 -200.085 280.325 -199.755 ;
        RECT 279.995 -201.445 280.325 -201.115 ;
        RECT 279.995 -202.805 280.325 -202.475 ;
        RECT 279.995 -204.165 280.325 -203.835 ;
        RECT 279.995 -205.525 280.325 -205.195 ;
        RECT 279.995 -206.885 280.325 -206.555 ;
        RECT 279.995 -208.245 280.325 -207.915 ;
        RECT 279.995 -209.605 280.325 -209.275 ;
        RECT 279.995 -210.965 280.325 -210.635 ;
        RECT 279.995 -212.325 280.325 -211.995 ;
        RECT 279.995 -213.685 280.325 -213.355 ;
        RECT 279.995 -215.045 280.325 -214.715 ;
        RECT 279.995 -216.405 280.325 -216.075 ;
        RECT 279.995 -217.765 280.325 -217.435 ;
        RECT 279.995 -219.125 280.325 -218.795 ;
        RECT 279.995 -220.485 280.325 -220.155 ;
        RECT 279.995 -221.845 280.325 -221.515 ;
        RECT 279.995 -223.205 280.325 -222.875 ;
        RECT 279.995 -224.565 280.325 -224.235 ;
        RECT 279.995 -225.925 280.325 -225.595 ;
        RECT 279.995 -227.285 280.325 -226.955 ;
        RECT 279.995 -228.645 280.325 -228.315 ;
        RECT 279.995 -230.005 280.325 -229.675 ;
        RECT 279.995 -231.365 280.325 -231.035 ;
        RECT 279.995 -232.725 280.325 -232.395 ;
        RECT 279.995 -234.085 280.325 -233.755 ;
        RECT 279.995 -235.445 280.325 -235.115 ;
        RECT 279.995 -236.805 280.325 -236.475 ;
        RECT 279.995 -238.165 280.325 -237.835 ;
        RECT 279.995 -243.81 280.325 -242.68 ;
        RECT 280 -243.925 280.32 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 246.76 281.685 247.89 ;
        RECT 281.355 241.915 281.685 242.245 ;
        RECT 281.355 240.555 281.685 240.885 ;
        RECT 281.355 239.195 281.685 239.525 ;
        RECT 281.355 237.835 281.685 238.165 ;
        RECT 281.36 237.16 281.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 -1.525 281.685 -1.195 ;
        RECT 281.355 -2.885 281.685 -2.555 ;
        RECT 281.36 -3.56 281.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 -238.165 281.685 -237.835 ;
        RECT 281.355 -243.81 281.685 -242.68 ;
        RECT 281.36 -243.925 281.68 -122.235 ;
        RECT 281.355 -122.565 281.685 -122.235 ;
        RECT 281.355 -123.925 281.685 -123.595 ;
        RECT 281.355 -125.285 281.685 -124.955 ;
        RECT 281.355 -126.645 281.685 -126.315 ;
        RECT 281.355 -128.005 281.685 -127.675 ;
        RECT 281.355 -129.365 281.685 -129.035 ;
        RECT 281.355 -130.725 281.685 -130.395 ;
        RECT 281.355 -132.085 281.685 -131.755 ;
        RECT 281.355 -133.445 281.685 -133.115 ;
        RECT 281.355 -134.805 281.685 -134.475 ;
        RECT 281.355 -136.165 281.685 -135.835 ;
        RECT 281.355 -137.525 281.685 -137.195 ;
        RECT 281.355 -138.885 281.685 -138.555 ;
        RECT 281.355 -140.245 281.685 -139.915 ;
        RECT 281.355 -141.605 281.685 -141.275 ;
        RECT 281.355 -142.965 281.685 -142.635 ;
        RECT 281.355 -144.325 281.685 -143.995 ;
        RECT 281.355 -145.685 281.685 -145.355 ;
        RECT 281.355 -147.045 281.685 -146.715 ;
        RECT 281.355 -148.405 281.685 -148.075 ;
        RECT 281.355 -149.765 281.685 -149.435 ;
        RECT 281.355 -151.125 281.685 -150.795 ;
        RECT 281.355 -152.485 281.685 -152.155 ;
        RECT 281.355 -153.845 281.685 -153.515 ;
        RECT 281.355 -155.205 281.685 -154.875 ;
        RECT 281.355 -156.565 281.685 -156.235 ;
        RECT 281.355 -157.925 281.685 -157.595 ;
        RECT 281.355 -159.285 281.685 -158.955 ;
        RECT 281.355 -160.645 281.685 -160.315 ;
        RECT 281.355 -162.005 281.685 -161.675 ;
        RECT 281.355 -163.365 281.685 -163.035 ;
        RECT 281.355 -164.725 281.685 -164.395 ;
        RECT 281.355 -166.085 281.685 -165.755 ;
        RECT 281.355 -167.445 281.685 -167.115 ;
        RECT 281.355 -168.805 281.685 -168.475 ;
        RECT 281.355 -170.165 281.685 -169.835 ;
        RECT 281.355 -171.525 281.685 -171.195 ;
        RECT 281.355 -172.885 281.685 -172.555 ;
        RECT 281.355 -174.245 281.685 -173.915 ;
        RECT 281.355 -175.605 281.685 -175.275 ;
        RECT 281.355 -176.965 281.685 -176.635 ;
        RECT 281.355 -178.325 281.685 -177.995 ;
        RECT 281.355 -179.685 281.685 -179.355 ;
        RECT 281.355 -181.045 281.685 -180.715 ;
        RECT 281.355 -182.405 281.685 -182.075 ;
        RECT 281.355 -183.765 281.685 -183.435 ;
        RECT 281.355 -185.125 281.685 -184.795 ;
        RECT 281.355 -186.485 281.685 -186.155 ;
        RECT 281.355 -187.845 281.685 -187.515 ;
        RECT 281.355 -189.205 281.685 -188.875 ;
        RECT 281.355 -190.565 281.685 -190.235 ;
        RECT 281.355 -191.925 281.685 -191.595 ;
        RECT 281.355 -193.285 281.685 -192.955 ;
        RECT 281.355 -194.645 281.685 -194.315 ;
        RECT 281.355 -196.005 281.685 -195.675 ;
        RECT 281.355 -197.365 281.685 -197.035 ;
        RECT 281.355 -198.725 281.685 -198.395 ;
        RECT 281.355 -200.085 281.685 -199.755 ;
        RECT 281.355 -201.445 281.685 -201.115 ;
        RECT 281.355 -202.805 281.685 -202.475 ;
        RECT 281.355 -204.165 281.685 -203.835 ;
        RECT 281.355 -205.525 281.685 -205.195 ;
        RECT 281.355 -206.885 281.685 -206.555 ;
        RECT 281.355 -208.245 281.685 -207.915 ;
        RECT 281.355 -209.605 281.685 -209.275 ;
        RECT 281.355 -210.965 281.685 -210.635 ;
        RECT 281.355 -212.325 281.685 -211.995 ;
        RECT 281.355 -213.685 281.685 -213.355 ;
        RECT 281.355 -215.045 281.685 -214.715 ;
        RECT 281.355 -216.405 281.685 -216.075 ;
        RECT 281.355 -217.765 281.685 -217.435 ;
        RECT 281.355 -219.125 281.685 -218.795 ;
        RECT 281.355 -220.485 281.685 -220.155 ;
        RECT 281.355 -221.845 281.685 -221.515 ;
        RECT 281.355 -223.205 281.685 -222.875 ;
        RECT 281.355 -224.565 281.685 -224.235 ;
        RECT 281.355 -225.925 281.685 -225.595 ;
        RECT 281.355 -227.285 281.685 -226.955 ;
        RECT 281.355 -228.645 281.685 -228.315 ;
        RECT 281.355 -230.005 281.685 -229.675 ;
        RECT 281.355 -231.365 281.685 -231.035 ;
        RECT 281.355 -232.725 281.685 -232.395 ;
        RECT 281.355 -234.085 281.685 -233.755 ;
        RECT 281.355 -235.445 281.685 -235.115 ;
        RECT 281.355 -236.805 281.685 -236.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.46 -125.535 242.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.275 246.76 243.605 247.89 ;
        RECT 243.275 241.915 243.605 242.245 ;
        RECT 243.275 240.555 243.605 240.885 ;
        RECT 243.275 239.195 243.605 239.525 ;
        RECT 243.275 237.835 243.605 238.165 ;
        RECT 243.28 237.16 243.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 246.76 244.965 247.89 ;
        RECT 244.635 241.915 244.965 242.245 ;
        RECT 244.635 240.555 244.965 240.885 ;
        RECT 244.635 239.195 244.965 239.525 ;
        RECT 244.635 237.835 244.965 238.165 ;
        RECT 244.64 237.16 244.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 -1.525 244.965 -1.195 ;
        RECT 244.635 -2.885 244.965 -2.555 ;
        RECT 244.64 -3.56 244.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 -122.565 244.965 -122.235 ;
        RECT 244.635 -123.925 244.965 -123.595 ;
        RECT 244.635 -125.285 244.965 -124.955 ;
        RECT 244.635 -126.645 244.965 -126.315 ;
        RECT 244.635 -128.005 244.965 -127.675 ;
        RECT 244.635 -129.365 244.965 -129.035 ;
        RECT 244.635 -130.725 244.965 -130.395 ;
        RECT 244.635 -132.085 244.965 -131.755 ;
        RECT 244.635 -133.445 244.965 -133.115 ;
        RECT 244.635 -134.805 244.965 -134.475 ;
        RECT 244.635 -136.165 244.965 -135.835 ;
        RECT 244.635 -137.525 244.965 -137.195 ;
        RECT 244.635 -138.885 244.965 -138.555 ;
        RECT 244.635 -140.245 244.965 -139.915 ;
        RECT 244.635 -141.605 244.965 -141.275 ;
        RECT 244.635 -142.965 244.965 -142.635 ;
        RECT 244.635 -144.325 244.965 -143.995 ;
        RECT 244.635 -145.685 244.965 -145.355 ;
        RECT 244.635 -147.045 244.965 -146.715 ;
        RECT 244.635 -148.405 244.965 -148.075 ;
        RECT 244.635 -149.765 244.965 -149.435 ;
        RECT 244.635 -151.125 244.965 -150.795 ;
        RECT 244.635 -152.485 244.965 -152.155 ;
        RECT 244.635 -153.845 244.965 -153.515 ;
        RECT 244.635 -155.205 244.965 -154.875 ;
        RECT 244.635 -156.565 244.965 -156.235 ;
        RECT 244.635 -157.925 244.965 -157.595 ;
        RECT 244.635 -159.285 244.965 -158.955 ;
        RECT 244.635 -160.645 244.965 -160.315 ;
        RECT 244.635 -162.005 244.965 -161.675 ;
        RECT 244.635 -163.365 244.965 -163.035 ;
        RECT 244.635 -164.725 244.965 -164.395 ;
        RECT 244.635 -166.085 244.965 -165.755 ;
        RECT 244.635 -167.445 244.965 -167.115 ;
        RECT 244.635 -168.805 244.965 -168.475 ;
        RECT 244.635 -170.165 244.965 -169.835 ;
        RECT 244.635 -171.525 244.965 -171.195 ;
        RECT 244.635 -172.885 244.965 -172.555 ;
        RECT 244.635 -174.245 244.965 -173.915 ;
        RECT 244.635 -175.605 244.965 -175.275 ;
        RECT 244.635 -176.965 244.965 -176.635 ;
        RECT 244.635 -178.325 244.965 -177.995 ;
        RECT 244.635 -179.685 244.965 -179.355 ;
        RECT 244.635 -181.045 244.965 -180.715 ;
        RECT 244.635 -182.405 244.965 -182.075 ;
        RECT 244.635 -183.765 244.965 -183.435 ;
        RECT 244.635 -185.125 244.965 -184.795 ;
        RECT 244.635 -186.485 244.965 -186.155 ;
        RECT 244.635 -187.845 244.965 -187.515 ;
        RECT 244.635 -189.205 244.965 -188.875 ;
        RECT 244.635 -190.565 244.965 -190.235 ;
        RECT 244.635 -191.925 244.965 -191.595 ;
        RECT 244.635 -193.285 244.965 -192.955 ;
        RECT 244.635 -194.645 244.965 -194.315 ;
        RECT 244.635 -196.005 244.965 -195.675 ;
        RECT 244.635 -197.365 244.965 -197.035 ;
        RECT 244.635 -198.725 244.965 -198.395 ;
        RECT 244.635 -200.085 244.965 -199.755 ;
        RECT 244.635 -201.445 244.965 -201.115 ;
        RECT 244.635 -202.805 244.965 -202.475 ;
        RECT 244.635 -204.165 244.965 -203.835 ;
        RECT 244.635 -205.525 244.965 -205.195 ;
        RECT 244.635 -206.885 244.965 -206.555 ;
        RECT 244.635 -208.245 244.965 -207.915 ;
        RECT 244.635 -209.605 244.965 -209.275 ;
        RECT 244.635 -210.965 244.965 -210.635 ;
        RECT 244.635 -212.325 244.965 -211.995 ;
        RECT 244.635 -213.685 244.965 -213.355 ;
        RECT 244.635 -215.045 244.965 -214.715 ;
        RECT 244.635 -216.405 244.965 -216.075 ;
        RECT 244.635 -217.765 244.965 -217.435 ;
        RECT 244.635 -219.125 244.965 -218.795 ;
        RECT 244.635 -220.485 244.965 -220.155 ;
        RECT 244.635 -221.845 244.965 -221.515 ;
        RECT 244.635 -223.205 244.965 -222.875 ;
        RECT 244.635 -224.565 244.965 -224.235 ;
        RECT 244.635 -225.925 244.965 -225.595 ;
        RECT 244.635 -227.285 244.965 -226.955 ;
        RECT 244.635 -228.645 244.965 -228.315 ;
        RECT 244.635 -230.005 244.965 -229.675 ;
        RECT 244.635 -231.365 244.965 -231.035 ;
        RECT 244.635 -232.725 244.965 -232.395 ;
        RECT 244.635 -234.085 244.965 -233.755 ;
        RECT 244.635 -235.445 244.965 -235.115 ;
        RECT 244.635 -236.805 244.965 -236.475 ;
        RECT 244.635 -238.165 244.965 -237.835 ;
        RECT 244.635 -243.81 244.965 -242.68 ;
        RECT 244.64 -243.925 244.96 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 246.76 246.325 247.89 ;
        RECT 245.995 241.915 246.325 242.245 ;
        RECT 245.995 240.555 246.325 240.885 ;
        RECT 245.995 239.195 246.325 239.525 ;
        RECT 245.995 237.835 246.325 238.165 ;
        RECT 246 237.16 246.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 -1.525 246.325 -1.195 ;
        RECT 245.995 -2.885 246.325 -2.555 ;
        RECT 246 -3.56 246.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 246.76 247.685 247.89 ;
        RECT 247.355 241.915 247.685 242.245 ;
        RECT 247.355 240.555 247.685 240.885 ;
        RECT 247.355 239.195 247.685 239.525 ;
        RECT 247.355 237.835 247.685 238.165 ;
        RECT 247.36 237.16 247.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 -1.525 247.685 -1.195 ;
        RECT 247.355 -2.885 247.685 -2.555 ;
        RECT 247.36 -3.56 247.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 -122.565 247.685 -122.235 ;
        RECT 247.355 -123.925 247.685 -123.595 ;
        RECT 247.355 -125.285 247.685 -124.955 ;
        RECT 247.355 -126.645 247.685 -126.315 ;
        RECT 247.355 -128.005 247.685 -127.675 ;
        RECT 247.355 -129.365 247.685 -129.035 ;
        RECT 247.355 -130.725 247.685 -130.395 ;
        RECT 247.355 -132.085 247.685 -131.755 ;
        RECT 247.355 -133.445 247.685 -133.115 ;
        RECT 247.355 -134.805 247.685 -134.475 ;
        RECT 247.355 -136.165 247.685 -135.835 ;
        RECT 247.355 -137.525 247.685 -137.195 ;
        RECT 247.355 -138.885 247.685 -138.555 ;
        RECT 247.355 -140.245 247.685 -139.915 ;
        RECT 247.355 -141.605 247.685 -141.275 ;
        RECT 247.355 -142.965 247.685 -142.635 ;
        RECT 247.355 -144.325 247.685 -143.995 ;
        RECT 247.355 -145.685 247.685 -145.355 ;
        RECT 247.355 -147.045 247.685 -146.715 ;
        RECT 247.355 -148.405 247.685 -148.075 ;
        RECT 247.355 -149.765 247.685 -149.435 ;
        RECT 247.355 -151.125 247.685 -150.795 ;
        RECT 247.355 -152.485 247.685 -152.155 ;
        RECT 247.355 -153.845 247.685 -153.515 ;
        RECT 247.355 -155.205 247.685 -154.875 ;
        RECT 247.355 -156.565 247.685 -156.235 ;
        RECT 247.355 -157.925 247.685 -157.595 ;
        RECT 247.355 -159.285 247.685 -158.955 ;
        RECT 247.355 -160.645 247.685 -160.315 ;
        RECT 247.355 -162.005 247.685 -161.675 ;
        RECT 247.355 -163.365 247.685 -163.035 ;
        RECT 247.355 -164.725 247.685 -164.395 ;
        RECT 247.355 -166.085 247.685 -165.755 ;
        RECT 247.355 -167.445 247.685 -167.115 ;
        RECT 247.355 -168.805 247.685 -168.475 ;
        RECT 247.355 -170.165 247.685 -169.835 ;
        RECT 247.355 -171.525 247.685 -171.195 ;
        RECT 247.355 -172.885 247.685 -172.555 ;
        RECT 247.355 -174.245 247.685 -173.915 ;
        RECT 247.355 -175.605 247.685 -175.275 ;
        RECT 247.355 -176.965 247.685 -176.635 ;
        RECT 247.355 -178.325 247.685 -177.995 ;
        RECT 247.355 -179.685 247.685 -179.355 ;
        RECT 247.355 -181.045 247.685 -180.715 ;
        RECT 247.355 -182.405 247.685 -182.075 ;
        RECT 247.355 -183.765 247.685 -183.435 ;
        RECT 247.355 -185.125 247.685 -184.795 ;
        RECT 247.355 -186.485 247.685 -186.155 ;
        RECT 247.355 -187.845 247.685 -187.515 ;
        RECT 247.355 -189.205 247.685 -188.875 ;
        RECT 247.355 -190.565 247.685 -190.235 ;
        RECT 247.355 -191.925 247.685 -191.595 ;
        RECT 247.355 -193.285 247.685 -192.955 ;
        RECT 247.355 -194.645 247.685 -194.315 ;
        RECT 247.355 -196.005 247.685 -195.675 ;
        RECT 247.355 -197.365 247.685 -197.035 ;
        RECT 247.355 -198.725 247.685 -198.395 ;
        RECT 247.355 -200.085 247.685 -199.755 ;
        RECT 247.355 -201.445 247.685 -201.115 ;
        RECT 247.355 -202.805 247.685 -202.475 ;
        RECT 247.355 -204.165 247.685 -203.835 ;
        RECT 247.355 -205.525 247.685 -205.195 ;
        RECT 247.355 -206.885 247.685 -206.555 ;
        RECT 247.355 -208.245 247.685 -207.915 ;
        RECT 247.355 -209.605 247.685 -209.275 ;
        RECT 247.355 -210.965 247.685 -210.635 ;
        RECT 247.355 -212.325 247.685 -211.995 ;
        RECT 247.355 -213.685 247.685 -213.355 ;
        RECT 247.355 -215.045 247.685 -214.715 ;
        RECT 247.355 -216.405 247.685 -216.075 ;
        RECT 247.355 -217.765 247.685 -217.435 ;
        RECT 247.355 -219.125 247.685 -218.795 ;
        RECT 247.355 -220.485 247.685 -220.155 ;
        RECT 247.355 -221.845 247.685 -221.515 ;
        RECT 247.355 -223.205 247.685 -222.875 ;
        RECT 247.355 -224.565 247.685 -224.235 ;
        RECT 247.355 -225.925 247.685 -225.595 ;
        RECT 247.355 -227.285 247.685 -226.955 ;
        RECT 247.355 -228.645 247.685 -228.315 ;
        RECT 247.355 -230.005 247.685 -229.675 ;
        RECT 247.355 -231.365 247.685 -231.035 ;
        RECT 247.355 -232.725 247.685 -232.395 ;
        RECT 247.355 -234.085 247.685 -233.755 ;
        RECT 247.355 -235.445 247.685 -235.115 ;
        RECT 247.355 -236.805 247.685 -236.475 ;
        RECT 247.355 -238.165 247.685 -237.835 ;
        RECT 247.355 -243.81 247.685 -242.68 ;
        RECT 247.36 -243.925 247.68 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 246.76 249.045 247.89 ;
        RECT 248.715 241.915 249.045 242.245 ;
        RECT 248.715 240.555 249.045 240.885 ;
        RECT 248.715 239.195 249.045 239.525 ;
        RECT 248.715 237.835 249.045 238.165 ;
        RECT 248.72 237.16 249.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 -1.525 249.045 -1.195 ;
        RECT 248.715 -2.885 249.045 -2.555 ;
        RECT 248.72 -3.56 249.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 -122.565 249.045 -122.235 ;
        RECT 248.715 -123.925 249.045 -123.595 ;
        RECT 248.715 -125.285 249.045 -124.955 ;
        RECT 248.715 -126.645 249.045 -126.315 ;
        RECT 248.715 -128.005 249.045 -127.675 ;
        RECT 248.715 -129.365 249.045 -129.035 ;
        RECT 248.715 -130.725 249.045 -130.395 ;
        RECT 248.715 -132.085 249.045 -131.755 ;
        RECT 248.715 -133.445 249.045 -133.115 ;
        RECT 248.715 -134.805 249.045 -134.475 ;
        RECT 248.715 -136.165 249.045 -135.835 ;
        RECT 248.715 -137.525 249.045 -137.195 ;
        RECT 248.715 -138.885 249.045 -138.555 ;
        RECT 248.715 -140.245 249.045 -139.915 ;
        RECT 248.715 -141.605 249.045 -141.275 ;
        RECT 248.715 -142.965 249.045 -142.635 ;
        RECT 248.715 -144.325 249.045 -143.995 ;
        RECT 248.715 -145.685 249.045 -145.355 ;
        RECT 248.715 -147.045 249.045 -146.715 ;
        RECT 248.715 -148.405 249.045 -148.075 ;
        RECT 248.715 -149.765 249.045 -149.435 ;
        RECT 248.715 -151.125 249.045 -150.795 ;
        RECT 248.715 -152.485 249.045 -152.155 ;
        RECT 248.715 -153.845 249.045 -153.515 ;
        RECT 248.715 -155.205 249.045 -154.875 ;
        RECT 248.715 -156.565 249.045 -156.235 ;
        RECT 248.715 -157.925 249.045 -157.595 ;
        RECT 248.715 -159.285 249.045 -158.955 ;
        RECT 248.715 -160.645 249.045 -160.315 ;
        RECT 248.715 -162.005 249.045 -161.675 ;
        RECT 248.715 -163.365 249.045 -163.035 ;
        RECT 248.715 -164.725 249.045 -164.395 ;
        RECT 248.715 -166.085 249.045 -165.755 ;
        RECT 248.715 -167.445 249.045 -167.115 ;
        RECT 248.715 -168.805 249.045 -168.475 ;
        RECT 248.715 -170.165 249.045 -169.835 ;
        RECT 248.715 -171.525 249.045 -171.195 ;
        RECT 248.715 -172.885 249.045 -172.555 ;
        RECT 248.715 -174.245 249.045 -173.915 ;
        RECT 248.715 -175.605 249.045 -175.275 ;
        RECT 248.715 -176.965 249.045 -176.635 ;
        RECT 248.715 -178.325 249.045 -177.995 ;
        RECT 248.715 -179.685 249.045 -179.355 ;
        RECT 248.715 -181.045 249.045 -180.715 ;
        RECT 248.715 -182.405 249.045 -182.075 ;
        RECT 248.715 -183.765 249.045 -183.435 ;
        RECT 248.715 -185.125 249.045 -184.795 ;
        RECT 248.715 -186.485 249.045 -186.155 ;
        RECT 248.715 -187.845 249.045 -187.515 ;
        RECT 248.715 -189.205 249.045 -188.875 ;
        RECT 248.715 -190.565 249.045 -190.235 ;
        RECT 248.715 -191.925 249.045 -191.595 ;
        RECT 248.715 -193.285 249.045 -192.955 ;
        RECT 248.715 -194.645 249.045 -194.315 ;
        RECT 248.715 -196.005 249.045 -195.675 ;
        RECT 248.715 -197.365 249.045 -197.035 ;
        RECT 248.715 -198.725 249.045 -198.395 ;
        RECT 248.715 -200.085 249.045 -199.755 ;
        RECT 248.715 -201.445 249.045 -201.115 ;
        RECT 248.715 -202.805 249.045 -202.475 ;
        RECT 248.715 -204.165 249.045 -203.835 ;
        RECT 248.715 -205.525 249.045 -205.195 ;
        RECT 248.715 -206.885 249.045 -206.555 ;
        RECT 248.715 -208.245 249.045 -207.915 ;
        RECT 248.715 -209.605 249.045 -209.275 ;
        RECT 248.715 -210.965 249.045 -210.635 ;
        RECT 248.715 -212.325 249.045 -211.995 ;
        RECT 248.715 -213.685 249.045 -213.355 ;
        RECT 248.715 -215.045 249.045 -214.715 ;
        RECT 248.715 -216.405 249.045 -216.075 ;
        RECT 248.715 -217.765 249.045 -217.435 ;
        RECT 248.715 -219.125 249.045 -218.795 ;
        RECT 248.715 -220.485 249.045 -220.155 ;
        RECT 248.715 -221.845 249.045 -221.515 ;
        RECT 248.715 -223.205 249.045 -222.875 ;
        RECT 248.715 -224.565 249.045 -224.235 ;
        RECT 248.715 -225.925 249.045 -225.595 ;
        RECT 248.715 -227.285 249.045 -226.955 ;
        RECT 248.715 -228.645 249.045 -228.315 ;
        RECT 248.715 -230.005 249.045 -229.675 ;
        RECT 248.715 -231.365 249.045 -231.035 ;
        RECT 248.715 -232.725 249.045 -232.395 ;
        RECT 248.715 -234.085 249.045 -233.755 ;
        RECT 248.715 -235.445 249.045 -235.115 ;
        RECT 248.715 -236.805 249.045 -236.475 ;
        RECT 248.715 -238.165 249.045 -237.835 ;
        RECT 248.715 -243.81 249.045 -242.68 ;
        RECT 248.72 -243.925 249.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 246.76 250.405 247.89 ;
        RECT 250.075 241.915 250.405 242.245 ;
        RECT 250.075 240.555 250.405 240.885 ;
        RECT 250.075 239.195 250.405 239.525 ;
        RECT 250.075 237.835 250.405 238.165 ;
        RECT 250.08 237.16 250.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 -1.525 250.405 -1.195 ;
        RECT 250.075 -2.885 250.405 -2.555 ;
        RECT 250.08 -3.56 250.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 -122.565 250.405 -122.235 ;
        RECT 250.075 -123.925 250.405 -123.595 ;
        RECT 250.075 -125.285 250.405 -124.955 ;
        RECT 250.075 -126.645 250.405 -126.315 ;
        RECT 250.075 -128.005 250.405 -127.675 ;
        RECT 250.075 -129.365 250.405 -129.035 ;
        RECT 250.075 -130.725 250.405 -130.395 ;
        RECT 250.075 -132.085 250.405 -131.755 ;
        RECT 250.075 -133.445 250.405 -133.115 ;
        RECT 250.075 -134.805 250.405 -134.475 ;
        RECT 250.075 -136.165 250.405 -135.835 ;
        RECT 250.075 -137.525 250.405 -137.195 ;
        RECT 250.075 -138.885 250.405 -138.555 ;
        RECT 250.075 -140.245 250.405 -139.915 ;
        RECT 250.075 -141.605 250.405 -141.275 ;
        RECT 250.075 -142.965 250.405 -142.635 ;
        RECT 250.075 -144.325 250.405 -143.995 ;
        RECT 250.075 -145.685 250.405 -145.355 ;
        RECT 250.075 -147.045 250.405 -146.715 ;
        RECT 250.075 -148.405 250.405 -148.075 ;
        RECT 250.075 -149.765 250.405 -149.435 ;
        RECT 250.075 -151.125 250.405 -150.795 ;
        RECT 250.075 -152.485 250.405 -152.155 ;
        RECT 250.075 -153.845 250.405 -153.515 ;
        RECT 250.075 -155.205 250.405 -154.875 ;
        RECT 250.075 -156.565 250.405 -156.235 ;
        RECT 250.075 -157.925 250.405 -157.595 ;
        RECT 250.075 -159.285 250.405 -158.955 ;
        RECT 250.075 -160.645 250.405 -160.315 ;
        RECT 250.075 -162.005 250.405 -161.675 ;
        RECT 250.075 -163.365 250.405 -163.035 ;
        RECT 250.075 -164.725 250.405 -164.395 ;
        RECT 250.075 -166.085 250.405 -165.755 ;
        RECT 250.075 -167.445 250.405 -167.115 ;
        RECT 250.075 -168.805 250.405 -168.475 ;
        RECT 250.075 -170.165 250.405 -169.835 ;
        RECT 250.075 -171.525 250.405 -171.195 ;
        RECT 250.075 -172.885 250.405 -172.555 ;
        RECT 250.075 -174.245 250.405 -173.915 ;
        RECT 250.075 -175.605 250.405 -175.275 ;
        RECT 250.075 -176.965 250.405 -176.635 ;
        RECT 250.075 -178.325 250.405 -177.995 ;
        RECT 250.075 -179.685 250.405 -179.355 ;
        RECT 250.075 -181.045 250.405 -180.715 ;
        RECT 250.075 -182.405 250.405 -182.075 ;
        RECT 250.075 -183.765 250.405 -183.435 ;
        RECT 250.075 -185.125 250.405 -184.795 ;
        RECT 250.075 -186.485 250.405 -186.155 ;
        RECT 250.075 -187.845 250.405 -187.515 ;
        RECT 250.075 -189.205 250.405 -188.875 ;
        RECT 250.075 -190.565 250.405 -190.235 ;
        RECT 250.075 -191.925 250.405 -191.595 ;
        RECT 250.075 -193.285 250.405 -192.955 ;
        RECT 250.075 -194.645 250.405 -194.315 ;
        RECT 250.075 -196.005 250.405 -195.675 ;
        RECT 250.075 -197.365 250.405 -197.035 ;
        RECT 250.075 -198.725 250.405 -198.395 ;
        RECT 250.075 -200.085 250.405 -199.755 ;
        RECT 250.075 -201.445 250.405 -201.115 ;
        RECT 250.075 -202.805 250.405 -202.475 ;
        RECT 250.075 -204.165 250.405 -203.835 ;
        RECT 250.075 -205.525 250.405 -205.195 ;
        RECT 250.075 -206.885 250.405 -206.555 ;
        RECT 250.075 -208.245 250.405 -207.915 ;
        RECT 250.075 -209.605 250.405 -209.275 ;
        RECT 250.075 -210.965 250.405 -210.635 ;
        RECT 250.075 -212.325 250.405 -211.995 ;
        RECT 250.075 -213.685 250.405 -213.355 ;
        RECT 250.075 -215.045 250.405 -214.715 ;
        RECT 250.075 -216.405 250.405 -216.075 ;
        RECT 250.075 -217.765 250.405 -217.435 ;
        RECT 250.075 -219.125 250.405 -218.795 ;
        RECT 250.075 -220.485 250.405 -220.155 ;
        RECT 250.075 -221.845 250.405 -221.515 ;
        RECT 250.075 -223.205 250.405 -222.875 ;
        RECT 250.075 -224.565 250.405 -224.235 ;
        RECT 250.075 -225.925 250.405 -225.595 ;
        RECT 250.075 -227.285 250.405 -226.955 ;
        RECT 250.075 -228.645 250.405 -228.315 ;
        RECT 250.075 -230.005 250.405 -229.675 ;
        RECT 250.075 -231.365 250.405 -231.035 ;
        RECT 250.075 -232.725 250.405 -232.395 ;
        RECT 250.075 -234.085 250.405 -233.755 ;
        RECT 250.075 -235.445 250.405 -235.115 ;
        RECT 250.075 -236.805 250.405 -236.475 ;
        RECT 250.075 -238.165 250.405 -237.835 ;
        RECT 250.075 -243.81 250.405 -242.68 ;
        RECT 250.08 -243.925 250.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 246.76 251.765 247.89 ;
        RECT 251.435 241.915 251.765 242.245 ;
        RECT 251.435 240.555 251.765 240.885 ;
        RECT 251.435 239.195 251.765 239.525 ;
        RECT 251.435 237.835 251.765 238.165 ;
        RECT 251.44 237.16 251.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 -1.525 251.765 -1.195 ;
        RECT 251.435 -2.885 251.765 -2.555 ;
        RECT 251.44 -3.56 251.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 -122.565 251.765 -122.235 ;
        RECT 251.435 -123.925 251.765 -123.595 ;
        RECT 251.435 -125.285 251.765 -124.955 ;
        RECT 251.435 -126.645 251.765 -126.315 ;
        RECT 251.435 -128.005 251.765 -127.675 ;
        RECT 251.435 -129.365 251.765 -129.035 ;
        RECT 251.435 -130.725 251.765 -130.395 ;
        RECT 251.435 -132.085 251.765 -131.755 ;
        RECT 251.435 -133.445 251.765 -133.115 ;
        RECT 251.435 -134.805 251.765 -134.475 ;
        RECT 251.435 -136.165 251.765 -135.835 ;
        RECT 251.435 -137.525 251.765 -137.195 ;
        RECT 251.435 -138.885 251.765 -138.555 ;
        RECT 251.435 -140.245 251.765 -139.915 ;
        RECT 251.435 -141.605 251.765 -141.275 ;
        RECT 251.435 -142.965 251.765 -142.635 ;
        RECT 251.435 -144.325 251.765 -143.995 ;
        RECT 251.435 -145.685 251.765 -145.355 ;
        RECT 251.435 -147.045 251.765 -146.715 ;
        RECT 251.435 -148.405 251.765 -148.075 ;
        RECT 251.435 -149.765 251.765 -149.435 ;
        RECT 251.435 -151.125 251.765 -150.795 ;
        RECT 251.435 -152.485 251.765 -152.155 ;
        RECT 251.435 -153.845 251.765 -153.515 ;
        RECT 251.435 -155.205 251.765 -154.875 ;
        RECT 251.435 -156.565 251.765 -156.235 ;
        RECT 251.435 -157.925 251.765 -157.595 ;
        RECT 251.435 -159.285 251.765 -158.955 ;
        RECT 251.435 -160.645 251.765 -160.315 ;
        RECT 251.435 -162.005 251.765 -161.675 ;
        RECT 251.435 -163.365 251.765 -163.035 ;
        RECT 251.435 -164.725 251.765 -164.395 ;
        RECT 251.435 -166.085 251.765 -165.755 ;
        RECT 251.435 -167.445 251.765 -167.115 ;
        RECT 251.435 -168.805 251.765 -168.475 ;
        RECT 251.435 -170.165 251.765 -169.835 ;
        RECT 251.435 -171.525 251.765 -171.195 ;
        RECT 251.435 -172.885 251.765 -172.555 ;
        RECT 251.435 -174.245 251.765 -173.915 ;
        RECT 251.435 -175.605 251.765 -175.275 ;
        RECT 251.435 -176.965 251.765 -176.635 ;
        RECT 251.435 -178.325 251.765 -177.995 ;
        RECT 251.435 -179.685 251.765 -179.355 ;
        RECT 251.435 -181.045 251.765 -180.715 ;
        RECT 251.435 -182.405 251.765 -182.075 ;
        RECT 251.435 -183.765 251.765 -183.435 ;
        RECT 251.435 -185.125 251.765 -184.795 ;
        RECT 251.435 -186.485 251.765 -186.155 ;
        RECT 251.435 -187.845 251.765 -187.515 ;
        RECT 251.435 -189.205 251.765 -188.875 ;
        RECT 251.435 -190.565 251.765 -190.235 ;
        RECT 251.435 -191.925 251.765 -191.595 ;
        RECT 251.435 -193.285 251.765 -192.955 ;
        RECT 251.435 -194.645 251.765 -194.315 ;
        RECT 251.435 -196.005 251.765 -195.675 ;
        RECT 251.435 -197.365 251.765 -197.035 ;
        RECT 251.435 -198.725 251.765 -198.395 ;
        RECT 251.435 -200.085 251.765 -199.755 ;
        RECT 251.435 -201.445 251.765 -201.115 ;
        RECT 251.435 -202.805 251.765 -202.475 ;
        RECT 251.435 -204.165 251.765 -203.835 ;
        RECT 251.435 -205.525 251.765 -205.195 ;
        RECT 251.435 -206.885 251.765 -206.555 ;
        RECT 251.435 -208.245 251.765 -207.915 ;
        RECT 251.435 -209.605 251.765 -209.275 ;
        RECT 251.435 -210.965 251.765 -210.635 ;
        RECT 251.435 -212.325 251.765 -211.995 ;
        RECT 251.435 -213.685 251.765 -213.355 ;
        RECT 251.435 -215.045 251.765 -214.715 ;
        RECT 251.435 -216.405 251.765 -216.075 ;
        RECT 251.435 -217.765 251.765 -217.435 ;
        RECT 251.435 -219.125 251.765 -218.795 ;
        RECT 251.435 -220.485 251.765 -220.155 ;
        RECT 251.435 -221.845 251.765 -221.515 ;
        RECT 251.435 -223.205 251.765 -222.875 ;
        RECT 251.435 -224.565 251.765 -224.235 ;
        RECT 251.435 -225.925 251.765 -225.595 ;
        RECT 251.435 -227.285 251.765 -226.955 ;
        RECT 251.435 -228.645 251.765 -228.315 ;
        RECT 251.435 -230.005 251.765 -229.675 ;
        RECT 251.435 -231.365 251.765 -231.035 ;
        RECT 251.435 -232.725 251.765 -232.395 ;
        RECT 251.435 -234.085 251.765 -233.755 ;
        RECT 251.435 -235.445 251.765 -235.115 ;
        RECT 251.435 -236.805 251.765 -236.475 ;
        RECT 251.435 -238.165 251.765 -237.835 ;
        RECT 251.435 -243.81 251.765 -242.68 ;
        RECT 251.44 -243.925 251.76 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 246.76 253.125 247.89 ;
        RECT 252.795 241.915 253.125 242.245 ;
        RECT 252.795 240.555 253.125 240.885 ;
        RECT 252.795 239.195 253.125 239.525 ;
        RECT 252.795 237.835 253.125 238.165 ;
        RECT 252.8 237.16 253.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 -126.645 253.125 -126.315 ;
        RECT 252.795 -128.005 253.125 -127.675 ;
        RECT 252.795 -129.365 253.125 -129.035 ;
        RECT 252.795 -130.725 253.125 -130.395 ;
        RECT 252.795 -132.085 253.125 -131.755 ;
        RECT 252.795 -133.445 253.125 -133.115 ;
        RECT 252.795 -134.805 253.125 -134.475 ;
        RECT 252.795 -136.165 253.125 -135.835 ;
        RECT 252.795 -137.525 253.125 -137.195 ;
        RECT 252.795 -138.885 253.125 -138.555 ;
        RECT 252.795 -140.245 253.125 -139.915 ;
        RECT 252.795 -141.605 253.125 -141.275 ;
        RECT 252.795 -142.965 253.125 -142.635 ;
        RECT 252.795 -144.325 253.125 -143.995 ;
        RECT 252.795 -145.685 253.125 -145.355 ;
        RECT 252.795 -147.045 253.125 -146.715 ;
        RECT 252.795 -148.405 253.125 -148.075 ;
        RECT 252.795 -149.765 253.125 -149.435 ;
        RECT 252.795 -151.125 253.125 -150.795 ;
        RECT 252.795 -152.485 253.125 -152.155 ;
        RECT 252.795 -153.845 253.125 -153.515 ;
        RECT 252.795 -155.205 253.125 -154.875 ;
        RECT 252.795 -156.565 253.125 -156.235 ;
        RECT 252.795 -157.925 253.125 -157.595 ;
        RECT 252.795 -159.285 253.125 -158.955 ;
        RECT 252.795 -160.645 253.125 -160.315 ;
        RECT 252.795 -162.005 253.125 -161.675 ;
        RECT 252.795 -163.365 253.125 -163.035 ;
        RECT 252.795 -164.725 253.125 -164.395 ;
        RECT 252.795 -166.085 253.125 -165.755 ;
        RECT 252.795 -167.445 253.125 -167.115 ;
        RECT 252.795 -168.805 253.125 -168.475 ;
        RECT 252.795 -170.165 253.125 -169.835 ;
        RECT 252.795 -171.525 253.125 -171.195 ;
        RECT 252.795 -172.885 253.125 -172.555 ;
        RECT 252.795 -174.245 253.125 -173.915 ;
        RECT 252.795 -175.605 253.125 -175.275 ;
        RECT 252.795 -176.965 253.125 -176.635 ;
        RECT 252.795 -178.325 253.125 -177.995 ;
        RECT 252.795 -179.685 253.125 -179.355 ;
        RECT 252.795 -181.045 253.125 -180.715 ;
        RECT 252.795 -182.405 253.125 -182.075 ;
        RECT 252.795 -183.765 253.125 -183.435 ;
        RECT 252.795 -185.125 253.125 -184.795 ;
        RECT 252.795 -186.485 253.125 -186.155 ;
        RECT 252.795 -187.845 253.125 -187.515 ;
        RECT 252.795 -189.205 253.125 -188.875 ;
        RECT 252.795 -190.565 253.125 -190.235 ;
        RECT 252.795 -191.925 253.125 -191.595 ;
        RECT 252.795 -193.285 253.125 -192.955 ;
        RECT 252.795 -194.645 253.125 -194.315 ;
        RECT 252.795 -196.005 253.125 -195.675 ;
        RECT 252.795 -197.365 253.125 -197.035 ;
        RECT 252.795 -198.725 253.125 -198.395 ;
        RECT 252.795 -200.085 253.125 -199.755 ;
        RECT 252.795 -201.445 253.125 -201.115 ;
        RECT 252.795 -202.805 253.125 -202.475 ;
        RECT 252.795 -204.165 253.125 -203.835 ;
        RECT 252.795 -205.525 253.125 -205.195 ;
        RECT 252.795 -206.885 253.125 -206.555 ;
        RECT 252.795 -208.245 253.125 -207.915 ;
        RECT 252.795 -209.605 253.125 -209.275 ;
        RECT 252.795 -210.965 253.125 -210.635 ;
        RECT 252.795 -212.325 253.125 -211.995 ;
        RECT 252.795 -213.685 253.125 -213.355 ;
        RECT 252.795 -215.045 253.125 -214.715 ;
        RECT 252.795 -216.405 253.125 -216.075 ;
        RECT 252.795 -217.765 253.125 -217.435 ;
        RECT 252.795 -219.125 253.125 -218.795 ;
        RECT 252.795 -220.485 253.125 -220.155 ;
        RECT 252.795 -221.845 253.125 -221.515 ;
        RECT 252.795 -223.205 253.125 -222.875 ;
        RECT 252.795 -224.565 253.125 -224.235 ;
        RECT 252.795 -225.925 253.125 -225.595 ;
        RECT 252.795 -227.285 253.125 -226.955 ;
        RECT 252.795 -228.645 253.125 -228.315 ;
        RECT 252.795 -230.005 253.125 -229.675 ;
        RECT 252.795 -231.365 253.125 -231.035 ;
        RECT 252.795 -232.725 253.125 -232.395 ;
        RECT 252.795 -234.085 253.125 -233.755 ;
        RECT 252.795 -235.445 253.125 -235.115 ;
        RECT 252.795 -236.805 253.125 -236.475 ;
        RECT 252.795 -238.165 253.125 -237.835 ;
        RECT 252.795 -243.81 253.125 -242.68 ;
        RECT 252.8 -243.925 253.12 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.36 -125.535 253.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.155 246.76 254.485 247.89 ;
        RECT 254.155 241.915 254.485 242.245 ;
        RECT 254.155 240.555 254.485 240.885 ;
        RECT 254.155 239.195 254.485 239.525 ;
        RECT 254.155 237.835 254.485 238.165 ;
        RECT 254.16 237.16 254.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 246.76 255.845 247.89 ;
        RECT 255.515 241.915 255.845 242.245 ;
        RECT 255.515 240.555 255.845 240.885 ;
        RECT 255.515 239.195 255.845 239.525 ;
        RECT 255.515 237.835 255.845 238.165 ;
        RECT 255.52 237.16 255.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 -1.525 255.845 -1.195 ;
        RECT 255.515 -2.885 255.845 -2.555 ;
        RECT 255.52 -3.56 255.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 -122.565 255.845 -122.235 ;
        RECT 255.515 -123.925 255.845 -123.595 ;
        RECT 255.515 -125.285 255.845 -124.955 ;
        RECT 255.515 -126.645 255.845 -126.315 ;
        RECT 255.515 -128.005 255.845 -127.675 ;
        RECT 255.515 -129.365 255.845 -129.035 ;
        RECT 255.515 -130.725 255.845 -130.395 ;
        RECT 255.515 -132.085 255.845 -131.755 ;
        RECT 255.515 -133.445 255.845 -133.115 ;
        RECT 255.515 -134.805 255.845 -134.475 ;
        RECT 255.515 -136.165 255.845 -135.835 ;
        RECT 255.515 -137.525 255.845 -137.195 ;
        RECT 255.515 -138.885 255.845 -138.555 ;
        RECT 255.515 -140.245 255.845 -139.915 ;
        RECT 255.515 -141.605 255.845 -141.275 ;
        RECT 255.515 -142.965 255.845 -142.635 ;
        RECT 255.515 -144.325 255.845 -143.995 ;
        RECT 255.515 -145.685 255.845 -145.355 ;
        RECT 255.515 -147.045 255.845 -146.715 ;
        RECT 255.515 -148.405 255.845 -148.075 ;
        RECT 255.515 -149.765 255.845 -149.435 ;
        RECT 255.515 -151.125 255.845 -150.795 ;
        RECT 255.515 -152.485 255.845 -152.155 ;
        RECT 255.515 -153.845 255.845 -153.515 ;
        RECT 255.515 -155.205 255.845 -154.875 ;
        RECT 255.515 -156.565 255.845 -156.235 ;
        RECT 255.515 -157.925 255.845 -157.595 ;
        RECT 255.515 -159.285 255.845 -158.955 ;
        RECT 255.515 -160.645 255.845 -160.315 ;
        RECT 255.515 -162.005 255.845 -161.675 ;
        RECT 255.515 -163.365 255.845 -163.035 ;
        RECT 255.515 -164.725 255.845 -164.395 ;
        RECT 255.515 -166.085 255.845 -165.755 ;
        RECT 255.515 -167.445 255.845 -167.115 ;
        RECT 255.515 -168.805 255.845 -168.475 ;
        RECT 255.515 -170.165 255.845 -169.835 ;
        RECT 255.515 -171.525 255.845 -171.195 ;
        RECT 255.515 -172.885 255.845 -172.555 ;
        RECT 255.515 -174.245 255.845 -173.915 ;
        RECT 255.515 -175.605 255.845 -175.275 ;
        RECT 255.515 -176.965 255.845 -176.635 ;
        RECT 255.515 -178.325 255.845 -177.995 ;
        RECT 255.515 -179.685 255.845 -179.355 ;
        RECT 255.515 -181.045 255.845 -180.715 ;
        RECT 255.515 -182.405 255.845 -182.075 ;
        RECT 255.515 -183.765 255.845 -183.435 ;
        RECT 255.515 -185.125 255.845 -184.795 ;
        RECT 255.515 -186.485 255.845 -186.155 ;
        RECT 255.515 -187.845 255.845 -187.515 ;
        RECT 255.515 -189.205 255.845 -188.875 ;
        RECT 255.515 -190.565 255.845 -190.235 ;
        RECT 255.515 -191.925 255.845 -191.595 ;
        RECT 255.515 -193.285 255.845 -192.955 ;
        RECT 255.515 -194.645 255.845 -194.315 ;
        RECT 255.515 -196.005 255.845 -195.675 ;
        RECT 255.515 -197.365 255.845 -197.035 ;
        RECT 255.515 -198.725 255.845 -198.395 ;
        RECT 255.515 -200.085 255.845 -199.755 ;
        RECT 255.515 -201.445 255.845 -201.115 ;
        RECT 255.515 -202.805 255.845 -202.475 ;
        RECT 255.515 -204.165 255.845 -203.835 ;
        RECT 255.515 -205.525 255.845 -205.195 ;
        RECT 255.515 -206.885 255.845 -206.555 ;
        RECT 255.515 -208.245 255.845 -207.915 ;
        RECT 255.515 -209.605 255.845 -209.275 ;
        RECT 255.515 -210.965 255.845 -210.635 ;
        RECT 255.515 -212.325 255.845 -211.995 ;
        RECT 255.515 -213.685 255.845 -213.355 ;
        RECT 255.515 -215.045 255.845 -214.715 ;
        RECT 255.515 -216.405 255.845 -216.075 ;
        RECT 255.515 -217.765 255.845 -217.435 ;
        RECT 255.515 -219.125 255.845 -218.795 ;
        RECT 255.515 -220.485 255.845 -220.155 ;
        RECT 255.515 -221.845 255.845 -221.515 ;
        RECT 255.515 -223.205 255.845 -222.875 ;
        RECT 255.515 -224.565 255.845 -224.235 ;
        RECT 255.515 -225.925 255.845 -225.595 ;
        RECT 255.515 -227.285 255.845 -226.955 ;
        RECT 255.515 -228.645 255.845 -228.315 ;
        RECT 255.515 -230.005 255.845 -229.675 ;
        RECT 255.515 -231.365 255.845 -231.035 ;
        RECT 255.515 -232.725 255.845 -232.395 ;
        RECT 255.515 -234.085 255.845 -233.755 ;
        RECT 255.515 -235.445 255.845 -235.115 ;
        RECT 255.515 -236.805 255.845 -236.475 ;
        RECT 255.515 -238.165 255.845 -237.835 ;
        RECT 255.515 -243.81 255.845 -242.68 ;
        RECT 255.52 -243.925 255.84 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 246.76 257.205 247.89 ;
        RECT 256.875 241.915 257.205 242.245 ;
        RECT 256.875 240.555 257.205 240.885 ;
        RECT 256.875 239.195 257.205 239.525 ;
        RECT 256.875 237.835 257.205 238.165 ;
        RECT 256.88 237.16 257.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 -1.525 257.205 -1.195 ;
        RECT 256.875 -2.885 257.205 -2.555 ;
        RECT 256.88 -3.56 257.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 246.76 258.565 247.89 ;
        RECT 258.235 241.915 258.565 242.245 ;
        RECT 258.235 240.555 258.565 240.885 ;
        RECT 258.235 239.195 258.565 239.525 ;
        RECT 258.235 237.835 258.565 238.165 ;
        RECT 258.24 237.16 258.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 -1.525 258.565 -1.195 ;
        RECT 258.235 -2.885 258.565 -2.555 ;
        RECT 258.24 -3.56 258.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 -122.565 258.565 -122.235 ;
        RECT 258.235 -123.925 258.565 -123.595 ;
        RECT 258.235 -125.285 258.565 -124.955 ;
        RECT 258.235 -126.645 258.565 -126.315 ;
        RECT 258.235 -128.005 258.565 -127.675 ;
        RECT 258.235 -129.365 258.565 -129.035 ;
        RECT 258.235 -130.725 258.565 -130.395 ;
        RECT 258.235 -132.085 258.565 -131.755 ;
        RECT 258.235 -133.445 258.565 -133.115 ;
        RECT 258.235 -134.805 258.565 -134.475 ;
        RECT 258.235 -136.165 258.565 -135.835 ;
        RECT 258.235 -137.525 258.565 -137.195 ;
        RECT 258.235 -138.885 258.565 -138.555 ;
        RECT 258.235 -140.245 258.565 -139.915 ;
        RECT 258.235 -141.605 258.565 -141.275 ;
        RECT 258.235 -142.965 258.565 -142.635 ;
        RECT 258.235 -144.325 258.565 -143.995 ;
        RECT 258.235 -145.685 258.565 -145.355 ;
        RECT 258.235 -147.045 258.565 -146.715 ;
        RECT 258.235 -148.405 258.565 -148.075 ;
        RECT 258.235 -149.765 258.565 -149.435 ;
        RECT 258.235 -151.125 258.565 -150.795 ;
        RECT 258.235 -152.485 258.565 -152.155 ;
        RECT 258.235 -153.845 258.565 -153.515 ;
        RECT 258.235 -155.205 258.565 -154.875 ;
        RECT 258.235 -156.565 258.565 -156.235 ;
        RECT 258.235 -157.925 258.565 -157.595 ;
        RECT 258.235 -159.285 258.565 -158.955 ;
        RECT 258.235 -160.645 258.565 -160.315 ;
        RECT 258.235 -162.005 258.565 -161.675 ;
        RECT 258.235 -163.365 258.565 -163.035 ;
        RECT 258.235 -164.725 258.565 -164.395 ;
        RECT 258.235 -166.085 258.565 -165.755 ;
        RECT 258.235 -167.445 258.565 -167.115 ;
        RECT 258.235 -168.805 258.565 -168.475 ;
        RECT 258.235 -170.165 258.565 -169.835 ;
        RECT 258.235 -171.525 258.565 -171.195 ;
        RECT 258.235 -172.885 258.565 -172.555 ;
        RECT 258.235 -174.245 258.565 -173.915 ;
        RECT 258.235 -175.605 258.565 -175.275 ;
        RECT 258.235 -176.965 258.565 -176.635 ;
        RECT 258.235 -178.325 258.565 -177.995 ;
        RECT 258.235 -179.685 258.565 -179.355 ;
        RECT 258.235 -181.045 258.565 -180.715 ;
        RECT 258.235 -182.405 258.565 -182.075 ;
        RECT 258.235 -183.765 258.565 -183.435 ;
        RECT 258.235 -185.125 258.565 -184.795 ;
        RECT 258.235 -186.485 258.565 -186.155 ;
        RECT 258.235 -187.845 258.565 -187.515 ;
        RECT 258.235 -189.205 258.565 -188.875 ;
        RECT 258.235 -190.565 258.565 -190.235 ;
        RECT 258.235 -191.925 258.565 -191.595 ;
        RECT 258.235 -193.285 258.565 -192.955 ;
        RECT 258.235 -194.645 258.565 -194.315 ;
        RECT 258.235 -196.005 258.565 -195.675 ;
        RECT 258.235 -197.365 258.565 -197.035 ;
        RECT 258.235 -198.725 258.565 -198.395 ;
        RECT 258.235 -200.085 258.565 -199.755 ;
        RECT 258.235 -201.445 258.565 -201.115 ;
        RECT 258.235 -202.805 258.565 -202.475 ;
        RECT 258.235 -204.165 258.565 -203.835 ;
        RECT 258.235 -205.525 258.565 -205.195 ;
        RECT 258.235 -206.885 258.565 -206.555 ;
        RECT 258.235 -208.245 258.565 -207.915 ;
        RECT 258.235 -209.605 258.565 -209.275 ;
        RECT 258.235 -210.965 258.565 -210.635 ;
        RECT 258.235 -212.325 258.565 -211.995 ;
        RECT 258.235 -213.685 258.565 -213.355 ;
        RECT 258.235 -215.045 258.565 -214.715 ;
        RECT 258.235 -216.405 258.565 -216.075 ;
        RECT 258.235 -217.765 258.565 -217.435 ;
        RECT 258.235 -219.125 258.565 -218.795 ;
        RECT 258.235 -220.485 258.565 -220.155 ;
        RECT 258.235 -221.845 258.565 -221.515 ;
        RECT 258.235 -223.205 258.565 -222.875 ;
        RECT 258.235 -224.565 258.565 -224.235 ;
        RECT 258.235 -225.925 258.565 -225.595 ;
        RECT 258.235 -227.285 258.565 -226.955 ;
        RECT 258.235 -228.645 258.565 -228.315 ;
        RECT 258.235 -230.005 258.565 -229.675 ;
        RECT 258.235 -231.365 258.565 -231.035 ;
        RECT 258.235 -232.725 258.565 -232.395 ;
        RECT 258.235 -234.085 258.565 -233.755 ;
        RECT 258.235 -235.445 258.565 -235.115 ;
        RECT 258.235 -236.805 258.565 -236.475 ;
        RECT 258.235 -238.165 258.565 -237.835 ;
        RECT 258.235 -243.81 258.565 -242.68 ;
        RECT 258.24 -243.925 258.56 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 246.76 259.925 247.89 ;
        RECT 259.595 241.915 259.925 242.245 ;
        RECT 259.595 240.555 259.925 240.885 ;
        RECT 259.595 239.195 259.925 239.525 ;
        RECT 259.595 237.835 259.925 238.165 ;
        RECT 259.6 237.16 259.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 -1.525 259.925 -1.195 ;
        RECT 259.595 -2.885 259.925 -2.555 ;
        RECT 259.6 -3.56 259.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 -122.565 259.925 -122.235 ;
        RECT 259.595 -123.925 259.925 -123.595 ;
        RECT 259.595 -125.285 259.925 -124.955 ;
        RECT 259.595 -126.645 259.925 -126.315 ;
        RECT 259.595 -128.005 259.925 -127.675 ;
        RECT 259.595 -129.365 259.925 -129.035 ;
        RECT 259.595 -130.725 259.925 -130.395 ;
        RECT 259.595 -132.085 259.925 -131.755 ;
        RECT 259.595 -133.445 259.925 -133.115 ;
        RECT 259.595 -134.805 259.925 -134.475 ;
        RECT 259.595 -136.165 259.925 -135.835 ;
        RECT 259.595 -137.525 259.925 -137.195 ;
        RECT 259.595 -138.885 259.925 -138.555 ;
        RECT 259.595 -140.245 259.925 -139.915 ;
        RECT 259.595 -141.605 259.925 -141.275 ;
        RECT 259.595 -142.965 259.925 -142.635 ;
        RECT 259.595 -144.325 259.925 -143.995 ;
        RECT 259.595 -145.685 259.925 -145.355 ;
        RECT 259.595 -147.045 259.925 -146.715 ;
        RECT 259.595 -148.405 259.925 -148.075 ;
        RECT 259.595 -149.765 259.925 -149.435 ;
        RECT 259.595 -151.125 259.925 -150.795 ;
        RECT 259.595 -152.485 259.925 -152.155 ;
        RECT 259.595 -153.845 259.925 -153.515 ;
        RECT 259.595 -155.205 259.925 -154.875 ;
        RECT 259.595 -156.565 259.925 -156.235 ;
        RECT 259.595 -157.925 259.925 -157.595 ;
        RECT 259.595 -159.285 259.925 -158.955 ;
        RECT 259.595 -160.645 259.925 -160.315 ;
        RECT 259.595 -162.005 259.925 -161.675 ;
        RECT 259.595 -163.365 259.925 -163.035 ;
        RECT 259.595 -164.725 259.925 -164.395 ;
        RECT 259.595 -166.085 259.925 -165.755 ;
        RECT 259.595 -167.445 259.925 -167.115 ;
        RECT 259.595 -168.805 259.925 -168.475 ;
        RECT 259.595 -170.165 259.925 -169.835 ;
        RECT 259.595 -171.525 259.925 -171.195 ;
        RECT 259.595 -172.885 259.925 -172.555 ;
        RECT 259.595 -174.245 259.925 -173.915 ;
        RECT 259.595 -175.605 259.925 -175.275 ;
        RECT 259.595 -176.965 259.925 -176.635 ;
        RECT 259.595 -178.325 259.925 -177.995 ;
        RECT 259.595 -179.685 259.925 -179.355 ;
        RECT 259.595 -181.045 259.925 -180.715 ;
        RECT 259.595 -182.405 259.925 -182.075 ;
        RECT 259.595 -183.765 259.925 -183.435 ;
        RECT 259.595 -185.125 259.925 -184.795 ;
        RECT 259.595 -186.485 259.925 -186.155 ;
        RECT 259.595 -187.845 259.925 -187.515 ;
        RECT 259.595 -189.205 259.925 -188.875 ;
        RECT 259.595 -190.565 259.925 -190.235 ;
        RECT 259.595 -191.925 259.925 -191.595 ;
        RECT 259.595 -193.285 259.925 -192.955 ;
        RECT 259.595 -194.645 259.925 -194.315 ;
        RECT 259.595 -196.005 259.925 -195.675 ;
        RECT 259.595 -197.365 259.925 -197.035 ;
        RECT 259.595 -198.725 259.925 -198.395 ;
        RECT 259.595 -200.085 259.925 -199.755 ;
        RECT 259.595 -201.445 259.925 -201.115 ;
        RECT 259.595 -202.805 259.925 -202.475 ;
        RECT 259.595 -204.165 259.925 -203.835 ;
        RECT 259.595 -205.525 259.925 -205.195 ;
        RECT 259.595 -206.885 259.925 -206.555 ;
        RECT 259.595 -208.245 259.925 -207.915 ;
        RECT 259.595 -209.605 259.925 -209.275 ;
        RECT 259.595 -210.965 259.925 -210.635 ;
        RECT 259.595 -212.325 259.925 -211.995 ;
        RECT 259.595 -213.685 259.925 -213.355 ;
        RECT 259.595 -215.045 259.925 -214.715 ;
        RECT 259.595 -216.405 259.925 -216.075 ;
        RECT 259.595 -217.765 259.925 -217.435 ;
        RECT 259.595 -219.125 259.925 -218.795 ;
        RECT 259.595 -220.485 259.925 -220.155 ;
        RECT 259.595 -221.845 259.925 -221.515 ;
        RECT 259.595 -223.205 259.925 -222.875 ;
        RECT 259.595 -224.565 259.925 -224.235 ;
        RECT 259.595 -225.925 259.925 -225.595 ;
        RECT 259.595 -227.285 259.925 -226.955 ;
        RECT 259.595 -228.645 259.925 -228.315 ;
        RECT 259.595 -230.005 259.925 -229.675 ;
        RECT 259.595 -231.365 259.925 -231.035 ;
        RECT 259.595 -232.725 259.925 -232.395 ;
        RECT 259.595 -234.085 259.925 -233.755 ;
        RECT 259.595 -235.445 259.925 -235.115 ;
        RECT 259.595 -236.805 259.925 -236.475 ;
        RECT 259.595 -238.165 259.925 -237.835 ;
        RECT 259.595 -243.81 259.925 -242.68 ;
        RECT 259.6 -243.925 259.92 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 246.76 261.285 247.89 ;
        RECT 260.955 241.915 261.285 242.245 ;
        RECT 260.955 240.555 261.285 240.885 ;
        RECT 260.955 239.195 261.285 239.525 ;
        RECT 260.955 237.835 261.285 238.165 ;
        RECT 260.96 237.16 261.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 -1.525 261.285 -1.195 ;
        RECT 260.955 -2.885 261.285 -2.555 ;
        RECT 260.96 -3.56 261.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 -122.565 261.285 -122.235 ;
        RECT 260.955 -123.925 261.285 -123.595 ;
        RECT 260.955 -125.285 261.285 -124.955 ;
        RECT 260.955 -126.645 261.285 -126.315 ;
        RECT 260.955 -128.005 261.285 -127.675 ;
        RECT 260.955 -129.365 261.285 -129.035 ;
        RECT 260.955 -130.725 261.285 -130.395 ;
        RECT 260.955 -132.085 261.285 -131.755 ;
        RECT 260.955 -133.445 261.285 -133.115 ;
        RECT 260.955 -134.805 261.285 -134.475 ;
        RECT 260.955 -136.165 261.285 -135.835 ;
        RECT 260.955 -137.525 261.285 -137.195 ;
        RECT 260.955 -138.885 261.285 -138.555 ;
        RECT 260.955 -140.245 261.285 -139.915 ;
        RECT 260.955 -141.605 261.285 -141.275 ;
        RECT 260.955 -142.965 261.285 -142.635 ;
        RECT 260.955 -144.325 261.285 -143.995 ;
        RECT 260.955 -145.685 261.285 -145.355 ;
        RECT 260.955 -147.045 261.285 -146.715 ;
        RECT 260.955 -148.405 261.285 -148.075 ;
        RECT 260.955 -149.765 261.285 -149.435 ;
        RECT 260.955 -151.125 261.285 -150.795 ;
        RECT 260.955 -152.485 261.285 -152.155 ;
        RECT 260.955 -153.845 261.285 -153.515 ;
        RECT 260.955 -155.205 261.285 -154.875 ;
        RECT 260.955 -156.565 261.285 -156.235 ;
        RECT 260.955 -157.925 261.285 -157.595 ;
        RECT 260.955 -159.285 261.285 -158.955 ;
        RECT 260.955 -160.645 261.285 -160.315 ;
        RECT 260.955 -162.005 261.285 -161.675 ;
        RECT 260.955 -163.365 261.285 -163.035 ;
        RECT 260.955 -164.725 261.285 -164.395 ;
        RECT 260.955 -166.085 261.285 -165.755 ;
        RECT 260.955 -167.445 261.285 -167.115 ;
        RECT 260.955 -168.805 261.285 -168.475 ;
        RECT 260.955 -170.165 261.285 -169.835 ;
        RECT 260.955 -171.525 261.285 -171.195 ;
        RECT 260.955 -172.885 261.285 -172.555 ;
        RECT 260.955 -174.245 261.285 -173.915 ;
        RECT 260.955 -175.605 261.285 -175.275 ;
        RECT 260.955 -176.965 261.285 -176.635 ;
        RECT 260.955 -178.325 261.285 -177.995 ;
        RECT 260.955 -179.685 261.285 -179.355 ;
        RECT 260.955 -181.045 261.285 -180.715 ;
        RECT 260.955 -182.405 261.285 -182.075 ;
        RECT 260.955 -183.765 261.285 -183.435 ;
        RECT 260.955 -185.125 261.285 -184.795 ;
        RECT 260.955 -186.485 261.285 -186.155 ;
        RECT 260.955 -187.845 261.285 -187.515 ;
        RECT 260.955 -189.205 261.285 -188.875 ;
        RECT 260.955 -190.565 261.285 -190.235 ;
        RECT 260.955 -191.925 261.285 -191.595 ;
        RECT 260.955 -193.285 261.285 -192.955 ;
        RECT 260.955 -194.645 261.285 -194.315 ;
        RECT 260.955 -196.005 261.285 -195.675 ;
        RECT 260.955 -197.365 261.285 -197.035 ;
        RECT 260.955 -198.725 261.285 -198.395 ;
        RECT 260.955 -200.085 261.285 -199.755 ;
        RECT 260.955 -201.445 261.285 -201.115 ;
        RECT 260.955 -202.805 261.285 -202.475 ;
        RECT 260.955 -204.165 261.285 -203.835 ;
        RECT 260.955 -205.525 261.285 -205.195 ;
        RECT 260.955 -206.885 261.285 -206.555 ;
        RECT 260.955 -208.245 261.285 -207.915 ;
        RECT 260.955 -209.605 261.285 -209.275 ;
        RECT 260.955 -210.965 261.285 -210.635 ;
        RECT 260.955 -212.325 261.285 -211.995 ;
        RECT 260.955 -213.685 261.285 -213.355 ;
        RECT 260.955 -215.045 261.285 -214.715 ;
        RECT 260.955 -216.405 261.285 -216.075 ;
        RECT 260.955 -217.765 261.285 -217.435 ;
        RECT 260.955 -219.125 261.285 -218.795 ;
        RECT 260.955 -220.485 261.285 -220.155 ;
        RECT 260.955 -221.845 261.285 -221.515 ;
        RECT 260.955 -223.205 261.285 -222.875 ;
        RECT 260.955 -224.565 261.285 -224.235 ;
        RECT 260.955 -225.925 261.285 -225.595 ;
        RECT 260.955 -227.285 261.285 -226.955 ;
        RECT 260.955 -228.645 261.285 -228.315 ;
        RECT 260.955 -230.005 261.285 -229.675 ;
        RECT 260.955 -231.365 261.285 -231.035 ;
        RECT 260.955 -232.725 261.285 -232.395 ;
        RECT 260.955 -234.085 261.285 -233.755 ;
        RECT 260.955 -235.445 261.285 -235.115 ;
        RECT 260.955 -236.805 261.285 -236.475 ;
        RECT 260.955 -238.165 261.285 -237.835 ;
        RECT 260.955 -243.81 261.285 -242.68 ;
        RECT 260.96 -243.925 261.28 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 237.835 262.645 238.165 ;
        RECT 262.32 237.16 262.64 248.005 ;
        RECT 262.315 246.76 262.645 247.89 ;
        RECT 262.315 241.915 262.645 242.245 ;
        RECT 262.315 240.555 262.645 240.885 ;
        RECT 262.315 239.195 262.645 239.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 246.76 227.285 247.89 ;
        RECT 226.955 241.915 227.285 242.245 ;
        RECT 226.955 240.555 227.285 240.885 ;
        RECT 226.955 239.195 227.285 239.525 ;
        RECT 226.955 237.835 227.285 238.165 ;
        RECT 226.96 237.16 227.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 -1.525 227.285 -1.195 ;
        RECT 226.955 -2.885 227.285 -2.555 ;
        RECT 226.96 -3.56 227.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 -122.565 227.285 -122.235 ;
        RECT 226.955 -123.925 227.285 -123.595 ;
        RECT 226.955 -125.285 227.285 -124.955 ;
        RECT 226.955 -126.645 227.285 -126.315 ;
        RECT 226.955 -128.005 227.285 -127.675 ;
        RECT 226.955 -129.365 227.285 -129.035 ;
        RECT 226.955 -130.725 227.285 -130.395 ;
        RECT 226.955 -132.085 227.285 -131.755 ;
        RECT 226.955 -133.445 227.285 -133.115 ;
        RECT 226.955 -134.805 227.285 -134.475 ;
        RECT 226.955 -136.165 227.285 -135.835 ;
        RECT 226.955 -137.525 227.285 -137.195 ;
        RECT 226.955 -138.885 227.285 -138.555 ;
        RECT 226.955 -140.245 227.285 -139.915 ;
        RECT 226.955 -141.605 227.285 -141.275 ;
        RECT 226.955 -142.965 227.285 -142.635 ;
        RECT 226.955 -144.325 227.285 -143.995 ;
        RECT 226.955 -145.685 227.285 -145.355 ;
        RECT 226.955 -147.045 227.285 -146.715 ;
        RECT 226.955 -148.405 227.285 -148.075 ;
        RECT 226.955 -149.765 227.285 -149.435 ;
        RECT 226.955 -151.125 227.285 -150.795 ;
        RECT 226.955 -152.485 227.285 -152.155 ;
        RECT 226.955 -153.845 227.285 -153.515 ;
        RECT 226.955 -155.205 227.285 -154.875 ;
        RECT 226.955 -156.565 227.285 -156.235 ;
        RECT 226.955 -157.925 227.285 -157.595 ;
        RECT 226.955 -159.285 227.285 -158.955 ;
        RECT 226.955 -160.645 227.285 -160.315 ;
        RECT 226.955 -162.005 227.285 -161.675 ;
        RECT 226.955 -163.365 227.285 -163.035 ;
        RECT 226.955 -164.725 227.285 -164.395 ;
        RECT 226.955 -166.085 227.285 -165.755 ;
        RECT 226.955 -167.445 227.285 -167.115 ;
        RECT 226.955 -168.805 227.285 -168.475 ;
        RECT 226.955 -170.165 227.285 -169.835 ;
        RECT 226.955 -171.525 227.285 -171.195 ;
        RECT 226.955 -172.885 227.285 -172.555 ;
        RECT 226.955 -174.245 227.285 -173.915 ;
        RECT 226.955 -175.605 227.285 -175.275 ;
        RECT 226.955 -176.965 227.285 -176.635 ;
        RECT 226.955 -178.325 227.285 -177.995 ;
        RECT 226.955 -179.685 227.285 -179.355 ;
        RECT 226.955 -181.045 227.285 -180.715 ;
        RECT 226.955 -182.405 227.285 -182.075 ;
        RECT 226.955 -183.765 227.285 -183.435 ;
        RECT 226.955 -185.125 227.285 -184.795 ;
        RECT 226.955 -186.485 227.285 -186.155 ;
        RECT 226.955 -187.845 227.285 -187.515 ;
        RECT 226.955 -189.205 227.285 -188.875 ;
        RECT 226.955 -190.565 227.285 -190.235 ;
        RECT 226.955 -191.925 227.285 -191.595 ;
        RECT 226.955 -193.285 227.285 -192.955 ;
        RECT 226.955 -194.645 227.285 -194.315 ;
        RECT 226.955 -196.005 227.285 -195.675 ;
        RECT 226.955 -197.365 227.285 -197.035 ;
        RECT 226.955 -198.725 227.285 -198.395 ;
        RECT 226.955 -200.085 227.285 -199.755 ;
        RECT 226.955 -201.445 227.285 -201.115 ;
        RECT 226.955 -202.805 227.285 -202.475 ;
        RECT 226.955 -204.165 227.285 -203.835 ;
        RECT 226.955 -205.525 227.285 -205.195 ;
        RECT 226.955 -206.885 227.285 -206.555 ;
        RECT 226.955 -208.245 227.285 -207.915 ;
        RECT 226.955 -209.605 227.285 -209.275 ;
        RECT 226.955 -210.965 227.285 -210.635 ;
        RECT 226.955 -212.325 227.285 -211.995 ;
        RECT 226.955 -213.685 227.285 -213.355 ;
        RECT 226.955 -215.045 227.285 -214.715 ;
        RECT 226.955 -216.405 227.285 -216.075 ;
        RECT 226.955 -217.765 227.285 -217.435 ;
        RECT 226.955 -219.125 227.285 -218.795 ;
        RECT 226.955 -220.485 227.285 -220.155 ;
        RECT 226.955 -221.845 227.285 -221.515 ;
        RECT 226.955 -223.205 227.285 -222.875 ;
        RECT 226.955 -224.565 227.285 -224.235 ;
        RECT 226.955 -225.925 227.285 -225.595 ;
        RECT 226.955 -227.285 227.285 -226.955 ;
        RECT 226.955 -228.645 227.285 -228.315 ;
        RECT 226.955 -230.005 227.285 -229.675 ;
        RECT 226.955 -231.365 227.285 -231.035 ;
        RECT 226.955 -232.725 227.285 -232.395 ;
        RECT 226.955 -234.085 227.285 -233.755 ;
        RECT 226.955 -235.445 227.285 -235.115 ;
        RECT 226.955 -236.805 227.285 -236.475 ;
        RECT 226.955 -238.165 227.285 -237.835 ;
        RECT 226.955 -243.81 227.285 -242.68 ;
        RECT 226.96 -243.925 227.28 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 246.76 228.645 247.89 ;
        RECT 228.315 241.915 228.645 242.245 ;
        RECT 228.315 240.555 228.645 240.885 ;
        RECT 228.315 239.195 228.645 239.525 ;
        RECT 228.315 237.835 228.645 238.165 ;
        RECT 228.32 237.16 228.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 -1.525 228.645 -1.195 ;
        RECT 228.315 -2.885 228.645 -2.555 ;
        RECT 228.32 -3.56 228.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 -122.565 228.645 -122.235 ;
        RECT 228.315 -123.925 228.645 -123.595 ;
        RECT 228.315 -125.285 228.645 -124.955 ;
        RECT 228.315 -126.645 228.645 -126.315 ;
        RECT 228.315 -128.005 228.645 -127.675 ;
        RECT 228.315 -129.365 228.645 -129.035 ;
        RECT 228.315 -130.725 228.645 -130.395 ;
        RECT 228.315 -132.085 228.645 -131.755 ;
        RECT 228.315 -133.445 228.645 -133.115 ;
        RECT 228.315 -134.805 228.645 -134.475 ;
        RECT 228.315 -136.165 228.645 -135.835 ;
        RECT 228.315 -137.525 228.645 -137.195 ;
        RECT 228.315 -138.885 228.645 -138.555 ;
        RECT 228.315 -140.245 228.645 -139.915 ;
        RECT 228.315 -141.605 228.645 -141.275 ;
        RECT 228.315 -142.965 228.645 -142.635 ;
        RECT 228.315 -144.325 228.645 -143.995 ;
        RECT 228.315 -145.685 228.645 -145.355 ;
        RECT 228.315 -147.045 228.645 -146.715 ;
        RECT 228.315 -148.405 228.645 -148.075 ;
        RECT 228.315 -149.765 228.645 -149.435 ;
        RECT 228.315 -151.125 228.645 -150.795 ;
        RECT 228.315 -152.485 228.645 -152.155 ;
        RECT 228.315 -153.845 228.645 -153.515 ;
        RECT 228.315 -155.205 228.645 -154.875 ;
        RECT 228.315 -156.565 228.645 -156.235 ;
        RECT 228.315 -157.925 228.645 -157.595 ;
        RECT 228.315 -159.285 228.645 -158.955 ;
        RECT 228.315 -160.645 228.645 -160.315 ;
        RECT 228.315 -162.005 228.645 -161.675 ;
        RECT 228.315 -163.365 228.645 -163.035 ;
        RECT 228.315 -164.725 228.645 -164.395 ;
        RECT 228.315 -166.085 228.645 -165.755 ;
        RECT 228.315 -167.445 228.645 -167.115 ;
        RECT 228.315 -168.805 228.645 -168.475 ;
        RECT 228.315 -170.165 228.645 -169.835 ;
        RECT 228.315 -171.525 228.645 -171.195 ;
        RECT 228.315 -172.885 228.645 -172.555 ;
        RECT 228.315 -174.245 228.645 -173.915 ;
        RECT 228.315 -175.605 228.645 -175.275 ;
        RECT 228.315 -176.965 228.645 -176.635 ;
        RECT 228.315 -178.325 228.645 -177.995 ;
        RECT 228.315 -179.685 228.645 -179.355 ;
        RECT 228.315 -181.045 228.645 -180.715 ;
        RECT 228.315 -182.405 228.645 -182.075 ;
        RECT 228.315 -183.765 228.645 -183.435 ;
        RECT 228.315 -185.125 228.645 -184.795 ;
        RECT 228.315 -186.485 228.645 -186.155 ;
        RECT 228.315 -187.845 228.645 -187.515 ;
        RECT 228.315 -189.205 228.645 -188.875 ;
        RECT 228.315 -190.565 228.645 -190.235 ;
        RECT 228.315 -191.925 228.645 -191.595 ;
        RECT 228.315 -193.285 228.645 -192.955 ;
        RECT 228.315 -194.645 228.645 -194.315 ;
        RECT 228.315 -196.005 228.645 -195.675 ;
        RECT 228.315 -197.365 228.645 -197.035 ;
        RECT 228.315 -198.725 228.645 -198.395 ;
        RECT 228.315 -200.085 228.645 -199.755 ;
        RECT 228.315 -201.445 228.645 -201.115 ;
        RECT 228.315 -202.805 228.645 -202.475 ;
        RECT 228.315 -204.165 228.645 -203.835 ;
        RECT 228.315 -205.525 228.645 -205.195 ;
        RECT 228.315 -206.885 228.645 -206.555 ;
        RECT 228.315 -208.245 228.645 -207.915 ;
        RECT 228.315 -209.605 228.645 -209.275 ;
        RECT 228.315 -210.965 228.645 -210.635 ;
        RECT 228.315 -212.325 228.645 -211.995 ;
        RECT 228.315 -213.685 228.645 -213.355 ;
        RECT 228.315 -215.045 228.645 -214.715 ;
        RECT 228.315 -216.405 228.645 -216.075 ;
        RECT 228.315 -217.765 228.645 -217.435 ;
        RECT 228.315 -219.125 228.645 -218.795 ;
        RECT 228.315 -220.485 228.645 -220.155 ;
        RECT 228.315 -221.845 228.645 -221.515 ;
        RECT 228.315 -223.205 228.645 -222.875 ;
        RECT 228.315 -224.565 228.645 -224.235 ;
        RECT 228.315 -225.925 228.645 -225.595 ;
        RECT 228.315 -227.285 228.645 -226.955 ;
        RECT 228.315 -228.645 228.645 -228.315 ;
        RECT 228.315 -230.005 228.645 -229.675 ;
        RECT 228.315 -231.365 228.645 -231.035 ;
        RECT 228.315 -232.725 228.645 -232.395 ;
        RECT 228.315 -234.085 228.645 -233.755 ;
        RECT 228.315 -235.445 228.645 -235.115 ;
        RECT 228.315 -236.805 228.645 -236.475 ;
        RECT 228.315 -238.165 228.645 -237.835 ;
        RECT 228.315 -243.81 228.645 -242.68 ;
        RECT 228.32 -243.925 228.64 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 246.76 230.005 247.89 ;
        RECT 229.675 241.915 230.005 242.245 ;
        RECT 229.675 240.555 230.005 240.885 ;
        RECT 229.675 239.195 230.005 239.525 ;
        RECT 229.675 237.835 230.005 238.165 ;
        RECT 229.68 237.16 230 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 -1.525 230.005 -1.195 ;
        RECT 229.675 -2.885 230.005 -2.555 ;
        RECT 229.68 -3.56 230 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 -122.565 230.005 -122.235 ;
        RECT 229.675 -123.925 230.005 -123.595 ;
        RECT 229.675 -125.285 230.005 -124.955 ;
        RECT 229.675 -126.645 230.005 -126.315 ;
        RECT 229.675 -128.005 230.005 -127.675 ;
        RECT 229.675 -129.365 230.005 -129.035 ;
        RECT 229.675 -130.725 230.005 -130.395 ;
        RECT 229.675 -132.085 230.005 -131.755 ;
        RECT 229.675 -133.445 230.005 -133.115 ;
        RECT 229.675 -134.805 230.005 -134.475 ;
        RECT 229.675 -136.165 230.005 -135.835 ;
        RECT 229.675 -137.525 230.005 -137.195 ;
        RECT 229.675 -138.885 230.005 -138.555 ;
        RECT 229.675 -140.245 230.005 -139.915 ;
        RECT 229.675 -141.605 230.005 -141.275 ;
        RECT 229.675 -142.965 230.005 -142.635 ;
        RECT 229.675 -144.325 230.005 -143.995 ;
        RECT 229.675 -145.685 230.005 -145.355 ;
        RECT 229.675 -147.045 230.005 -146.715 ;
        RECT 229.675 -148.405 230.005 -148.075 ;
        RECT 229.675 -149.765 230.005 -149.435 ;
        RECT 229.675 -151.125 230.005 -150.795 ;
        RECT 229.675 -152.485 230.005 -152.155 ;
        RECT 229.675 -153.845 230.005 -153.515 ;
        RECT 229.675 -155.205 230.005 -154.875 ;
        RECT 229.675 -156.565 230.005 -156.235 ;
        RECT 229.675 -157.925 230.005 -157.595 ;
        RECT 229.675 -159.285 230.005 -158.955 ;
        RECT 229.675 -160.645 230.005 -160.315 ;
        RECT 229.675 -162.005 230.005 -161.675 ;
        RECT 229.675 -163.365 230.005 -163.035 ;
        RECT 229.675 -164.725 230.005 -164.395 ;
        RECT 229.675 -166.085 230.005 -165.755 ;
        RECT 229.675 -167.445 230.005 -167.115 ;
        RECT 229.675 -168.805 230.005 -168.475 ;
        RECT 229.675 -170.165 230.005 -169.835 ;
        RECT 229.675 -171.525 230.005 -171.195 ;
        RECT 229.675 -172.885 230.005 -172.555 ;
        RECT 229.675 -174.245 230.005 -173.915 ;
        RECT 229.675 -175.605 230.005 -175.275 ;
        RECT 229.675 -176.965 230.005 -176.635 ;
        RECT 229.675 -178.325 230.005 -177.995 ;
        RECT 229.675 -179.685 230.005 -179.355 ;
        RECT 229.675 -181.045 230.005 -180.715 ;
        RECT 229.675 -182.405 230.005 -182.075 ;
        RECT 229.675 -183.765 230.005 -183.435 ;
        RECT 229.675 -185.125 230.005 -184.795 ;
        RECT 229.675 -186.485 230.005 -186.155 ;
        RECT 229.675 -187.845 230.005 -187.515 ;
        RECT 229.675 -189.205 230.005 -188.875 ;
        RECT 229.675 -190.565 230.005 -190.235 ;
        RECT 229.675 -191.925 230.005 -191.595 ;
        RECT 229.675 -193.285 230.005 -192.955 ;
        RECT 229.675 -194.645 230.005 -194.315 ;
        RECT 229.675 -196.005 230.005 -195.675 ;
        RECT 229.675 -197.365 230.005 -197.035 ;
        RECT 229.675 -198.725 230.005 -198.395 ;
        RECT 229.675 -200.085 230.005 -199.755 ;
        RECT 229.675 -201.445 230.005 -201.115 ;
        RECT 229.675 -202.805 230.005 -202.475 ;
        RECT 229.675 -204.165 230.005 -203.835 ;
        RECT 229.675 -205.525 230.005 -205.195 ;
        RECT 229.675 -206.885 230.005 -206.555 ;
        RECT 229.675 -208.245 230.005 -207.915 ;
        RECT 229.675 -209.605 230.005 -209.275 ;
        RECT 229.675 -210.965 230.005 -210.635 ;
        RECT 229.675 -212.325 230.005 -211.995 ;
        RECT 229.675 -213.685 230.005 -213.355 ;
        RECT 229.675 -215.045 230.005 -214.715 ;
        RECT 229.675 -216.405 230.005 -216.075 ;
        RECT 229.675 -217.765 230.005 -217.435 ;
        RECT 229.675 -219.125 230.005 -218.795 ;
        RECT 229.675 -220.485 230.005 -220.155 ;
        RECT 229.675 -221.845 230.005 -221.515 ;
        RECT 229.675 -223.205 230.005 -222.875 ;
        RECT 229.675 -224.565 230.005 -224.235 ;
        RECT 229.675 -225.925 230.005 -225.595 ;
        RECT 229.675 -227.285 230.005 -226.955 ;
        RECT 229.675 -228.645 230.005 -228.315 ;
        RECT 229.675 -230.005 230.005 -229.675 ;
        RECT 229.675 -231.365 230.005 -231.035 ;
        RECT 229.675 -232.725 230.005 -232.395 ;
        RECT 229.675 -234.085 230.005 -233.755 ;
        RECT 229.675 -235.445 230.005 -235.115 ;
        RECT 229.675 -236.805 230.005 -236.475 ;
        RECT 229.675 -238.165 230.005 -237.835 ;
        RECT 229.675 -243.81 230.005 -242.68 ;
        RECT 229.68 -243.925 230 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 246.76 231.365 247.89 ;
        RECT 231.035 241.915 231.365 242.245 ;
        RECT 231.035 240.555 231.365 240.885 ;
        RECT 231.035 239.195 231.365 239.525 ;
        RECT 231.035 237.835 231.365 238.165 ;
        RECT 231.04 237.16 231.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 -126.645 231.365 -126.315 ;
        RECT 231.035 -128.005 231.365 -127.675 ;
        RECT 231.035 -129.365 231.365 -129.035 ;
        RECT 231.035 -130.725 231.365 -130.395 ;
        RECT 231.035 -132.085 231.365 -131.755 ;
        RECT 231.035 -133.445 231.365 -133.115 ;
        RECT 231.035 -134.805 231.365 -134.475 ;
        RECT 231.035 -136.165 231.365 -135.835 ;
        RECT 231.035 -137.525 231.365 -137.195 ;
        RECT 231.035 -138.885 231.365 -138.555 ;
        RECT 231.035 -140.245 231.365 -139.915 ;
        RECT 231.035 -141.605 231.365 -141.275 ;
        RECT 231.035 -142.965 231.365 -142.635 ;
        RECT 231.035 -144.325 231.365 -143.995 ;
        RECT 231.035 -145.685 231.365 -145.355 ;
        RECT 231.035 -147.045 231.365 -146.715 ;
        RECT 231.035 -148.405 231.365 -148.075 ;
        RECT 231.035 -149.765 231.365 -149.435 ;
        RECT 231.035 -151.125 231.365 -150.795 ;
        RECT 231.035 -152.485 231.365 -152.155 ;
        RECT 231.035 -153.845 231.365 -153.515 ;
        RECT 231.035 -155.205 231.365 -154.875 ;
        RECT 231.035 -156.565 231.365 -156.235 ;
        RECT 231.035 -157.925 231.365 -157.595 ;
        RECT 231.035 -159.285 231.365 -158.955 ;
        RECT 231.035 -160.645 231.365 -160.315 ;
        RECT 231.035 -162.005 231.365 -161.675 ;
        RECT 231.035 -163.365 231.365 -163.035 ;
        RECT 231.035 -164.725 231.365 -164.395 ;
        RECT 231.035 -166.085 231.365 -165.755 ;
        RECT 231.035 -167.445 231.365 -167.115 ;
        RECT 231.035 -168.805 231.365 -168.475 ;
        RECT 231.035 -170.165 231.365 -169.835 ;
        RECT 231.035 -171.525 231.365 -171.195 ;
        RECT 231.035 -172.885 231.365 -172.555 ;
        RECT 231.035 -174.245 231.365 -173.915 ;
        RECT 231.035 -175.605 231.365 -175.275 ;
        RECT 231.035 -176.965 231.365 -176.635 ;
        RECT 231.035 -178.325 231.365 -177.995 ;
        RECT 231.035 -179.685 231.365 -179.355 ;
        RECT 231.035 -181.045 231.365 -180.715 ;
        RECT 231.035 -182.405 231.365 -182.075 ;
        RECT 231.035 -183.765 231.365 -183.435 ;
        RECT 231.035 -185.125 231.365 -184.795 ;
        RECT 231.035 -186.485 231.365 -186.155 ;
        RECT 231.035 -187.845 231.365 -187.515 ;
        RECT 231.035 -189.205 231.365 -188.875 ;
        RECT 231.035 -190.565 231.365 -190.235 ;
        RECT 231.035 -191.925 231.365 -191.595 ;
        RECT 231.035 -193.285 231.365 -192.955 ;
        RECT 231.035 -194.645 231.365 -194.315 ;
        RECT 231.035 -196.005 231.365 -195.675 ;
        RECT 231.035 -197.365 231.365 -197.035 ;
        RECT 231.035 -198.725 231.365 -198.395 ;
        RECT 231.035 -200.085 231.365 -199.755 ;
        RECT 231.035 -201.445 231.365 -201.115 ;
        RECT 231.035 -202.805 231.365 -202.475 ;
        RECT 231.035 -204.165 231.365 -203.835 ;
        RECT 231.035 -205.525 231.365 -205.195 ;
        RECT 231.035 -206.885 231.365 -206.555 ;
        RECT 231.035 -208.245 231.365 -207.915 ;
        RECT 231.035 -209.605 231.365 -209.275 ;
        RECT 231.035 -210.965 231.365 -210.635 ;
        RECT 231.035 -212.325 231.365 -211.995 ;
        RECT 231.035 -213.685 231.365 -213.355 ;
        RECT 231.035 -215.045 231.365 -214.715 ;
        RECT 231.035 -216.405 231.365 -216.075 ;
        RECT 231.035 -217.765 231.365 -217.435 ;
        RECT 231.035 -219.125 231.365 -218.795 ;
        RECT 231.035 -220.485 231.365 -220.155 ;
        RECT 231.035 -221.845 231.365 -221.515 ;
        RECT 231.035 -223.205 231.365 -222.875 ;
        RECT 231.035 -224.565 231.365 -224.235 ;
        RECT 231.035 -225.925 231.365 -225.595 ;
        RECT 231.035 -227.285 231.365 -226.955 ;
        RECT 231.035 -228.645 231.365 -228.315 ;
        RECT 231.035 -230.005 231.365 -229.675 ;
        RECT 231.035 -231.365 231.365 -231.035 ;
        RECT 231.035 -232.725 231.365 -232.395 ;
        RECT 231.035 -234.085 231.365 -233.755 ;
        RECT 231.035 -235.445 231.365 -235.115 ;
        RECT 231.035 -236.805 231.365 -236.475 ;
        RECT 231.035 -238.165 231.365 -237.835 ;
        RECT 231.035 -243.81 231.365 -242.68 ;
        RECT 231.04 -243.925 231.36 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.56 -125.535 231.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.395 246.76 232.725 247.89 ;
        RECT 232.395 241.915 232.725 242.245 ;
        RECT 232.395 240.555 232.725 240.885 ;
        RECT 232.395 239.195 232.725 239.525 ;
        RECT 232.395 237.835 232.725 238.165 ;
        RECT 232.4 237.16 232.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 246.76 234.085 247.89 ;
        RECT 233.755 241.915 234.085 242.245 ;
        RECT 233.755 240.555 234.085 240.885 ;
        RECT 233.755 239.195 234.085 239.525 ;
        RECT 233.755 237.835 234.085 238.165 ;
        RECT 233.76 237.16 234.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 -1.525 234.085 -1.195 ;
        RECT 233.755 -2.885 234.085 -2.555 ;
        RECT 233.76 -3.56 234.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 -122.565 234.085 -122.235 ;
        RECT 233.755 -123.925 234.085 -123.595 ;
        RECT 233.755 -125.285 234.085 -124.955 ;
        RECT 233.755 -126.645 234.085 -126.315 ;
        RECT 233.755 -128.005 234.085 -127.675 ;
        RECT 233.755 -129.365 234.085 -129.035 ;
        RECT 233.755 -130.725 234.085 -130.395 ;
        RECT 233.755 -132.085 234.085 -131.755 ;
        RECT 233.755 -133.445 234.085 -133.115 ;
        RECT 233.755 -134.805 234.085 -134.475 ;
        RECT 233.755 -136.165 234.085 -135.835 ;
        RECT 233.755 -137.525 234.085 -137.195 ;
        RECT 233.755 -138.885 234.085 -138.555 ;
        RECT 233.755 -140.245 234.085 -139.915 ;
        RECT 233.755 -141.605 234.085 -141.275 ;
        RECT 233.755 -142.965 234.085 -142.635 ;
        RECT 233.755 -144.325 234.085 -143.995 ;
        RECT 233.755 -145.685 234.085 -145.355 ;
        RECT 233.755 -147.045 234.085 -146.715 ;
        RECT 233.755 -148.405 234.085 -148.075 ;
        RECT 233.755 -149.765 234.085 -149.435 ;
        RECT 233.755 -151.125 234.085 -150.795 ;
        RECT 233.755 -152.485 234.085 -152.155 ;
        RECT 233.755 -153.845 234.085 -153.515 ;
        RECT 233.755 -155.205 234.085 -154.875 ;
        RECT 233.755 -156.565 234.085 -156.235 ;
        RECT 233.755 -157.925 234.085 -157.595 ;
        RECT 233.755 -159.285 234.085 -158.955 ;
        RECT 233.755 -160.645 234.085 -160.315 ;
        RECT 233.755 -162.005 234.085 -161.675 ;
        RECT 233.755 -163.365 234.085 -163.035 ;
        RECT 233.755 -164.725 234.085 -164.395 ;
        RECT 233.755 -166.085 234.085 -165.755 ;
        RECT 233.755 -167.445 234.085 -167.115 ;
        RECT 233.755 -168.805 234.085 -168.475 ;
        RECT 233.755 -170.165 234.085 -169.835 ;
        RECT 233.755 -171.525 234.085 -171.195 ;
        RECT 233.755 -172.885 234.085 -172.555 ;
        RECT 233.755 -174.245 234.085 -173.915 ;
        RECT 233.755 -175.605 234.085 -175.275 ;
        RECT 233.755 -176.965 234.085 -176.635 ;
        RECT 233.755 -178.325 234.085 -177.995 ;
        RECT 233.755 -179.685 234.085 -179.355 ;
        RECT 233.755 -181.045 234.085 -180.715 ;
        RECT 233.755 -182.405 234.085 -182.075 ;
        RECT 233.755 -183.765 234.085 -183.435 ;
        RECT 233.755 -185.125 234.085 -184.795 ;
        RECT 233.755 -186.485 234.085 -186.155 ;
        RECT 233.755 -187.845 234.085 -187.515 ;
        RECT 233.755 -189.205 234.085 -188.875 ;
        RECT 233.755 -190.565 234.085 -190.235 ;
        RECT 233.755 -191.925 234.085 -191.595 ;
        RECT 233.755 -193.285 234.085 -192.955 ;
        RECT 233.755 -194.645 234.085 -194.315 ;
        RECT 233.755 -196.005 234.085 -195.675 ;
        RECT 233.755 -197.365 234.085 -197.035 ;
        RECT 233.755 -198.725 234.085 -198.395 ;
        RECT 233.755 -200.085 234.085 -199.755 ;
        RECT 233.755 -201.445 234.085 -201.115 ;
        RECT 233.755 -202.805 234.085 -202.475 ;
        RECT 233.755 -204.165 234.085 -203.835 ;
        RECT 233.755 -205.525 234.085 -205.195 ;
        RECT 233.755 -206.885 234.085 -206.555 ;
        RECT 233.755 -208.245 234.085 -207.915 ;
        RECT 233.755 -209.605 234.085 -209.275 ;
        RECT 233.755 -210.965 234.085 -210.635 ;
        RECT 233.755 -212.325 234.085 -211.995 ;
        RECT 233.755 -213.685 234.085 -213.355 ;
        RECT 233.755 -215.045 234.085 -214.715 ;
        RECT 233.755 -216.405 234.085 -216.075 ;
        RECT 233.755 -217.765 234.085 -217.435 ;
        RECT 233.755 -219.125 234.085 -218.795 ;
        RECT 233.755 -220.485 234.085 -220.155 ;
        RECT 233.755 -221.845 234.085 -221.515 ;
        RECT 233.755 -223.205 234.085 -222.875 ;
        RECT 233.755 -224.565 234.085 -224.235 ;
        RECT 233.755 -225.925 234.085 -225.595 ;
        RECT 233.755 -227.285 234.085 -226.955 ;
        RECT 233.755 -228.645 234.085 -228.315 ;
        RECT 233.755 -230.005 234.085 -229.675 ;
        RECT 233.755 -231.365 234.085 -231.035 ;
        RECT 233.755 -232.725 234.085 -232.395 ;
        RECT 233.755 -234.085 234.085 -233.755 ;
        RECT 233.755 -235.445 234.085 -235.115 ;
        RECT 233.755 -236.805 234.085 -236.475 ;
        RECT 233.755 -238.165 234.085 -237.835 ;
        RECT 233.755 -243.81 234.085 -242.68 ;
        RECT 233.76 -243.925 234.08 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 246.76 235.445 247.89 ;
        RECT 235.115 241.915 235.445 242.245 ;
        RECT 235.115 240.555 235.445 240.885 ;
        RECT 235.115 239.195 235.445 239.525 ;
        RECT 235.115 237.835 235.445 238.165 ;
        RECT 235.12 237.16 235.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 -1.525 235.445 -1.195 ;
        RECT 235.115 -2.885 235.445 -2.555 ;
        RECT 235.12 -3.56 235.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 246.76 236.805 247.89 ;
        RECT 236.475 241.915 236.805 242.245 ;
        RECT 236.475 240.555 236.805 240.885 ;
        RECT 236.475 239.195 236.805 239.525 ;
        RECT 236.475 237.835 236.805 238.165 ;
        RECT 236.48 237.16 236.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 -1.525 236.805 -1.195 ;
        RECT 236.475 -2.885 236.805 -2.555 ;
        RECT 236.48 -3.56 236.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 -122.565 236.805 -122.235 ;
        RECT 236.475 -123.925 236.805 -123.595 ;
        RECT 236.475 -125.285 236.805 -124.955 ;
        RECT 236.475 -126.645 236.805 -126.315 ;
        RECT 236.475 -128.005 236.805 -127.675 ;
        RECT 236.475 -129.365 236.805 -129.035 ;
        RECT 236.475 -130.725 236.805 -130.395 ;
        RECT 236.475 -132.085 236.805 -131.755 ;
        RECT 236.475 -133.445 236.805 -133.115 ;
        RECT 236.475 -134.805 236.805 -134.475 ;
        RECT 236.475 -136.165 236.805 -135.835 ;
        RECT 236.475 -137.525 236.805 -137.195 ;
        RECT 236.475 -138.885 236.805 -138.555 ;
        RECT 236.475 -140.245 236.805 -139.915 ;
        RECT 236.475 -141.605 236.805 -141.275 ;
        RECT 236.475 -142.965 236.805 -142.635 ;
        RECT 236.475 -144.325 236.805 -143.995 ;
        RECT 236.475 -145.685 236.805 -145.355 ;
        RECT 236.475 -147.045 236.805 -146.715 ;
        RECT 236.475 -148.405 236.805 -148.075 ;
        RECT 236.475 -149.765 236.805 -149.435 ;
        RECT 236.475 -151.125 236.805 -150.795 ;
        RECT 236.475 -152.485 236.805 -152.155 ;
        RECT 236.475 -153.845 236.805 -153.515 ;
        RECT 236.475 -155.205 236.805 -154.875 ;
        RECT 236.475 -156.565 236.805 -156.235 ;
        RECT 236.475 -157.925 236.805 -157.595 ;
        RECT 236.475 -159.285 236.805 -158.955 ;
        RECT 236.475 -160.645 236.805 -160.315 ;
        RECT 236.475 -162.005 236.805 -161.675 ;
        RECT 236.475 -163.365 236.805 -163.035 ;
        RECT 236.475 -164.725 236.805 -164.395 ;
        RECT 236.475 -166.085 236.805 -165.755 ;
        RECT 236.475 -167.445 236.805 -167.115 ;
        RECT 236.475 -168.805 236.805 -168.475 ;
        RECT 236.475 -170.165 236.805 -169.835 ;
        RECT 236.475 -171.525 236.805 -171.195 ;
        RECT 236.475 -172.885 236.805 -172.555 ;
        RECT 236.475 -174.245 236.805 -173.915 ;
        RECT 236.475 -175.605 236.805 -175.275 ;
        RECT 236.475 -176.965 236.805 -176.635 ;
        RECT 236.475 -178.325 236.805 -177.995 ;
        RECT 236.475 -179.685 236.805 -179.355 ;
        RECT 236.475 -181.045 236.805 -180.715 ;
        RECT 236.475 -182.405 236.805 -182.075 ;
        RECT 236.475 -183.765 236.805 -183.435 ;
        RECT 236.475 -185.125 236.805 -184.795 ;
        RECT 236.475 -186.485 236.805 -186.155 ;
        RECT 236.475 -187.845 236.805 -187.515 ;
        RECT 236.475 -189.205 236.805 -188.875 ;
        RECT 236.475 -190.565 236.805 -190.235 ;
        RECT 236.475 -191.925 236.805 -191.595 ;
        RECT 236.475 -193.285 236.805 -192.955 ;
        RECT 236.475 -194.645 236.805 -194.315 ;
        RECT 236.475 -196.005 236.805 -195.675 ;
        RECT 236.475 -197.365 236.805 -197.035 ;
        RECT 236.475 -198.725 236.805 -198.395 ;
        RECT 236.475 -200.085 236.805 -199.755 ;
        RECT 236.475 -201.445 236.805 -201.115 ;
        RECT 236.475 -202.805 236.805 -202.475 ;
        RECT 236.475 -204.165 236.805 -203.835 ;
        RECT 236.475 -205.525 236.805 -205.195 ;
        RECT 236.475 -206.885 236.805 -206.555 ;
        RECT 236.475 -208.245 236.805 -207.915 ;
        RECT 236.475 -209.605 236.805 -209.275 ;
        RECT 236.475 -210.965 236.805 -210.635 ;
        RECT 236.475 -212.325 236.805 -211.995 ;
        RECT 236.475 -213.685 236.805 -213.355 ;
        RECT 236.475 -215.045 236.805 -214.715 ;
        RECT 236.475 -216.405 236.805 -216.075 ;
        RECT 236.475 -217.765 236.805 -217.435 ;
        RECT 236.475 -219.125 236.805 -218.795 ;
        RECT 236.475 -220.485 236.805 -220.155 ;
        RECT 236.475 -221.845 236.805 -221.515 ;
        RECT 236.475 -223.205 236.805 -222.875 ;
        RECT 236.475 -224.565 236.805 -224.235 ;
        RECT 236.475 -225.925 236.805 -225.595 ;
        RECT 236.475 -227.285 236.805 -226.955 ;
        RECT 236.475 -228.645 236.805 -228.315 ;
        RECT 236.475 -230.005 236.805 -229.675 ;
        RECT 236.475 -231.365 236.805 -231.035 ;
        RECT 236.475 -232.725 236.805 -232.395 ;
        RECT 236.475 -234.085 236.805 -233.755 ;
        RECT 236.475 -235.445 236.805 -235.115 ;
        RECT 236.475 -236.805 236.805 -236.475 ;
        RECT 236.475 -238.165 236.805 -237.835 ;
        RECT 236.475 -243.81 236.805 -242.68 ;
        RECT 236.48 -243.925 236.8 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 246.76 238.165 247.89 ;
        RECT 237.835 241.915 238.165 242.245 ;
        RECT 237.835 240.555 238.165 240.885 ;
        RECT 237.835 239.195 238.165 239.525 ;
        RECT 237.835 237.835 238.165 238.165 ;
        RECT 237.84 237.16 238.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 -1.525 238.165 -1.195 ;
        RECT 237.835 -2.885 238.165 -2.555 ;
        RECT 237.84 -3.56 238.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 -122.565 238.165 -122.235 ;
        RECT 237.835 -123.925 238.165 -123.595 ;
        RECT 237.835 -125.285 238.165 -124.955 ;
        RECT 237.835 -126.645 238.165 -126.315 ;
        RECT 237.835 -128.005 238.165 -127.675 ;
        RECT 237.835 -129.365 238.165 -129.035 ;
        RECT 237.835 -130.725 238.165 -130.395 ;
        RECT 237.835 -132.085 238.165 -131.755 ;
        RECT 237.835 -133.445 238.165 -133.115 ;
        RECT 237.835 -134.805 238.165 -134.475 ;
        RECT 237.835 -136.165 238.165 -135.835 ;
        RECT 237.835 -137.525 238.165 -137.195 ;
        RECT 237.835 -138.885 238.165 -138.555 ;
        RECT 237.835 -140.245 238.165 -139.915 ;
        RECT 237.835 -141.605 238.165 -141.275 ;
        RECT 237.835 -142.965 238.165 -142.635 ;
        RECT 237.835 -144.325 238.165 -143.995 ;
        RECT 237.835 -145.685 238.165 -145.355 ;
        RECT 237.835 -147.045 238.165 -146.715 ;
        RECT 237.835 -148.405 238.165 -148.075 ;
        RECT 237.835 -149.765 238.165 -149.435 ;
        RECT 237.835 -151.125 238.165 -150.795 ;
        RECT 237.835 -152.485 238.165 -152.155 ;
        RECT 237.835 -153.845 238.165 -153.515 ;
        RECT 237.835 -155.205 238.165 -154.875 ;
        RECT 237.835 -156.565 238.165 -156.235 ;
        RECT 237.835 -157.925 238.165 -157.595 ;
        RECT 237.835 -159.285 238.165 -158.955 ;
        RECT 237.835 -160.645 238.165 -160.315 ;
        RECT 237.835 -162.005 238.165 -161.675 ;
        RECT 237.835 -163.365 238.165 -163.035 ;
        RECT 237.835 -164.725 238.165 -164.395 ;
        RECT 237.835 -166.085 238.165 -165.755 ;
        RECT 237.835 -167.445 238.165 -167.115 ;
        RECT 237.835 -168.805 238.165 -168.475 ;
        RECT 237.835 -170.165 238.165 -169.835 ;
        RECT 237.835 -171.525 238.165 -171.195 ;
        RECT 237.835 -172.885 238.165 -172.555 ;
        RECT 237.835 -174.245 238.165 -173.915 ;
        RECT 237.835 -175.605 238.165 -175.275 ;
        RECT 237.835 -176.965 238.165 -176.635 ;
        RECT 237.835 -178.325 238.165 -177.995 ;
        RECT 237.835 -179.685 238.165 -179.355 ;
        RECT 237.835 -181.045 238.165 -180.715 ;
        RECT 237.835 -182.405 238.165 -182.075 ;
        RECT 237.835 -183.765 238.165 -183.435 ;
        RECT 237.835 -185.125 238.165 -184.795 ;
        RECT 237.835 -186.485 238.165 -186.155 ;
        RECT 237.835 -187.845 238.165 -187.515 ;
        RECT 237.835 -189.205 238.165 -188.875 ;
        RECT 237.835 -190.565 238.165 -190.235 ;
        RECT 237.835 -191.925 238.165 -191.595 ;
        RECT 237.835 -193.285 238.165 -192.955 ;
        RECT 237.835 -194.645 238.165 -194.315 ;
        RECT 237.835 -196.005 238.165 -195.675 ;
        RECT 237.835 -197.365 238.165 -197.035 ;
        RECT 237.835 -198.725 238.165 -198.395 ;
        RECT 237.835 -200.085 238.165 -199.755 ;
        RECT 237.835 -201.445 238.165 -201.115 ;
        RECT 237.835 -202.805 238.165 -202.475 ;
        RECT 237.835 -204.165 238.165 -203.835 ;
        RECT 237.835 -205.525 238.165 -205.195 ;
        RECT 237.835 -206.885 238.165 -206.555 ;
        RECT 237.835 -208.245 238.165 -207.915 ;
        RECT 237.835 -209.605 238.165 -209.275 ;
        RECT 237.835 -210.965 238.165 -210.635 ;
        RECT 237.835 -212.325 238.165 -211.995 ;
        RECT 237.835 -213.685 238.165 -213.355 ;
        RECT 237.835 -215.045 238.165 -214.715 ;
        RECT 237.835 -216.405 238.165 -216.075 ;
        RECT 237.835 -217.765 238.165 -217.435 ;
        RECT 237.835 -219.125 238.165 -218.795 ;
        RECT 237.835 -220.485 238.165 -220.155 ;
        RECT 237.835 -221.845 238.165 -221.515 ;
        RECT 237.835 -223.205 238.165 -222.875 ;
        RECT 237.835 -224.565 238.165 -224.235 ;
        RECT 237.835 -225.925 238.165 -225.595 ;
        RECT 237.835 -227.285 238.165 -226.955 ;
        RECT 237.835 -228.645 238.165 -228.315 ;
        RECT 237.835 -230.005 238.165 -229.675 ;
        RECT 237.835 -231.365 238.165 -231.035 ;
        RECT 237.835 -232.725 238.165 -232.395 ;
        RECT 237.835 -234.085 238.165 -233.755 ;
        RECT 237.835 -235.445 238.165 -235.115 ;
        RECT 237.835 -236.805 238.165 -236.475 ;
        RECT 237.835 -238.165 238.165 -237.835 ;
        RECT 237.835 -243.81 238.165 -242.68 ;
        RECT 237.84 -243.925 238.16 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 246.76 239.525 247.89 ;
        RECT 239.195 241.915 239.525 242.245 ;
        RECT 239.195 240.555 239.525 240.885 ;
        RECT 239.195 239.195 239.525 239.525 ;
        RECT 239.195 237.835 239.525 238.165 ;
        RECT 239.2 237.16 239.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 -1.525 239.525 -1.195 ;
        RECT 239.195 -2.885 239.525 -2.555 ;
        RECT 239.2 -3.56 239.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 -122.565 239.525 -122.235 ;
        RECT 239.195 -123.925 239.525 -123.595 ;
        RECT 239.195 -125.285 239.525 -124.955 ;
        RECT 239.195 -126.645 239.525 -126.315 ;
        RECT 239.195 -128.005 239.525 -127.675 ;
        RECT 239.195 -129.365 239.525 -129.035 ;
        RECT 239.195 -130.725 239.525 -130.395 ;
        RECT 239.195 -132.085 239.525 -131.755 ;
        RECT 239.195 -133.445 239.525 -133.115 ;
        RECT 239.195 -134.805 239.525 -134.475 ;
        RECT 239.195 -136.165 239.525 -135.835 ;
        RECT 239.195 -137.525 239.525 -137.195 ;
        RECT 239.195 -138.885 239.525 -138.555 ;
        RECT 239.195 -140.245 239.525 -139.915 ;
        RECT 239.195 -141.605 239.525 -141.275 ;
        RECT 239.195 -142.965 239.525 -142.635 ;
        RECT 239.195 -144.325 239.525 -143.995 ;
        RECT 239.195 -145.685 239.525 -145.355 ;
        RECT 239.195 -147.045 239.525 -146.715 ;
        RECT 239.195 -148.405 239.525 -148.075 ;
        RECT 239.195 -149.765 239.525 -149.435 ;
        RECT 239.195 -151.125 239.525 -150.795 ;
        RECT 239.195 -152.485 239.525 -152.155 ;
        RECT 239.195 -153.845 239.525 -153.515 ;
        RECT 239.195 -155.205 239.525 -154.875 ;
        RECT 239.195 -156.565 239.525 -156.235 ;
        RECT 239.195 -157.925 239.525 -157.595 ;
        RECT 239.195 -159.285 239.525 -158.955 ;
        RECT 239.195 -160.645 239.525 -160.315 ;
        RECT 239.195 -162.005 239.525 -161.675 ;
        RECT 239.195 -163.365 239.525 -163.035 ;
        RECT 239.195 -164.725 239.525 -164.395 ;
        RECT 239.195 -166.085 239.525 -165.755 ;
        RECT 239.195 -167.445 239.525 -167.115 ;
        RECT 239.195 -168.805 239.525 -168.475 ;
        RECT 239.195 -170.165 239.525 -169.835 ;
        RECT 239.195 -171.525 239.525 -171.195 ;
        RECT 239.195 -172.885 239.525 -172.555 ;
        RECT 239.195 -174.245 239.525 -173.915 ;
        RECT 239.195 -175.605 239.525 -175.275 ;
        RECT 239.195 -176.965 239.525 -176.635 ;
        RECT 239.195 -178.325 239.525 -177.995 ;
        RECT 239.195 -179.685 239.525 -179.355 ;
        RECT 239.195 -181.045 239.525 -180.715 ;
        RECT 239.195 -182.405 239.525 -182.075 ;
        RECT 239.195 -183.765 239.525 -183.435 ;
        RECT 239.195 -185.125 239.525 -184.795 ;
        RECT 239.195 -186.485 239.525 -186.155 ;
        RECT 239.195 -187.845 239.525 -187.515 ;
        RECT 239.195 -189.205 239.525 -188.875 ;
        RECT 239.195 -190.565 239.525 -190.235 ;
        RECT 239.195 -191.925 239.525 -191.595 ;
        RECT 239.195 -193.285 239.525 -192.955 ;
        RECT 239.195 -194.645 239.525 -194.315 ;
        RECT 239.195 -196.005 239.525 -195.675 ;
        RECT 239.195 -197.365 239.525 -197.035 ;
        RECT 239.195 -198.725 239.525 -198.395 ;
        RECT 239.195 -200.085 239.525 -199.755 ;
        RECT 239.195 -201.445 239.525 -201.115 ;
        RECT 239.195 -202.805 239.525 -202.475 ;
        RECT 239.195 -204.165 239.525 -203.835 ;
        RECT 239.195 -205.525 239.525 -205.195 ;
        RECT 239.195 -206.885 239.525 -206.555 ;
        RECT 239.195 -208.245 239.525 -207.915 ;
        RECT 239.195 -209.605 239.525 -209.275 ;
        RECT 239.195 -210.965 239.525 -210.635 ;
        RECT 239.195 -212.325 239.525 -211.995 ;
        RECT 239.195 -213.685 239.525 -213.355 ;
        RECT 239.195 -215.045 239.525 -214.715 ;
        RECT 239.195 -216.405 239.525 -216.075 ;
        RECT 239.195 -217.765 239.525 -217.435 ;
        RECT 239.195 -219.125 239.525 -218.795 ;
        RECT 239.195 -220.485 239.525 -220.155 ;
        RECT 239.195 -221.845 239.525 -221.515 ;
        RECT 239.195 -223.205 239.525 -222.875 ;
        RECT 239.195 -224.565 239.525 -224.235 ;
        RECT 239.195 -225.925 239.525 -225.595 ;
        RECT 239.195 -227.285 239.525 -226.955 ;
        RECT 239.195 -228.645 239.525 -228.315 ;
        RECT 239.195 -230.005 239.525 -229.675 ;
        RECT 239.195 -231.365 239.525 -231.035 ;
        RECT 239.195 -232.725 239.525 -232.395 ;
        RECT 239.195 -234.085 239.525 -233.755 ;
        RECT 239.195 -235.445 239.525 -235.115 ;
        RECT 239.195 -236.805 239.525 -236.475 ;
        RECT 239.195 -238.165 239.525 -237.835 ;
        RECT 239.195 -243.81 239.525 -242.68 ;
        RECT 239.2 -243.925 239.52 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 246.76 240.885 247.89 ;
        RECT 240.555 241.915 240.885 242.245 ;
        RECT 240.555 240.555 240.885 240.885 ;
        RECT 240.555 239.195 240.885 239.525 ;
        RECT 240.555 237.835 240.885 238.165 ;
        RECT 240.56 237.16 240.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 -1.525 240.885 -1.195 ;
        RECT 240.555 -2.885 240.885 -2.555 ;
        RECT 240.56 -3.56 240.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 -122.565 240.885 -122.235 ;
        RECT 240.555 -123.925 240.885 -123.595 ;
        RECT 240.555 -125.285 240.885 -124.955 ;
        RECT 240.555 -126.645 240.885 -126.315 ;
        RECT 240.555 -128.005 240.885 -127.675 ;
        RECT 240.555 -129.365 240.885 -129.035 ;
        RECT 240.555 -130.725 240.885 -130.395 ;
        RECT 240.555 -132.085 240.885 -131.755 ;
        RECT 240.555 -133.445 240.885 -133.115 ;
        RECT 240.555 -134.805 240.885 -134.475 ;
        RECT 240.555 -136.165 240.885 -135.835 ;
        RECT 240.555 -137.525 240.885 -137.195 ;
        RECT 240.555 -138.885 240.885 -138.555 ;
        RECT 240.555 -140.245 240.885 -139.915 ;
        RECT 240.555 -141.605 240.885 -141.275 ;
        RECT 240.555 -142.965 240.885 -142.635 ;
        RECT 240.555 -144.325 240.885 -143.995 ;
        RECT 240.555 -145.685 240.885 -145.355 ;
        RECT 240.555 -147.045 240.885 -146.715 ;
        RECT 240.555 -148.405 240.885 -148.075 ;
        RECT 240.555 -149.765 240.885 -149.435 ;
        RECT 240.555 -151.125 240.885 -150.795 ;
        RECT 240.555 -152.485 240.885 -152.155 ;
        RECT 240.555 -153.845 240.885 -153.515 ;
        RECT 240.555 -155.205 240.885 -154.875 ;
        RECT 240.555 -156.565 240.885 -156.235 ;
        RECT 240.555 -157.925 240.885 -157.595 ;
        RECT 240.555 -159.285 240.885 -158.955 ;
        RECT 240.555 -160.645 240.885 -160.315 ;
        RECT 240.555 -162.005 240.885 -161.675 ;
        RECT 240.555 -163.365 240.885 -163.035 ;
        RECT 240.555 -164.725 240.885 -164.395 ;
        RECT 240.555 -166.085 240.885 -165.755 ;
        RECT 240.555 -167.445 240.885 -167.115 ;
        RECT 240.555 -168.805 240.885 -168.475 ;
        RECT 240.555 -170.165 240.885 -169.835 ;
        RECT 240.555 -171.525 240.885 -171.195 ;
        RECT 240.555 -172.885 240.885 -172.555 ;
        RECT 240.555 -174.245 240.885 -173.915 ;
        RECT 240.555 -175.605 240.885 -175.275 ;
        RECT 240.555 -176.965 240.885 -176.635 ;
        RECT 240.555 -178.325 240.885 -177.995 ;
        RECT 240.555 -179.685 240.885 -179.355 ;
        RECT 240.555 -181.045 240.885 -180.715 ;
        RECT 240.555 -182.405 240.885 -182.075 ;
        RECT 240.555 -183.765 240.885 -183.435 ;
        RECT 240.555 -185.125 240.885 -184.795 ;
        RECT 240.555 -186.485 240.885 -186.155 ;
        RECT 240.555 -187.845 240.885 -187.515 ;
        RECT 240.555 -189.205 240.885 -188.875 ;
        RECT 240.555 -190.565 240.885 -190.235 ;
        RECT 240.555 -191.925 240.885 -191.595 ;
        RECT 240.555 -193.285 240.885 -192.955 ;
        RECT 240.555 -194.645 240.885 -194.315 ;
        RECT 240.555 -196.005 240.885 -195.675 ;
        RECT 240.555 -197.365 240.885 -197.035 ;
        RECT 240.555 -198.725 240.885 -198.395 ;
        RECT 240.555 -200.085 240.885 -199.755 ;
        RECT 240.555 -201.445 240.885 -201.115 ;
        RECT 240.555 -202.805 240.885 -202.475 ;
        RECT 240.555 -204.165 240.885 -203.835 ;
        RECT 240.555 -205.525 240.885 -205.195 ;
        RECT 240.555 -206.885 240.885 -206.555 ;
        RECT 240.555 -208.245 240.885 -207.915 ;
        RECT 240.555 -209.605 240.885 -209.275 ;
        RECT 240.555 -210.965 240.885 -210.635 ;
        RECT 240.555 -212.325 240.885 -211.995 ;
        RECT 240.555 -213.685 240.885 -213.355 ;
        RECT 240.555 -215.045 240.885 -214.715 ;
        RECT 240.555 -216.405 240.885 -216.075 ;
        RECT 240.555 -217.765 240.885 -217.435 ;
        RECT 240.555 -219.125 240.885 -218.795 ;
        RECT 240.555 -220.485 240.885 -220.155 ;
        RECT 240.555 -221.845 240.885 -221.515 ;
        RECT 240.555 -223.205 240.885 -222.875 ;
        RECT 240.555 -224.565 240.885 -224.235 ;
        RECT 240.555 -225.925 240.885 -225.595 ;
        RECT 240.555 -227.285 240.885 -226.955 ;
        RECT 240.555 -228.645 240.885 -228.315 ;
        RECT 240.555 -230.005 240.885 -229.675 ;
        RECT 240.555 -231.365 240.885 -231.035 ;
        RECT 240.555 -232.725 240.885 -232.395 ;
        RECT 240.555 -234.085 240.885 -233.755 ;
        RECT 240.555 -235.445 240.885 -235.115 ;
        RECT 240.555 -236.805 240.885 -236.475 ;
        RECT 240.555 -238.165 240.885 -237.835 ;
        RECT 240.555 -243.81 240.885 -242.68 ;
        RECT 240.56 -243.925 240.88 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 246.76 242.245 247.89 ;
        RECT 241.915 241.915 242.245 242.245 ;
        RECT 241.915 240.555 242.245 240.885 ;
        RECT 241.915 239.195 242.245 239.525 ;
        RECT 241.915 237.835 242.245 238.165 ;
        RECT 241.92 237.16 242.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 -129.365 242.245 -129.035 ;
        RECT 241.915 -130.725 242.245 -130.395 ;
        RECT 241.915 -132.085 242.245 -131.755 ;
        RECT 241.915 -133.445 242.245 -133.115 ;
        RECT 241.915 -134.805 242.245 -134.475 ;
        RECT 241.915 -136.165 242.245 -135.835 ;
        RECT 241.915 -137.525 242.245 -137.195 ;
        RECT 241.915 -138.885 242.245 -138.555 ;
        RECT 241.915 -140.245 242.245 -139.915 ;
        RECT 241.915 -141.605 242.245 -141.275 ;
        RECT 241.915 -142.965 242.245 -142.635 ;
        RECT 241.915 -144.325 242.245 -143.995 ;
        RECT 241.915 -145.685 242.245 -145.355 ;
        RECT 241.915 -147.045 242.245 -146.715 ;
        RECT 241.915 -148.405 242.245 -148.075 ;
        RECT 241.915 -149.765 242.245 -149.435 ;
        RECT 241.915 -151.125 242.245 -150.795 ;
        RECT 241.915 -152.485 242.245 -152.155 ;
        RECT 241.915 -153.845 242.245 -153.515 ;
        RECT 241.915 -155.205 242.245 -154.875 ;
        RECT 241.915 -156.565 242.245 -156.235 ;
        RECT 241.915 -157.925 242.245 -157.595 ;
        RECT 241.915 -159.285 242.245 -158.955 ;
        RECT 241.915 -160.645 242.245 -160.315 ;
        RECT 241.915 -162.005 242.245 -161.675 ;
        RECT 241.915 -163.365 242.245 -163.035 ;
        RECT 241.915 -164.725 242.245 -164.395 ;
        RECT 241.915 -166.085 242.245 -165.755 ;
        RECT 241.915 -167.445 242.245 -167.115 ;
        RECT 241.915 -168.805 242.245 -168.475 ;
        RECT 241.915 -170.165 242.245 -169.835 ;
        RECT 241.915 -171.525 242.245 -171.195 ;
        RECT 241.915 -172.885 242.245 -172.555 ;
        RECT 241.915 -174.245 242.245 -173.915 ;
        RECT 241.915 -175.605 242.245 -175.275 ;
        RECT 241.915 -176.965 242.245 -176.635 ;
        RECT 241.915 -178.325 242.245 -177.995 ;
        RECT 241.915 -179.685 242.245 -179.355 ;
        RECT 241.915 -181.045 242.245 -180.715 ;
        RECT 241.915 -182.405 242.245 -182.075 ;
        RECT 241.915 -183.765 242.245 -183.435 ;
        RECT 241.915 -185.125 242.245 -184.795 ;
        RECT 241.915 -186.485 242.245 -186.155 ;
        RECT 241.915 -187.845 242.245 -187.515 ;
        RECT 241.915 -189.205 242.245 -188.875 ;
        RECT 241.915 -190.565 242.245 -190.235 ;
        RECT 241.915 -191.925 242.245 -191.595 ;
        RECT 241.915 -193.285 242.245 -192.955 ;
        RECT 241.915 -194.645 242.245 -194.315 ;
        RECT 241.915 -196.005 242.245 -195.675 ;
        RECT 241.915 -197.365 242.245 -197.035 ;
        RECT 241.915 -198.725 242.245 -198.395 ;
        RECT 241.915 -200.085 242.245 -199.755 ;
        RECT 241.915 -201.445 242.245 -201.115 ;
        RECT 241.915 -202.805 242.245 -202.475 ;
        RECT 241.915 -204.165 242.245 -203.835 ;
        RECT 241.915 -205.525 242.245 -205.195 ;
        RECT 241.915 -206.885 242.245 -206.555 ;
        RECT 241.915 -208.245 242.245 -207.915 ;
        RECT 241.915 -209.605 242.245 -209.275 ;
        RECT 241.915 -210.965 242.245 -210.635 ;
        RECT 241.915 -212.325 242.245 -211.995 ;
        RECT 241.915 -213.685 242.245 -213.355 ;
        RECT 241.915 -215.045 242.245 -214.715 ;
        RECT 241.915 -216.405 242.245 -216.075 ;
        RECT 241.915 -217.765 242.245 -217.435 ;
        RECT 241.915 -219.125 242.245 -218.795 ;
        RECT 241.915 -220.485 242.245 -220.155 ;
        RECT 241.915 -221.845 242.245 -221.515 ;
        RECT 241.915 -223.205 242.245 -222.875 ;
        RECT 241.915 -224.565 242.245 -224.235 ;
        RECT 241.915 -225.925 242.245 -225.595 ;
        RECT 241.915 -227.285 242.245 -226.955 ;
        RECT 241.915 -228.645 242.245 -228.315 ;
        RECT 241.915 -230.005 242.245 -229.675 ;
        RECT 241.915 -231.365 242.245 -231.035 ;
        RECT 241.915 -232.725 242.245 -232.395 ;
        RECT 241.915 -234.085 242.245 -233.755 ;
        RECT 241.915 -235.445 242.245 -235.115 ;
        RECT 241.915 -236.805 242.245 -236.475 ;
        RECT 241.915 -238.165 242.245 -237.835 ;
        RECT 241.915 -243.81 242.245 -242.68 ;
        RECT 241.92 -243.925 242.24 -126.315 ;
        RECT 241.915 -126.645 242.245 -126.315 ;
        RECT 241.915 -128.005 242.245 -127.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 246.76 208.245 247.89 ;
        RECT 207.915 241.915 208.245 242.245 ;
        RECT 207.915 240.555 208.245 240.885 ;
        RECT 207.915 239.195 208.245 239.525 ;
        RECT 207.915 237.835 208.245 238.165 ;
        RECT 207.92 237.16 208.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 -1.525 208.245 -1.195 ;
        RECT 207.915 -2.885 208.245 -2.555 ;
        RECT 207.92 -3.56 208.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 -122.565 208.245 -122.235 ;
        RECT 207.915 -123.925 208.245 -123.595 ;
        RECT 207.915 -125.285 208.245 -124.955 ;
        RECT 207.915 -126.645 208.245 -126.315 ;
        RECT 207.915 -128.005 208.245 -127.675 ;
        RECT 207.915 -129.365 208.245 -129.035 ;
        RECT 207.915 -130.725 208.245 -130.395 ;
        RECT 207.915 -132.085 208.245 -131.755 ;
        RECT 207.915 -133.445 208.245 -133.115 ;
        RECT 207.915 -134.805 208.245 -134.475 ;
        RECT 207.915 -136.165 208.245 -135.835 ;
        RECT 207.915 -137.525 208.245 -137.195 ;
        RECT 207.915 -138.885 208.245 -138.555 ;
        RECT 207.915 -140.245 208.245 -139.915 ;
        RECT 207.915 -141.605 208.245 -141.275 ;
        RECT 207.915 -142.965 208.245 -142.635 ;
        RECT 207.915 -144.325 208.245 -143.995 ;
        RECT 207.915 -145.685 208.245 -145.355 ;
        RECT 207.915 -147.045 208.245 -146.715 ;
        RECT 207.915 -148.405 208.245 -148.075 ;
        RECT 207.915 -149.765 208.245 -149.435 ;
        RECT 207.915 -151.125 208.245 -150.795 ;
        RECT 207.915 -152.485 208.245 -152.155 ;
        RECT 207.915 -153.845 208.245 -153.515 ;
        RECT 207.915 -155.205 208.245 -154.875 ;
        RECT 207.915 -156.565 208.245 -156.235 ;
        RECT 207.915 -157.925 208.245 -157.595 ;
        RECT 207.915 -159.285 208.245 -158.955 ;
        RECT 207.915 -160.645 208.245 -160.315 ;
        RECT 207.915 -162.005 208.245 -161.675 ;
        RECT 207.915 -163.365 208.245 -163.035 ;
        RECT 207.915 -164.725 208.245 -164.395 ;
        RECT 207.915 -166.085 208.245 -165.755 ;
        RECT 207.915 -167.445 208.245 -167.115 ;
        RECT 207.915 -168.805 208.245 -168.475 ;
        RECT 207.915 -170.165 208.245 -169.835 ;
        RECT 207.915 -171.525 208.245 -171.195 ;
        RECT 207.915 -172.885 208.245 -172.555 ;
        RECT 207.915 -174.245 208.245 -173.915 ;
        RECT 207.915 -175.605 208.245 -175.275 ;
        RECT 207.915 -176.965 208.245 -176.635 ;
        RECT 207.915 -178.325 208.245 -177.995 ;
        RECT 207.915 -179.685 208.245 -179.355 ;
        RECT 207.915 -181.045 208.245 -180.715 ;
        RECT 207.915 -182.405 208.245 -182.075 ;
        RECT 207.915 -183.765 208.245 -183.435 ;
        RECT 207.915 -185.125 208.245 -184.795 ;
        RECT 207.915 -186.485 208.245 -186.155 ;
        RECT 207.915 -187.845 208.245 -187.515 ;
        RECT 207.915 -189.205 208.245 -188.875 ;
        RECT 207.915 -190.565 208.245 -190.235 ;
        RECT 207.915 -191.925 208.245 -191.595 ;
        RECT 207.915 -193.285 208.245 -192.955 ;
        RECT 207.915 -194.645 208.245 -194.315 ;
        RECT 207.915 -196.005 208.245 -195.675 ;
        RECT 207.915 -197.365 208.245 -197.035 ;
        RECT 207.915 -198.725 208.245 -198.395 ;
        RECT 207.915 -200.085 208.245 -199.755 ;
        RECT 207.915 -201.445 208.245 -201.115 ;
        RECT 207.915 -202.805 208.245 -202.475 ;
        RECT 207.915 -204.165 208.245 -203.835 ;
        RECT 207.915 -205.525 208.245 -205.195 ;
        RECT 207.915 -206.885 208.245 -206.555 ;
        RECT 207.915 -208.245 208.245 -207.915 ;
        RECT 207.915 -209.605 208.245 -209.275 ;
        RECT 207.915 -210.965 208.245 -210.635 ;
        RECT 207.915 -212.325 208.245 -211.995 ;
        RECT 207.915 -213.685 208.245 -213.355 ;
        RECT 207.915 -215.045 208.245 -214.715 ;
        RECT 207.915 -216.405 208.245 -216.075 ;
        RECT 207.915 -217.765 208.245 -217.435 ;
        RECT 207.915 -219.125 208.245 -218.795 ;
        RECT 207.915 -220.485 208.245 -220.155 ;
        RECT 207.915 -221.845 208.245 -221.515 ;
        RECT 207.915 -223.205 208.245 -222.875 ;
        RECT 207.915 -224.565 208.245 -224.235 ;
        RECT 207.915 -225.925 208.245 -225.595 ;
        RECT 207.915 -227.285 208.245 -226.955 ;
        RECT 207.915 -228.645 208.245 -228.315 ;
        RECT 207.915 -230.005 208.245 -229.675 ;
        RECT 207.915 -231.365 208.245 -231.035 ;
        RECT 207.915 -232.725 208.245 -232.395 ;
        RECT 207.915 -234.085 208.245 -233.755 ;
        RECT 207.915 -235.445 208.245 -235.115 ;
        RECT 207.915 -236.805 208.245 -236.475 ;
        RECT 207.915 -238.165 208.245 -237.835 ;
        RECT 207.915 -243.81 208.245 -242.68 ;
        RECT 207.92 -243.925 208.24 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 246.76 209.605 247.89 ;
        RECT 209.275 241.915 209.605 242.245 ;
        RECT 209.275 240.555 209.605 240.885 ;
        RECT 209.275 239.195 209.605 239.525 ;
        RECT 209.275 237.835 209.605 238.165 ;
        RECT 209.28 237.16 209.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 -126.645 209.605 -126.315 ;
        RECT 209.275 -128.005 209.605 -127.675 ;
        RECT 209.275 -129.365 209.605 -129.035 ;
        RECT 209.275 -130.725 209.605 -130.395 ;
        RECT 209.275 -132.085 209.605 -131.755 ;
        RECT 209.275 -133.445 209.605 -133.115 ;
        RECT 209.275 -134.805 209.605 -134.475 ;
        RECT 209.275 -136.165 209.605 -135.835 ;
        RECT 209.275 -137.525 209.605 -137.195 ;
        RECT 209.275 -138.885 209.605 -138.555 ;
        RECT 209.275 -140.245 209.605 -139.915 ;
        RECT 209.275 -141.605 209.605 -141.275 ;
        RECT 209.275 -142.965 209.605 -142.635 ;
        RECT 209.275 -144.325 209.605 -143.995 ;
        RECT 209.275 -145.685 209.605 -145.355 ;
        RECT 209.275 -147.045 209.605 -146.715 ;
        RECT 209.275 -148.405 209.605 -148.075 ;
        RECT 209.275 -149.765 209.605 -149.435 ;
        RECT 209.275 -151.125 209.605 -150.795 ;
        RECT 209.275 -152.485 209.605 -152.155 ;
        RECT 209.275 -153.845 209.605 -153.515 ;
        RECT 209.275 -155.205 209.605 -154.875 ;
        RECT 209.275 -156.565 209.605 -156.235 ;
        RECT 209.275 -157.925 209.605 -157.595 ;
        RECT 209.275 -159.285 209.605 -158.955 ;
        RECT 209.275 -160.645 209.605 -160.315 ;
        RECT 209.275 -162.005 209.605 -161.675 ;
        RECT 209.275 -163.365 209.605 -163.035 ;
        RECT 209.275 -164.725 209.605 -164.395 ;
        RECT 209.275 -166.085 209.605 -165.755 ;
        RECT 209.275 -167.445 209.605 -167.115 ;
        RECT 209.275 -168.805 209.605 -168.475 ;
        RECT 209.275 -170.165 209.605 -169.835 ;
        RECT 209.275 -171.525 209.605 -171.195 ;
        RECT 209.275 -172.885 209.605 -172.555 ;
        RECT 209.275 -174.245 209.605 -173.915 ;
        RECT 209.275 -175.605 209.605 -175.275 ;
        RECT 209.275 -176.965 209.605 -176.635 ;
        RECT 209.275 -178.325 209.605 -177.995 ;
        RECT 209.275 -179.685 209.605 -179.355 ;
        RECT 209.275 -181.045 209.605 -180.715 ;
        RECT 209.275 -182.405 209.605 -182.075 ;
        RECT 209.275 -183.765 209.605 -183.435 ;
        RECT 209.275 -185.125 209.605 -184.795 ;
        RECT 209.275 -186.485 209.605 -186.155 ;
        RECT 209.275 -187.845 209.605 -187.515 ;
        RECT 209.275 -189.205 209.605 -188.875 ;
        RECT 209.275 -190.565 209.605 -190.235 ;
        RECT 209.275 -191.925 209.605 -191.595 ;
        RECT 209.275 -193.285 209.605 -192.955 ;
        RECT 209.275 -194.645 209.605 -194.315 ;
        RECT 209.275 -196.005 209.605 -195.675 ;
        RECT 209.275 -197.365 209.605 -197.035 ;
        RECT 209.275 -198.725 209.605 -198.395 ;
        RECT 209.275 -200.085 209.605 -199.755 ;
        RECT 209.275 -201.445 209.605 -201.115 ;
        RECT 209.275 -202.805 209.605 -202.475 ;
        RECT 209.275 -204.165 209.605 -203.835 ;
        RECT 209.275 -205.525 209.605 -205.195 ;
        RECT 209.275 -206.885 209.605 -206.555 ;
        RECT 209.275 -208.245 209.605 -207.915 ;
        RECT 209.275 -209.605 209.605 -209.275 ;
        RECT 209.275 -210.965 209.605 -210.635 ;
        RECT 209.275 -212.325 209.605 -211.995 ;
        RECT 209.275 -213.685 209.605 -213.355 ;
        RECT 209.275 -215.045 209.605 -214.715 ;
        RECT 209.275 -216.405 209.605 -216.075 ;
        RECT 209.275 -217.765 209.605 -217.435 ;
        RECT 209.275 -219.125 209.605 -218.795 ;
        RECT 209.275 -220.485 209.605 -220.155 ;
        RECT 209.275 -221.845 209.605 -221.515 ;
        RECT 209.275 -223.205 209.605 -222.875 ;
        RECT 209.275 -224.565 209.605 -224.235 ;
        RECT 209.275 -225.925 209.605 -225.595 ;
        RECT 209.275 -227.285 209.605 -226.955 ;
        RECT 209.275 -228.645 209.605 -228.315 ;
        RECT 209.275 -230.005 209.605 -229.675 ;
        RECT 209.275 -231.365 209.605 -231.035 ;
        RECT 209.275 -232.725 209.605 -232.395 ;
        RECT 209.275 -234.085 209.605 -233.755 ;
        RECT 209.275 -235.445 209.605 -235.115 ;
        RECT 209.275 -236.805 209.605 -236.475 ;
        RECT 209.275 -238.165 209.605 -237.835 ;
        RECT 209.275 -243.81 209.605 -242.68 ;
        RECT 209.28 -243.925 209.6 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.76 -125.535 210.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.635 246.76 210.965 247.89 ;
        RECT 210.635 241.915 210.965 242.245 ;
        RECT 210.635 240.555 210.965 240.885 ;
        RECT 210.635 239.195 210.965 239.525 ;
        RECT 210.635 237.835 210.965 238.165 ;
        RECT 210.64 237.16 210.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 246.76 212.325 247.89 ;
        RECT 211.995 241.915 212.325 242.245 ;
        RECT 211.995 240.555 212.325 240.885 ;
        RECT 211.995 239.195 212.325 239.525 ;
        RECT 211.995 237.835 212.325 238.165 ;
        RECT 212 237.16 212.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 -1.525 212.325 -1.195 ;
        RECT 211.995 -2.885 212.325 -2.555 ;
        RECT 212 -3.56 212.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 -122.565 212.325 -122.235 ;
        RECT 211.995 -123.925 212.325 -123.595 ;
        RECT 211.995 -125.285 212.325 -124.955 ;
        RECT 211.995 -126.645 212.325 -126.315 ;
        RECT 211.995 -128.005 212.325 -127.675 ;
        RECT 211.995 -129.365 212.325 -129.035 ;
        RECT 211.995 -130.725 212.325 -130.395 ;
        RECT 211.995 -132.085 212.325 -131.755 ;
        RECT 211.995 -133.445 212.325 -133.115 ;
        RECT 211.995 -134.805 212.325 -134.475 ;
        RECT 211.995 -136.165 212.325 -135.835 ;
        RECT 211.995 -137.525 212.325 -137.195 ;
        RECT 211.995 -138.885 212.325 -138.555 ;
        RECT 211.995 -140.245 212.325 -139.915 ;
        RECT 211.995 -141.605 212.325 -141.275 ;
        RECT 211.995 -142.965 212.325 -142.635 ;
        RECT 211.995 -144.325 212.325 -143.995 ;
        RECT 211.995 -145.685 212.325 -145.355 ;
        RECT 211.995 -147.045 212.325 -146.715 ;
        RECT 211.995 -148.405 212.325 -148.075 ;
        RECT 211.995 -149.765 212.325 -149.435 ;
        RECT 211.995 -151.125 212.325 -150.795 ;
        RECT 211.995 -152.485 212.325 -152.155 ;
        RECT 211.995 -153.845 212.325 -153.515 ;
        RECT 211.995 -155.205 212.325 -154.875 ;
        RECT 211.995 -156.565 212.325 -156.235 ;
        RECT 211.995 -157.925 212.325 -157.595 ;
        RECT 211.995 -159.285 212.325 -158.955 ;
        RECT 211.995 -160.645 212.325 -160.315 ;
        RECT 211.995 -162.005 212.325 -161.675 ;
        RECT 211.995 -163.365 212.325 -163.035 ;
        RECT 211.995 -164.725 212.325 -164.395 ;
        RECT 211.995 -166.085 212.325 -165.755 ;
        RECT 211.995 -167.445 212.325 -167.115 ;
        RECT 211.995 -168.805 212.325 -168.475 ;
        RECT 211.995 -170.165 212.325 -169.835 ;
        RECT 211.995 -171.525 212.325 -171.195 ;
        RECT 211.995 -172.885 212.325 -172.555 ;
        RECT 211.995 -174.245 212.325 -173.915 ;
        RECT 211.995 -175.605 212.325 -175.275 ;
        RECT 211.995 -176.965 212.325 -176.635 ;
        RECT 211.995 -178.325 212.325 -177.995 ;
        RECT 211.995 -179.685 212.325 -179.355 ;
        RECT 211.995 -181.045 212.325 -180.715 ;
        RECT 211.995 -182.405 212.325 -182.075 ;
        RECT 211.995 -183.765 212.325 -183.435 ;
        RECT 211.995 -185.125 212.325 -184.795 ;
        RECT 211.995 -186.485 212.325 -186.155 ;
        RECT 211.995 -187.845 212.325 -187.515 ;
        RECT 211.995 -189.205 212.325 -188.875 ;
        RECT 211.995 -190.565 212.325 -190.235 ;
        RECT 211.995 -191.925 212.325 -191.595 ;
        RECT 211.995 -193.285 212.325 -192.955 ;
        RECT 211.995 -194.645 212.325 -194.315 ;
        RECT 211.995 -196.005 212.325 -195.675 ;
        RECT 211.995 -197.365 212.325 -197.035 ;
        RECT 211.995 -198.725 212.325 -198.395 ;
        RECT 211.995 -200.085 212.325 -199.755 ;
        RECT 211.995 -201.445 212.325 -201.115 ;
        RECT 211.995 -202.805 212.325 -202.475 ;
        RECT 211.995 -204.165 212.325 -203.835 ;
        RECT 211.995 -205.525 212.325 -205.195 ;
        RECT 211.995 -206.885 212.325 -206.555 ;
        RECT 211.995 -208.245 212.325 -207.915 ;
        RECT 211.995 -209.605 212.325 -209.275 ;
        RECT 211.995 -210.965 212.325 -210.635 ;
        RECT 211.995 -212.325 212.325 -211.995 ;
        RECT 211.995 -213.685 212.325 -213.355 ;
        RECT 211.995 -215.045 212.325 -214.715 ;
        RECT 211.995 -216.405 212.325 -216.075 ;
        RECT 211.995 -217.765 212.325 -217.435 ;
        RECT 211.995 -219.125 212.325 -218.795 ;
        RECT 211.995 -220.485 212.325 -220.155 ;
        RECT 211.995 -221.845 212.325 -221.515 ;
        RECT 211.995 -223.205 212.325 -222.875 ;
        RECT 211.995 -224.565 212.325 -224.235 ;
        RECT 211.995 -225.925 212.325 -225.595 ;
        RECT 211.995 -227.285 212.325 -226.955 ;
        RECT 211.995 -228.645 212.325 -228.315 ;
        RECT 211.995 -230.005 212.325 -229.675 ;
        RECT 211.995 -231.365 212.325 -231.035 ;
        RECT 211.995 -232.725 212.325 -232.395 ;
        RECT 211.995 -234.085 212.325 -233.755 ;
        RECT 211.995 -235.445 212.325 -235.115 ;
        RECT 211.995 -236.805 212.325 -236.475 ;
        RECT 211.995 -238.165 212.325 -237.835 ;
        RECT 211.995 -243.81 212.325 -242.68 ;
        RECT 212 -243.925 212.32 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 246.76 213.685 247.89 ;
        RECT 213.355 241.915 213.685 242.245 ;
        RECT 213.355 240.555 213.685 240.885 ;
        RECT 213.355 239.195 213.685 239.525 ;
        RECT 213.355 237.835 213.685 238.165 ;
        RECT 213.36 237.16 213.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 -1.525 213.685 -1.195 ;
        RECT 213.355 -2.885 213.685 -2.555 ;
        RECT 213.36 -3.56 213.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 246.76 215.045 247.89 ;
        RECT 214.715 241.915 215.045 242.245 ;
        RECT 214.715 240.555 215.045 240.885 ;
        RECT 214.715 239.195 215.045 239.525 ;
        RECT 214.715 237.835 215.045 238.165 ;
        RECT 214.72 237.16 215.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 -1.525 215.045 -1.195 ;
        RECT 214.715 -2.885 215.045 -2.555 ;
        RECT 214.72 -3.56 215.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 -122.565 215.045 -122.235 ;
        RECT 214.715 -123.925 215.045 -123.595 ;
        RECT 214.715 -125.285 215.045 -124.955 ;
        RECT 214.715 -126.645 215.045 -126.315 ;
        RECT 214.715 -128.005 215.045 -127.675 ;
        RECT 214.715 -129.365 215.045 -129.035 ;
        RECT 214.715 -130.725 215.045 -130.395 ;
        RECT 214.715 -132.085 215.045 -131.755 ;
        RECT 214.715 -133.445 215.045 -133.115 ;
        RECT 214.715 -134.805 215.045 -134.475 ;
        RECT 214.715 -136.165 215.045 -135.835 ;
        RECT 214.715 -137.525 215.045 -137.195 ;
        RECT 214.715 -138.885 215.045 -138.555 ;
        RECT 214.715 -140.245 215.045 -139.915 ;
        RECT 214.715 -141.605 215.045 -141.275 ;
        RECT 214.715 -142.965 215.045 -142.635 ;
        RECT 214.715 -144.325 215.045 -143.995 ;
        RECT 214.715 -145.685 215.045 -145.355 ;
        RECT 214.715 -147.045 215.045 -146.715 ;
        RECT 214.715 -148.405 215.045 -148.075 ;
        RECT 214.715 -149.765 215.045 -149.435 ;
        RECT 214.715 -151.125 215.045 -150.795 ;
        RECT 214.715 -152.485 215.045 -152.155 ;
        RECT 214.715 -153.845 215.045 -153.515 ;
        RECT 214.715 -155.205 215.045 -154.875 ;
        RECT 214.715 -156.565 215.045 -156.235 ;
        RECT 214.715 -157.925 215.045 -157.595 ;
        RECT 214.715 -159.285 215.045 -158.955 ;
        RECT 214.715 -160.645 215.045 -160.315 ;
        RECT 214.715 -162.005 215.045 -161.675 ;
        RECT 214.715 -163.365 215.045 -163.035 ;
        RECT 214.715 -164.725 215.045 -164.395 ;
        RECT 214.715 -166.085 215.045 -165.755 ;
        RECT 214.715 -167.445 215.045 -167.115 ;
        RECT 214.715 -168.805 215.045 -168.475 ;
        RECT 214.715 -170.165 215.045 -169.835 ;
        RECT 214.715 -171.525 215.045 -171.195 ;
        RECT 214.715 -172.885 215.045 -172.555 ;
        RECT 214.715 -174.245 215.045 -173.915 ;
        RECT 214.715 -175.605 215.045 -175.275 ;
        RECT 214.715 -176.965 215.045 -176.635 ;
        RECT 214.715 -178.325 215.045 -177.995 ;
        RECT 214.715 -179.685 215.045 -179.355 ;
        RECT 214.715 -181.045 215.045 -180.715 ;
        RECT 214.715 -182.405 215.045 -182.075 ;
        RECT 214.715 -183.765 215.045 -183.435 ;
        RECT 214.715 -185.125 215.045 -184.795 ;
        RECT 214.715 -186.485 215.045 -186.155 ;
        RECT 214.715 -187.845 215.045 -187.515 ;
        RECT 214.715 -189.205 215.045 -188.875 ;
        RECT 214.715 -190.565 215.045 -190.235 ;
        RECT 214.715 -191.925 215.045 -191.595 ;
        RECT 214.715 -193.285 215.045 -192.955 ;
        RECT 214.715 -194.645 215.045 -194.315 ;
        RECT 214.715 -196.005 215.045 -195.675 ;
        RECT 214.715 -197.365 215.045 -197.035 ;
        RECT 214.715 -198.725 215.045 -198.395 ;
        RECT 214.715 -200.085 215.045 -199.755 ;
        RECT 214.715 -201.445 215.045 -201.115 ;
        RECT 214.715 -202.805 215.045 -202.475 ;
        RECT 214.715 -204.165 215.045 -203.835 ;
        RECT 214.715 -205.525 215.045 -205.195 ;
        RECT 214.715 -206.885 215.045 -206.555 ;
        RECT 214.715 -208.245 215.045 -207.915 ;
        RECT 214.715 -209.605 215.045 -209.275 ;
        RECT 214.715 -210.965 215.045 -210.635 ;
        RECT 214.715 -212.325 215.045 -211.995 ;
        RECT 214.715 -213.685 215.045 -213.355 ;
        RECT 214.715 -215.045 215.045 -214.715 ;
        RECT 214.715 -216.405 215.045 -216.075 ;
        RECT 214.715 -217.765 215.045 -217.435 ;
        RECT 214.715 -219.125 215.045 -218.795 ;
        RECT 214.715 -220.485 215.045 -220.155 ;
        RECT 214.715 -221.845 215.045 -221.515 ;
        RECT 214.715 -223.205 215.045 -222.875 ;
        RECT 214.715 -224.565 215.045 -224.235 ;
        RECT 214.715 -225.925 215.045 -225.595 ;
        RECT 214.715 -227.285 215.045 -226.955 ;
        RECT 214.715 -228.645 215.045 -228.315 ;
        RECT 214.715 -230.005 215.045 -229.675 ;
        RECT 214.715 -231.365 215.045 -231.035 ;
        RECT 214.715 -232.725 215.045 -232.395 ;
        RECT 214.715 -234.085 215.045 -233.755 ;
        RECT 214.715 -235.445 215.045 -235.115 ;
        RECT 214.715 -236.805 215.045 -236.475 ;
        RECT 214.715 -238.165 215.045 -237.835 ;
        RECT 214.715 -243.81 215.045 -242.68 ;
        RECT 214.72 -243.925 215.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 246.76 216.405 247.89 ;
        RECT 216.075 241.915 216.405 242.245 ;
        RECT 216.075 240.555 216.405 240.885 ;
        RECT 216.075 239.195 216.405 239.525 ;
        RECT 216.075 237.835 216.405 238.165 ;
        RECT 216.08 237.16 216.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 -1.525 216.405 -1.195 ;
        RECT 216.075 -2.885 216.405 -2.555 ;
        RECT 216.08 -3.56 216.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 -122.565 216.405 -122.235 ;
        RECT 216.075 -123.925 216.405 -123.595 ;
        RECT 216.075 -125.285 216.405 -124.955 ;
        RECT 216.075 -126.645 216.405 -126.315 ;
        RECT 216.075 -128.005 216.405 -127.675 ;
        RECT 216.075 -129.365 216.405 -129.035 ;
        RECT 216.075 -130.725 216.405 -130.395 ;
        RECT 216.075 -132.085 216.405 -131.755 ;
        RECT 216.075 -133.445 216.405 -133.115 ;
        RECT 216.075 -134.805 216.405 -134.475 ;
        RECT 216.075 -136.165 216.405 -135.835 ;
        RECT 216.075 -137.525 216.405 -137.195 ;
        RECT 216.075 -138.885 216.405 -138.555 ;
        RECT 216.075 -140.245 216.405 -139.915 ;
        RECT 216.075 -141.605 216.405 -141.275 ;
        RECT 216.075 -142.965 216.405 -142.635 ;
        RECT 216.075 -144.325 216.405 -143.995 ;
        RECT 216.075 -145.685 216.405 -145.355 ;
        RECT 216.075 -147.045 216.405 -146.715 ;
        RECT 216.075 -148.405 216.405 -148.075 ;
        RECT 216.075 -149.765 216.405 -149.435 ;
        RECT 216.075 -151.125 216.405 -150.795 ;
        RECT 216.075 -152.485 216.405 -152.155 ;
        RECT 216.075 -153.845 216.405 -153.515 ;
        RECT 216.075 -155.205 216.405 -154.875 ;
        RECT 216.075 -156.565 216.405 -156.235 ;
        RECT 216.075 -157.925 216.405 -157.595 ;
        RECT 216.075 -159.285 216.405 -158.955 ;
        RECT 216.075 -160.645 216.405 -160.315 ;
        RECT 216.075 -162.005 216.405 -161.675 ;
        RECT 216.075 -163.365 216.405 -163.035 ;
        RECT 216.075 -164.725 216.405 -164.395 ;
        RECT 216.075 -166.085 216.405 -165.755 ;
        RECT 216.075 -167.445 216.405 -167.115 ;
        RECT 216.075 -168.805 216.405 -168.475 ;
        RECT 216.075 -170.165 216.405 -169.835 ;
        RECT 216.075 -171.525 216.405 -171.195 ;
        RECT 216.075 -172.885 216.405 -172.555 ;
        RECT 216.075 -174.245 216.405 -173.915 ;
        RECT 216.075 -175.605 216.405 -175.275 ;
        RECT 216.075 -176.965 216.405 -176.635 ;
        RECT 216.075 -178.325 216.405 -177.995 ;
        RECT 216.075 -179.685 216.405 -179.355 ;
        RECT 216.075 -181.045 216.405 -180.715 ;
        RECT 216.075 -182.405 216.405 -182.075 ;
        RECT 216.075 -183.765 216.405 -183.435 ;
        RECT 216.075 -185.125 216.405 -184.795 ;
        RECT 216.075 -186.485 216.405 -186.155 ;
        RECT 216.075 -187.845 216.405 -187.515 ;
        RECT 216.075 -189.205 216.405 -188.875 ;
        RECT 216.075 -190.565 216.405 -190.235 ;
        RECT 216.075 -191.925 216.405 -191.595 ;
        RECT 216.075 -193.285 216.405 -192.955 ;
        RECT 216.075 -194.645 216.405 -194.315 ;
        RECT 216.075 -196.005 216.405 -195.675 ;
        RECT 216.075 -197.365 216.405 -197.035 ;
        RECT 216.075 -198.725 216.405 -198.395 ;
        RECT 216.075 -200.085 216.405 -199.755 ;
        RECT 216.075 -201.445 216.405 -201.115 ;
        RECT 216.075 -202.805 216.405 -202.475 ;
        RECT 216.075 -204.165 216.405 -203.835 ;
        RECT 216.075 -205.525 216.405 -205.195 ;
        RECT 216.075 -206.885 216.405 -206.555 ;
        RECT 216.075 -208.245 216.405 -207.915 ;
        RECT 216.075 -209.605 216.405 -209.275 ;
        RECT 216.075 -210.965 216.405 -210.635 ;
        RECT 216.075 -212.325 216.405 -211.995 ;
        RECT 216.075 -213.685 216.405 -213.355 ;
        RECT 216.075 -215.045 216.405 -214.715 ;
        RECT 216.075 -216.405 216.405 -216.075 ;
        RECT 216.075 -217.765 216.405 -217.435 ;
        RECT 216.075 -219.125 216.405 -218.795 ;
        RECT 216.075 -220.485 216.405 -220.155 ;
        RECT 216.075 -221.845 216.405 -221.515 ;
        RECT 216.075 -223.205 216.405 -222.875 ;
        RECT 216.075 -224.565 216.405 -224.235 ;
        RECT 216.075 -225.925 216.405 -225.595 ;
        RECT 216.075 -227.285 216.405 -226.955 ;
        RECT 216.075 -228.645 216.405 -228.315 ;
        RECT 216.075 -230.005 216.405 -229.675 ;
        RECT 216.075 -231.365 216.405 -231.035 ;
        RECT 216.075 -232.725 216.405 -232.395 ;
        RECT 216.075 -234.085 216.405 -233.755 ;
        RECT 216.075 -235.445 216.405 -235.115 ;
        RECT 216.075 -236.805 216.405 -236.475 ;
        RECT 216.075 -238.165 216.405 -237.835 ;
        RECT 216.075 -243.81 216.405 -242.68 ;
        RECT 216.08 -243.925 216.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 246.76 217.765 247.89 ;
        RECT 217.435 241.915 217.765 242.245 ;
        RECT 217.435 240.555 217.765 240.885 ;
        RECT 217.435 239.195 217.765 239.525 ;
        RECT 217.435 237.835 217.765 238.165 ;
        RECT 217.44 237.16 217.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 -1.525 217.765 -1.195 ;
        RECT 217.435 -2.885 217.765 -2.555 ;
        RECT 217.44 -3.56 217.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 -122.565 217.765 -122.235 ;
        RECT 217.435 -123.925 217.765 -123.595 ;
        RECT 217.435 -125.285 217.765 -124.955 ;
        RECT 217.435 -126.645 217.765 -126.315 ;
        RECT 217.435 -128.005 217.765 -127.675 ;
        RECT 217.435 -129.365 217.765 -129.035 ;
        RECT 217.435 -130.725 217.765 -130.395 ;
        RECT 217.435 -132.085 217.765 -131.755 ;
        RECT 217.435 -133.445 217.765 -133.115 ;
        RECT 217.435 -134.805 217.765 -134.475 ;
        RECT 217.435 -136.165 217.765 -135.835 ;
        RECT 217.435 -137.525 217.765 -137.195 ;
        RECT 217.435 -138.885 217.765 -138.555 ;
        RECT 217.435 -140.245 217.765 -139.915 ;
        RECT 217.435 -141.605 217.765 -141.275 ;
        RECT 217.435 -142.965 217.765 -142.635 ;
        RECT 217.435 -144.325 217.765 -143.995 ;
        RECT 217.435 -145.685 217.765 -145.355 ;
        RECT 217.435 -147.045 217.765 -146.715 ;
        RECT 217.435 -148.405 217.765 -148.075 ;
        RECT 217.435 -149.765 217.765 -149.435 ;
        RECT 217.435 -151.125 217.765 -150.795 ;
        RECT 217.435 -152.485 217.765 -152.155 ;
        RECT 217.435 -153.845 217.765 -153.515 ;
        RECT 217.435 -155.205 217.765 -154.875 ;
        RECT 217.435 -156.565 217.765 -156.235 ;
        RECT 217.435 -157.925 217.765 -157.595 ;
        RECT 217.435 -159.285 217.765 -158.955 ;
        RECT 217.435 -160.645 217.765 -160.315 ;
        RECT 217.435 -162.005 217.765 -161.675 ;
        RECT 217.435 -163.365 217.765 -163.035 ;
        RECT 217.435 -164.725 217.765 -164.395 ;
        RECT 217.435 -166.085 217.765 -165.755 ;
        RECT 217.435 -167.445 217.765 -167.115 ;
        RECT 217.435 -168.805 217.765 -168.475 ;
        RECT 217.435 -170.165 217.765 -169.835 ;
        RECT 217.435 -171.525 217.765 -171.195 ;
        RECT 217.435 -172.885 217.765 -172.555 ;
        RECT 217.435 -174.245 217.765 -173.915 ;
        RECT 217.435 -175.605 217.765 -175.275 ;
        RECT 217.435 -176.965 217.765 -176.635 ;
        RECT 217.435 -178.325 217.765 -177.995 ;
        RECT 217.435 -179.685 217.765 -179.355 ;
        RECT 217.435 -181.045 217.765 -180.715 ;
        RECT 217.435 -182.405 217.765 -182.075 ;
        RECT 217.435 -183.765 217.765 -183.435 ;
        RECT 217.435 -185.125 217.765 -184.795 ;
        RECT 217.435 -186.485 217.765 -186.155 ;
        RECT 217.435 -187.845 217.765 -187.515 ;
        RECT 217.435 -189.205 217.765 -188.875 ;
        RECT 217.435 -190.565 217.765 -190.235 ;
        RECT 217.435 -191.925 217.765 -191.595 ;
        RECT 217.435 -193.285 217.765 -192.955 ;
        RECT 217.435 -194.645 217.765 -194.315 ;
        RECT 217.435 -196.005 217.765 -195.675 ;
        RECT 217.435 -197.365 217.765 -197.035 ;
        RECT 217.435 -198.725 217.765 -198.395 ;
        RECT 217.435 -200.085 217.765 -199.755 ;
        RECT 217.435 -201.445 217.765 -201.115 ;
        RECT 217.435 -202.805 217.765 -202.475 ;
        RECT 217.435 -204.165 217.765 -203.835 ;
        RECT 217.435 -205.525 217.765 -205.195 ;
        RECT 217.435 -206.885 217.765 -206.555 ;
        RECT 217.435 -208.245 217.765 -207.915 ;
        RECT 217.435 -209.605 217.765 -209.275 ;
        RECT 217.435 -210.965 217.765 -210.635 ;
        RECT 217.435 -212.325 217.765 -211.995 ;
        RECT 217.435 -213.685 217.765 -213.355 ;
        RECT 217.435 -215.045 217.765 -214.715 ;
        RECT 217.435 -216.405 217.765 -216.075 ;
        RECT 217.435 -217.765 217.765 -217.435 ;
        RECT 217.435 -219.125 217.765 -218.795 ;
        RECT 217.435 -220.485 217.765 -220.155 ;
        RECT 217.435 -221.845 217.765 -221.515 ;
        RECT 217.435 -223.205 217.765 -222.875 ;
        RECT 217.435 -224.565 217.765 -224.235 ;
        RECT 217.435 -225.925 217.765 -225.595 ;
        RECT 217.435 -227.285 217.765 -226.955 ;
        RECT 217.435 -228.645 217.765 -228.315 ;
        RECT 217.435 -230.005 217.765 -229.675 ;
        RECT 217.435 -231.365 217.765 -231.035 ;
        RECT 217.435 -232.725 217.765 -232.395 ;
        RECT 217.435 -234.085 217.765 -233.755 ;
        RECT 217.435 -235.445 217.765 -235.115 ;
        RECT 217.435 -236.805 217.765 -236.475 ;
        RECT 217.435 -238.165 217.765 -237.835 ;
        RECT 217.435 -243.81 217.765 -242.68 ;
        RECT 217.44 -243.925 217.76 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 246.76 219.125 247.89 ;
        RECT 218.795 241.915 219.125 242.245 ;
        RECT 218.795 240.555 219.125 240.885 ;
        RECT 218.795 239.195 219.125 239.525 ;
        RECT 218.795 237.835 219.125 238.165 ;
        RECT 218.8 237.16 219.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 -1.525 219.125 -1.195 ;
        RECT 218.795 -2.885 219.125 -2.555 ;
        RECT 218.8 -3.56 219.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 -122.565 219.125 -122.235 ;
        RECT 218.795 -123.925 219.125 -123.595 ;
        RECT 218.795 -125.285 219.125 -124.955 ;
        RECT 218.795 -126.645 219.125 -126.315 ;
        RECT 218.795 -128.005 219.125 -127.675 ;
        RECT 218.795 -129.365 219.125 -129.035 ;
        RECT 218.795 -130.725 219.125 -130.395 ;
        RECT 218.795 -132.085 219.125 -131.755 ;
        RECT 218.795 -133.445 219.125 -133.115 ;
        RECT 218.795 -134.805 219.125 -134.475 ;
        RECT 218.795 -136.165 219.125 -135.835 ;
        RECT 218.795 -137.525 219.125 -137.195 ;
        RECT 218.795 -138.885 219.125 -138.555 ;
        RECT 218.795 -140.245 219.125 -139.915 ;
        RECT 218.795 -141.605 219.125 -141.275 ;
        RECT 218.795 -142.965 219.125 -142.635 ;
        RECT 218.795 -144.325 219.125 -143.995 ;
        RECT 218.795 -145.685 219.125 -145.355 ;
        RECT 218.795 -147.045 219.125 -146.715 ;
        RECT 218.795 -148.405 219.125 -148.075 ;
        RECT 218.795 -149.765 219.125 -149.435 ;
        RECT 218.795 -151.125 219.125 -150.795 ;
        RECT 218.795 -152.485 219.125 -152.155 ;
        RECT 218.795 -153.845 219.125 -153.515 ;
        RECT 218.795 -155.205 219.125 -154.875 ;
        RECT 218.795 -156.565 219.125 -156.235 ;
        RECT 218.795 -157.925 219.125 -157.595 ;
        RECT 218.795 -159.285 219.125 -158.955 ;
        RECT 218.795 -160.645 219.125 -160.315 ;
        RECT 218.795 -162.005 219.125 -161.675 ;
        RECT 218.795 -163.365 219.125 -163.035 ;
        RECT 218.795 -164.725 219.125 -164.395 ;
        RECT 218.795 -166.085 219.125 -165.755 ;
        RECT 218.795 -167.445 219.125 -167.115 ;
        RECT 218.795 -168.805 219.125 -168.475 ;
        RECT 218.795 -170.165 219.125 -169.835 ;
        RECT 218.795 -171.525 219.125 -171.195 ;
        RECT 218.795 -172.885 219.125 -172.555 ;
        RECT 218.795 -174.245 219.125 -173.915 ;
        RECT 218.795 -175.605 219.125 -175.275 ;
        RECT 218.795 -176.965 219.125 -176.635 ;
        RECT 218.795 -178.325 219.125 -177.995 ;
        RECT 218.795 -179.685 219.125 -179.355 ;
        RECT 218.795 -181.045 219.125 -180.715 ;
        RECT 218.795 -182.405 219.125 -182.075 ;
        RECT 218.795 -183.765 219.125 -183.435 ;
        RECT 218.795 -185.125 219.125 -184.795 ;
        RECT 218.795 -186.485 219.125 -186.155 ;
        RECT 218.795 -187.845 219.125 -187.515 ;
        RECT 218.795 -189.205 219.125 -188.875 ;
        RECT 218.795 -190.565 219.125 -190.235 ;
        RECT 218.795 -191.925 219.125 -191.595 ;
        RECT 218.795 -193.285 219.125 -192.955 ;
        RECT 218.795 -194.645 219.125 -194.315 ;
        RECT 218.795 -196.005 219.125 -195.675 ;
        RECT 218.795 -197.365 219.125 -197.035 ;
        RECT 218.795 -198.725 219.125 -198.395 ;
        RECT 218.795 -200.085 219.125 -199.755 ;
        RECT 218.795 -201.445 219.125 -201.115 ;
        RECT 218.795 -202.805 219.125 -202.475 ;
        RECT 218.795 -204.165 219.125 -203.835 ;
        RECT 218.795 -205.525 219.125 -205.195 ;
        RECT 218.795 -206.885 219.125 -206.555 ;
        RECT 218.795 -208.245 219.125 -207.915 ;
        RECT 218.795 -209.605 219.125 -209.275 ;
        RECT 218.795 -210.965 219.125 -210.635 ;
        RECT 218.795 -212.325 219.125 -211.995 ;
        RECT 218.795 -213.685 219.125 -213.355 ;
        RECT 218.795 -215.045 219.125 -214.715 ;
        RECT 218.795 -216.405 219.125 -216.075 ;
        RECT 218.795 -217.765 219.125 -217.435 ;
        RECT 218.795 -219.125 219.125 -218.795 ;
        RECT 218.795 -220.485 219.125 -220.155 ;
        RECT 218.795 -221.845 219.125 -221.515 ;
        RECT 218.795 -223.205 219.125 -222.875 ;
        RECT 218.795 -224.565 219.125 -224.235 ;
        RECT 218.795 -225.925 219.125 -225.595 ;
        RECT 218.795 -227.285 219.125 -226.955 ;
        RECT 218.795 -228.645 219.125 -228.315 ;
        RECT 218.795 -230.005 219.125 -229.675 ;
        RECT 218.795 -231.365 219.125 -231.035 ;
        RECT 218.795 -232.725 219.125 -232.395 ;
        RECT 218.795 -234.085 219.125 -233.755 ;
        RECT 218.795 -235.445 219.125 -235.115 ;
        RECT 218.795 -236.805 219.125 -236.475 ;
        RECT 218.795 -238.165 219.125 -237.835 ;
        RECT 218.795 -243.81 219.125 -242.68 ;
        RECT 218.8 -243.925 219.12 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 246.76 220.485 247.89 ;
        RECT 220.155 241.915 220.485 242.245 ;
        RECT 220.155 240.555 220.485 240.885 ;
        RECT 220.155 239.195 220.485 239.525 ;
        RECT 220.155 237.835 220.485 238.165 ;
        RECT 220.16 237.16 220.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 -126.645 220.485 -126.315 ;
        RECT 220.155 -128.005 220.485 -127.675 ;
        RECT 220.155 -129.365 220.485 -129.035 ;
        RECT 220.155 -130.725 220.485 -130.395 ;
        RECT 220.155 -132.085 220.485 -131.755 ;
        RECT 220.155 -133.445 220.485 -133.115 ;
        RECT 220.155 -134.805 220.485 -134.475 ;
        RECT 220.155 -136.165 220.485 -135.835 ;
        RECT 220.155 -137.525 220.485 -137.195 ;
        RECT 220.155 -138.885 220.485 -138.555 ;
        RECT 220.155 -140.245 220.485 -139.915 ;
        RECT 220.155 -141.605 220.485 -141.275 ;
        RECT 220.155 -142.965 220.485 -142.635 ;
        RECT 220.155 -144.325 220.485 -143.995 ;
        RECT 220.155 -145.685 220.485 -145.355 ;
        RECT 220.155 -147.045 220.485 -146.715 ;
        RECT 220.155 -148.405 220.485 -148.075 ;
        RECT 220.155 -149.765 220.485 -149.435 ;
        RECT 220.155 -151.125 220.485 -150.795 ;
        RECT 220.155 -152.485 220.485 -152.155 ;
        RECT 220.155 -153.845 220.485 -153.515 ;
        RECT 220.155 -155.205 220.485 -154.875 ;
        RECT 220.155 -156.565 220.485 -156.235 ;
        RECT 220.155 -157.925 220.485 -157.595 ;
        RECT 220.155 -159.285 220.485 -158.955 ;
        RECT 220.155 -160.645 220.485 -160.315 ;
        RECT 220.155 -162.005 220.485 -161.675 ;
        RECT 220.155 -163.365 220.485 -163.035 ;
        RECT 220.155 -164.725 220.485 -164.395 ;
        RECT 220.155 -166.085 220.485 -165.755 ;
        RECT 220.155 -167.445 220.485 -167.115 ;
        RECT 220.155 -168.805 220.485 -168.475 ;
        RECT 220.155 -170.165 220.485 -169.835 ;
        RECT 220.155 -171.525 220.485 -171.195 ;
        RECT 220.155 -172.885 220.485 -172.555 ;
        RECT 220.155 -174.245 220.485 -173.915 ;
        RECT 220.155 -175.605 220.485 -175.275 ;
        RECT 220.155 -176.965 220.485 -176.635 ;
        RECT 220.155 -178.325 220.485 -177.995 ;
        RECT 220.155 -179.685 220.485 -179.355 ;
        RECT 220.155 -181.045 220.485 -180.715 ;
        RECT 220.155 -182.405 220.485 -182.075 ;
        RECT 220.155 -183.765 220.485 -183.435 ;
        RECT 220.155 -185.125 220.485 -184.795 ;
        RECT 220.155 -186.485 220.485 -186.155 ;
        RECT 220.155 -187.845 220.485 -187.515 ;
        RECT 220.155 -189.205 220.485 -188.875 ;
        RECT 220.155 -190.565 220.485 -190.235 ;
        RECT 220.155 -191.925 220.485 -191.595 ;
        RECT 220.155 -193.285 220.485 -192.955 ;
        RECT 220.155 -194.645 220.485 -194.315 ;
        RECT 220.155 -196.005 220.485 -195.675 ;
        RECT 220.155 -197.365 220.485 -197.035 ;
        RECT 220.155 -198.725 220.485 -198.395 ;
        RECT 220.155 -200.085 220.485 -199.755 ;
        RECT 220.155 -201.445 220.485 -201.115 ;
        RECT 220.155 -202.805 220.485 -202.475 ;
        RECT 220.155 -204.165 220.485 -203.835 ;
        RECT 220.155 -205.525 220.485 -205.195 ;
        RECT 220.155 -206.885 220.485 -206.555 ;
        RECT 220.155 -208.245 220.485 -207.915 ;
        RECT 220.155 -209.605 220.485 -209.275 ;
        RECT 220.155 -210.965 220.485 -210.635 ;
        RECT 220.155 -212.325 220.485 -211.995 ;
        RECT 220.155 -213.685 220.485 -213.355 ;
        RECT 220.155 -215.045 220.485 -214.715 ;
        RECT 220.155 -216.405 220.485 -216.075 ;
        RECT 220.155 -217.765 220.485 -217.435 ;
        RECT 220.155 -219.125 220.485 -218.795 ;
        RECT 220.155 -220.485 220.485 -220.155 ;
        RECT 220.155 -221.845 220.485 -221.515 ;
        RECT 220.155 -223.205 220.485 -222.875 ;
        RECT 220.155 -224.565 220.485 -224.235 ;
        RECT 220.155 -225.925 220.485 -225.595 ;
        RECT 220.155 -227.285 220.485 -226.955 ;
        RECT 220.155 -228.645 220.485 -228.315 ;
        RECT 220.155 -230.005 220.485 -229.675 ;
        RECT 220.155 -231.365 220.485 -231.035 ;
        RECT 220.155 -232.725 220.485 -232.395 ;
        RECT 220.155 -234.085 220.485 -233.755 ;
        RECT 220.155 -235.445 220.485 -235.115 ;
        RECT 220.155 -236.805 220.485 -236.475 ;
        RECT 220.155 -238.165 220.485 -237.835 ;
        RECT 220.155 -243.81 220.485 -242.68 ;
        RECT 220.16 -243.925 220.48 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.66 -125.535 220.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.515 246.76 221.845 247.89 ;
        RECT 221.515 241.915 221.845 242.245 ;
        RECT 221.515 240.555 221.845 240.885 ;
        RECT 221.515 239.195 221.845 239.525 ;
        RECT 221.515 237.835 221.845 238.165 ;
        RECT 221.52 237.16 221.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 246.76 223.205 247.89 ;
        RECT 222.875 241.915 223.205 242.245 ;
        RECT 222.875 240.555 223.205 240.885 ;
        RECT 222.875 239.195 223.205 239.525 ;
        RECT 222.875 237.835 223.205 238.165 ;
        RECT 222.88 237.16 223.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 -1.525 223.205 -1.195 ;
        RECT 222.875 -2.885 223.205 -2.555 ;
        RECT 222.88 -3.56 223.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 -122.565 223.205 -122.235 ;
        RECT 222.875 -123.925 223.205 -123.595 ;
        RECT 222.875 -125.285 223.205 -124.955 ;
        RECT 222.875 -126.645 223.205 -126.315 ;
        RECT 222.875 -128.005 223.205 -127.675 ;
        RECT 222.875 -129.365 223.205 -129.035 ;
        RECT 222.875 -130.725 223.205 -130.395 ;
        RECT 222.875 -132.085 223.205 -131.755 ;
        RECT 222.875 -133.445 223.205 -133.115 ;
        RECT 222.875 -134.805 223.205 -134.475 ;
        RECT 222.875 -136.165 223.205 -135.835 ;
        RECT 222.875 -137.525 223.205 -137.195 ;
        RECT 222.875 -138.885 223.205 -138.555 ;
        RECT 222.875 -140.245 223.205 -139.915 ;
        RECT 222.875 -141.605 223.205 -141.275 ;
        RECT 222.875 -142.965 223.205 -142.635 ;
        RECT 222.875 -144.325 223.205 -143.995 ;
        RECT 222.875 -145.685 223.205 -145.355 ;
        RECT 222.875 -147.045 223.205 -146.715 ;
        RECT 222.875 -148.405 223.205 -148.075 ;
        RECT 222.875 -149.765 223.205 -149.435 ;
        RECT 222.875 -151.125 223.205 -150.795 ;
        RECT 222.875 -152.485 223.205 -152.155 ;
        RECT 222.875 -153.845 223.205 -153.515 ;
        RECT 222.875 -155.205 223.205 -154.875 ;
        RECT 222.875 -156.565 223.205 -156.235 ;
        RECT 222.875 -157.925 223.205 -157.595 ;
        RECT 222.875 -159.285 223.205 -158.955 ;
        RECT 222.875 -160.645 223.205 -160.315 ;
        RECT 222.875 -162.005 223.205 -161.675 ;
        RECT 222.875 -163.365 223.205 -163.035 ;
        RECT 222.875 -164.725 223.205 -164.395 ;
        RECT 222.875 -166.085 223.205 -165.755 ;
        RECT 222.875 -167.445 223.205 -167.115 ;
        RECT 222.875 -168.805 223.205 -168.475 ;
        RECT 222.875 -170.165 223.205 -169.835 ;
        RECT 222.875 -171.525 223.205 -171.195 ;
        RECT 222.875 -172.885 223.205 -172.555 ;
        RECT 222.875 -174.245 223.205 -173.915 ;
        RECT 222.875 -175.605 223.205 -175.275 ;
        RECT 222.875 -176.965 223.205 -176.635 ;
        RECT 222.875 -178.325 223.205 -177.995 ;
        RECT 222.875 -179.685 223.205 -179.355 ;
        RECT 222.875 -181.045 223.205 -180.715 ;
        RECT 222.875 -182.405 223.205 -182.075 ;
        RECT 222.875 -183.765 223.205 -183.435 ;
        RECT 222.875 -185.125 223.205 -184.795 ;
        RECT 222.875 -186.485 223.205 -186.155 ;
        RECT 222.875 -187.845 223.205 -187.515 ;
        RECT 222.875 -189.205 223.205 -188.875 ;
        RECT 222.875 -190.565 223.205 -190.235 ;
        RECT 222.875 -191.925 223.205 -191.595 ;
        RECT 222.875 -193.285 223.205 -192.955 ;
        RECT 222.875 -194.645 223.205 -194.315 ;
        RECT 222.875 -196.005 223.205 -195.675 ;
        RECT 222.875 -197.365 223.205 -197.035 ;
        RECT 222.875 -198.725 223.205 -198.395 ;
        RECT 222.875 -200.085 223.205 -199.755 ;
        RECT 222.875 -201.445 223.205 -201.115 ;
        RECT 222.875 -202.805 223.205 -202.475 ;
        RECT 222.875 -204.165 223.205 -203.835 ;
        RECT 222.875 -205.525 223.205 -205.195 ;
        RECT 222.875 -206.885 223.205 -206.555 ;
        RECT 222.875 -208.245 223.205 -207.915 ;
        RECT 222.875 -209.605 223.205 -209.275 ;
        RECT 222.875 -210.965 223.205 -210.635 ;
        RECT 222.875 -212.325 223.205 -211.995 ;
        RECT 222.875 -213.685 223.205 -213.355 ;
        RECT 222.875 -215.045 223.205 -214.715 ;
        RECT 222.875 -216.405 223.205 -216.075 ;
        RECT 222.875 -217.765 223.205 -217.435 ;
        RECT 222.875 -219.125 223.205 -218.795 ;
        RECT 222.875 -220.485 223.205 -220.155 ;
        RECT 222.875 -221.845 223.205 -221.515 ;
        RECT 222.875 -223.205 223.205 -222.875 ;
        RECT 222.875 -224.565 223.205 -224.235 ;
        RECT 222.875 -225.925 223.205 -225.595 ;
        RECT 222.875 -227.285 223.205 -226.955 ;
        RECT 222.875 -228.645 223.205 -228.315 ;
        RECT 222.875 -230.005 223.205 -229.675 ;
        RECT 222.875 -231.365 223.205 -231.035 ;
        RECT 222.875 -232.725 223.205 -232.395 ;
        RECT 222.875 -234.085 223.205 -233.755 ;
        RECT 222.875 -235.445 223.205 -235.115 ;
        RECT 222.875 -236.805 223.205 -236.475 ;
        RECT 222.875 -238.165 223.205 -237.835 ;
        RECT 222.875 -243.81 223.205 -242.68 ;
        RECT 222.88 -243.925 223.2 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 246.76 224.565 247.89 ;
        RECT 224.235 241.915 224.565 242.245 ;
        RECT 224.235 240.555 224.565 240.885 ;
        RECT 224.235 239.195 224.565 239.525 ;
        RECT 224.235 237.835 224.565 238.165 ;
        RECT 224.24 237.16 224.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 -1.525 224.565 -1.195 ;
        RECT 224.235 -2.885 224.565 -2.555 ;
        RECT 224.24 -3.56 224.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 246.76 225.925 247.89 ;
        RECT 225.595 241.915 225.925 242.245 ;
        RECT 225.595 240.555 225.925 240.885 ;
        RECT 225.595 239.195 225.925 239.525 ;
        RECT 225.595 237.835 225.925 238.165 ;
        RECT 225.6 237.16 225.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 -1.525 225.925 -1.195 ;
        RECT 225.595 -2.885 225.925 -2.555 ;
        RECT 225.6 -3.56 225.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 -160.645 225.925 -160.315 ;
        RECT 225.595 -162.005 225.925 -161.675 ;
        RECT 225.595 -163.365 225.925 -163.035 ;
        RECT 225.595 -164.725 225.925 -164.395 ;
        RECT 225.595 -166.085 225.925 -165.755 ;
        RECT 225.595 -167.445 225.925 -167.115 ;
        RECT 225.595 -168.805 225.925 -168.475 ;
        RECT 225.595 -170.165 225.925 -169.835 ;
        RECT 225.595 -171.525 225.925 -171.195 ;
        RECT 225.595 -172.885 225.925 -172.555 ;
        RECT 225.595 -174.245 225.925 -173.915 ;
        RECT 225.595 -175.605 225.925 -175.275 ;
        RECT 225.595 -176.965 225.925 -176.635 ;
        RECT 225.595 -178.325 225.925 -177.995 ;
        RECT 225.595 -179.685 225.925 -179.355 ;
        RECT 225.595 -181.045 225.925 -180.715 ;
        RECT 225.595 -182.405 225.925 -182.075 ;
        RECT 225.595 -183.765 225.925 -183.435 ;
        RECT 225.595 -185.125 225.925 -184.795 ;
        RECT 225.595 -186.485 225.925 -186.155 ;
        RECT 225.595 -187.845 225.925 -187.515 ;
        RECT 225.595 -189.205 225.925 -188.875 ;
        RECT 225.595 -190.565 225.925 -190.235 ;
        RECT 225.595 -191.925 225.925 -191.595 ;
        RECT 225.595 -193.285 225.925 -192.955 ;
        RECT 225.595 -194.645 225.925 -194.315 ;
        RECT 225.595 -196.005 225.925 -195.675 ;
        RECT 225.595 -197.365 225.925 -197.035 ;
        RECT 225.595 -198.725 225.925 -198.395 ;
        RECT 225.595 -200.085 225.925 -199.755 ;
        RECT 225.595 -201.445 225.925 -201.115 ;
        RECT 225.595 -202.805 225.925 -202.475 ;
        RECT 225.595 -204.165 225.925 -203.835 ;
        RECT 225.595 -205.525 225.925 -205.195 ;
        RECT 225.595 -206.885 225.925 -206.555 ;
        RECT 225.595 -208.245 225.925 -207.915 ;
        RECT 225.595 -209.605 225.925 -209.275 ;
        RECT 225.595 -210.965 225.925 -210.635 ;
        RECT 225.595 -212.325 225.925 -211.995 ;
        RECT 225.595 -213.685 225.925 -213.355 ;
        RECT 225.595 -215.045 225.925 -214.715 ;
        RECT 225.595 -216.405 225.925 -216.075 ;
        RECT 225.595 -217.765 225.925 -217.435 ;
        RECT 225.595 -219.125 225.925 -218.795 ;
        RECT 225.595 -220.485 225.925 -220.155 ;
        RECT 225.595 -221.845 225.925 -221.515 ;
        RECT 225.595 -223.205 225.925 -222.875 ;
        RECT 225.595 -224.565 225.925 -224.235 ;
        RECT 225.595 -225.925 225.925 -225.595 ;
        RECT 225.595 -227.285 225.925 -226.955 ;
        RECT 225.595 -228.645 225.925 -228.315 ;
        RECT 225.595 -230.005 225.925 -229.675 ;
        RECT 225.595 -231.365 225.925 -231.035 ;
        RECT 225.595 -232.725 225.925 -232.395 ;
        RECT 225.595 -234.085 225.925 -233.755 ;
        RECT 225.595 -235.445 225.925 -235.115 ;
        RECT 225.595 -236.805 225.925 -236.475 ;
        RECT 225.595 -238.165 225.925 -237.835 ;
        RECT 225.595 -243.81 225.925 -242.68 ;
        RECT 225.6 -243.925 225.92 -122.235 ;
        RECT 225.595 -122.565 225.925 -122.235 ;
        RECT 225.595 -123.925 225.925 -123.595 ;
        RECT 225.595 -125.285 225.925 -124.955 ;
        RECT 225.595 -126.645 225.925 -126.315 ;
        RECT 225.595 -128.005 225.925 -127.675 ;
        RECT 225.595 -129.365 225.925 -129.035 ;
        RECT 225.595 -130.725 225.925 -130.395 ;
        RECT 225.595 -132.085 225.925 -131.755 ;
        RECT 225.595 -133.445 225.925 -133.115 ;
        RECT 225.595 -134.805 225.925 -134.475 ;
        RECT 225.595 -136.165 225.925 -135.835 ;
        RECT 225.595 -137.525 225.925 -137.195 ;
        RECT 225.595 -138.885 225.925 -138.555 ;
        RECT 225.595 -140.245 225.925 -139.915 ;
        RECT 225.595 -141.605 225.925 -141.275 ;
        RECT 225.595 -142.965 225.925 -142.635 ;
        RECT 225.595 -144.325 225.925 -143.995 ;
        RECT 225.595 -145.685 225.925 -145.355 ;
        RECT 225.595 -147.045 225.925 -146.715 ;
        RECT 225.595 -148.405 225.925 -148.075 ;
        RECT 225.595 -149.765 225.925 -149.435 ;
        RECT 225.595 -151.125 225.925 -150.795 ;
        RECT 225.595 -152.485 225.925 -152.155 ;
        RECT 225.595 -153.845 225.925 -153.515 ;
        RECT 225.595 -155.205 225.925 -154.875 ;
        RECT 225.595 -156.565 225.925 -156.235 ;
        RECT 225.595 -157.925 225.925 -157.595 ;
        RECT 225.595 -159.285 225.925 -158.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 246.76 187.845 247.89 ;
        RECT 187.515 241.915 187.845 242.245 ;
        RECT 187.515 240.555 187.845 240.885 ;
        RECT 187.515 239.195 187.845 239.525 ;
        RECT 187.515 237.835 187.845 238.165 ;
        RECT 187.52 237.16 187.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 -126.645 187.845 -126.315 ;
        RECT 187.515 -128.005 187.845 -127.675 ;
        RECT 187.515 -129.365 187.845 -129.035 ;
        RECT 187.515 -130.725 187.845 -130.395 ;
        RECT 187.515 -132.085 187.845 -131.755 ;
        RECT 187.515 -133.445 187.845 -133.115 ;
        RECT 187.515 -134.805 187.845 -134.475 ;
        RECT 187.515 -136.165 187.845 -135.835 ;
        RECT 187.515 -137.525 187.845 -137.195 ;
        RECT 187.515 -138.885 187.845 -138.555 ;
        RECT 187.515 -140.245 187.845 -139.915 ;
        RECT 187.515 -141.605 187.845 -141.275 ;
        RECT 187.515 -142.965 187.845 -142.635 ;
        RECT 187.515 -144.325 187.845 -143.995 ;
        RECT 187.515 -145.685 187.845 -145.355 ;
        RECT 187.515 -147.045 187.845 -146.715 ;
        RECT 187.515 -148.405 187.845 -148.075 ;
        RECT 187.515 -149.765 187.845 -149.435 ;
        RECT 187.515 -151.125 187.845 -150.795 ;
        RECT 187.515 -152.485 187.845 -152.155 ;
        RECT 187.515 -153.845 187.845 -153.515 ;
        RECT 187.515 -155.205 187.845 -154.875 ;
        RECT 187.515 -156.565 187.845 -156.235 ;
        RECT 187.515 -157.925 187.845 -157.595 ;
        RECT 187.515 -159.285 187.845 -158.955 ;
        RECT 187.515 -160.645 187.845 -160.315 ;
        RECT 187.515 -162.005 187.845 -161.675 ;
        RECT 187.515 -163.365 187.845 -163.035 ;
        RECT 187.515 -164.725 187.845 -164.395 ;
        RECT 187.515 -166.085 187.845 -165.755 ;
        RECT 187.515 -167.445 187.845 -167.115 ;
        RECT 187.515 -168.805 187.845 -168.475 ;
        RECT 187.515 -170.165 187.845 -169.835 ;
        RECT 187.515 -171.525 187.845 -171.195 ;
        RECT 187.515 -172.885 187.845 -172.555 ;
        RECT 187.515 -174.245 187.845 -173.915 ;
        RECT 187.515 -175.605 187.845 -175.275 ;
        RECT 187.515 -176.965 187.845 -176.635 ;
        RECT 187.515 -178.325 187.845 -177.995 ;
        RECT 187.515 -179.685 187.845 -179.355 ;
        RECT 187.515 -181.045 187.845 -180.715 ;
        RECT 187.515 -182.405 187.845 -182.075 ;
        RECT 187.515 -183.765 187.845 -183.435 ;
        RECT 187.515 -185.125 187.845 -184.795 ;
        RECT 187.515 -186.485 187.845 -186.155 ;
        RECT 187.515 -187.845 187.845 -187.515 ;
        RECT 187.515 -189.205 187.845 -188.875 ;
        RECT 187.515 -190.565 187.845 -190.235 ;
        RECT 187.515 -191.925 187.845 -191.595 ;
        RECT 187.515 -193.285 187.845 -192.955 ;
        RECT 187.515 -194.645 187.845 -194.315 ;
        RECT 187.515 -196.005 187.845 -195.675 ;
        RECT 187.515 -197.365 187.845 -197.035 ;
        RECT 187.515 -198.725 187.845 -198.395 ;
        RECT 187.515 -200.085 187.845 -199.755 ;
        RECT 187.515 -201.445 187.845 -201.115 ;
        RECT 187.515 -202.805 187.845 -202.475 ;
        RECT 187.515 -204.165 187.845 -203.835 ;
        RECT 187.515 -205.525 187.845 -205.195 ;
        RECT 187.515 -206.885 187.845 -206.555 ;
        RECT 187.515 -208.245 187.845 -207.915 ;
        RECT 187.515 -209.605 187.845 -209.275 ;
        RECT 187.515 -210.965 187.845 -210.635 ;
        RECT 187.515 -212.325 187.845 -211.995 ;
        RECT 187.515 -213.685 187.845 -213.355 ;
        RECT 187.515 -215.045 187.845 -214.715 ;
        RECT 187.515 -216.405 187.845 -216.075 ;
        RECT 187.515 -217.765 187.845 -217.435 ;
        RECT 187.515 -219.125 187.845 -218.795 ;
        RECT 187.515 -220.485 187.845 -220.155 ;
        RECT 187.515 -221.845 187.845 -221.515 ;
        RECT 187.515 -223.205 187.845 -222.875 ;
        RECT 187.515 -224.565 187.845 -224.235 ;
        RECT 187.515 -225.925 187.845 -225.595 ;
        RECT 187.515 -227.285 187.845 -226.955 ;
        RECT 187.515 -228.645 187.845 -228.315 ;
        RECT 187.515 -230.005 187.845 -229.675 ;
        RECT 187.515 -231.365 187.845 -231.035 ;
        RECT 187.515 -232.725 187.845 -232.395 ;
        RECT 187.515 -234.085 187.845 -233.755 ;
        RECT 187.515 -235.445 187.845 -235.115 ;
        RECT 187.515 -236.805 187.845 -236.475 ;
        RECT 187.515 -238.165 187.845 -237.835 ;
        RECT 187.515 -243.81 187.845 -242.68 ;
        RECT 187.52 -243.925 187.84 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.96 -125.535 188.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 246.76 189.205 247.89 ;
        RECT 188.875 241.915 189.205 242.245 ;
        RECT 188.875 240.555 189.205 240.885 ;
        RECT 188.875 239.195 189.205 239.525 ;
        RECT 188.875 237.835 189.205 238.165 ;
        RECT 188.88 237.16 189.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 246.76 190.565 247.89 ;
        RECT 190.235 241.915 190.565 242.245 ;
        RECT 190.235 240.555 190.565 240.885 ;
        RECT 190.235 239.195 190.565 239.525 ;
        RECT 190.235 237.835 190.565 238.165 ;
        RECT 190.24 237.16 190.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 -1.525 190.565 -1.195 ;
        RECT 190.235 -2.885 190.565 -2.555 ;
        RECT 190.24 -3.56 190.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 246.76 191.925 247.89 ;
        RECT 191.595 241.915 191.925 242.245 ;
        RECT 191.595 240.555 191.925 240.885 ;
        RECT 191.595 239.195 191.925 239.525 ;
        RECT 191.595 237.835 191.925 238.165 ;
        RECT 191.6 237.16 191.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 -1.525 191.925 -1.195 ;
        RECT 191.595 -2.885 191.925 -2.555 ;
        RECT 191.6 -3.56 191.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 246.76 193.285 247.89 ;
        RECT 192.955 241.915 193.285 242.245 ;
        RECT 192.955 240.555 193.285 240.885 ;
        RECT 192.955 239.195 193.285 239.525 ;
        RECT 192.955 237.835 193.285 238.165 ;
        RECT 192.96 237.16 193.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 -1.525 193.285 -1.195 ;
        RECT 192.955 -2.885 193.285 -2.555 ;
        RECT 192.96 -3.56 193.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 -122.565 193.285 -122.235 ;
        RECT 192.955 -123.925 193.285 -123.595 ;
        RECT 192.955 -125.285 193.285 -124.955 ;
        RECT 192.955 -126.645 193.285 -126.315 ;
        RECT 192.955 -128.005 193.285 -127.675 ;
        RECT 192.955 -129.365 193.285 -129.035 ;
        RECT 192.955 -130.725 193.285 -130.395 ;
        RECT 192.955 -132.085 193.285 -131.755 ;
        RECT 192.955 -133.445 193.285 -133.115 ;
        RECT 192.955 -134.805 193.285 -134.475 ;
        RECT 192.955 -136.165 193.285 -135.835 ;
        RECT 192.955 -137.525 193.285 -137.195 ;
        RECT 192.955 -138.885 193.285 -138.555 ;
        RECT 192.955 -140.245 193.285 -139.915 ;
        RECT 192.955 -141.605 193.285 -141.275 ;
        RECT 192.955 -142.965 193.285 -142.635 ;
        RECT 192.955 -144.325 193.285 -143.995 ;
        RECT 192.955 -145.685 193.285 -145.355 ;
        RECT 192.955 -147.045 193.285 -146.715 ;
        RECT 192.955 -148.405 193.285 -148.075 ;
        RECT 192.955 -149.765 193.285 -149.435 ;
        RECT 192.955 -151.125 193.285 -150.795 ;
        RECT 192.955 -152.485 193.285 -152.155 ;
        RECT 192.955 -153.845 193.285 -153.515 ;
        RECT 192.955 -155.205 193.285 -154.875 ;
        RECT 192.955 -156.565 193.285 -156.235 ;
        RECT 192.955 -157.925 193.285 -157.595 ;
        RECT 192.955 -159.285 193.285 -158.955 ;
        RECT 192.955 -160.645 193.285 -160.315 ;
        RECT 192.955 -162.005 193.285 -161.675 ;
        RECT 192.955 -163.365 193.285 -163.035 ;
        RECT 192.955 -164.725 193.285 -164.395 ;
        RECT 192.955 -166.085 193.285 -165.755 ;
        RECT 192.955 -167.445 193.285 -167.115 ;
        RECT 192.955 -168.805 193.285 -168.475 ;
        RECT 192.955 -170.165 193.285 -169.835 ;
        RECT 192.955 -171.525 193.285 -171.195 ;
        RECT 192.955 -172.885 193.285 -172.555 ;
        RECT 192.955 -174.245 193.285 -173.915 ;
        RECT 192.955 -175.605 193.285 -175.275 ;
        RECT 192.955 -176.965 193.285 -176.635 ;
        RECT 192.955 -178.325 193.285 -177.995 ;
        RECT 192.955 -179.685 193.285 -179.355 ;
        RECT 192.955 -181.045 193.285 -180.715 ;
        RECT 192.955 -182.405 193.285 -182.075 ;
        RECT 192.955 -183.765 193.285 -183.435 ;
        RECT 192.955 -185.125 193.285 -184.795 ;
        RECT 192.955 -186.485 193.285 -186.155 ;
        RECT 192.955 -187.845 193.285 -187.515 ;
        RECT 192.955 -189.205 193.285 -188.875 ;
        RECT 192.955 -190.565 193.285 -190.235 ;
        RECT 192.955 -191.925 193.285 -191.595 ;
        RECT 192.955 -193.285 193.285 -192.955 ;
        RECT 192.955 -194.645 193.285 -194.315 ;
        RECT 192.955 -196.005 193.285 -195.675 ;
        RECT 192.955 -197.365 193.285 -197.035 ;
        RECT 192.955 -198.725 193.285 -198.395 ;
        RECT 192.955 -200.085 193.285 -199.755 ;
        RECT 192.955 -201.445 193.285 -201.115 ;
        RECT 192.955 -202.805 193.285 -202.475 ;
        RECT 192.955 -204.165 193.285 -203.835 ;
        RECT 192.955 -205.525 193.285 -205.195 ;
        RECT 192.955 -206.885 193.285 -206.555 ;
        RECT 192.955 -208.245 193.285 -207.915 ;
        RECT 192.955 -209.605 193.285 -209.275 ;
        RECT 192.955 -210.965 193.285 -210.635 ;
        RECT 192.955 -212.325 193.285 -211.995 ;
        RECT 192.955 -213.685 193.285 -213.355 ;
        RECT 192.955 -215.045 193.285 -214.715 ;
        RECT 192.955 -216.405 193.285 -216.075 ;
        RECT 192.955 -217.765 193.285 -217.435 ;
        RECT 192.955 -219.125 193.285 -218.795 ;
        RECT 192.955 -220.485 193.285 -220.155 ;
        RECT 192.955 -221.845 193.285 -221.515 ;
        RECT 192.955 -223.205 193.285 -222.875 ;
        RECT 192.955 -224.565 193.285 -224.235 ;
        RECT 192.955 -225.925 193.285 -225.595 ;
        RECT 192.955 -227.285 193.285 -226.955 ;
        RECT 192.955 -228.645 193.285 -228.315 ;
        RECT 192.955 -230.005 193.285 -229.675 ;
        RECT 192.955 -231.365 193.285 -231.035 ;
        RECT 192.955 -232.725 193.285 -232.395 ;
        RECT 192.955 -234.085 193.285 -233.755 ;
        RECT 192.955 -235.445 193.285 -235.115 ;
        RECT 192.955 -236.805 193.285 -236.475 ;
        RECT 192.955 -238.165 193.285 -237.835 ;
        RECT 192.955 -243.81 193.285 -242.68 ;
        RECT 192.96 -243.925 193.28 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 246.76 194.645 247.89 ;
        RECT 194.315 241.915 194.645 242.245 ;
        RECT 194.315 240.555 194.645 240.885 ;
        RECT 194.315 239.195 194.645 239.525 ;
        RECT 194.315 237.835 194.645 238.165 ;
        RECT 194.32 237.16 194.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 -1.525 194.645 -1.195 ;
        RECT 194.315 -2.885 194.645 -2.555 ;
        RECT 194.32 -3.56 194.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 -122.565 194.645 -122.235 ;
        RECT 194.315 -123.925 194.645 -123.595 ;
        RECT 194.315 -125.285 194.645 -124.955 ;
        RECT 194.315 -126.645 194.645 -126.315 ;
        RECT 194.315 -128.005 194.645 -127.675 ;
        RECT 194.315 -129.365 194.645 -129.035 ;
        RECT 194.315 -130.725 194.645 -130.395 ;
        RECT 194.315 -132.085 194.645 -131.755 ;
        RECT 194.315 -133.445 194.645 -133.115 ;
        RECT 194.315 -134.805 194.645 -134.475 ;
        RECT 194.315 -136.165 194.645 -135.835 ;
        RECT 194.315 -137.525 194.645 -137.195 ;
        RECT 194.315 -138.885 194.645 -138.555 ;
        RECT 194.315 -140.245 194.645 -139.915 ;
        RECT 194.315 -141.605 194.645 -141.275 ;
        RECT 194.315 -142.965 194.645 -142.635 ;
        RECT 194.315 -144.325 194.645 -143.995 ;
        RECT 194.315 -145.685 194.645 -145.355 ;
        RECT 194.315 -147.045 194.645 -146.715 ;
        RECT 194.315 -148.405 194.645 -148.075 ;
        RECT 194.315 -149.765 194.645 -149.435 ;
        RECT 194.315 -151.125 194.645 -150.795 ;
        RECT 194.315 -152.485 194.645 -152.155 ;
        RECT 194.315 -153.845 194.645 -153.515 ;
        RECT 194.315 -155.205 194.645 -154.875 ;
        RECT 194.315 -156.565 194.645 -156.235 ;
        RECT 194.315 -157.925 194.645 -157.595 ;
        RECT 194.315 -159.285 194.645 -158.955 ;
        RECT 194.315 -160.645 194.645 -160.315 ;
        RECT 194.315 -162.005 194.645 -161.675 ;
        RECT 194.315 -163.365 194.645 -163.035 ;
        RECT 194.315 -164.725 194.645 -164.395 ;
        RECT 194.315 -166.085 194.645 -165.755 ;
        RECT 194.315 -167.445 194.645 -167.115 ;
        RECT 194.315 -168.805 194.645 -168.475 ;
        RECT 194.315 -170.165 194.645 -169.835 ;
        RECT 194.315 -171.525 194.645 -171.195 ;
        RECT 194.315 -172.885 194.645 -172.555 ;
        RECT 194.315 -174.245 194.645 -173.915 ;
        RECT 194.315 -175.605 194.645 -175.275 ;
        RECT 194.315 -176.965 194.645 -176.635 ;
        RECT 194.315 -178.325 194.645 -177.995 ;
        RECT 194.315 -179.685 194.645 -179.355 ;
        RECT 194.315 -181.045 194.645 -180.715 ;
        RECT 194.315 -182.405 194.645 -182.075 ;
        RECT 194.315 -183.765 194.645 -183.435 ;
        RECT 194.315 -185.125 194.645 -184.795 ;
        RECT 194.315 -186.485 194.645 -186.155 ;
        RECT 194.315 -187.845 194.645 -187.515 ;
        RECT 194.315 -189.205 194.645 -188.875 ;
        RECT 194.315 -190.565 194.645 -190.235 ;
        RECT 194.315 -191.925 194.645 -191.595 ;
        RECT 194.315 -193.285 194.645 -192.955 ;
        RECT 194.315 -194.645 194.645 -194.315 ;
        RECT 194.315 -196.005 194.645 -195.675 ;
        RECT 194.315 -197.365 194.645 -197.035 ;
        RECT 194.315 -198.725 194.645 -198.395 ;
        RECT 194.315 -200.085 194.645 -199.755 ;
        RECT 194.315 -201.445 194.645 -201.115 ;
        RECT 194.315 -202.805 194.645 -202.475 ;
        RECT 194.315 -204.165 194.645 -203.835 ;
        RECT 194.315 -205.525 194.645 -205.195 ;
        RECT 194.315 -206.885 194.645 -206.555 ;
        RECT 194.315 -208.245 194.645 -207.915 ;
        RECT 194.315 -209.605 194.645 -209.275 ;
        RECT 194.315 -210.965 194.645 -210.635 ;
        RECT 194.315 -212.325 194.645 -211.995 ;
        RECT 194.315 -213.685 194.645 -213.355 ;
        RECT 194.315 -215.045 194.645 -214.715 ;
        RECT 194.315 -216.405 194.645 -216.075 ;
        RECT 194.315 -217.765 194.645 -217.435 ;
        RECT 194.315 -219.125 194.645 -218.795 ;
        RECT 194.315 -220.485 194.645 -220.155 ;
        RECT 194.315 -221.845 194.645 -221.515 ;
        RECT 194.315 -223.205 194.645 -222.875 ;
        RECT 194.315 -224.565 194.645 -224.235 ;
        RECT 194.315 -225.925 194.645 -225.595 ;
        RECT 194.315 -227.285 194.645 -226.955 ;
        RECT 194.315 -228.645 194.645 -228.315 ;
        RECT 194.315 -230.005 194.645 -229.675 ;
        RECT 194.315 -231.365 194.645 -231.035 ;
        RECT 194.315 -232.725 194.645 -232.395 ;
        RECT 194.315 -234.085 194.645 -233.755 ;
        RECT 194.315 -235.445 194.645 -235.115 ;
        RECT 194.315 -236.805 194.645 -236.475 ;
        RECT 194.315 -238.165 194.645 -237.835 ;
        RECT 194.315 -243.81 194.645 -242.68 ;
        RECT 194.32 -243.925 194.64 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 246.76 196.005 247.89 ;
        RECT 195.675 241.915 196.005 242.245 ;
        RECT 195.675 240.555 196.005 240.885 ;
        RECT 195.675 239.195 196.005 239.525 ;
        RECT 195.675 237.835 196.005 238.165 ;
        RECT 195.68 237.16 196 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -1.525 196.005 -1.195 ;
        RECT 195.675 -2.885 196.005 -2.555 ;
        RECT 195.68 -3.56 196 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -122.565 196.005 -122.235 ;
        RECT 195.675 -123.925 196.005 -123.595 ;
        RECT 195.675 -125.285 196.005 -124.955 ;
        RECT 195.675 -126.645 196.005 -126.315 ;
        RECT 195.675 -128.005 196.005 -127.675 ;
        RECT 195.675 -129.365 196.005 -129.035 ;
        RECT 195.675 -130.725 196.005 -130.395 ;
        RECT 195.675 -132.085 196.005 -131.755 ;
        RECT 195.675 -133.445 196.005 -133.115 ;
        RECT 195.675 -134.805 196.005 -134.475 ;
        RECT 195.675 -136.165 196.005 -135.835 ;
        RECT 195.675 -137.525 196.005 -137.195 ;
        RECT 195.675 -138.885 196.005 -138.555 ;
        RECT 195.675 -140.245 196.005 -139.915 ;
        RECT 195.675 -141.605 196.005 -141.275 ;
        RECT 195.675 -142.965 196.005 -142.635 ;
        RECT 195.675 -144.325 196.005 -143.995 ;
        RECT 195.675 -145.685 196.005 -145.355 ;
        RECT 195.675 -147.045 196.005 -146.715 ;
        RECT 195.675 -148.405 196.005 -148.075 ;
        RECT 195.675 -149.765 196.005 -149.435 ;
        RECT 195.675 -151.125 196.005 -150.795 ;
        RECT 195.675 -152.485 196.005 -152.155 ;
        RECT 195.675 -153.845 196.005 -153.515 ;
        RECT 195.675 -155.205 196.005 -154.875 ;
        RECT 195.675 -156.565 196.005 -156.235 ;
        RECT 195.675 -157.925 196.005 -157.595 ;
        RECT 195.675 -159.285 196.005 -158.955 ;
        RECT 195.675 -160.645 196.005 -160.315 ;
        RECT 195.675 -162.005 196.005 -161.675 ;
        RECT 195.675 -163.365 196.005 -163.035 ;
        RECT 195.675 -164.725 196.005 -164.395 ;
        RECT 195.675 -166.085 196.005 -165.755 ;
        RECT 195.675 -167.445 196.005 -167.115 ;
        RECT 195.675 -168.805 196.005 -168.475 ;
        RECT 195.675 -170.165 196.005 -169.835 ;
        RECT 195.675 -171.525 196.005 -171.195 ;
        RECT 195.675 -172.885 196.005 -172.555 ;
        RECT 195.675 -174.245 196.005 -173.915 ;
        RECT 195.675 -175.605 196.005 -175.275 ;
        RECT 195.675 -176.965 196.005 -176.635 ;
        RECT 195.675 -178.325 196.005 -177.995 ;
        RECT 195.675 -179.685 196.005 -179.355 ;
        RECT 195.675 -181.045 196.005 -180.715 ;
        RECT 195.675 -182.405 196.005 -182.075 ;
        RECT 195.675 -183.765 196.005 -183.435 ;
        RECT 195.675 -185.125 196.005 -184.795 ;
        RECT 195.675 -186.485 196.005 -186.155 ;
        RECT 195.675 -187.845 196.005 -187.515 ;
        RECT 195.675 -189.205 196.005 -188.875 ;
        RECT 195.675 -190.565 196.005 -190.235 ;
        RECT 195.675 -191.925 196.005 -191.595 ;
        RECT 195.675 -193.285 196.005 -192.955 ;
        RECT 195.675 -194.645 196.005 -194.315 ;
        RECT 195.675 -196.005 196.005 -195.675 ;
        RECT 195.675 -197.365 196.005 -197.035 ;
        RECT 195.675 -198.725 196.005 -198.395 ;
        RECT 195.675 -200.085 196.005 -199.755 ;
        RECT 195.675 -201.445 196.005 -201.115 ;
        RECT 195.675 -202.805 196.005 -202.475 ;
        RECT 195.675 -204.165 196.005 -203.835 ;
        RECT 195.675 -205.525 196.005 -205.195 ;
        RECT 195.675 -206.885 196.005 -206.555 ;
        RECT 195.675 -208.245 196.005 -207.915 ;
        RECT 195.675 -209.605 196.005 -209.275 ;
        RECT 195.675 -210.965 196.005 -210.635 ;
        RECT 195.675 -212.325 196.005 -211.995 ;
        RECT 195.675 -213.685 196.005 -213.355 ;
        RECT 195.675 -215.045 196.005 -214.715 ;
        RECT 195.675 -216.405 196.005 -216.075 ;
        RECT 195.675 -217.765 196.005 -217.435 ;
        RECT 195.675 -219.125 196.005 -218.795 ;
        RECT 195.675 -220.485 196.005 -220.155 ;
        RECT 195.675 -221.845 196.005 -221.515 ;
        RECT 195.675 -223.205 196.005 -222.875 ;
        RECT 195.675 -224.565 196.005 -224.235 ;
        RECT 195.675 -225.925 196.005 -225.595 ;
        RECT 195.675 -227.285 196.005 -226.955 ;
        RECT 195.675 -228.645 196.005 -228.315 ;
        RECT 195.675 -230.005 196.005 -229.675 ;
        RECT 195.675 -231.365 196.005 -231.035 ;
        RECT 195.675 -232.725 196.005 -232.395 ;
        RECT 195.675 -234.085 196.005 -233.755 ;
        RECT 195.675 -235.445 196.005 -235.115 ;
        RECT 195.675 -236.805 196.005 -236.475 ;
        RECT 195.675 -238.165 196.005 -237.835 ;
        RECT 195.675 -243.81 196.005 -242.68 ;
        RECT 195.68 -243.925 196 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 246.76 197.365 247.89 ;
        RECT 197.035 241.915 197.365 242.245 ;
        RECT 197.035 240.555 197.365 240.885 ;
        RECT 197.035 239.195 197.365 239.525 ;
        RECT 197.035 237.835 197.365 238.165 ;
        RECT 197.04 237.16 197.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -1.525 197.365 -1.195 ;
        RECT 197.035 -2.885 197.365 -2.555 ;
        RECT 197.04 -3.56 197.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -122.565 197.365 -122.235 ;
        RECT 197.035 -123.925 197.365 -123.595 ;
        RECT 197.035 -125.285 197.365 -124.955 ;
        RECT 197.035 -126.645 197.365 -126.315 ;
        RECT 197.035 -128.005 197.365 -127.675 ;
        RECT 197.035 -129.365 197.365 -129.035 ;
        RECT 197.035 -130.725 197.365 -130.395 ;
        RECT 197.035 -132.085 197.365 -131.755 ;
        RECT 197.035 -133.445 197.365 -133.115 ;
        RECT 197.035 -134.805 197.365 -134.475 ;
        RECT 197.035 -136.165 197.365 -135.835 ;
        RECT 197.035 -137.525 197.365 -137.195 ;
        RECT 197.035 -138.885 197.365 -138.555 ;
        RECT 197.035 -140.245 197.365 -139.915 ;
        RECT 197.035 -141.605 197.365 -141.275 ;
        RECT 197.035 -142.965 197.365 -142.635 ;
        RECT 197.035 -144.325 197.365 -143.995 ;
        RECT 197.035 -145.685 197.365 -145.355 ;
        RECT 197.035 -147.045 197.365 -146.715 ;
        RECT 197.035 -148.405 197.365 -148.075 ;
        RECT 197.035 -149.765 197.365 -149.435 ;
        RECT 197.035 -151.125 197.365 -150.795 ;
        RECT 197.035 -152.485 197.365 -152.155 ;
        RECT 197.035 -153.845 197.365 -153.515 ;
        RECT 197.035 -155.205 197.365 -154.875 ;
        RECT 197.035 -156.565 197.365 -156.235 ;
        RECT 197.035 -157.925 197.365 -157.595 ;
        RECT 197.035 -159.285 197.365 -158.955 ;
        RECT 197.035 -160.645 197.365 -160.315 ;
        RECT 197.035 -162.005 197.365 -161.675 ;
        RECT 197.035 -163.365 197.365 -163.035 ;
        RECT 197.035 -164.725 197.365 -164.395 ;
        RECT 197.035 -166.085 197.365 -165.755 ;
        RECT 197.035 -167.445 197.365 -167.115 ;
        RECT 197.035 -168.805 197.365 -168.475 ;
        RECT 197.035 -170.165 197.365 -169.835 ;
        RECT 197.035 -171.525 197.365 -171.195 ;
        RECT 197.035 -172.885 197.365 -172.555 ;
        RECT 197.035 -174.245 197.365 -173.915 ;
        RECT 197.035 -175.605 197.365 -175.275 ;
        RECT 197.035 -176.965 197.365 -176.635 ;
        RECT 197.035 -178.325 197.365 -177.995 ;
        RECT 197.035 -179.685 197.365 -179.355 ;
        RECT 197.035 -181.045 197.365 -180.715 ;
        RECT 197.035 -182.405 197.365 -182.075 ;
        RECT 197.035 -183.765 197.365 -183.435 ;
        RECT 197.035 -185.125 197.365 -184.795 ;
        RECT 197.035 -186.485 197.365 -186.155 ;
        RECT 197.035 -187.845 197.365 -187.515 ;
        RECT 197.035 -189.205 197.365 -188.875 ;
        RECT 197.035 -190.565 197.365 -190.235 ;
        RECT 197.035 -191.925 197.365 -191.595 ;
        RECT 197.035 -193.285 197.365 -192.955 ;
        RECT 197.035 -194.645 197.365 -194.315 ;
        RECT 197.035 -196.005 197.365 -195.675 ;
        RECT 197.035 -197.365 197.365 -197.035 ;
        RECT 197.035 -198.725 197.365 -198.395 ;
        RECT 197.035 -200.085 197.365 -199.755 ;
        RECT 197.035 -201.445 197.365 -201.115 ;
        RECT 197.035 -202.805 197.365 -202.475 ;
        RECT 197.035 -204.165 197.365 -203.835 ;
        RECT 197.035 -205.525 197.365 -205.195 ;
        RECT 197.035 -206.885 197.365 -206.555 ;
        RECT 197.035 -208.245 197.365 -207.915 ;
        RECT 197.035 -209.605 197.365 -209.275 ;
        RECT 197.035 -210.965 197.365 -210.635 ;
        RECT 197.035 -212.325 197.365 -211.995 ;
        RECT 197.035 -213.685 197.365 -213.355 ;
        RECT 197.035 -215.045 197.365 -214.715 ;
        RECT 197.035 -216.405 197.365 -216.075 ;
        RECT 197.035 -217.765 197.365 -217.435 ;
        RECT 197.035 -219.125 197.365 -218.795 ;
        RECT 197.035 -220.485 197.365 -220.155 ;
        RECT 197.035 -221.845 197.365 -221.515 ;
        RECT 197.035 -223.205 197.365 -222.875 ;
        RECT 197.035 -224.565 197.365 -224.235 ;
        RECT 197.035 -225.925 197.365 -225.595 ;
        RECT 197.035 -227.285 197.365 -226.955 ;
        RECT 197.035 -228.645 197.365 -228.315 ;
        RECT 197.035 -230.005 197.365 -229.675 ;
        RECT 197.035 -231.365 197.365 -231.035 ;
        RECT 197.035 -232.725 197.365 -232.395 ;
        RECT 197.035 -234.085 197.365 -233.755 ;
        RECT 197.035 -235.445 197.365 -235.115 ;
        RECT 197.035 -236.805 197.365 -236.475 ;
        RECT 197.035 -238.165 197.365 -237.835 ;
        RECT 197.035 -243.81 197.365 -242.68 ;
        RECT 197.04 -243.925 197.36 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 246.76 198.725 247.89 ;
        RECT 198.395 241.915 198.725 242.245 ;
        RECT 198.395 240.555 198.725 240.885 ;
        RECT 198.395 239.195 198.725 239.525 ;
        RECT 198.395 237.835 198.725 238.165 ;
        RECT 198.4 237.16 198.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 -126.645 198.725 -126.315 ;
        RECT 198.395 -128.005 198.725 -127.675 ;
        RECT 198.395 -129.365 198.725 -129.035 ;
        RECT 198.395 -130.725 198.725 -130.395 ;
        RECT 198.395 -132.085 198.725 -131.755 ;
        RECT 198.395 -133.445 198.725 -133.115 ;
        RECT 198.395 -134.805 198.725 -134.475 ;
        RECT 198.395 -136.165 198.725 -135.835 ;
        RECT 198.395 -137.525 198.725 -137.195 ;
        RECT 198.395 -138.885 198.725 -138.555 ;
        RECT 198.395 -140.245 198.725 -139.915 ;
        RECT 198.395 -141.605 198.725 -141.275 ;
        RECT 198.395 -142.965 198.725 -142.635 ;
        RECT 198.395 -144.325 198.725 -143.995 ;
        RECT 198.395 -145.685 198.725 -145.355 ;
        RECT 198.395 -147.045 198.725 -146.715 ;
        RECT 198.395 -148.405 198.725 -148.075 ;
        RECT 198.395 -149.765 198.725 -149.435 ;
        RECT 198.395 -151.125 198.725 -150.795 ;
        RECT 198.395 -152.485 198.725 -152.155 ;
        RECT 198.395 -153.845 198.725 -153.515 ;
        RECT 198.395 -155.205 198.725 -154.875 ;
        RECT 198.395 -156.565 198.725 -156.235 ;
        RECT 198.395 -157.925 198.725 -157.595 ;
        RECT 198.395 -159.285 198.725 -158.955 ;
        RECT 198.395 -160.645 198.725 -160.315 ;
        RECT 198.395 -162.005 198.725 -161.675 ;
        RECT 198.395 -163.365 198.725 -163.035 ;
        RECT 198.395 -164.725 198.725 -164.395 ;
        RECT 198.395 -166.085 198.725 -165.755 ;
        RECT 198.395 -167.445 198.725 -167.115 ;
        RECT 198.395 -168.805 198.725 -168.475 ;
        RECT 198.395 -170.165 198.725 -169.835 ;
        RECT 198.395 -171.525 198.725 -171.195 ;
        RECT 198.395 -172.885 198.725 -172.555 ;
        RECT 198.395 -174.245 198.725 -173.915 ;
        RECT 198.395 -175.605 198.725 -175.275 ;
        RECT 198.395 -176.965 198.725 -176.635 ;
        RECT 198.395 -178.325 198.725 -177.995 ;
        RECT 198.395 -179.685 198.725 -179.355 ;
        RECT 198.395 -181.045 198.725 -180.715 ;
        RECT 198.395 -182.405 198.725 -182.075 ;
        RECT 198.395 -183.765 198.725 -183.435 ;
        RECT 198.395 -185.125 198.725 -184.795 ;
        RECT 198.395 -186.485 198.725 -186.155 ;
        RECT 198.395 -187.845 198.725 -187.515 ;
        RECT 198.395 -189.205 198.725 -188.875 ;
        RECT 198.395 -190.565 198.725 -190.235 ;
        RECT 198.395 -191.925 198.725 -191.595 ;
        RECT 198.395 -193.285 198.725 -192.955 ;
        RECT 198.395 -194.645 198.725 -194.315 ;
        RECT 198.395 -196.005 198.725 -195.675 ;
        RECT 198.395 -197.365 198.725 -197.035 ;
        RECT 198.395 -198.725 198.725 -198.395 ;
        RECT 198.395 -200.085 198.725 -199.755 ;
        RECT 198.395 -201.445 198.725 -201.115 ;
        RECT 198.395 -202.805 198.725 -202.475 ;
        RECT 198.395 -204.165 198.725 -203.835 ;
        RECT 198.395 -205.525 198.725 -205.195 ;
        RECT 198.395 -206.885 198.725 -206.555 ;
        RECT 198.395 -208.245 198.725 -207.915 ;
        RECT 198.395 -209.605 198.725 -209.275 ;
        RECT 198.395 -210.965 198.725 -210.635 ;
        RECT 198.395 -212.325 198.725 -211.995 ;
        RECT 198.395 -213.685 198.725 -213.355 ;
        RECT 198.395 -215.045 198.725 -214.715 ;
        RECT 198.395 -216.405 198.725 -216.075 ;
        RECT 198.395 -217.765 198.725 -217.435 ;
        RECT 198.395 -219.125 198.725 -218.795 ;
        RECT 198.395 -220.485 198.725 -220.155 ;
        RECT 198.395 -221.845 198.725 -221.515 ;
        RECT 198.395 -223.205 198.725 -222.875 ;
        RECT 198.395 -224.565 198.725 -224.235 ;
        RECT 198.395 -225.925 198.725 -225.595 ;
        RECT 198.395 -227.285 198.725 -226.955 ;
        RECT 198.395 -228.645 198.725 -228.315 ;
        RECT 198.395 -230.005 198.725 -229.675 ;
        RECT 198.395 -231.365 198.725 -231.035 ;
        RECT 198.395 -232.725 198.725 -232.395 ;
        RECT 198.395 -234.085 198.725 -233.755 ;
        RECT 198.395 -235.445 198.725 -235.115 ;
        RECT 198.395 -236.805 198.725 -236.475 ;
        RECT 198.395 -238.165 198.725 -237.835 ;
        RECT 198.395 -243.81 198.725 -242.68 ;
        RECT 198.4 -243.925 198.72 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.86 -125.535 199.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 246.76 200.085 247.89 ;
        RECT 199.755 241.915 200.085 242.245 ;
        RECT 199.755 240.555 200.085 240.885 ;
        RECT 199.755 239.195 200.085 239.525 ;
        RECT 199.755 237.835 200.085 238.165 ;
        RECT 199.76 237.16 200.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 246.76 201.445 247.89 ;
        RECT 201.115 241.915 201.445 242.245 ;
        RECT 201.115 240.555 201.445 240.885 ;
        RECT 201.115 239.195 201.445 239.525 ;
        RECT 201.115 237.835 201.445 238.165 ;
        RECT 201.12 237.16 201.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -1.525 201.445 -1.195 ;
        RECT 201.115 -2.885 201.445 -2.555 ;
        RECT 201.12 -3.56 201.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -122.565 201.445 -122.235 ;
        RECT 201.115 -123.925 201.445 -123.595 ;
        RECT 201.115 -125.285 201.445 -124.955 ;
        RECT 201.115 -126.645 201.445 -126.315 ;
        RECT 201.115 -128.005 201.445 -127.675 ;
        RECT 201.115 -129.365 201.445 -129.035 ;
        RECT 201.115 -130.725 201.445 -130.395 ;
        RECT 201.115 -132.085 201.445 -131.755 ;
        RECT 201.115 -133.445 201.445 -133.115 ;
        RECT 201.115 -134.805 201.445 -134.475 ;
        RECT 201.115 -136.165 201.445 -135.835 ;
        RECT 201.115 -137.525 201.445 -137.195 ;
        RECT 201.115 -138.885 201.445 -138.555 ;
        RECT 201.115 -140.245 201.445 -139.915 ;
        RECT 201.115 -141.605 201.445 -141.275 ;
        RECT 201.115 -142.965 201.445 -142.635 ;
        RECT 201.115 -144.325 201.445 -143.995 ;
        RECT 201.115 -145.685 201.445 -145.355 ;
        RECT 201.115 -147.045 201.445 -146.715 ;
        RECT 201.115 -148.405 201.445 -148.075 ;
        RECT 201.115 -149.765 201.445 -149.435 ;
        RECT 201.115 -151.125 201.445 -150.795 ;
        RECT 201.115 -152.485 201.445 -152.155 ;
        RECT 201.115 -153.845 201.445 -153.515 ;
        RECT 201.115 -155.205 201.445 -154.875 ;
        RECT 201.115 -156.565 201.445 -156.235 ;
        RECT 201.115 -157.925 201.445 -157.595 ;
        RECT 201.115 -159.285 201.445 -158.955 ;
        RECT 201.115 -160.645 201.445 -160.315 ;
        RECT 201.115 -162.005 201.445 -161.675 ;
        RECT 201.115 -163.365 201.445 -163.035 ;
        RECT 201.115 -164.725 201.445 -164.395 ;
        RECT 201.115 -166.085 201.445 -165.755 ;
        RECT 201.115 -167.445 201.445 -167.115 ;
        RECT 201.115 -168.805 201.445 -168.475 ;
        RECT 201.115 -170.165 201.445 -169.835 ;
        RECT 201.115 -171.525 201.445 -171.195 ;
        RECT 201.115 -172.885 201.445 -172.555 ;
        RECT 201.115 -174.245 201.445 -173.915 ;
        RECT 201.115 -175.605 201.445 -175.275 ;
        RECT 201.115 -176.965 201.445 -176.635 ;
        RECT 201.115 -178.325 201.445 -177.995 ;
        RECT 201.115 -179.685 201.445 -179.355 ;
        RECT 201.115 -181.045 201.445 -180.715 ;
        RECT 201.115 -182.405 201.445 -182.075 ;
        RECT 201.115 -183.765 201.445 -183.435 ;
        RECT 201.115 -185.125 201.445 -184.795 ;
        RECT 201.115 -186.485 201.445 -186.155 ;
        RECT 201.115 -187.845 201.445 -187.515 ;
        RECT 201.115 -189.205 201.445 -188.875 ;
        RECT 201.115 -190.565 201.445 -190.235 ;
        RECT 201.115 -191.925 201.445 -191.595 ;
        RECT 201.115 -193.285 201.445 -192.955 ;
        RECT 201.115 -194.645 201.445 -194.315 ;
        RECT 201.115 -196.005 201.445 -195.675 ;
        RECT 201.115 -197.365 201.445 -197.035 ;
        RECT 201.115 -198.725 201.445 -198.395 ;
        RECT 201.115 -200.085 201.445 -199.755 ;
        RECT 201.115 -201.445 201.445 -201.115 ;
        RECT 201.115 -202.805 201.445 -202.475 ;
        RECT 201.115 -204.165 201.445 -203.835 ;
        RECT 201.115 -205.525 201.445 -205.195 ;
        RECT 201.115 -206.885 201.445 -206.555 ;
        RECT 201.115 -208.245 201.445 -207.915 ;
        RECT 201.115 -209.605 201.445 -209.275 ;
        RECT 201.115 -210.965 201.445 -210.635 ;
        RECT 201.115 -212.325 201.445 -211.995 ;
        RECT 201.115 -213.685 201.445 -213.355 ;
        RECT 201.115 -215.045 201.445 -214.715 ;
        RECT 201.115 -216.405 201.445 -216.075 ;
        RECT 201.115 -217.765 201.445 -217.435 ;
        RECT 201.115 -219.125 201.445 -218.795 ;
        RECT 201.115 -220.485 201.445 -220.155 ;
        RECT 201.115 -221.845 201.445 -221.515 ;
        RECT 201.115 -223.205 201.445 -222.875 ;
        RECT 201.115 -224.565 201.445 -224.235 ;
        RECT 201.115 -225.925 201.445 -225.595 ;
        RECT 201.115 -227.285 201.445 -226.955 ;
        RECT 201.115 -228.645 201.445 -228.315 ;
        RECT 201.115 -230.005 201.445 -229.675 ;
        RECT 201.115 -231.365 201.445 -231.035 ;
        RECT 201.115 -232.725 201.445 -232.395 ;
        RECT 201.115 -234.085 201.445 -233.755 ;
        RECT 201.115 -235.445 201.445 -235.115 ;
        RECT 201.115 -236.805 201.445 -236.475 ;
        RECT 201.115 -238.165 201.445 -237.835 ;
        RECT 201.115 -243.81 201.445 -242.68 ;
        RECT 201.12 -243.925 201.44 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 246.76 202.805 247.89 ;
        RECT 202.475 241.915 202.805 242.245 ;
        RECT 202.475 240.555 202.805 240.885 ;
        RECT 202.475 239.195 202.805 239.525 ;
        RECT 202.475 237.835 202.805 238.165 ;
        RECT 202.48 237.16 202.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 -1.525 202.805 -1.195 ;
        RECT 202.475 -2.885 202.805 -2.555 ;
        RECT 202.48 -3.56 202.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 246.76 204.165 247.89 ;
        RECT 203.835 241.915 204.165 242.245 ;
        RECT 203.835 240.555 204.165 240.885 ;
        RECT 203.835 239.195 204.165 239.525 ;
        RECT 203.835 237.835 204.165 238.165 ;
        RECT 203.84 237.16 204.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 -1.525 204.165 -1.195 ;
        RECT 203.835 -2.885 204.165 -2.555 ;
        RECT 203.84 -3.56 204.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 -122.565 204.165 -122.235 ;
        RECT 203.835 -123.925 204.165 -123.595 ;
        RECT 203.835 -125.285 204.165 -124.955 ;
        RECT 203.835 -126.645 204.165 -126.315 ;
        RECT 203.835 -128.005 204.165 -127.675 ;
        RECT 203.835 -129.365 204.165 -129.035 ;
        RECT 203.835 -130.725 204.165 -130.395 ;
        RECT 203.835 -132.085 204.165 -131.755 ;
        RECT 203.835 -133.445 204.165 -133.115 ;
        RECT 203.835 -134.805 204.165 -134.475 ;
        RECT 203.835 -136.165 204.165 -135.835 ;
        RECT 203.835 -137.525 204.165 -137.195 ;
        RECT 203.835 -138.885 204.165 -138.555 ;
        RECT 203.835 -140.245 204.165 -139.915 ;
        RECT 203.835 -141.605 204.165 -141.275 ;
        RECT 203.835 -142.965 204.165 -142.635 ;
        RECT 203.835 -144.325 204.165 -143.995 ;
        RECT 203.835 -145.685 204.165 -145.355 ;
        RECT 203.835 -147.045 204.165 -146.715 ;
        RECT 203.835 -148.405 204.165 -148.075 ;
        RECT 203.835 -149.765 204.165 -149.435 ;
        RECT 203.835 -151.125 204.165 -150.795 ;
        RECT 203.835 -152.485 204.165 -152.155 ;
        RECT 203.835 -153.845 204.165 -153.515 ;
        RECT 203.835 -155.205 204.165 -154.875 ;
        RECT 203.835 -156.565 204.165 -156.235 ;
        RECT 203.835 -157.925 204.165 -157.595 ;
        RECT 203.835 -159.285 204.165 -158.955 ;
        RECT 203.835 -160.645 204.165 -160.315 ;
        RECT 203.835 -162.005 204.165 -161.675 ;
        RECT 203.835 -163.365 204.165 -163.035 ;
        RECT 203.835 -164.725 204.165 -164.395 ;
        RECT 203.835 -166.085 204.165 -165.755 ;
        RECT 203.835 -167.445 204.165 -167.115 ;
        RECT 203.835 -168.805 204.165 -168.475 ;
        RECT 203.835 -170.165 204.165 -169.835 ;
        RECT 203.835 -171.525 204.165 -171.195 ;
        RECT 203.835 -172.885 204.165 -172.555 ;
        RECT 203.835 -174.245 204.165 -173.915 ;
        RECT 203.835 -175.605 204.165 -175.275 ;
        RECT 203.835 -176.965 204.165 -176.635 ;
        RECT 203.835 -178.325 204.165 -177.995 ;
        RECT 203.835 -179.685 204.165 -179.355 ;
        RECT 203.835 -181.045 204.165 -180.715 ;
        RECT 203.835 -182.405 204.165 -182.075 ;
        RECT 203.835 -183.765 204.165 -183.435 ;
        RECT 203.835 -185.125 204.165 -184.795 ;
        RECT 203.835 -186.485 204.165 -186.155 ;
        RECT 203.835 -187.845 204.165 -187.515 ;
        RECT 203.835 -189.205 204.165 -188.875 ;
        RECT 203.835 -190.565 204.165 -190.235 ;
        RECT 203.835 -191.925 204.165 -191.595 ;
        RECT 203.835 -193.285 204.165 -192.955 ;
        RECT 203.835 -194.645 204.165 -194.315 ;
        RECT 203.835 -196.005 204.165 -195.675 ;
        RECT 203.835 -197.365 204.165 -197.035 ;
        RECT 203.835 -198.725 204.165 -198.395 ;
        RECT 203.835 -200.085 204.165 -199.755 ;
        RECT 203.835 -201.445 204.165 -201.115 ;
        RECT 203.835 -202.805 204.165 -202.475 ;
        RECT 203.835 -204.165 204.165 -203.835 ;
        RECT 203.835 -205.525 204.165 -205.195 ;
        RECT 203.835 -206.885 204.165 -206.555 ;
        RECT 203.835 -208.245 204.165 -207.915 ;
        RECT 203.835 -209.605 204.165 -209.275 ;
        RECT 203.835 -210.965 204.165 -210.635 ;
        RECT 203.835 -212.325 204.165 -211.995 ;
        RECT 203.835 -213.685 204.165 -213.355 ;
        RECT 203.835 -215.045 204.165 -214.715 ;
        RECT 203.835 -216.405 204.165 -216.075 ;
        RECT 203.835 -217.765 204.165 -217.435 ;
        RECT 203.835 -219.125 204.165 -218.795 ;
        RECT 203.835 -220.485 204.165 -220.155 ;
        RECT 203.835 -221.845 204.165 -221.515 ;
        RECT 203.835 -223.205 204.165 -222.875 ;
        RECT 203.835 -224.565 204.165 -224.235 ;
        RECT 203.835 -225.925 204.165 -225.595 ;
        RECT 203.835 -227.285 204.165 -226.955 ;
        RECT 203.835 -228.645 204.165 -228.315 ;
        RECT 203.835 -230.005 204.165 -229.675 ;
        RECT 203.835 -231.365 204.165 -231.035 ;
        RECT 203.835 -232.725 204.165 -232.395 ;
        RECT 203.835 -234.085 204.165 -233.755 ;
        RECT 203.835 -235.445 204.165 -235.115 ;
        RECT 203.835 -236.805 204.165 -236.475 ;
        RECT 203.835 -238.165 204.165 -237.835 ;
        RECT 203.835 -243.81 204.165 -242.68 ;
        RECT 203.84 -243.925 204.16 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 246.76 205.525 247.89 ;
        RECT 205.195 241.915 205.525 242.245 ;
        RECT 205.195 240.555 205.525 240.885 ;
        RECT 205.195 239.195 205.525 239.525 ;
        RECT 205.195 237.835 205.525 238.165 ;
        RECT 205.2 237.16 205.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 -1.525 205.525 -1.195 ;
        RECT 205.195 -2.885 205.525 -2.555 ;
        RECT 205.2 -3.56 205.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 -122.565 205.525 -122.235 ;
        RECT 205.195 -123.925 205.525 -123.595 ;
        RECT 205.195 -125.285 205.525 -124.955 ;
        RECT 205.195 -126.645 205.525 -126.315 ;
        RECT 205.195 -128.005 205.525 -127.675 ;
        RECT 205.195 -129.365 205.525 -129.035 ;
        RECT 205.195 -130.725 205.525 -130.395 ;
        RECT 205.195 -132.085 205.525 -131.755 ;
        RECT 205.195 -133.445 205.525 -133.115 ;
        RECT 205.195 -134.805 205.525 -134.475 ;
        RECT 205.195 -136.165 205.525 -135.835 ;
        RECT 205.195 -137.525 205.525 -137.195 ;
        RECT 205.195 -138.885 205.525 -138.555 ;
        RECT 205.195 -140.245 205.525 -139.915 ;
        RECT 205.195 -141.605 205.525 -141.275 ;
        RECT 205.195 -142.965 205.525 -142.635 ;
        RECT 205.195 -144.325 205.525 -143.995 ;
        RECT 205.195 -145.685 205.525 -145.355 ;
        RECT 205.195 -147.045 205.525 -146.715 ;
        RECT 205.195 -148.405 205.525 -148.075 ;
        RECT 205.195 -149.765 205.525 -149.435 ;
        RECT 205.195 -151.125 205.525 -150.795 ;
        RECT 205.195 -152.485 205.525 -152.155 ;
        RECT 205.195 -153.845 205.525 -153.515 ;
        RECT 205.195 -155.205 205.525 -154.875 ;
        RECT 205.195 -156.565 205.525 -156.235 ;
        RECT 205.195 -157.925 205.525 -157.595 ;
        RECT 205.195 -159.285 205.525 -158.955 ;
        RECT 205.195 -160.645 205.525 -160.315 ;
        RECT 205.195 -162.005 205.525 -161.675 ;
        RECT 205.195 -163.365 205.525 -163.035 ;
        RECT 205.195 -164.725 205.525 -164.395 ;
        RECT 205.195 -166.085 205.525 -165.755 ;
        RECT 205.195 -167.445 205.525 -167.115 ;
        RECT 205.195 -168.805 205.525 -168.475 ;
        RECT 205.195 -170.165 205.525 -169.835 ;
        RECT 205.195 -171.525 205.525 -171.195 ;
        RECT 205.195 -172.885 205.525 -172.555 ;
        RECT 205.195 -174.245 205.525 -173.915 ;
        RECT 205.195 -175.605 205.525 -175.275 ;
        RECT 205.195 -176.965 205.525 -176.635 ;
        RECT 205.195 -178.325 205.525 -177.995 ;
        RECT 205.195 -179.685 205.525 -179.355 ;
        RECT 205.195 -181.045 205.525 -180.715 ;
        RECT 205.195 -182.405 205.525 -182.075 ;
        RECT 205.195 -183.765 205.525 -183.435 ;
        RECT 205.195 -185.125 205.525 -184.795 ;
        RECT 205.195 -186.485 205.525 -186.155 ;
        RECT 205.195 -187.845 205.525 -187.515 ;
        RECT 205.195 -189.205 205.525 -188.875 ;
        RECT 205.195 -190.565 205.525 -190.235 ;
        RECT 205.195 -191.925 205.525 -191.595 ;
        RECT 205.195 -193.285 205.525 -192.955 ;
        RECT 205.195 -194.645 205.525 -194.315 ;
        RECT 205.195 -196.005 205.525 -195.675 ;
        RECT 205.195 -197.365 205.525 -197.035 ;
        RECT 205.195 -198.725 205.525 -198.395 ;
        RECT 205.195 -200.085 205.525 -199.755 ;
        RECT 205.195 -201.445 205.525 -201.115 ;
        RECT 205.195 -202.805 205.525 -202.475 ;
        RECT 205.195 -204.165 205.525 -203.835 ;
        RECT 205.195 -205.525 205.525 -205.195 ;
        RECT 205.195 -206.885 205.525 -206.555 ;
        RECT 205.195 -208.245 205.525 -207.915 ;
        RECT 205.195 -209.605 205.525 -209.275 ;
        RECT 205.195 -210.965 205.525 -210.635 ;
        RECT 205.195 -212.325 205.525 -211.995 ;
        RECT 205.195 -213.685 205.525 -213.355 ;
        RECT 205.195 -215.045 205.525 -214.715 ;
        RECT 205.195 -216.405 205.525 -216.075 ;
        RECT 205.195 -217.765 205.525 -217.435 ;
        RECT 205.195 -219.125 205.525 -218.795 ;
        RECT 205.195 -220.485 205.525 -220.155 ;
        RECT 205.195 -221.845 205.525 -221.515 ;
        RECT 205.195 -223.205 205.525 -222.875 ;
        RECT 205.195 -224.565 205.525 -224.235 ;
        RECT 205.195 -225.925 205.525 -225.595 ;
        RECT 205.195 -227.285 205.525 -226.955 ;
        RECT 205.195 -228.645 205.525 -228.315 ;
        RECT 205.195 -230.005 205.525 -229.675 ;
        RECT 205.195 -231.365 205.525 -231.035 ;
        RECT 205.195 -232.725 205.525 -232.395 ;
        RECT 205.195 -234.085 205.525 -233.755 ;
        RECT 205.195 -235.445 205.525 -235.115 ;
        RECT 205.195 -236.805 205.525 -236.475 ;
        RECT 205.195 -238.165 205.525 -237.835 ;
        RECT 205.195 -243.81 205.525 -242.68 ;
        RECT 205.2 -243.925 205.52 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 246.76 206.885 247.89 ;
        RECT 206.555 241.915 206.885 242.245 ;
        RECT 206.555 240.555 206.885 240.885 ;
        RECT 206.555 239.195 206.885 239.525 ;
        RECT 206.555 237.835 206.885 238.165 ;
        RECT 206.56 237.16 206.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 -1.525 206.885 -1.195 ;
        RECT 206.555 -2.885 206.885 -2.555 ;
        RECT 206.56 -3.56 206.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 -174.245 206.885 -173.915 ;
        RECT 206.555 -175.605 206.885 -175.275 ;
        RECT 206.555 -176.965 206.885 -176.635 ;
        RECT 206.555 -178.325 206.885 -177.995 ;
        RECT 206.555 -179.685 206.885 -179.355 ;
        RECT 206.555 -181.045 206.885 -180.715 ;
        RECT 206.555 -182.405 206.885 -182.075 ;
        RECT 206.555 -183.765 206.885 -183.435 ;
        RECT 206.555 -185.125 206.885 -184.795 ;
        RECT 206.555 -186.485 206.885 -186.155 ;
        RECT 206.555 -187.845 206.885 -187.515 ;
        RECT 206.555 -189.205 206.885 -188.875 ;
        RECT 206.555 -190.565 206.885 -190.235 ;
        RECT 206.555 -191.925 206.885 -191.595 ;
        RECT 206.555 -193.285 206.885 -192.955 ;
        RECT 206.555 -194.645 206.885 -194.315 ;
        RECT 206.555 -196.005 206.885 -195.675 ;
        RECT 206.555 -197.365 206.885 -197.035 ;
        RECT 206.555 -198.725 206.885 -198.395 ;
        RECT 206.555 -200.085 206.885 -199.755 ;
        RECT 206.555 -201.445 206.885 -201.115 ;
        RECT 206.555 -202.805 206.885 -202.475 ;
        RECT 206.555 -204.165 206.885 -203.835 ;
        RECT 206.555 -205.525 206.885 -205.195 ;
        RECT 206.555 -206.885 206.885 -206.555 ;
        RECT 206.555 -208.245 206.885 -207.915 ;
        RECT 206.555 -209.605 206.885 -209.275 ;
        RECT 206.555 -210.965 206.885 -210.635 ;
        RECT 206.555 -212.325 206.885 -211.995 ;
        RECT 206.555 -213.685 206.885 -213.355 ;
        RECT 206.555 -215.045 206.885 -214.715 ;
        RECT 206.555 -216.405 206.885 -216.075 ;
        RECT 206.555 -217.765 206.885 -217.435 ;
        RECT 206.555 -219.125 206.885 -218.795 ;
        RECT 206.555 -220.485 206.885 -220.155 ;
        RECT 206.555 -221.845 206.885 -221.515 ;
        RECT 206.555 -223.205 206.885 -222.875 ;
        RECT 206.555 -224.565 206.885 -224.235 ;
        RECT 206.555 -225.925 206.885 -225.595 ;
        RECT 206.555 -227.285 206.885 -226.955 ;
        RECT 206.555 -228.645 206.885 -228.315 ;
        RECT 206.555 -230.005 206.885 -229.675 ;
        RECT 206.555 -231.365 206.885 -231.035 ;
        RECT 206.555 -232.725 206.885 -232.395 ;
        RECT 206.555 -234.085 206.885 -233.755 ;
        RECT 206.555 -235.445 206.885 -235.115 ;
        RECT 206.555 -236.805 206.885 -236.475 ;
        RECT 206.555 -238.165 206.885 -237.835 ;
        RECT 206.555 -243.81 206.885 -242.68 ;
        RECT 206.56 -243.925 206.88 -122.235 ;
        RECT 206.555 -122.565 206.885 -122.235 ;
        RECT 206.555 -123.925 206.885 -123.595 ;
        RECT 206.555 -125.285 206.885 -124.955 ;
        RECT 206.555 -126.645 206.885 -126.315 ;
        RECT 206.555 -128.005 206.885 -127.675 ;
        RECT 206.555 -129.365 206.885 -129.035 ;
        RECT 206.555 -130.725 206.885 -130.395 ;
        RECT 206.555 -132.085 206.885 -131.755 ;
        RECT 206.555 -133.445 206.885 -133.115 ;
        RECT 206.555 -134.805 206.885 -134.475 ;
        RECT 206.555 -136.165 206.885 -135.835 ;
        RECT 206.555 -137.525 206.885 -137.195 ;
        RECT 206.555 -138.885 206.885 -138.555 ;
        RECT 206.555 -140.245 206.885 -139.915 ;
        RECT 206.555 -141.605 206.885 -141.275 ;
        RECT 206.555 -142.965 206.885 -142.635 ;
        RECT 206.555 -144.325 206.885 -143.995 ;
        RECT 206.555 -145.685 206.885 -145.355 ;
        RECT 206.555 -147.045 206.885 -146.715 ;
        RECT 206.555 -148.405 206.885 -148.075 ;
        RECT 206.555 -149.765 206.885 -149.435 ;
        RECT 206.555 -151.125 206.885 -150.795 ;
        RECT 206.555 -152.485 206.885 -152.155 ;
        RECT 206.555 -153.845 206.885 -153.515 ;
        RECT 206.555 -155.205 206.885 -154.875 ;
        RECT 206.555 -156.565 206.885 -156.235 ;
        RECT 206.555 -157.925 206.885 -157.595 ;
        RECT 206.555 -159.285 206.885 -158.955 ;
        RECT 206.555 -160.645 206.885 -160.315 ;
        RECT 206.555 -162.005 206.885 -161.675 ;
        RECT 206.555 -163.365 206.885 -163.035 ;
        RECT 206.555 -164.725 206.885 -164.395 ;
        RECT 206.555 -166.085 206.885 -165.755 ;
        RECT 206.555 -167.445 206.885 -167.115 ;
        RECT 206.555 -168.805 206.885 -168.475 ;
        RECT 206.555 -170.165 206.885 -169.835 ;
        RECT 206.555 -171.525 206.885 -171.195 ;
        RECT 206.555 -172.885 206.885 -172.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 246.76 166.085 247.89 ;
        RECT 165.755 241.915 166.085 242.245 ;
        RECT 165.755 240.555 166.085 240.885 ;
        RECT 165.755 239.195 166.085 239.525 ;
        RECT 165.755 237.835 166.085 238.165 ;
        RECT 165.76 237.16 166.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 -126.645 166.085 -126.315 ;
        RECT 165.755 -128.005 166.085 -127.675 ;
        RECT 165.755 -129.365 166.085 -129.035 ;
        RECT 165.755 -130.725 166.085 -130.395 ;
        RECT 165.755 -132.085 166.085 -131.755 ;
        RECT 165.755 -133.445 166.085 -133.115 ;
        RECT 165.755 -134.805 166.085 -134.475 ;
        RECT 165.755 -136.165 166.085 -135.835 ;
        RECT 165.755 -137.525 166.085 -137.195 ;
        RECT 165.755 -138.885 166.085 -138.555 ;
        RECT 165.755 -140.245 166.085 -139.915 ;
        RECT 165.755 -141.605 166.085 -141.275 ;
        RECT 165.755 -142.965 166.085 -142.635 ;
        RECT 165.755 -144.325 166.085 -143.995 ;
        RECT 165.755 -145.685 166.085 -145.355 ;
        RECT 165.755 -147.045 166.085 -146.715 ;
        RECT 165.755 -148.405 166.085 -148.075 ;
        RECT 165.755 -149.765 166.085 -149.435 ;
        RECT 165.755 -151.125 166.085 -150.795 ;
        RECT 165.755 -152.485 166.085 -152.155 ;
        RECT 165.755 -153.845 166.085 -153.515 ;
        RECT 165.755 -155.205 166.085 -154.875 ;
        RECT 165.755 -156.565 166.085 -156.235 ;
        RECT 165.755 -157.925 166.085 -157.595 ;
        RECT 165.755 -159.285 166.085 -158.955 ;
        RECT 165.755 -160.645 166.085 -160.315 ;
        RECT 165.755 -162.005 166.085 -161.675 ;
        RECT 165.755 -163.365 166.085 -163.035 ;
        RECT 165.755 -164.725 166.085 -164.395 ;
        RECT 165.755 -166.085 166.085 -165.755 ;
        RECT 165.755 -167.445 166.085 -167.115 ;
        RECT 165.755 -168.805 166.085 -168.475 ;
        RECT 165.755 -170.165 166.085 -169.835 ;
        RECT 165.755 -171.525 166.085 -171.195 ;
        RECT 165.755 -172.885 166.085 -172.555 ;
        RECT 165.755 -174.245 166.085 -173.915 ;
        RECT 165.755 -175.605 166.085 -175.275 ;
        RECT 165.755 -176.965 166.085 -176.635 ;
        RECT 165.755 -178.325 166.085 -177.995 ;
        RECT 165.755 -179.685 166.085 -179.355 ;
        RECT 165.755 -181.045 166.085 -180.715 ;
        RECT 165.755 -182.405 166.085 -182.075 ;
        RECT 165.755 -183.765 166.085 -183.435 ;
        RECT 165.755 -185.125 166.085 -184.795 ;
        RECT 165.755 -186.485 166.085 -186.155 ;
        RECT 165.755 -187.845 166.085 -187.515 ;
        RECT 165.755 -189.205 166.085 -188.875 ;
        RECT 165.755 -190.565 166.085 -190.235 ;
        RECT 165.755 -191.925 166.085 -191.595 ;
        RECT 165.755 -193.285 166.085 -192.955 ;
        RECT 165.755 -194.645 166.085 -194.315 ;
        RECT 165.755 -196.005 166.085 -195.675 ;
        RECT 165.755 -197.365 166.085 -197.035 ;
        RECT 165.755 -198.725 166.085 -198.395 ;
        RECT 165.755 -200.085 166.085 -199.755 ;
        RECT 165.755 -201.445 166.085 -201.115 ;
        RECT 165.755 -202.805 166.085 -202.475 ;
        RECT 165.755 -204.165 166.085 -203.835 ;
        RECT 165.755 -205.525 166.085 -205.195 ;
        RECT 165.755 -206.885 166.085 -206.555 ;
        RECT 165.755 -208.245 166.085 -207.915 ;
        RECT 165.755 -209.605 166.085 -209.275 ;
        RECT 165.755 -210.965 166.085 -210.635 ;
        RECT 165.755 -212.325 166.085 -211.995 ;
        RECT 165.755 -213.685 166.085 -213.355 ;
        RECT 165.755 -215.045 166.085 -214.715 ;
        RECT 165.755 -216.405 166.085 -216.075 ;
        RECT 165.755 -217.765 166.085 -217.435 ;
        RECT 165.755 -219.125 166.085 -218.795 ;
        RECT 165.755 -220.485 166.085 -220.155 ;
        RECT 165.755 -221.845 166.085 -221.515 ;
        RECT 165.755 -223.205 166.085 -222.875 ;
        RECT 165.755 -224.565 166.085 -224.235 ;
        RECT 165.755 -225.925 166.085 -225.595 ;
        RECT 165.755 -227.285 166.085 -226.955 ;
        RECT 165.755 -228.645 166.085 -228.315 ;
        RECT 165.755 -230.005 166.085 -229.675 ;
        RECT 165.755 -231.365 166.085 -231.035 ;
        RECT 165.755 -232.725 166.085 -232.395 ;
        RECT 165.755 -234.085 166.085 -233.755 ;
        RECT 165.755 -235.445 166.085 -235.115 ;
        RECT 165.755 -236.805 166.085 -236.475 ;
        RECT 165.755 -238.165 166.085 -237.835 ;
        RECT 165.755 -243.81 166.085 -242.68 ;
        RECT 165.76 -243.925 166.08 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.16 -125.535 166.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 246.76 167.445 247.89 ;
        RECT 167.115 241.915 167.445 242.245 ;
        RECT 167.115 240.555 167.445 240.885 ;
        RECT 167.115 239.195 167.445 239.525 ;
        RECT 167.115 237.835 167.445 238.165 ;
        RECT 167.12 237.16 167.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 246.76 168.805 247.89 ;
        RECT 168.475 241.915 168.805 242.245 ;
        RECT 168.475 240.555 168.805 240.885 ;
        RECT 168.475 239.195 168.805 239.525 ;
        RECT 168.475 237.835 168.805 238.165 ;
        RECT 168.48 237.16 168.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 -1.525 168.805 -1.195 ;
        RECT 168.475 -2.885 168.805 -2.555 ;
        RECT 168.48 -3.56 168.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 246.76 170.165 247.89 ;
        RECT 169.835 241.915 170.165 242.245 ;
        RECT 169.835 240.555 170.165 240.885 ;
        RECT 169.835 239.195 170.165 239.525 ;
        RECT 169.835 237.835 170.165 238.165 ;
        RECT 169.84 237.16 170.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 -1.525 170.165 -1.195 ;
        RECT 169.835 -2.885 170.165 -2.555 ;
        RECT 169.84 -3.56 170.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 246.76 171.525 247.89 ;
        RECT 171.195 241.915 171.525 242.245 ;
        RECT 171.195 240.555 171.525 240.885 ;
        RECT 171.195 239.195 171.525 239.525 ;
        RECT 171.195 237.835 171.525 238.165 ;
        RECT 171.2 237.16 171.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -1.525 171.525 -1.195 ;
        RECT 171.195 -2.885 171.525 -2.555 ;
        RECT 171.2 -3.56 171.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -122.565 171.525 -122.235 ;
        RECT 171.195 -123.925 171.525 -123.595 ;
        RECT 171.195 -125.285 171.525 -124.955 ;
        RECT 171.195 -126.645 171.525 -126.315 ;
        RECT 171.195 -128.005 171.525 -127.675 ;
        RECT 171.195 -129.365 171.525 -129.035 ;
        RECT 171.195 -130.725 171.525 -130.395 ;
        RECT 171.195 -132.085 171.525 -131.755 ;
        RECT 171.195 -133.445 171.525 -133.115 ;
        RECT 171.195 -134.805 171.525 -134.475 ;
        RECT 171.195 -136.165 171.525 -135.835 ;
        RECT 171.195 -137.525 171.525 -137.195 ;
        RECT 171.195 -138.885 171.525 -138.555 ;
        RECT 171.195 -140.245 171.525 -139.915 ;
        RECT 171.195 -141.605 171.525 -141.275 ;
        RECT 171.195 -142.965 171.525 -142.635 ;
        RECT 171.195 -144.325 171.525 -143.995 ;
        RECT 171.195 -145.685 171.525 -145.355 ;
        RECT 171.195 -147.045 171.525 -146.715 ;
        RECT 171.195 -148.405 171.525 -148.075 ;
        RECT 171.195 -149.765 171.525 -149.435 ;
        RECT 171.195 -151.125 171.525 -150.795 ;
        RECT 171.195 -152.485 171.525 -152.155 ;
        RECT 171.195 -153.845 171.525 -153.515 ;
        RECT 171.195 -155.205 171.525 -154.875 ;
        RECT 171.195 -156.565 171.525 -156.235 ;
        RECT 171.195 -157.925 171.525 -157.595 ;
        RECT 171.195 -159.285 171.525 -158.955 ;
        RECT 171.195 -160.645 171.525 -160.315 ;
        RECT 171.195 -162.005 171.525 -161.675 ;
        RECT 171.195 -163.365 171.525 -163.035 ;
        RECT 171.195 -164.725 171.525 -164.395 ;
        RECT 171.195 -166.085 171.525 -165.755 ;
        RECT 171.195 -167.445 171.525 -167.115 ;
        RECT 171.195 -168.805 171.525 -168.475 ;
        RECT 171.195 -170.165 171.525 -169.835 ;
        RECT 171.195 -171.525 171.525 -171.195 ;
        RECT 171.195 -172.885 171.525 -172.555 ;
        RECT 171.195 -174.245 171.525 -173.915 ;
        RECT 171.195 -175.605 171.525 -175.275 ;
        RECT 171.195 -176.965 171.525 -176.635 ;
        RECT 171.195 -178.325 171.525 -177.995 ;
        RECT 171.195 -179.685 171.525 -179.355 ;
        RECT 171.195 -181.045 171.525 -180.715 ;
        RECT 171.195 -182.405 171.525 -182.075 ;
        RECT 171.195 -183.765 171.525 -183.435 ;
        RECT 171.195 -185.125 171.525 -184.795 ;
        RECT 171.195 -186.485 171.525 -186.155 ;
        RECT 171.195 -187.845 171.525 -187.515 ;
        RECT 171.195 -189.205 171.525 -188.875 ;
        RECT 171.195 -190.565 171.525 -190.235 ;
        RECT 171.195 -191.925 171.525 -191.595 ;
        RECT 171.195 -193.285 171.525 -192.955 ;
        RECT 171.195 -194.645 171.525 -194.315 ;
        RECT 171.195 -196.005 171.525 -195.675 ;
        RECT 171.195 -197.365 171.525 -197.035 ;
        RECT 171.195 -198.725 171.525 -198.395 ;
        RECT 171.195 -200.085 171.525 -199.755 ;
        RECT 171.195 -201.445 171.525 -201.115 ;
        RECT 171.195 -202.805 171.525 -202.475 ;
        RECT 171.195 -204.165 171.525 -203.835 ;
        RECT 171.195 -205.525 171.525 -205.195 ;
        RECT 171.195 -206.885 171.525 -206.555 ;
        RECT 171.195 -208.245 171.525 -207.915 ;
        RECT 171.195 -209.605 171.525 -209.275 ;
        RECT 171.195 -210.965 171.525 -210.635 ;
        RECT 171.195 -212.325 171.525 -211.995 ;
        RECT 171.195 -213.685 171.525 -213.355 ;
        RECT 171.195 -215.045 171.525 -214.715 ;
        RECT 171.195 -216.405 171.525 -216.075 ;
        RECT 171.195 -217.765 171.525 -217.435 ;
        RECT 171.195 -219.125 171.525 -218.795 ;
        RECT 171.195 -220.485 171.525 -220.155 ;
        RECT 171.195 -221.845 171.525 -221.515 ;
        RECT 171.195 -223.205 171.525 -222.875 ;
        RECT 171.195 -224.565 171.525 -224.235 ;
        RECT 171.195 -225.925 171.525 -225.595 ;
        RECT 171.195 -227.285 171.525 -226.955 ;
        RECT 171.195 -228.645 171.525 -228.315 ;
        RECT 171.195 -230.005 171.525 -229.675 ;
        RECT 171.195 -231.365 171.525 -231.035 ;
        RECT 171.195 -232.725 171.525 -232.395 ;
        RECT 171.195 -234.085 171.525 -233.755 ;
        RECT 171.195 -235.445 171.525 -235.115 ;
        RECT 171.195 -236.805 171.525 -236.475 ;
        RECT 171.195 -238.165 171.525 -237.835 ;
        RECT 171.195 -243.81 171.525 -242.68 ;
        RECT 171.2 -243.925 171.52 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 246.76 172.885 247.89 ;
        RECT 172.555 241.915 172.885 242.245 ;
        RECT 172.555 240.555 172.885 240.885 ;
        RECT 172.555 239.195 172.885 239.525 ;
        RECT 172.555 237.835 172.885 238.165 ;
        RECT 172.56 237.16 172.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -1.525 172.885 -1.195 ;
        RECT 172.555 -2.885 172.885 -2.555 ;
        RECT 172.56 -3.56 172.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -122.565 172.885 -122.235 ;
        RECT 172.555 -123.925 172.885 -123.595 ;
        RECT 172.555 -125.285 172.885 -124.955 ;
        RECT 172.555 -126.645 172.885 -126.315 ;
        RECT 172.555 -128.005 172.885 -127.675 ;
        RECT 172.555 -129.365 172.885 -129.035 ;
        RECT 172.555 -130.725 172.885 -130.395 ;
        RECT 172.555 -132.085 172.885 -131.755 ;
        RECT 172.555 -133.445 172.885 -133.115 ;
        RECT 172.555 -134.805 172.885 -134.475 ;
        RECT 172.555 -136.165 172.885 -135.835 ;
        RECT 172.555 -137.525 172.885 -137.195 ;
        RECT 172.555 -138.885 172.885 -138.555 ;
        RECT 172.555 -140.245 172.885 -139.915 ;
        RECT 172.555 -141.605 172.885 -141.275 ;
        RECT 172.555 -142.965 172.885 -142.635 ;
        RECT 172.555 -144.325 172.885 -143.995 ;
        RECT 172.555 -145.685 172.885 -145.355 ;
        RECT 172.555 -147.045 172.885 -146.715 ;
        RECT 172.555 -148.405 172.885 -148.075 ;
        RECT 172.555 -149.765 172.885 -149.435 ;
        RECT 172.555 -151.125 172.885 -150.795 ;
        RECT 172.555 -152.485 172.885 -152.155 ;
        RECT 172.555 -153.845 172.885 -153.515 ;
        RECT 172.555 -155.205 172.885 -154.875 ;
        RECT 172.555 -156.565 172.885 -156.235 ;
        RECT 172.555 -157.925 172.885 -157.595 ;
        RECT 172.555 -159.285 172.885 -158.955 ;
        RECT 172.555 -160.645 172.885 -160.315 ;
        RECT 172.555 -162.005 172.885 -161.675 ;
        RECT 172.555 -163.365 172.885 -163.035 ;
        RECT 172.555 -164.725 172.885 -164.395 ;
        RECT 172.555 -166.085 172.885 -165.755 ;
        RECT 172.555 -167.445 172.885 -167.115 ;
        RECT 172.555 -168.805 172.885 -168.475 ;
        RECT 172.555 -170.165 172.885 -169.835 ;
        RECT 172.555 -171.525 172.885 -171.195 ;
        RECT 172.555 -172.885 172.885 -172.555 ;
        RECT 172.555 -174.245 172.885 -173.915 ;
        RECT 172.555 -175.605 172.885 -175.275 ;
        RECT 172.555 -176.965 172.885 -176.635 ;
        RECT 172.555 -178.325 172.885 -177.995 ;
        RECT 172.555 -179.685 172.885 -179.355 ;
        RECT 172.555 -181.045 172.885 -180.715 ;
        RECT 172.555 -182.405 172.885 -182.075 ;
        RECT 172.555 -183.765 172.885 -183.435 ;
        RECT 172.555 -185.125 172.885 -184.795 ;
        RECT 172.555 -186.485 172.885 -186.155 ;
        RECT 172.555 -187.845 172.885 -187.515 ;
        RECT 172.555 -189.205 172.885 -188.875 ;
        RECT 172.555 -190.565 172.885 -190.235 ;
        RECT 172.555 -191.925 172.885 -191.595 ;
        RECT 172.555 -193.285 172.885 -192.955 ;
        RECT 172.555 -194.645 172.885 -194.315 ;
        RECT 172.555 -196.005 172.885 -195.675 ;
        RECT 172.555 -197.365 172.885 -197.035 ;
        RECT 172.555 -198.725 172.885 -198.395 ;
        RECT 172.555 -200.085 172.885 -199.755 ;
        RECT 172.555 -201.445 172.885 -201.115 ;
        RECT 172.555 -202.805 172.885 -202.475 ;
        RECT 172.555 -204.165 172.885 -203.835 ;
        RECT 172.555 -205.525 172.885 -205.195 ;
        RECT 172.555 -206.885 172.885 -206.555 ;
        RECT 172.555 -208.245 172.885 -207.915 ;
        RECT 172.555 -209.605 172.885 -209.275 ;
        RECT 172.555 -210.965 172.885 -210.635 ;
        RECT 172.555 -212.325 172.885 -211.995 ;
        RECT 172.555 -213.685 172.885 -213.355 ;
        RECT 172.555 -215.045 172.885 -214.715 ;
        RECT 172.555 -216.405 172.885 -216.075 ;
        RECT 172.555 -217.765 172.885 -217.435 ;
        RECT 172.555 -219.125 172.885 -218.795 ;
        RECT 172.555 -220.485 172.885 -220.155 ;
        RECT 172.555 -221.845 172.885 -221.515 ;
        RECT 172.555 -223.205 172.885 -222.875 ;
        RECT 172.555 -224.565 172.885 -224.235 ;
        RECT 172.555 -225.925 172.885 -225.595 ;
        RECT 172.555 -227.285 172.885 -226.955 ;
        RECT 172.555 -228.645 172.885 -228.315 ;
        RECT 172.555 -230.005 172.885 -229.675 ;
        RECT 172.555 -231.365 172.885 -231.035 ;
        RECT 172.555 -232.725 172.885 -232.395 ;
        RECT 172.555 -234.085 172.885 -233.755 ;
        RECT 172.555 -235.445 172.885 -235.115 ;
        RECT 172.555 -236.805 172.885 -236.475 ;
        RECT 172.555 -238.165 172.885 -237.835 ;
        RECT 172.555 -243.81 172.885 -242.68 ;
        RECT 172.56 -243.925 172.88 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 246.76 174.245 247.89 ;
        RECT 173.915 241.915 174.245 242.245 ;
        RECT 173.915 240.555 174.245 240.885 ;
        RECT 173.915 239.195 174.245 239.525 ;
        RECT 173.915 237.835 174.245 238.165 ;
        RECT 173.92 237.16 174.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 -1.525 174.245 -1.195 ;
        RECT 173.915 -2.885 174.245 -2.555 ;
        RECT 173.92 -3.56 174.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 -122.565 174.245 -122.235 ;
        RECT 173.915 -123.925 174.245 -123.595 ;
        RECT 173.915 -125.285 174.245 -124.955 ;
        RECT 173.915 -126.645 174.245 -126.315 ;
        RECT 173.915 -128.005 174.245 -127.675 ;
        RECT 173.915 -129.365 174.245 -129.035 ;
        RECT 173.915 -130.725 174.245 -130.395 ;
        RECT 173.915 -132.085 174.245 -131.755 ;
        RECT 173.915 -133.445 174.245 -133.115 ;
        RECT 173.915 -134.805 174.245 -134.475 ;
        RECT 173.915 -136.165 174.245 -135.835 ;
        RECT 173.915 -137.525 174.245 -137.195 ;
        RECT 173.915 -138.885 174.245 -138.555 ;
        RECT 173.915 -140.245 174.245 -139.915 ;
        RECT 173.915 -141.605 174.245 -141.275 ;
        RECT 173.915 -142.965 174.245 -142.635 ;
        RECT 173.915 -144.325 174.245 -143.995 ;
        RECT 173.915 -145.685 174.245 -145.355 ;
        RECT 173.915 -147.045 174.245 -146.715 ;
        RECT 173.915 -148.405 174.245 -148.075 ;
        RECT 173.915 -149.765 174.245 -149.435 ;
        RECT 173.915 -151.125 174.245 -150.795 ;
        RECT 173.915 -152.485 174.245 -152.155 ;
        RECT 173.915 -153.845 174.245 -153.515 ;
        RECT 173.915 -155.205 174.245 -154.875 ;
        RECT 173.915 -156.565 174.245 -156.235 ;
        RECT 173.915 -157.925 174.245 -157.595 ;
        RECT 173.915 -159.285 174.245 -158.955 ;
        RECT 173.915 -160.645 174.245 -160.315 ;
        RECT 173.915 -162.005 174.245 -161.675 ;
        RECT 173.915 -163.365 174.245 -163.035 ;
        RECT 173.915 -164.725 174.245 -164.395 ;
        RECT 173.915 -166.085 174.245 -165.755 ;
        RECT 173.915 -167.445 174.245 -167.115 ;
        RECT 173.915 -168.805 174.245 -168.475 ;
        RECT 173.915 -170.165 174.245 -169.835 ;
        RECT 173.915 -171.525 174.245 -171.195 ;
        RECT 173.915 -172.885 174.245 -172.555 ;
        RECT 173.915 -174.245 174.245 -173.915 ;
        RECT 173.915 -175.605 174.245 -175.275 ;
        RECT 173.915 -176.965 174.245 -176.635 ;
        RECT 173.915 -178.325 174.245 -177.995 ;
        RECT 173.915 -179.685 174.245 -179.355 ;
        RECT 173.915 -181.045 174.245 -180.715 ;
        RECT 173.915 -182.405 174.245 -182.075 ;
        RECT 173.915 -183.765 174.245 -183.435 ;
        RECT 173.915 -185.125 174.245 -184.795 ;
        RECT 173.915 -186.485 174.245 -186.155 ;
        RECT 173.915 -187.845 174.245 -187.515 ;
        RECT 173.915 -189.205 174.245 -188.875 ;
        RECT 173.915 -190.565 174.245 -190.235 ;
        RECT 173.915 -191.925 174.245 -191.595 ;
        RECT 173.915 -193.285 174.245 -192.955 ;
        RECT 173.915 -194.645 174.245 -194.315 ;
        RECT 173.915 -196.005 174.245 -195.675 ;
        RECT 173.915 -197.365 174.245 -197.035 ;
        RECT 173.915 -198.725 174.245 -198.395 ;
        RECT 173.915 -200.085 174.245 -199.755 ;
        RECT 173.915 -201.445 174.245 -201.115 ;
        RECT 173.915 -202.805 174.245 -202.475 ;
        RECT 173.915 -204.165 174.245 -203.835 ;
        RECT 173.915 -205.525 174.245 -205.195 ;
        RECT 173.915 -206.885 174.245 -206.555 ;
        RECT 173.915 -208.245 174.245 -207.915 ;
        RECT 173.915 -209.605 174.245 -209.275 ;
        RECT 173.915 -210.965 174.245 -210.635 ;
        RECT 173.915 -212.325 174.245 -211.995 ;
        RECT 173.915 -213.685 174.245 -213.355 ;
        RECT 173.915 -215.045 174.245 -214.715 ;
        RECT 173.915 -216.405 174.245 -216.075 ;
        RECT 173.915 -217.765 174.245 -217.435 ;
        RECT 173.915 -219.125 174.245 -218.795 ;
        RECT 173.915 -220.485 174.245 -220.155 ;
        RECT 173.915 -221.845 174.245 -221.515 ;
        RECT 173.915 -223.205 174.245 -222.875 ;
        RECT 173.915 -224.565 174.245 -224.235 ;
        RECT 173.915 -225.925 174.245 -225.595 ;
        RECT 173.915 -227.285 174.245 -226.955 ;
        RECT 173.915 -228.645 174.245 -228.315 ;
        RECT 173.915 -230.005 174.245 -229.675 ;
        RECT 173.915 -231.365 174.245 -231.035 ;
        RECT 173.915 -232.725 174.245 -232.395 ;
        RECT 173.915 -234.085 174.245 -233.755 ;
        RECT 173.915 -235.445 174.245 -235.115 ;
        RECT 173.915 -236.805 174.245 -236.475 ;
        RECT 173.915 -238.165 174.245 -237.835 ;
        RECT 173.915 -243.81 174.245 -242.68 ;
        RECT 173.92 -243.925 174.24 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 246.76 175.605 247.89 ;
        RECT 175.275 241.915 175.605 242.245 ;
        RECT 175.275 240.555 175.605 240.885 ;
        RECT 175.275 239.195 175.605 239.525 ;
        RECT 175.275 237.835 175.605 238.165 ;
        RECT 175.28 237.16 175.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -1.525 175.605 -1.195 ;
        RECT 175.275 -2.885 175.605 -2.555 ;
        RECT 175.28 -3.56 175.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -122.565 175.605 -122.235 ;
        RECT 175.275 -123.925 175.605 -123.595 ;
        RECT 175.275 -125.285 175.605 -124.955 ;
        RECT 175.275 -126.645 175.605 -126.315 ;
        RECT 175.275 -128.005 175.605 -127.675 ;
        RECT 175.275 -129.365 175.605 -129.035 ;
        RECT 175.275 -130.725 175.605 -130.395 ;
        RECT 175.275 -132.085 175.605 -131.755 ;
        RECT 175.275 -133.445 175.605 -133.115 ;
        RECT 175.275 -134.805 175.605 -134.475 ;
        RECT 175.275 -136.165 175.605 -135.835 ;
        RECT 175.275 -137.525 175.605 -137.195 ;
        RECT 175.275 -138.885 175.605 -138.555 ;
        RECT 175.275 -140.245 175.605 -139.915 ;
        RECT 175.275 -141.605 175.605 -141.275 ;
        RECT 175.275 -142.965 175.605 -142.635 ;
        RECT 175.275 -144.325 175.605 -143.995 ;
        RECT 175.275 -145.685 175.605 -145.355 ;
        RECT 175.275 -147.045 175.605 -146.715 ;
        RECT 175.275 -148.405 175.605 -148.075 ;
        RECT 175.275 -149.765 175.605 -149.435 ;
        RECT 175.275 -151.125 175.605 -150.795 ;
        RECT 175.275 -152.485 175.605 -152.155 ;
        RECT 175.275 -153.845 175.605 -153.515 ;
        RECT 175.275 -155.205 175.605 -154.875 ;
        RECT 175.275 -156.565 175.605 -156.235 ;
        RECT 175.275 -157.925 175.605 -157.595 ;
        RECT 175.275 -159.285 175.605 -158.955 ;
        RECT 175.275 -160.645 175.605 -160.315 ;
        RECT 175.275 -162.005 175.605 -161.675 ;
        RECT 175.275 -163.365 175.605 -163.035 ;
        RECT 175.275 -164.725 175.605 -164.395 ;
        RECT 175.275 -166.085 175.605 -165.755 ;
        RECT 175.275 -167.445 175.605 -167.115 ;
        RECT 175.275 -168.805 175.605 -168.475 ;
        RECT 175.275 -170.165 175.605 -169.835 ;
        RECT 175.275 -171.525 175.605 -171.195 ;
        RECT 175.275 -172.885 175.605 -172.555 ;
        RECT 175.275 -174.245 175.605 -173.915 ;
        RECT 175.275 -175.605 175.605 -175.275 ;
        RECT 175.275 -176.965 175.605 -176.635 ;
        RECT 175.275 -178.325 175.605 -177.995 ;
        RECT 175.275 -179.685 175.605 -179.355 ;
        RECT 175.275 -181.045 175.605 -180.715 ;
        RECT 175.275 -182.405 175.605 -182.075 ;
        RECT 175.275 -183.765 175.605 -183.435 ;
        RECT 175.275 -185.125 175.605 -184.795 ;
        RECT 175.275 -186.485 175.605 -186.155 ;
        RECT 175.275 -187.845 175.605 -187.515 ;
        RECT 175.275 -189.205 175.605 -188.875 ;
        RECT 175.275 -190.565 175.605 -190.235 ;
        RECT 175.275 -191.925 175.605 -191.595 ;
        RECT 175.275 -193.285 175.605 -192.955 ;
        RECT 175.275 -194.645 175.605 -194.315 ;
        RECT 175.275 -196.005 175.605 -195.675 ;
        RECT 175.275 -197.365 175.605 -197.035 ;
        RECT 175.275 -198.725 175.605 -198.395 ;
        RECT 175.275 -200.085 175.605 -199.755 ;
        RECT 175.275 -201.445 175.605 -201.115 ;
        RECT 175.275 -202.805 175.605 -202.475 ;
        RECT 175.275 -204.165 175.605 -203.835 ;
        RECT 175.275 -205.525 175.605 -205.195 ;
        RECT 175.275 -206.885 175.605 -206.555 ;
        RECT 175.275 -208.245 175.605 -207.915 ;
        RECT 175.275 -209.605 175.605 -209.275 ;
        RECT 175.275 -210.965 175.605 -210.635 ;
        RECT 175.275 -212.325 175.605 -211.995 ;
        RECT 175.275 -213.685 175.605 -213.355 ;
        RECT 175.275 -215.045 175.605 -214.715 ;
        RECT 175.275 -216.405 175.605 -216.075 ;
        RECT 175.275 -217.765 175.605 -217.435 ;
        RECT 175.275 -219.125 175.605 -218.795 ;
        RECT 175.275 -220.485 175.605 -220.155 ;
        RECT 175.275 -221.845 175.605 -221.515 ;
        RECT 175.275 -223.205 175.605 -222.875 ;
        RECT 175.275 -224.565 175.605 -224.235 ;
        RECT 175.275 -225.925 175.605 -225.595 ;
        RECT 175.275 -227.285 175.605 -226.955 ;
        RECT 175.275 -228.645 175.605 -228.315 ;
        RECT 175.275 -230.005 175.605 -229.675 ;
        RECT 175.275 -231.365 175.605 -231.035 ;
        RECT 175.275 -232.725 175.605 -232.395 ;
        RECT 175.275 -234.085 175.605 -233.755 ;
        RECT 175.275 -235.445 175.605 -235.115 ;
        RECT 175.275 -236.805 175.605 -236.475 ;
        RECT 175.275 -238.165 175.605 -237.835 ;
        RECT 175.275 -243.81 175.605 -242.68 ;
        RECT 175.28 -243.925 175.6 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 246.76 176.965 247.89 ;
        RECT 176.635 241.915 176.965 242.245 ;
        RECT 176.635 240.555 176.965 240.885 ;
        RECT 176.635 239.195 176.965 239.525 ;
        RECT 176.635 237.835 176.965 238.165 ;
        RECT 176.64 237.16 176.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 -126.645 176.965 -126.315 ;
        RECT 176.635 -128.005 176.965 -127.675 ;
        RECT 176.635 -129.365 176.965 -129.035 ;
        RECT 176.635 -130.725 176.965 -130.395 ;
        RECT 176.635 -132.085 176.965 -131.755 ;
        RECT 176.635 -133.445 176.965 -133.115 ;
        RECT 176.635 -134.805 176.965 -134.475 ;
        RECT 176.635 -136.165 176.965 -135.835 ;
        RECT 176.635 -137.525 176.965 -137.195 ;
        RECT 176.635 -138.885 176.965 -138.555 ;
        RECT 176.635 -140.245 176.965 -139.915 ;
        RECT 176.635 -141.605 176.965 -141.275 ;
        RECT 176.635 -142.965 176.965 -142.635 ;
        RECT 176.635 -144.325 176.965 -143.995 ;
        RECT 176.635 -145.685 176.965 -145.355 ;
        RECT 176.635 -147.045 176.965 -146.715 ;
        RECT 176.635 -148.405 176.965 -148.075 ;
        RECT 176.635 -149.765 176.965 -149.435 ;
        RECT 176.635 -151.125 176.965 -150.795 ;
        RECT 176.635 -152.485 176.965 -152.155 ;
        RECT 176.635 -153.845 176.965 -153.515 ;
        RECT 176.635 -155.205 176.965 -154.875 ;
        RECT 176.635 -156.565 176.965 -156.235 ;
        RECT 176.635 -157.925 176.965 -157.595 ;
        RECT 176.635 -159.285 176.965 -158.955 ;
        RECT 176.635 -160.645 176.965 -160.315 ;
        RECT 176.635 -162.005 176.965 -161.675 ;
        RECT 176.635 -163.365 176.965 -163.035 ;
        RECT 176.635 -164.725 176.965 -164.395 ;
        RECT 176.635 -166.085 176.965 -165.755 ;
        RECT 176.635 -167.445 176.965 -167.115 ;
        RECT 176.635 -168.805 176.965 -168.475 ;
        RECT 176.635 -170.165 176.965 -169.835 ;
        RECT 176.635 -171.525 176.965 -171.195 ;
        RECT 176.635 -172.885 176.965 -172.555 ;
        RECT 176.635 -174.245 176.965 -173.915 ;
        RECT 176.635 -175.605 176.965 -175.275 ;
        RECT 176.635 -176.965 176.965 -176.635 ;
        RECT 176.635 -178.325 176.965 -177.995 ;
        RECT 176.635 -179.685 176.965 -179.355 ;
        RECT 176.635 -181.045 176.965 -180.715 ;
        RECT 176.635 -182.405 176.965 -182.075 ;
        RECT 176.635 -183.765 176.965 -183.435 ;
        RECT 176.635 -185.125 176.965 -184.795 ;
        RECT 176.635 -186.485 176.965 -186.155 ;
        RECT 176.635 -187.845 176.965 -187.515 ;
        RECT 176.635 -189.205 176.965 -188.875 ;
        RECT 176.635 -190.565 176.965 -190.235 ;
        RECT 176.635 -191.925 176.965 -191.595 ;
        RECT 176.635 -193.285 176.965 -192.955 ;
        RECT 176.635 -194.645 176.965 -194.315 ;
        RECT 176.635 -196.005 176.965 -195.675 ;
        RECT 176.635 -197.365 176.965 -197.035 ;
        RECT 176.635 -198.725 176.965 -198.395 ;
        RECT 176.635 -200.085 176.965 -199.755 ;
        RECT 176.635 -201.445 176.965 -201.115 ;
        RECT 176.635 -202.805 176.965 -202.475 ;
        RECT 176.635 -204.165 176.965 -203.835 ;
        RECT 176.635 -205.525 176.965 -205.195 ;
        RECT 176.635 -206.885 176.965 -206.555 ;
        RECT 176.635 -208.245 176.965 -207.915 ;
        RECT 176.635 -209.605 176.965 -209.275 ;
        RECT 176.635 -210.965 176.965 -210.635 ;
        RECT 176.635 -212.325 176.965 -211.995 ;
        RECT 176.635 -213.685 176.965 -213.355 ;
        RECT 176.635 -215.045 176.965 -214.715 ;
        RECT 176.635 -216.405 176.965 -216.075 ;
        RECT 176.635 -217.765 176.965 -217.435 ;
        RECT 176.635 -219.125 176.965 -218.795 ;
        RECT 176.635 -220.485 176.965 -220.155 ;
        RECT 176.635 -221.845 176.965 -221.515 ;
        RECT 176.635 -223.205 176.965 -222.875 ;
        RECT 176.635 -224.565 176.965 -224.235 ;
        RECT 176.635 -225.925 176.965 -225.595 ;
        RECT 176.635 -227.285 176.965 -226.955 ;
        RECT 176.635 -228.645 176.965 -228.315 ;
        RECT 176.635 -230.005 176.965 -229.675 ;
        RECT 176.635 -231.365 176.965 -231.035 ;
        RECT 176.635 -232.725 176.965 -232.395 ;
        RECT 176.635 -234.085 176.965 -233.755 ;
        RECT 176.635 -235.445 176.965 -235.115 ;
        RECT 176.635 -236.805 176.965 -236.475 ;
        RECT 176.635 -238.165 176.965 -237.835 ;
        RECT 176.635 -243.81 176.965 -242.68 ;
        RECT 176.64 -243.925 176.96 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.06 -125.535 177.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 246.76 178.325 247.89 ;
        RECT 177.995 241.915 178.325 242.245 ;
        RECT 177.995 240.555 178.325 240.885 ;
        RECT 177.995 239.195 178.325 239.525 ;
        RECT 177.995 237.835 178.325 238.165 ;
        RECT 178 237.16 178.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 246.76 179.685 247.89 ;
        RECT 179.355 241.915 179.685 242.245 ;
        RECT 179.355 240.555 179.685 240.885 ;
        RECT 179.355 239.195 179.685 239.525 ;
        RECT 179.355 237.835 179.685 238.165 ;
        RECT 179.36 237.16 179.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 -1.525 179.685 -1.195 ;
        RECT 179.355 -2.885 179.685 -2.555 ;
        RECT 179.36 -3.56 179.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 246.76 181.045 247.89 ;
        RECT 180.715 241.915 181.045 242.245 ;
        RECT 180.715 240.555 181.045 240.885 ;
        RECT 180.715 239.195 181.045 239.525 ;
        RECT 180.715 237.835 181.045 238.165 ;
        RECT 180.72 237.16 181.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 -1.525 181.045 -1.195 ;
        RECT 180.715 -2.885 181.045 -2.555 ;
        RECT 180.72 -3.56 181.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 246.76 182.405 247.89 ;
        RECT 182.075 241.915 182.405 242.245 ;
        RECT 182.075 240.555 182.405 240.885 ;
        RECT 182.075 239.195 182.405 239.525 ;
        RECT 182.075 237.835 182.405 238.165 ;
        RECT 182.08 237.16 182.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 -1.525 182.405 -1.195 ;
        RECT 182.075 -2.885 182.405 -2.555 ;
        RECT 182.08 -3.56 182.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 -122.565 182.405 -122.235 ;
        RECT 182.075 -123.925 182.405 -123.595 ;
        RECT 182.075 -125.285 182.405 -124.955 ;
        RECT 182.075 -126.645 182.405 -126.315 ;
        RECT 182.075 -128.005 182.405 -127.675 ;
        RECT 182.075 -129.365 182.405 -129.035 ;
        RECT 182.075 -130.725 182.405 -130.395 ;
        RECT 182.075 -132.085 182.405 -131.755 ;
        RECT 182.075 -133.445 182.405 -133.115 ;
        RECT 182.075 -134.805 182.405 -134.475 ;
        RECT 182.075 -136.165 182.405 -135.835 ;
        RECT 182.075 -137.525 182.405 -137.195 ;
        RECT 182.075 -138.885 182.405 -138.555 ;
        RECT 182.075 -140.245 182.405 -139.915 ;
        RECT 182.075 -141.605 182.405 -141.275 ;
        RECT 182.075 -142.965 182.405 -142.635 ;
        RECT 182.075 -144.325 182.405 -143.995 ;
        RECT 182.075 -145.685 182.405 -145.355 ;
        RECT 182.075 -147.045 182.405 -146.715 ;
        RECT 182.075 -148.405 182.405 -148.075 ;
        RECT 182.075 -149.765 182.405 -149.435 ;
        RECT 182.075 -151.125 182.405 -150.795 ;
        RECT 182.075 -152.485 182.405 -152.155 ;
        RECT 182.075 -153.845 182.405 -153.515 ;
        RECT 182.075 -155.205 182.405 -154.875 ;
        RECT 182.075 -156.565 182.405 -156.235 ;
        RECT 182.075 -157.925 182.405 -157.595 ;
        RECT 182.075 -159.285 182.405 -158.955 ;
        RECT 182.075 -160.645 182.405 -160.315 ;
        RECT 182.075 -162.005 182.405 -161.675 ;
        RECT 182.075 -163.365 182.405 -163.035 ;
        RECT 182.075 -164.725 182.405 -164.395 ;
        RECT 182.075 -166.085 182.405 -165.755 ;
        RECT 182.075 -167.445 182.405 -167.115 ;
        RECT 182.075 -168.805 182.405 -168.475 ;
        RECT 182.075 -170.165 182.405 -169.835 ;
        RECT 182.075 -171.525 182.405 -171.195 ;
        RECT 182.075 -172.885 182.405 -172.555 ;
        RECT 182.075 -174.245 182.405 -173.915 ;
        RECT 182.075 -175.605 182.405 -175.275 ;
        RECT 182.075 -176.965 182.405 -176.635 ;
        RECT 182.075 -178.325 182.405 -177.995 ;
        RECT 182.075 -179.685 182.405 -179.355 ;
        RECT 182.075 -181.045 182.405 -180.715 ;
        RECT 182.075 -182.405 182.405 -182.075 ;
        RECT 182.075 -183.765 182.405 -183.435 ;
        RECT 182.075 -185.125 182.405 -184.795 ;
        RECT 182.075 -186.485 182.405 -186.155 ;
        RECT 182.075 -187.845 182.405 -187.515 ;
        RECT 182.075 -189.205 182.405 -188.875 ;
        RECT 182.075 -190.565 182.405 -190.235 ;
        RECT 182.075 -191.925 182.405 -191.595 ;
        RECT 182.075 -193.285 182.405 -192.955 ;
        RECT 182.075 -194.645 182.405 -194.315 ;
        RECT 182.075 -196.005 182.405 -195.675 ;
        RECT 182.075 -197.365 182.405 -197.035 ;
        RECT 182.075 -198.725 182.405 -198.395 ;
        RECT 182.075 -200.085 182.405 -199.755 ;
        RECT 182.075 -201.445 182.405 -201.115 ;
        RECT 182.075 -202.805 182.405 -202.475 ;
        RECT 182.075 -204.165 182.405 -203.835 ;
        RECT 182.075 -205.525 182.405 -205.195 ;
        RECT 182.075 -206.885 182.405 -206.555 ;
        RECT 182.075 -208.245 182.405 -207.915 ;
        RECT 182.075 -209.605 182.405 -209.275 ;
        RECT 182.075 -210.965 182.405 -210.635 ;
        RECT 182.075 -212.325 182.405 -211.995 ;
        RECT 182.075 -213.685 182.405 -213.355 ;
        RECT 182.075 -215.045 182.405 -214.715 ;
        RECT 182.075 -216.405 182.405 -216.075 ;
        RECT 182.075 -217.765 182.405 -217.435 ;
        RECT 182.075 -219.125 182.405 -218.795 ;
        RECT 182.075 -220.485 182.405 -220.155 ;
        RECT 182.075 -221.845 182.405 -221.515 ;
        RECT 182.075 -223.205 182.405 -222.875 ;
        RECT 182.075 -224.565 182.405 -224.235 ;
        RECT 182.075 -225.925 182.405 -225.595 ;
        RECT 182.075 -227.285 182.405 -226.955 ;
        RECT 182.075 -228.645 182.405 -228.315 ;
        RECT 182.075 -230.005 182.405 -229.675 ;
        RECT 182.075 -231.365 182.405 -231.035 ;
        RECT 182.075 -232.725 182.405 -232.395 ;
        RECT 182.075 -234.085 182.405 -233.755 ;
        RECT 182.075 -235.445 182.405 -235.115 ;
        RECT 182.075 -236.805 182.405 -236.475 ;
        RECT 182.075 -238.165 182.405 -237.835 ;
        RECT 182.075 -243.81 182.405 -242.68 ;
        RECT 182.08 -243.925 182.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 246.76 183.765 247.89 ;
        RECT 183.435 241.915 183.765 242.245 ;
        RECT 183.435 240.555 183.765 240.885 ;
        RECT 183.435 239.195 183.765 239.525 ;
        RECT 183.435 237.835 183.765 238.165 ;
        RECT 183.44 237.16 183.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -1.525 183.765 -1.195 ;
        RECT 183.435 -2.885 183.765 -2.555 ;
        RECT 183.44 -3.56 183.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -122.565 183.765 -122.235 ;
        RECT 183.435 -123.925 183.765 -123.595 ;
        RECT 183.435 -125.285 183.765 -124.955 ;
        RECT 183.435 -126.645 183.765 -126.315 ;
        RECT 183.435 -128.005 183.765 -127.675 ;
        RECT 183.435 -129.365 183.765 -129.035 ;
        RECT 183.435 -130.725 183.765 -130.395 ;
        RECT 183.435 -132.085 183.765 -131.755 ;
        RECT 183.435 -133.445 183.765 -133.115 ;
        RECT 183.435 -134.805 183.765 -134.475 ;
        RECT 183.435 -136.165 183.765 -135.835 ;
        RECT 183.435 -137.525 183.765 -137.195 ;
        RECT 183.435 -138.885 183.765 -138.555 ;
        RECT 183.435 -140.245 183.765 -139.915 ;
        RECT 183.435 -141.605 183.765 -141.275 ;
        RECT 183.435 -142.965 183.765 -142.635 ;
        RECT 183.435 -144.325 183.765 -143.995 ;
        RECT 183.435 -145.685 183.765 -145.355 ;
        RECT 183.435 -147.045 183.765 -146.715 ;
        RECT 183.435 -148.405 183.765 -148.075 ;
        RECT 183.435 -149.765 183.765 -149.435 ;
        RECT 183.435 -151.125 183.765 -150.795 ;
        RECT 183.435 -152.485 183.765 -152.155 ;
        RECT 183.435 -153.845 183.765 -153.515 ;
        RECT 183.435 -155.205 183.765 -154.875 ;
        RECT 183.435 -156.565 183.765 -156.235 ;
        RECT 183.435 -157.925 183.765 -157.595 ;
        RECT 183.435 -159.285 183.765 -158.955 ;
        RECT 183.435 -160.645 183.765 -160.315 ;
        RECT 183.435 -162.005 183.765 -161.675 ;
        RECT 183.435 -163.365 183.765 -163.035 ;
        RECT 183.435 -164.725 183.765 -164.395 ;
        RECT 183.435 -166.085 183.765 -165.755 ;
        RECT 183.435 -167.445 183.765 -167.115 ;
        RECT 183.435 -168.805 183.765 -168.475 ;
        RECT 183.435 -170.165 183.765 -169.835 ;
        RECT 183.435 -171.525 183.765 -171.195 ;
        RECT 183.435 -172.885 183.765 -172.555 ;
        RECT 183.435 -174.245 183.765 -173.915 ;
        RECT 183.435 -175.605 183.765 -175.275 ;
        RECT 183.435 -176.965 183.765 -176.635 ;
        RECT 183.435 -178.325 183.765 -177.995 ;
        RECT 183.435 -179.685 183.765 -179.355 ;
        RECT 183.435 -181.045 183.765 -180.715 ;
        RECT 183.435 -182.405 183.765 -182.075 ;
        RECT 183.435 -183.765 183.765 -183.435 ;
        RECT 183.435 -185.125 183.765 -184.795 ;
        RECT 183.435 -186.485 183.765 -186.155 ;
        RECT 183.435 -187.845 183.765 -187.515 ;
        RECT 183.435 -189.205 183.765 -188.875 ;
        RECT 183.435 -190.565 183.765 -190.235 ;
        RECT 183.435 -191.925 183.765 -191.595 ;
        RECT 183.435 -193.285 183.765 -192.955 ;
        RECT 183.435 -194.645 183.765 -194.315 ;
        RECT 183.435 -196.005 183.765 -195.675 ;
        RECT 183.435 -197.365 183.765 -197.035 ;
        RECT 183.435 -198.725 183.765 -198.395 ;
        RECT 183.435 -200.085 183.765 -199.755 ;
        RECT 183.435 -201.445 183.765 -201.115 ;
        RECT 183.435 -202.805 183.765 -202.475 ;
        RECT 183.435 -204.165 183.765 -203.835 ;
        RECT 183.435 -205.525 183.765 -205.195 ;
        RECT 183.435 -206.885 183.765 -206.555 ;
        RECT 183.435 -208.245 183.765 -207.915 ;
        RECT 183.435 -209.605 183.765 -209.275 ;
        RECT 183.435 -210.965 183.765 -210.635 ;
        RECT 183.435 -212.325 183.765 -211.995 ;
        RECT 183.435 -213.685 183.765 -213.355 ;
        RECT 183.435 -215.045 183.765 -214.715 ;
        RECT 183.435 -216.405 183.765 -216.075 ;
        RECT 183.435 -217.765 183.765 -217.435 ;
        RECT 183.435 -219.125 183.765 -218.795 ;
        RECT 183.435 -220.485 183.765 -220.155 ;
        RECT 183.435 -221.845 183.765 -221.515 ;
        RECT 183.435 -223.205 183.765 -222.875 ;
        RECT 183.435 -224.565 183.765 -224.235 ;
        RECT 183.435 -225.925 183.765 -225.595 ;
        RECT 183.435 -227.285 183.765 -226.955 ;
        RECT 183.435 -228.645 183.765 -228.315 ;
        RECT 183.435 -230.005 183.765 -229.675 ;
        RECT 183.435 -231.365 183.765 -231.035 ;
        RECT 183.435 -232.725 183.765 -232.395 ;
        RECT 183.435 -234.085 183.765 -233.755 ;
        RECT 183.435 -235.445 183.765 -235.115 ;
        RECT 183.435 -236.805 183.765 -236.475 ;
        RECT 183.435 -238.165 183.765 -237.835 ;
        RECT 183.435 -243.81 183.765 -242.68 ;
        RECT 183.44 -243.925 183.76 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 246.76 185.125 247.89 ;
        RECT 184.795 241.915 185.125 242.245 ;
        RECT 184.795 240.555 185.125 240.885 ;
        RECT 184.795 239.195 185.125 239.525 ;
        RECT 184.795 237.835 185.125 238.165 ;
        RECT 184.8 237.16 185.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -1.525 185.125 -1.195 ;
        RECT 184.795 -2.885 185.125 -2.555 ;
        RECT 184.8 -3.56 185.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -122.565 185.125 -122.235 ;
        RECT 184.795 -123.925 185.125 -123.595 ;
        RECT 184.795 -125.285 185.125 -124.955 ;
        RECT 184.795 -126.645 185.125 -126.315 ;
        RECT 184.795 -128.005 185.125 -127.675 ;
        RECT 184.795 -129.365 185.125 -129.035 ;
        RECT 184.795 -130.725 185.125 -130.395 ;
        RECT 184.795 -132.085 185.125 -131.755 ;
        RECT 184.795 -133.445 185.125 -133.115 ;
        RECT 184.795 -134.805 185.125 -134.475 ;
        RECT 184.795 -136.165 185.125 -135.835 ;
        RECT 184.795 -137.525 185.125 -137.195 ;
        RECT 184.795 -138.885 185.125 -138.555 ;
        RECT 184.795 -140.245 185.125 -139.915 ;
        RECT 184.795 -141.605 185.125 -141.275 ;
        RECT 184.795 -142.965 185.125 -142.635 ;
        RECT 184.795 -144.325 185.125 -143.995 ;
        RECT 184.795 -145.685 185.125 -145.355 ;
        RECT 184.795 -147.045 185.125 -146.715 ;
        RECT 184.795 -148.405 185.125 -148.075 ;
        RECT 184.795 -149.765 185.125 -149.435 ;
        RECT 184.795 -151.125 185.125 -150.795 ;
        RECT 184.795 -152.485 185.125 -152.155 ;
        RECT 184.795 -153.845 185.125 -153.515 ;
        RECT 184.795 -155.205 185.125 -154.875 ;
        RECT 184.795 -156.565 185.125 -156.235 ;
        RECT 184.795 -157.925 185.125 -157.595 ;
        RECT 184.795 -159.285 185.125 -158.955 ;
        RECT 184.795 -160.645 185.125 -160.315 ;
        RECT 184.795 -162.005 185.125 -161.675 ;
        RECT 184.795 -163.365 185.125 -163.035 ;
        RECT 184.795 -164.725 185.125 -164.395 ;
        RECT 184.795 -166.085 185.125 -165.755 ;
        RECT 184.795 -167.445 185.125 -167.115 ;
        RECT 184.795 -168.805 185.125 -168.475 ;
        RECT 184.795 -170.165 185.125 -169.835 ;
        RECT 184.795 -171.525 185.125 -171.195 ;
        RECT 184.795 -172.885 185.125 -172.555 ;
        RECT 184.795 -174.245 185.125 -173.915 ;
        RECT 184.795 -175.605 185.125 -175.275 ;
        RECT 184.795 -176.965 185.125 -176.635 ;
        RECT 184.795 -178.325 185.125 -177.995 ;
        RECT 184.795 -179.685 185.125 -179.355 ;
        RECT 184.795 -181.045 185.125 -180.715 ;
        RECT 184.795 -182.405 185.125 -182.075 ;
        RECT 184.795 -183.765 185.125 -183.435 ;
        RECT 184.795 -185.125 185.125 -184.795 ;
        RECT 184.795 -186.485 185.125 -186.155 ;
        RECT 184.795 -187.845 185.125 -187.515 ;
        RECT 184.795 -189.205 185.125 -188.875 ;
        RECT 184.795 -190.565 185.125 -190.235 ;
        RECT 184.795 -191.925 185.125 -191.595 ;
        RECT 184.795 -193.285 185.125 -192.955 ;
        RECT 184.795 -194.645 185.125 -194.315 ;
        RECT 184.795 -196.005 185.125 -195.675 ;
        RECT 184.795 -197.365 185.125 -197.035 ;
        RECT 184.795 -198.725 185.125 -198.395 ;
        RECT 184.795 -200.085 185.125 -199.755 ;
        RECT 184.795 -201.445 185.125 -201.115 ;
        RECT 184.795 -202.805 185.125 -202.475 ;
        RECT 184.795 -204.165 185.125 -203.835 ;
        RECT 184.795 -205.525 185.125 -205.195 ;
        RECT 184.795 -206.885 185.125 -206.555 ;
        RECT 184.795 -208.245 185.125 -207.915 ;
        RECT 184.795 -209.605 185.125 -209.275 ;
        RECT 184.795 -210.965 185.125 -210.635 ;
        RECT 184.795 -212.325 185.125 -211.995 ;
        RECT 184.795 -213.685 185.125 -213.355 ;
        RECT 184.795 -215.045 185.125 -214.715 ;
        RECT 184.795 -216.405 185.125 -216.075 ;
        RECT 184.795 -217.765 185.125 -217.435 ;
        RECT 184.795 -219.125 185.125 -218.795 ;
        RECT 184.795 -220.485 185.125 -220.155 ;
        RECT 184.795 -221.845 185.125 -221.515 ;
        RECT 184.795 -223.205 185.125 -222.875 ;
        RECT 184.795 -224.565 185.125 -224.235 ;
        RECT 184.795 -225.925 185.125 -225.595 ;
        RECT 184.795 -227.285 185.125 -226.955 ;
        RECT 184.795 -228.645 185.125 -228.315 ;
        RECT 184.795 -230.005 185.125 -229.675 ;
        RECT 184.795 -231.365 185.125 -231.035 ;
        RECT 184.795 -232.725 185.125 -232.395 ;
        RECT 184.795 -234.085 185.125 -233.755 ;
        RECT 184.795 -235.445 185.125 -235.115 ;
        RECT 184.795 -236.805 185.125 -236.475 ;
        RECT 184.795 -238.165 185.125 -237.835 ;
        RECT 184.795 -243.81 185.125 -242.68 ;
        RECT 184.8 -243.925 185.12 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 246.76 186.485 247.89 ;
        RECT 186.155 241.915 186.485 242.245 ;
        RECT 186.155 240.555 186.485 240.885 ;
        RECT 186.155 239.195 186.485 239.525 ;
        RECT 186.155 237.835 186.485 238.165 ;
        RECT 186.16 237.16 186.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 -1.525 186.485 -1.195 ;
        RECT 186.155 -2.885 186.485 -2.555 ;
        RECT 186.16 -3.56 186.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 -175.605 186.485 -175.275 ;
        RECT 186.155 -176.965 186.485 -176.635 ;
        RECT 186.155 -178.325 186.485 -177.995 ;
        RECT 186.155 -179.685 186.485 -179.355 ;
        RECT 186.155 -181.045 186.485 -180.715 ;
        RECT 186.155 -182.405 186.485 -182.075 ;
        RECT 186.155 -183.765 186.485 -183.435 ;
        RECT 186.155 -185.125 186.485 -184.795 ;
        RECT 186.155 -186.485 186.485 -186.155 ;
        RECT 186.155 -187.845 186.485 -187.515 ;
        RECT 186.155 -189.205 186.485 -188.875 ;
        RECT 186.155 -190.565 186.485 -190.235 ;
        RECT 186.155 -191.925 186.485 -191.595 ;
        RECT 186.155 -193.285 186.485 -192.955 ;
        RECT 186.155 -194.645 186.485 -194.315 ;
        RECT 186.155 -196.005 186.485 -195.675 ;
        RECT 186.155 -197.365 186.485 -197.035 ;
        RECT 186.155 -198.725 186.485 -198.395 ;
        RECT 186.155 -200.085 186.485 -199.755 ;
        RECT 186.155 -201.445 186.485 -201.115 ;
        RECT 186.155 -202.805 186.485 -202.475 ;
        RECT 186.155 -204.165 186.485 -203.835 ;
        RECT 186.155 -205.525 186.485 -205.195 ;
        RECT 186.155 -206.885 186.485 -206.555 ;
        RECT 186.155 -208.245 186.485 -207.915 ;
        RECT 186.155 -209.605 186.485 -209.275 ;
        RECT 186.155 -210.965 186.485 -210.635 ;
        RECT 186.155 -212.325 186.485 -211.995 ;
        RECT 186.155 -213.685 186.485 -213.355 ;
        RECT 186.155 -215.045 186.485 -214.715 ;
        RECT 186.155 -216.405 186.485 -216.075 ;
        RECT 186.155 -217.765 186.485 -217.435 ;
        RECT 186.155 -219.125 186.485 -218.795 ;
        RECT 186.155 -220.485 186.485 -220.155 ;
        RECT 186.155 -221.845 186.485 -221.515 ;
        RECT 186.155 -223.205 186.485 -222.875 ;
        RECT 186.155 -224.565 186.485 -224.235 ;
        RECT 186.155 -225.925 186.485 -225.595 ;
        RECT 186.155 -227.285 186.485 -226.955 ;
        RECT 186.155 -228.645 186.485 -228.315 ;
        RECT 186.155 -230.005 186.485 -229.675 ;
        RECT 186.155 -231.365 186.485 -231.035 ;
        RECT 186.155 -232.725 186.485 -232.395 ;
        RECT 186.155 -234.085 186.485 -233.755 ;
        RECT 186.155 -235.445 186.485 -235.115 ;
        RECT 186.155 -236.805 186.485 -236.475 ;
        RECT 186.155 -238.165 186.485 -237.835 ;
        RECT 186.155 -243.81 186.485 -242.68 ;
        RECT 186.16 -243.925 186.48 -122.235 ;
        RECT 186.155 -122.565 186.485 -122.235 ;
        RECT 186.155 -123.925 186.485 -123.595 ;
        RECT 186.155 -125.285 186.485 -124.955 ;
        RECT 186.155 -126.645 186.485 -126.315 ;
        RECT 186.155 -128.005 186.485 -127.675 ;
        RECT 186.155 -129.365 186.485 -129.035 ;
        RECT 186.155 -130.725 186.485 -130.395 ;
        RECT 186.155 -132.085 186.485 -131.755 ;
        RECT 186.155 -133.445 186.485 -133.115 ;
        RECT 186.155 -134.805 186.485 -134.475 ;
        RECT 186.155 -136.165 186.485 -135.835 ;
        RECT 186.155 -137.525 186.485 -137.195 ;
        RECT 186.155 -138.885 186.485 -138.555 ;
        RECT 186.155 -140.245 186.485 -139.915 ;
        RECT 186.155 -141.605 186.485 -141.275 ;
        RECT 186.155 -142.965 186.485 -142.635 ;
        RECT 186.155 -144.325 186.485 -143.995 ;
        RECT 186.155 -145.685 186.485 -145.355 ;
        RECT 186.155 -147.045 186.485 -146.715 ;
        RECT 186.155 -148.405 186.485 -148.075 ;
        RECT 186.155 -149.765 186.485 -149.435 ;
        RECT 186.155 -151.125 186.485 -150.795 ;
        RECT 186.155 -152.485 186.485 -152.155 ;
        RECT 186.155 -153.845 186.485 -153.515 ;
        RECT 186.155 -155.205 186.485 -154.875 ;
        RECT 186.155 -156.565 186.485 -156.235 ;
        RECT 186.155 -157.925 186.485 -157.595 ;
        RECT 186.155 -159.285 186.485 -158.955 ;
        RECT 186.155 -160.645 186.485 -160.315 ;
        RECT 186.155 -162.005 186.485 -161.675 ;
        RECT 186.155 -163.365 186.485 -163.035 ;
        RECT 186.155 -164.725 186.485 -164.395 ;
        RECT 186.155 -166.085 186.485 -165.755 ;
        RECT 186.155 -167.445 186.485 -167.115 ;
        RECT 186.155 -168.805 186.485 -168.475 ;
        RECT 186.155 -170.165 186.485 -169.835 ;
        RECT 186.155 -171.525 186.485 -171.195 ;
        RECT 186.155 -172.885 186.485 -172.555 ;
        RECT 186.155 -174.245 186.485 -173.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 246.76 149.765 247.89 ;
        RECT 149.435 241.915 149.765 242.245 ;
        RECT 149.435 240.555 149.765 240.885 ;
        RECT 149.435 239.195 149.765 239.525 ;
        RECT 149.435 237.835 149.765 238.165 ;
        RECT 149.44 237.16 149.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 -1.525 149.765 -1.195 ;
        RECT 149.435 -2.885 149.765 -2.555 ;
        RECT 149.44 -3.56 149.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 -122.565 149.765 -122.235 ;
        RECT 149.435 -123.925 149.765 -123.595 ;
        RECT 149.435 -125.285 149.765 -124.955 ;
        RECT 149.435 -126.645 149.765 -126.315 ;
        RECT 149.435 -128.005 149.765 -127.675 ;
        RECT 149.435 -129.365 149.765 -129.035 ;
        RECT 149.435 -130.725 149.765 -130.395 ;
        RECT 149.435 -132.085 149.765 -131.755 ;
        RECT 149.435 -133.445 149.765 -133.115 ;
        RECT 149.435 -134.805 149.765 -134.475 ;
        RECT 149.435 -136.165 149.765 -135.835 ;
        RECT 149.435 -137.525 149.765 -137.195 ;
        RECT 149.435 -138.885 149.765 -138.555 ;
        RECT 149.435 -140.245 149.765 -139.915 ;
        RECT 149.435 -141.605 149.765 -141.275 ;
        RECT 149.435 -142.965 149.765 -142.635 ;
        RECT 149.435 -144.325 149.765 -143.995 ;
        RECT 149.435 -145.685 149.765 -145.355 ;
        RECT 149.435 -147.045 149.765 -146.715 ;
        RECT 149.435 -148.405 149.765 -148.075 ;
        RECT 149.435 -149.765 149.765 -149.435 ;
        RECT 149.435 -151.125 149.765 -150.795 ;
        RECT 149.435 -152.485 149.765 -152.155 ;
        RECT 149.435 -153.845 149.765 -153.515 ;
        RECT 149.435 -155.205 149.765 -154.875 ;
        RECT 149.435 -156.565 149.765 -156.235 ;
        RECT 149.435 -157.925 149.765 -157.595 ;
        RECT 149.435 -159.285 149.765 -158.955 ;
        RECT 149.435 -160.645 149.765 -160.315 ;
        RECT 149.435 -162.005 149.765 -161.675 ;
        RECT 149.435 -163.365 149.765 -163.035 ;
        RECT 149.435 -164.725 149.765 -164.395 ;
        RECT 149.435 -166.085 149.765 -165.755 ;
        RECT 149.435 -167.445 149.765 -167.115 ;
        RECT 149.435 -168.805 149.765 -168.475 ;
        RECT 149.435 -170.165 149.765 -169.835 ;
        RECT 149.435 -171.525 149.765 -171.195 ;
        RECT 149.435 -172.885 149.765 -172.555 ;
        RECT 149.435 -174.245 149.765 -173.915 ;
        RECT 149.435 -175.605 149.765 -175.275 ;
        RECT 149.435 -176.965 149.765 -176.635 ;
        RECT 149.435 -178.325 149.765 -177.995 ;
        RECT 149.435 -179.685 149.765 -179.355 ;
        RECT 149.435 -181.045 149.765 -180.715 ;
        RECT 149.435 -182.405 149.765 -182.075 ;
        RECT 149.435 -183.765 149.765 -183.435 ;
        RECT 149.435 -185.125 149.765 -184.795 ;
        RECT 149.435 -186.485 149.765 -186.155 ;
        RECT 149.435 -187.845 149.765 -187.515 ;
        RECT 149.435 -189.205 149.765 -188.875 ;
        RECT 149.435 -190.565 149.765 -190.235 ;
        RECT 149.435 -191.925 149.765 -191.595 ;
        RECT 149.435 -193.285 149.765 -192.955 ;
        RECT 149.435 -194.645 149.765 -194.315 ;
        RECT 149.435 -196.005 149.765 -195.675 ;
        RECT 149.435 -197.365 149.765 -197.035 ;
        RECT 149.435 -198.725 149.765 -198.395 ;
        RECT 149.435 -200.085 149.765 -199.755 ;
        RECT 149.435 -201.445 149.765 -201.115 ;
        RECT 149.435 -202.805 149.765 -202.475 ;
        RECT 149.435 -204.165 149.765 -203.835 ;
        RECT 149.435 -205.525 149.765 -205.195 ;
        RECT 149.435 -206.885 149.765 -206.555 ;
        RECT 149.435 -208.245 149.765 -207.915 ;
        RECT 149.435 -209.605 149.765 -209.275 ;
        RECT 149.435 -210.965 149.765 -210.635 ;
        RECT 149.435 -212.325 149.765 -211.995 ;
        RECT 149.435 -213.685 149.765 -213.355 ;
        RECT 149.435 -215.045 149.765 -214.715 ;
        RECT 149.435 -216.405 149.765 -216.075 ;
        RECT 149.435 -217.765 149.765 -217.435 ;
        RECT 149.435 -219.125 149.765 -218.795 ;
        RECT 149.435 -220.485 149.765 -220.155 ;
        RECT 149.435 -221.845 149.765 -221.515 ;
        RECT 149.435 -223.205 149.765 -222.875 ;
        RECT 149.435 -224.565 149.765 -224.235 ;
        RECT 149.435 -225.925 149.765 -225.595 ;
        RECT 149.435 -227.285 149.765 -226.955 ;
        RECT 149.435 -228.645 149.765 -228.315 ;
        RECT 149.435 -230.005 149.765 -229.675 ;
        RECT 149.435 -231.365 149.765 -231.035 ;
        RECT 149.435 -232.725 149.765 -232.395 ;
        RECT 149.435 -234.085 149.765 -233.755 ;
        RECT 149.435 -235.445 149.765 -235.115 ;
        RECT 149.435 -236.805 149.765 -236.475 ;
        RECT 149.435 -238.165 149.765 -237.835 ;
        RECT 149.435 -243.81 149.765 -242.68 ;
        RECT 149.44 -243.925 149.76 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 246.76 151.125 247.89 ;
        RECT 150.795 241.915 151.125 242.245 ;
        RECT 150.795 240.555 151.125 240.885 ;
        RECT 150.795 239.195 151.125 239.525 ;
        RECT 150.795 237.835 151.125 238.165 ;
        RECT 150.8 237.16 151.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 -1.525 151.125 -1.195 ;
        RECT 150.795 -2.885 151.125 -2.555 ;
        RECT 150.8 -3.56 151.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 -122.565 151.125 -122.235 ;
        RECT 150.795 -123.925 151.125 -123.595 ;
        RECT 150.795 -125.285 151.125 -124.955 ;
        RECT 150.795 -126.645 151.125 -126.315 ;
        RECT 150.795 -128.005 151.125 -127.675 ;
        RECT 150.795 -129.365 151.125 -129.035 ;
        RECT 150.795 -130.725 151.125 -130.395 ;
        RECT 150.795 -132.085 151.125 -131.755 ;
        RECT 150.795 -133.445 151.125 -133.115 ;
        RECT 150.795 -134.805 151.125 -134.475 ;
        RECT 150.795 -136.165 151.125 -135.835 ;
        RECT 150.795 -137.525 151.125 -137.195 ;
        RECT 150.795 -138.885 151.125 -138.555 ;
        RECT 150.795 -140.245 151.125 -139.915 ;
        RECT 150.795 -141.605 151.125 -141.275 ;
        RECT 150.795 -142.965 151.125 -142.635 ;
        RECT 150.795 -144.325 151.125 -143.995 ;
        RECT 150.795 -145.685 151.125 -145.355 ;
        RECT 150.795 -147.045 151.125 -146.715 ;
        RECT 150.795 -148.405 151.125 -148.075 ;
        RECT 150.795 -149.765 151.125 -149.435 ;
        RECT 150.795 -151.125 151.125 -150.795 ;
        RECT 150.795 -152.485 151.125 -152.155 ;
        RECT 150.795 -153.845 151.125 -153.515 ;
        RECT 150.795 -155.205 151.125 -154.875 ;
        RECT 150.795 -156.565 151.125 -156.235 ;
        RECT 150.795 -157.925 151.125 -157.595 ;
        RECT 150.795 -159.285 151.125 -158.955 ;
        RECT 150.795 -160.645 151.125 -160.315 ;
        RECT 150.795 -162.005 151.125 -161.675 ;
        RECT 150.795 -163.365 151.125 -163.035 ;
        RECT 150.795 -164.725 151.125 -164.395 ;
        RECT 150.795 -166.085 151.125 -165.755 ;
        RECT 150.795 -167.445 151.125 -167.115 ;
        RECT 150.795 -168.805 151.125 -168.475 ;
        RECT 150.795 -170.165 151.125 -169.835 ;
        RECT 150.795 -171.525 151.125 -171.195 ;
        RECT 150.795 -172.885 151.125 -172.555 ;
        RECT 150.795 -174.245 151.125 -173.915 ;
        RECT 150.795 -175.605 151.125 -175.275 ;
        RECT 150.795 -176.965 151.125 -176.635 ;
        RECT 150.795 -178.325 151.125 -177.995 ;
        RECT 150.795 -179.685 151.125 -179.355 ;
        RECT 150.795 -181.045 151.125 -180.715 ;
        RECT 150.795 -182.405 151.125 -182.075 ;
        RECT 150.795 -183.765 151.125 -183.435 ;
        RECT 150.795 -185.125 151.125 -184.795 ;
        RECT 150.795 -186.485 151.125 -186.155 ;
        RECT 150.795 -187.845 151.125 -187.515 ;
        RECT 150.795 -189.205 151.125 -188.875 ;
        RECT 150.795 -190.565 151.125 -190.235 ;
        RECT 150.795 -191.925 151.125 -191.595 ;
        RECT 150.795 -193.285 151.125 -192.955 ;
        RECT 150.795 -194.645 151.125 -194.315 ;
        RECT 150.795 -196.005 151.125 -195.675 ;
        RECT 150.795 -197.365 151.125 -197.035 ;
        RECT 150.795 -198.725 151.125 -198.395 ;
        RECT 150.795 -200.085 151.125 -199.755 ;
        RECT 150.795 -201.445 151.125 -201.115 ;
        RECT 150.795 -202.805 151.125 -202.475 ;
        RECT 150.795 -204.165 151.125 -203.835 ;
        RECT 150.795 -205.525 151.125 -205.195 ;
        RECT 150.795 -206.885 151.125 -206.555 ;
        RECT 150.795 -208.245 151.125 -207.915 ;
        RECT 150.795 -209.605 151.125 -209.275 ;
        RECT 150.795 -210.965 151.125 -210.635 ;
        RECT 150.795 -212.325 151.125 -211.995 ;
        RECT 150.795 -213.685 151.125 -213.355 ;
        RECT 150.795 -215.045 151.125 -214.715 ;
        RECT 150.795 -216.405 151.125 -216.075 ;
        RECT 150.795 -217.765 151.125 -217.435 ;
        RECT 150.795 -219.125 151.125 -218.795 ;
        RECT 150.795 -220.485 151.125 -220.155 ;
        RECT 150.795 -221.845 151.125 -221.515 ;
        RECT 150.795 -223.205 151.125 -222.875 ;
        RECT 150.795 -224.565 151.125 -224.235 ;
        RECT 150.795 -225.925 151.125 -225.595 ;
        RECT 150.795 -227.285 151.125 -226.955 ;
        RECT 150.795 -228.645 151.125 -228.315 ;
        RECT 150.795 -230.005 151.125 -229.675 ;
        RECT 150.795 -231.365 151.125 -231.035 ;
        RECT 150.795 -232.725 151.125 -232.395 ;
        RECT 150.795 -234.085 151.125 -233.755 ;
        RECT 150.795 -235.445 151.125 -235.115 ;
        RECT 150.795 -236.805 151.125 -236.475 ;
        RECT 150.795 -238.165 151.125 -237.835 ;
        RECT 150.795 -243.81 151.125 -242.68 ;
        RECT 150.8 -243.925 151.12 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 246.76 152.485 247.89 ;
        RECT 152.155 241.915 152.485 242.245 ;
        RECT 152.155 240.555 152.485 240.885 ;
        RECT 152.155 239.195 152.485 239.525 ;
        RECT 152.155 237.835 152.485 238.165 ;
        RECT 152.16 237.16 152.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 -1.525 152.485 -1.195 ;
        RECT 152.155 -2.885 152.485 -2.555 ;
        RECT 152.16 -3.56 152.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 -122.565 152.485 -122.235 ;
        RECT 152.155 -123.925 152.485 -123.595 ;
        RECT 152.155 -125.285 152.485 -124.955 ;
        RECT 152.155 -126.645 152.485 -126.315 ;
        RECT 152.155 -128.005 152.485 -127.675 ;
        RECT 152.155 -129.365 152.485 -129.035 ;
        RECT 152.155 -130.725 152.485 -130.395 ;
        RECT 152.155 -132.085 152.485 -131.755 ;
        RECT 152.155 -133.445 152.485 -133.115 ;
        RECT 152.155 -134.805 152.485 -134.475 ;
        RECT 152.155 -136.165 152.485 -135.835 ;
        RECT 152.155 -137.525 152.485 -137.195 ;
        RECT 152.155 -138.885 152.485 -138.555 ;
        RECT 152.155 -140.245 152.485 -139.915 ;
        RECT 152.155 -141.605 152.485 -141.275 ;
        RECT 152.155 -142.965 152.485 -142.635 ;
        RECT 152.155 -144.325 152.485 -143.995 ;
        RECT 152.155 -145.685 152.485 -145.355 ;
        RECT 152.155 -147.045 152.485 -146.715 ;
        RECT 152.155 -148.405 152.485 -148.075 ;
        RECT 152.155 -149.765 152.485 -149.435 ;
        RECT 152.155 -151.125 152.485 -150.795 ;
        RECT 152.155 -152.485 152.485 -152.155 ;
        RECT 152.155 -153.845 152.485 -153.515 ;
        RECT 152.155 -155.205 152.485 -154.875 ;
        RECT 152.155 -156.565 152.485 -156.235 ;
        RECT 152.155 -157.925 152.485 -157.595 ;
        RECT 152.155 -159.285 152.485 -158.955 ;
        RECT 152.155 -160.645 152.485 -160.315 ;
        RECT 152.155 -162.005 152.485 -161.675 ;
        RECT 152.155 -163.365 152.485 -163.035 ;
        RECT 152.155 -164.725 152.485 -164.395 ;
        RECT 152.155 -166.085 152.485 -165.755 ;
        RECT 152.155 -167.445 152.485 -167.115 ;
        RECT 152.155 -168.805 152.485 -168.475 ;
        RECT 152.155 -170.165 152.485 -169.835 ;
        RECT 152.155 -171.525 152.485 -171.195 ;
        RECT 152.155 -172.885 152.485 -172.555 ;
        RECT 152.155 -174.245 152.485 -173.915 ;
        RECT 152.155 -175.605 152.485 -175.275 ;
        RECT 152.155 -176.965 152.485 -176.635 ;
        RECT 152.155 -178.325 152.485 -177.995 ;
        RECT 152.155 -179.685 152.485 -179.355 ;
        RECT 152.155 -181.045 152.485 -180.715 ;
        RECT 152.155 -182.405 152.485 -182.075 ;
        RECT 152.155 -183.765 152.485 -183.435 ;
        RECT 152.155 -185.125 152.485 -184.795 ;
        RECT 152.155 -186.485 152.485 -186.155 ;
        RECT 152.155 -187.845 152.485 -187.515 ;
        RECT 152.155 -189.205 152.485 -188.875 ;
        RECT 152.155 -190.565 152.485 -190.235 ;
        RECT 152.155 -191.925 152.485 -191.595 ;
        RECT 152.155 -193.285 152.485 -192.955 ;
        RECT 152.155 -194.645 152.485 -194.315 ;
        RECT 152.155 -196.005 152.485 -195.675 ;
        RECT 152.155 -197.365 152.485 -197.035 ;
        RECT 152.155 -198.725 152.485 -198.395 ;
        RECT 152.155 -200.085 152.485 -199.755 ;
        RECT 152.155 -201.445 152.485 -201.115 ;
        RECT 152.155 -202.805 152.485 -202.475 ;
        RECT 152.155 -204.165 152.485 -203.835 ;
        RECT 152.155 -205.525 152.485 -205.195 ;
        RECT 152.155 -206.885 152.485 -206.555 ;
        RECT 152.155 -208.245 152.485 -207.915 ;
        RECT 152.155 -209.605 152.485 -209.275 ;
        RECT 152.155 -210.965 152.485 -210.635 ;
        RECT 152.155 -212.325 152.485 -211.995 ;
        RECT 152.155 -213.685 152.485 -213.355 ;
        RECT 152.155 -215.045 152.485 -214.715 ;
        RECT 152.155 -216.405 152.485 -216.075 ;
        RECT 152.155 -217.765 152.485 -217.435 ;
        RECT 152.155 -219.125 152.485 -218.795 ;
        RECT 152.155 -220.485 152.485 -220.155 ;
        RECT 152.155 -221.845 152.485 -221.515 ;
        RECT 152.155 -223.205 152.485 -222.875 ;
        RECT 152.155 -224.565 152.485 -224.235 ;
        RECT 152.155 -225.925 152.485 -225.595 ;
        RECT 152.155 -227.285 152.485 -226.955 ;
        RECT 152.155 -228.645 152.485 -228.315 ;
        RECT 152.155 -230.005 152.485 -229.675 ;
        RECT 152.155 -231.365 152.485 -231.035 ;
        RECT 152.155 -232.725 152.485 -232.395 ;
        RECT 152.155 -234.085 152.485 -233.755 ;
        RECT 152.155 -235.445 152.485 -235.115 ;
        RECT 152.155 -236.805 152.485 -236.475 ;
        RECT 152.155 -238.165 152.485 -237.835 ;
        RECT 152.155 -243.81 152.485 -242.68 ;
        RECT 152.16 -243.925 152.48 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 246.76 153.845 247.89 ;
        RECT 153.515 241.915 153.845 242.245 ;
        RECT 153.515 240.555 153.845 240.885 ;
        RECT 153.515 239.195 153.845 239.525 ;
        RECT 153.515 237.835 153.845 238.165 ;
        RECT 153.52 237.16 153.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 -1.525 153.845 -1.195 ;
        RECT 153.515 -2.885 153.845 -2.555 ;
        RECT 153.52 -3.56 153.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 -122.565 153.845 -122.235 ;
        RECT 153.515 -123.925 153.845 -123.595 ;
        RECT 153.515 -125.285 153.845 -124.955 ;
        RECT 153.515 -126.645 153.845 -126.315 ;
        RECT 153.515 -128.005 153.845 -127.675 ;
        RECT 153.515 -129.365 153.845 -129.035 ;
        RECT 153.515 -130.725 153.845 -130.395 ;
        RECT 153.515 -132.085 153.845 -131.755 ;
        RECT 153.515 -133.445 153.845 -133.115 ;
        RECT 153.515 -134.805 153.845 -134.475 ;
        RECT 153.515 -136.165 153.845 -135.835 ;
        RECT 153.515 -137.525 153.845 -137.195 ;
        RECT 153.515 -138.885 153.845 -138.555 ;
        RECT 153.515 -140.245 153.845 -139.915 ;
        RECT 153.515 -141.605 153.845 -141.275 ;
        RECT 153.515 -142.965 153.845 -142.635 ;
        RECT 153.515 -144.325 153.845 -143.995 ;
        RECT 153.515 -145.685 153.845 -145.355 ;
        RECT 153.515 -147.045 153.845 -146.715 ;
        RECT 153.515 -148.405 153.845 -148.075 ;
        RECT 153.515 -149.765 153.845 -149.435 ;
        RECT 153.515 -151.125 153.845 -150.795 ;
        RECT 153.515 -152.485 153.845 -152.155 ;
        RECT 153.515 -153.845 153.845 -153.515 ;
        RECT 153.515 -155.205 153.845 -154.875 ;
        RECT 153.515 -156.565 153.845 -156.235 ;
        RECT 153.515 -157.925 153.845 -157.595 ;
        RECT 153.515 -159.285 153.845 -158.955 ;
        RECT 153.515 -160.645 153.845 -160.315 ;
        RECT 153.515 -162.005 153.845 -161.675 ;
        RECT 153.515 -163.365 153.845 -163.035 ;
        RECT 153.515 -164.725 153.845 -164.395 ;
        RECT 153.515 -166.085 153.845 -165.755 ;
        RECT 153.515 -167.445 153.845 -167.115 ;
        RECT 153.515 -168.805 153.845 -168.475 ;
        RECT 153.515 -170.165 153.845 -169.835 ;
        RECT 153.515 -171.525 153.845 -171.195 ;
        RECT 153.515 -172.885 153.845 -172.555 ;
        RECT 153.515 -174.245 153.845 -173.915 ;
        RECT 153.515 -175.605 153.845 -175.275 ;
        RECT 153.515 -176.965 153.845 -176.635 ;
        RECT 153.515 -178.325 153.845 -177.995 ;
        RECT 153.515 -179.685 153.845 -179.355 ;
        RECT 153.515 -181.045 153.845 -180.715 ;
        RECT 153.515 -182.405 153.845 -182.075 ;
        RECT 153.515 -183.765 153.845 -183.435 ;
        RECT 153.515 -185.125 153.845 -184.795 ;
        RECT 153.515 -186.485 153.845 -186.155 ;
        RECT 153.515 -187.845 153.845 -187.515 ;
        RECT 153.515 -189.205 153.845 -188.875 ;
        RECT 153.515 -190.565 153.845 -190.235 ;
        RECT 153.515 -191.925 153.845 -191.595 ;
        RECT 153.515 -193.285 153.845 -192.955 ;
        RECT 153.515 -194.645 153.845 -194.315 ;
        RECT 153.515 -196.005 153.845 -195.675 ;
        RECT 153.515 -197.365 153.845 -197.035 ;
        RECT 153.515 -198.725 153.845 -198.395 ;
        RECT 153.515 -200.085 153.845 -199.755 ;
        RECT 153.515 -201.445 153.845 -201.115 ;
        RECT 153.515 -202.805 153.845 -202.475 ;
        RECT 153.515 -204.165 153.845 -203.835 ;
        RECT 153.515 -205.525 153.845 -205.195 ;
        RECT 153.515 -206.885 153.845 -206.555 ;
        RECT 153.515 -208.245 153.845 -207.915 ;
        RECT 153.515 -209.605 153.845 -209.275 ;
        RECT 153.515 -210.965 153.845 -210.635 ;
        RECT 153.515 -212.325 153.845 -211.995 ;
        RECT 153.515 -213.685 153.845 -213.355 ;
        RECT 153.515 -215.045 153.845 -214.715 ;
        RECT 153.515 -216.405 153.845 -216.075 ;
        RECT 153.515 -217.765 153.845 -217.435 ;
        RECT 153.515 -219.125 153.845 -218.795 ;
        RECT 153.515 -220.485 153.845 -220.155 ;
        RECT 153.515 -221.845 153.845 -221.515 ;
        RECT 153.515 -223.205 153.845 -222.875 ;
        RECT 153.515 -224.565 153.845 -224.235 ;
        RECT 153.515 -225.925 153.845 -225.595 ;
        RECT 153.515 -227.285 153.845 -226.955 ;
        RECT 153.515 -228.645 153.845 -228.315 ;
        RECT 153.515 -230.005 153.845 -229.675 ;
        RECT 153.515 -231.365 153.845 -231.035 ;
        RECT 153.515 -232.725 153.845 -232.395 ;
        RECT 153.515 -234.085 153.845 -233.755 ;
        RECT 153.515 -235.445 153.845 -235.115 ;
        RECT 153.515 -236.805 153.845 -236.475 ;
        RECT 153.515 -238.165 153.845 -237.835 ;
        RECT 153.515 -243.81 153.845 -242.68 ;
        RECT 153.52 -243.925 153.84 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 246.76 155.205 247.89 ;
        RECT 154.875 241.915 155.205 242.245 ;
        RECT 154.875 240.555 155.205 240.885 ;
        RECT 154.875 239.195 155.205 239.525 ;
        RECT 154.875 237.835 155.205 238.165 ;
        RECT 154.88 237.16 155.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 -126.645 155.205 -126.315 ;
        RECT 154.875 -128.005 155.205 -127.675 ;
        RECT 154.875 -129.365 155.205 -129.035 ;
        RECT 154.875 -130.725 155.205 -130.395 ;
        RECT 154.875 -132.085 155.205 -131.755 ;
        RECT 154.875 -133.445 155.205 -133.115 ;
        RECT 154.875 -134.805 155.205 -134.475 ;
        RECT 154.875 -136.165 155.205 -135.835 ;
        RECT 154.875 -137.525 155.205 -137.195 ;
        RECT 154.875 -138.885 155.205 -138.555 ;
        RECT 154.875 -140.245 155.205 -139.915 ;
        RECT 154.875 -141.605 155.205 -141.275 ;
        RECT 154.875 -142.965 155.205 -142.635 ;
        RECT 154.875 -144.325 155.205 -143.995 ;
        RECT 154.875 -145.685 155.205 -145.355 ;
        RECT 154.875 -147.045 155.205 -146.715 ;
        RECT 154.875 -148.405 155.205 -148.075 ;
        RECT 154.875 -149.765 155.205 -149.435 ;
        RECT 154.875 -151.125 155.205 -150.795 ;
        RECT 154.875 -152.485 155.205 -152.155 ;
        RECT 154.875 -153.845 155.205 -153.515 ;
        RECT 154.875 -155.205 155.205 -154.875 ;
        RECT 154.875 -156.565 155.205 -156.235 ;
        RECT 154.875 -157.925 155.205 -157.595 ;
        RECT 154.875 -159.285 155.205 -158.955 ;
        RECT 154.875 -160.645 155.205 -160.315 ;
        RECT 154.875 -162.005 155.205 -161.675 ;
        RECT 154.875 -163.365 155.205 -163.035 ;
        RECT 154.875 -164.725 155.205 -164.395 ;
        RECT 154.875 -166.085 155.205 -165.755 ;
        RECT 154.875 -167.445 155.205 -167.115 ;
        RECT 154.875 -168.805 155.205 -168.475 ;
        RECT 154.875 -170.165 155.205 -169.835 ;
        RECT 154.875 -171.525 155.205 -171.195 ;
        RECT 154.875 -172.885 155.205 -172.555 ;
        RECT 154.875 -174.245 155.205 -173.915 ;
        RECT 154.875 -175.605 155.205 -175.275 ;
        RECT 154.875 -176.965 155.205 -176.635 ;
        RECT 154.875 -178.325 155.205 -177.995 ;
        RECT 154.875 -179.685 155.205 -179.355 ;
        RECT 154.875 -181.045 155.205 -180.715 ;
        RECT 154.875 -182.405 155.205 -182.075 ;
        RECT 154.875 -183.765 155.205 -183.435 ;
        RECT 154.875 -185.125 155.205 -184.795 ;
        RECT 154.875 -186.485 155.205 -186.155 ;
        RECT 154.875 -187.845 155.205 -187.515 ;
        RECT 154.875 -189.205 155.205 -188.875 ;
        RECT 154.875 -190.565 155.205 -190.235 ;
        RECT 154.875 -191.925 155.205 -191.595 ;
        RECT 154.875 -193.285 155.205 -192.955 ;
        RECT 154.875 -194.645 155.205 -194.315 ;
        RECT 154.875 -196.005 155.205 -195.675 ;
        RECT 154.875 -197.365 155.205 -197.035 ;
        RECT 154.875 -198.725 155.205 -198.395 ;
        RECT 154.875 -200.085 155.205 -199.755 ;
        RECT 154.875 -201.445 155.205 -201.115 ;
        RECT 154.875 -202.805 155.205 -202.475 ;
        RECT 154.875 -204.165 155.205 -203.835 ;
        RECT 154.875 -205.525 155.205 -205.195 ;
        RECT 154.875 -206.885 155.205 -206.555 ;
        RECT 154.875 -208.245 155.205 -207.915 ;
        RECT 154.875 -209.605 155.205 -209.275 ;
        RECT 154.875 -210.965 155.205 -210.635 ;
        RECT 154.875 -212.325 155.205 -211.995 ;
        RECT 154.875 -213.685 155.205 -213.355 ;
        RECT 154.875 -215.045 155.205 -214.715 ;
        RECT 154.875 -216.405 155.205 -216.075 ;
        RECT 154.875 -217.765 155.205 -217.435 ;
        RECT 154.875 -219.125 155.205 -218.795 ;
        RECT 154.875 -220.485 155.205 -220.155 ;
        RECT 154.875 -221.845 155.205 -221.515 ;
        RECT 154.875 -223.205 155.205 -222.875 ;
        RECT 154.875 -224.565 155.205 -224.235 ;
        RECT 154.875 -225.925 155.205 -225.595 ;
        RECT 154.875 -227.285 155.205 -226.955 ;
        RECT 154.875 -228.645 155.205 -228.315 ;
        RECT 154.875 -230.005 155.205 -229.675 ;
        RECT 154.875 -231.365 155.205 -231.035 ;
        RECT 154.875 -232.725 155.205 -232.395 ;
        RECT 154.875 -234.085 155.205 -233.755 ;
        RECT 154.875 -235.445 155.205 -235.115 ;
        RECT 154.875 -236.805 155.205 -236.475 ;
        RECT 154.875 -238.165 155.205 -237.835 ;
        RECT 154.875 -243.81 155.205 -242.68 ;
        RECT 154.88 -243.925 155.2 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.26 -125.535 155.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.235 246.76 156.565 247.89 ;
        RECT 156.235 241.915 156.565 242.245 ;
        RECT 156.235 240.555 156.565 240.885 ;
        RECT 156.235 239.195 156.565 239.525 ;
        RECT 156.235 237.835 156.565 238.165 ;
        RECT 156.24 237.16 156.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 246.76 157.925 247.89 ;
        RECT 157.595 241.915 157.925 242.245 ;
        RECT 157.595 240.555 157.925 240.885 ;
        RECT 157.595 239.195 157.925 239.525 ;
        RECT 157.595 237.835 157.925 238.165 ;
        RECT 157.6 237.16 157.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 -1.525 157.925 -1.195 ;
        RECT 157.595 -2.885 157.925 -2.555 ;
        RECT 157.6 -3.56 157.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 246.76 159.285 247.89 ;
        RECT 158.955 241.915 159.285 242.245 ;
        RECT 158.955 240.555 159.285 240.885 ;
        RECT 158.955 239.195 159.285 239.525 ;
        RECT 158.955 237.835 159.285 238.165 ;
        RECT 158.96 237.16 159.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -1.525 159.285 -1.195 ;
        RECT 158.955 -2.885 159.285 -2.555 ;
        RECT 158.96 -3.56 159.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -122.565 159.285 -122.235 ;
        RECT 158.955 -123.925 159.285 -123.595 ;
        RECT 158.955 -125.285 159.285 -124.955 ;
        RECT 158.955 -126.645 159.285 -126.315 ;
        RECT 158.955 -128.005 159.285 -127.675 ;
        RECT 158.955 -129.365 159.285 -129.035 ;
        RECT 158.955 -130.725 159.285 -130.395 ;
        RECT 158.955 -132.085 159.285 -131.755 ;
        RECT 158.955 -133.445 159.285 -133.115 ;
        RECT 158.955 -134.805 159.285 -134.475 ;
        RECT 158.955 -136.165 159.285 -135.835 ;
        RECT 158.955 -137.525 159.285 -137.195 ;
        RECT 158.955 -138.885 159.285 -138.555 ;
        RECT 158.955 -140.245 159.285 -139.915 ;
        RECT 158.955 -141.605 159.285 -141.275 ;
        RECT 158.955 -142.965 159.285 -142.635 ;
        RECT 158.955 -144.325 159.285 -143.995 ;
        RECT 158.955 -145.685 159.285 -145.355 ;
        RECT 158.955 -147.045 159.285 -146.715 ;
        RECT 158.955 -148.405 159.285 -148.075 ;
        RECT 158.955 -149.765 159.285 -149.435 ;
        RECT 158.955 -151.125 159.285 -150.795 ;
        RECT 158.955 -152.485 159.285 -152.155 ;
        RECT 158.955 -153.845 159.285 -153.515 ;
        RECT 158.955 -155.205 159.285 -154.875 ;
        RECT 158.955 -156.565 159.285 -156.235 ;
        RECT 158.955 -157.925 159.285 -157.595 ;
        RECT 158.955 -159.285 159.285 -158.955 ;
        RECT 158.955 -160.645 159.285 -160.315 ;
        RECT 158.955 -162.005 159.285 -161.675 ;
        RECT 158.955 -163.365 159.285 -163.035 ;
        RECT 158.955 -164.725 159.285 -164.395 ;
        RECT 158.955 -166.085 159.285 -165.755 ;
        RECT 158.955 -167.445 159.285 -167.115 ;
        RECT 158.955 -168.805 159.285 -168.475 ;
        RECT 158.955 -170.165 159.285 -169.835 ;
        RECT 158.955 -171.525 159.285 -171.195 ;
        RECT 158.955 -172.885 159.285 -172.555 ;
        RECT 158.955 -174.245 159.285 -173.915 ;
        RECT 158.955 -175.605 159.285 -175.275 ;
        RECT 158.955 -176.965 159.285 -176.635 ;
        RECT 158.955 -178.325 159.285 -177.995 ;
        RECT 158.955 -179.685 159.285 -179.355 ;
        RECT 158.955 -181.045 159.285 -180.715 ;
        RECT 158.955 -182.405 159.285 -182.075 ;
        RECT 158.955 -183.765 159.285 -183.435 ;
        RECT 158.955 -185.125 159.285 -184.795 ;
        RECT 158.955 -186.485 159.285 -186.155 ;
        RECT 158.955 -187.845 159.285 -187.515 ;
        RECT 158.955 -189.205 159.285 -188.875 ;
        RECT 158.955 -190.565 159.285 -190.235 ;
        RECT 158.955 -191.925 159.285 -191.595 ;
        RECT 158.955 -193.285 159.285 -192.955 ;
        RECT 158.955 -194.645 159.285 -194.315 ;
        RECT 158.955 -196.005 159.285 -195.675 ;
        RECT 158.955 -197.365 159.285 -197.035 ;
        RECT 158.955 -198.725 159.285 -198.395 ;
        RECT 158.955 -200.085 159.285 -199.755 ;
        RECT 158.955 -201.445 159.285 -201.115 ;
        RECT 158.955 -202.805 159.285 -202.475 ;
        RECT 158.955 -204.165 159.285 -203.835 ;
        RECT 158.955 -205.525 159.285 -205.195 ;
        RECT 158.955 -206.885 159.285 -206.555 ;
        RECT 158.955 -208.245 159.285 -207.915 ;
        RECT 158.955 -209.605 159.285 -209.275 ;
        RECT 158.955 -210.965 159.285 -210.635 ;
        RECT 158.955 -212.325 159.285 -211.995 ;
        RECT 158.955 -213.685 159.285 -213.355 ;
        RECT 158.955 -215.045 159.285 -214.715 ;
        RECT 158.955 -216.405 159.285 -216.075 ;
        RECT 158.955 -217.765 159.285 -217.435 ;
        RECT 158.955 -219.125 159.285 -218.795 ;
        RECT 158.955 -220.485 159.285 -220.155 ;
        RECT 158.955 -221.845 159.285 -221.515 ;
        RECT 158.955 -223.205 159.285 -222.875 ;
        RECT 158.955 -224.565 159.285 -224.235 ;
        RECT 158.955 -225.925 159.285 -225.595 ;
        RECT 158.955 -227.285 159.285 -226.955 ;
        RECT 158.955 -228.645 159.285 -228.315 ;
        RECT 158.955 -230.005 159.285 -229.675 ;
        RECT 158.955 -231.365 159.285 -231.035 ;
        RECT 158.955 -232.725 159.285 -232.395 ;
        RECT 158.955 -234.085 159.285 -233.755 ;
        RECT 158.955 -235.445 159.285 -235.115 ;
        RECT 158.955 -236.805 159.285 -236.475 ;
        RECT 158.955 -238.165 159.285 -237.835 ;
        RECT 158.955 -243.81 159.285 -242.68 ;
        RECT 158.96 -243.925 159.28 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 246.76 160.645 247.89 ;
        RECT 160.315 241.915 160.645 242.245 ;
        RECT 160.315 240.555 160.645 240.885 ;
        RECT 160.315 239.195 160.645 239.525 ;
        RECT 160.315 237.835 160.645 238.165 ;
        RECT 160.32 237.16 160.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -1.525 160.645 -1.195 ;
        RECT 160.315 -2.885 160.645 -2.555 ;
        RECT 160.32 -3.56 160.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -122.565 160.645 -122.235 ;
        RECT 160.315 -123.925 160.645 -123.595 ;
        RECT 160.315 -125.285 160.645 -124.955 ;
        RECT 160.315 -126.645 160.645 -126.315 ;
        RECT 160.315 -128.005 160.645 -127.675 ;
        RECT 160.315 -129.365 160.645 -129.035 ;
        RECT 160.315 -130.725 160.645 -130.395 ;
        RECT 160.315 -132.085 160.645 -131.755 ;
        RECT 160.315 -133.445 160.645 -133.115 ;
        RECT 160.315 -134.805 160.645 -134.475 ;
        RECT 160.315 -136.165 160.645 -135.835 ;
        RECT 160.315 -137.525 160.645 -137.195 ;
        RECT 160.315 -138.885 160.645 -138.555 ;
        RECT 160.315 -140.245 160.645 -139.915 ;
        RECT 160.315 -141.605 160.645 -141.275 ;
        RECT 160.315 -142.965 160.645 -142.635 ;
        RECT 160.315 -144.325 160.645 -143.995 ;
        RECT 160.315 -145.685 160.645 -145.355 ;
        RECT 160.315 -147.045 160.645 -146.715 ;
        RECT 160.315 -148.405 160.645 -148.075 ;
        RECT 160.315 -149.765 160.645 -149.435 ;
        RECT 160.315 -151.125 160.645 -150.795 ;
        RECT 160.315 -152.485 160.645 -152.155 ;
        RECT 160.315 -153.845 160.645 -153.515 ;
        RECT 160.315 -155.205 160.645 -154.875 ;
        RECT 160.315 -156.565 160.645 -156.235 ;
        RECT 160.315 -157.925 160.645 -157.595 ;
        RECT 160.315 -159.285 160.645 -158.955 ;
        RECT 160.315 -160.645 160.645 -160.315 ;
        RECT 160.315 -162.005 160.645 -161.675 ;
        RECT 160.315 -163.365 160.645 -163.035 ;
        RECT 160.315 -164.725 160.645 -164.395 ;
        RECT 160.315 -166.085 160.645 -165.755 ;
        RECT 160.315 -167.445 160.645 -167.115 ;
        RECT 160.315 -168.805 160.645 -168.475 ;
        RECT 160.315 -170.165 160.645 -169.835 ;
        RECT 160.315 -171.525 160.645 -171.195 ;
        RECT 160.315 -172.885 160.645 -172.555 ;
        RECT 160.315 -174.245 160.645 -173.915 ;
        RECT 160.315 -175.605 160.645 -175.275 ;
        RECT 160.315 -176.965 160.645 -176.635 ;
        RECT 160.315 -178.325 160.645 -177.995 ;
        RECT 160.315 -179.685 160.645 -179.355 ;
        RECT 160.315 -181.045 160.645 -180.715 ;
        RECT 160.315 -182.405 160.645 -182.075 ;
        RECT 160.315 -183.765 160.645 -183.435 ;
        RECT 160.315 -185.125 160.645 -184.795 ;
        RECT 160.315 -186.485 160.645 -186.155 ;
        RECT 160.315 -187.845 160.645 -187.515 ;
        RECT 160.315 -189.205 160.645 -188.875 ;
        RECT 160.315 -190.565 160.645 -190.235 ;
        RECT 160.315 -191.925 160.645 -191.595 ;
        RECT 160.315 -193.285 160.645 -192.955 ;
        RECT 160.315 -194.645 160.645 -194.315 ;
        RECT 160.315 -196.005 160.645 -195.675 ;
        RECT 160.315 -197.365 160.645 -197.035 ;
        RECT 160.315 -198.725 160.645 -198.395 ;
        RECT 160.315 -200.085 160.645 -199.755 ;
        RECT 160.315 -201.445 160.645 -201.115 ;
        RECT 160.315 -202.805 160.645 -202.475 ;
        RECT 160.315 -204.165 160.645 -203.835 ;
        RECT 160.315 -205.525 160.645 -205.195 ;
        RECT 160.315 -206.885 160.645 -206.555 ;
        RECT 160.315 -208.245 160.645 -207.915 ;
        RECT 160.315 -209.605 160.645 -209.275 ;
        RECT 160.315 -210.965 160.645 -210.635 ;
        RECT 160.315 -212.325 160.645 -211.995 ;
        RECT 160.315 -213.685 160.645 -213.355 ;
        RECT 160.315 -215.045 160.645 -214.715 ;
        RECT 160.315 -216.405 160.645 -216.075 ;
        RECT 160.315 -217.765 160.645 -217.435 ;
        RECT 160.315 -219.125 160.645 -218.795 ;
        RECT 160.315 -220.485 160.645 -220.155 ;
        RECT 160.315 -221.845 160.645 -221.515 ;
        RECT 160.315 -223.205 160.645 -222.875 ;
        RECT 160.315 -224.565 160.645 -224.235 ;
        RECT 160.315 -225.925 160.645 -225.595 ;
        RECT 160.315 -227.285 160.645 -226.955 ;
        RECT 160.315 -228.645 160.645 -228.315 ;
        RECT 160.315 -230.005 160.645 -229.675 ;
        RECT 160.315 -231.365 160.645 -231.035 ;
        RECT 160.315 -232.725 160.645 -232.395 ;
        RECT 160.315 -234.085 160.645 -233.755 ;
        RECT 160.315 -235.445 160.645 -235.115 ;
        RECT 160.315 -236.805 160.645 -236.475 ;
        RECT 160.315 -238.165 160.645 -237.835 ;
        RECT 160.315 -243.81 160.645 -242.68 ;
        RECT 160.32 -243.925 160.64 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 246.76 162.005 247.89 ;
        RECT 161.675 241.915 162.005 242.245 ;
        RECT 161.675 240.555 162.005 240.885 ;
        RECT 161.675 239.195 162.005 239.525 ;
        RECT 161.675 237.835 162.005 238.165 ;
        RECT 161.68 237.16 162 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 -1.525 162.005 -1.195 ;
        RECT 161.675 -2.885 162.005 -2.555 ;
        RECT 161.68 -3.56 162 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 -122.565 162.005 -122.235 ;
        RECT 161.675 -123.925 162.005 -123.595 ;
        RECT 161.675 -125.285 162.005 -124.955 ;
        RECT 161.675 -126.645 162.005 -126.315 ;
        RECT 161.675 -128.005 162.005 -127.675 ;
        RECT 161.675 -129.365 162.005 -129.035 ;
        RECT 161.675 -130.725 162.005 -130.395 ;
        RECT 161.675 -132.085 162.005 -131.755 ;
        RECT 161.675 -133.445 162.005 -133.115 ;
        RECT 161.675 -134.805 162.005 -134.475 ;
        RECT 161.675 -136.165 162.005 -135.835 ;
        RECT 161.675 -137.525 162.005 -137.195 ;
        RECT 161.675 -138.885 162.005 -138.555 ;
        RECT 161.675 -140.245 162.005 -139.915 ;
        RECT 161.675 -141.605 162.005 -141.275 ;
        RECT 161.675 -142.965 162.005 -142.635 ;
        RECT 161.675 -144.325 162.005 -143.995 ;
        RECT 161.675 -145.685 162.005 -145.355 ;
        RECT 161.675 -147.045 162.005 -146.715 ;
        RECT 161.675 -148.405 162.005 -148.075 ;
        RECT 161.675 -149.765 162.005 -149.435 ;
        RECT 161.675 -151.125 162.005 -150.795 ;
        RECT 161.675 -152.485 162.005 -152.155 ;
        RECT 161.675 -153.845 162.005 -153.515 ;
        RECT 161.675 -155.205 162.005 -154.875 ;
        RECT 161.675 -156.565 162.005 -156.235 ;
        RECT 161.675 -157.925 162.005 -157.595 ;
        RECT 161.675 -159.285 162.005 -158.955 ;
        RECT 161.675 -160.645 162.005 -160.315 ;
        RECT 161.675 -162.005 162.005 -161.675 ;
        RECT 161.675 -163.365 162.005 -163.035 ;
        RECT 161.675 -164.725 162.005 -164.395 ;
        RECT 161.675 -166.085 162.005 -165.755 ;
        RECT 161.675 -167.445 162.005 -167.115 ;
        RECT 161.675 -168.805 162.005 -168.475 ;
        RECT 161.675 -170.165 162.005 -169.835 ;
        RECT 161.675 -171.525 162.005 -171.195 ;
        RECT 161.675 -172.885 162.005 -172.555 ;
        RECT 161.675 -174.245 162.005 -173.915 ;
        RECT 161.675 -175.605 162.005 -175.275 ;
        RECT 161.675 -176.965 162.005 -176.635 ;
        RECT 161.675 -178.325 162.005 -177.995 ;
        RECT 161.675 -179.685 162.005 -179.355 ;
        RECT 161.675 -181.045 162.005 -180.715 ;
        RECT 161.675 -182.405 162.005 -182.075 ;
        RECT 161.675 -183.765 162.005 -183.435 ;
        RECT 161.675 -185.125 162.005 -184.795 ;
        RECT 161.675 -186.485 162.005 -186.155 ;
        RECT 161.675 -187.845 162.005 -187.515 ;
        RECT 161.675 -189.205 162.005 -188.875 ;
        RECT 161.675 -190.565 162.005 -190.235 ;
        RECT 161.675 -191.925 162.005 -191.595 ;
        RECT 161.675 -193.285 162.005 -192.955 ;
        RECT 161.675 -194.645 162.005 -194.315 ;
        RECT 161.675 -196.005 162.005 -195.675 ;
        RECT 161.675 -197.365 162.005 -197.035 ;
        RECT 161.675 -198.725 162.005 -198.395 ;
        RECT 161.675 -200.085 162.005 -199.755 ;
        RECT 161.675 -201.445 162.005 -201.115 ;
        RECT 161.675 -202.805 162.005 -202.475 ;
        RECT 161.675 -204.165 162.005 -203.835 ;
        RECT 161.675 -205.525 162.005 -205.195 ;
        RECT 161.675 -206.885 162.005 -206.555 ;
        RECT 161.675 -208.245 162.005 -207.915 ;
        RECT 161.675 -209.605 162.005 -209.275 ;
        RECT 161.675 -210.965 162.005 -210.635 ;
        RECT 161.675 -212.325 162.005 -211.995 ;
        RECT 161.675 -213.685 162.005 -213.355 ;
        RECT 161.675 -215.045 162.005 -214.715 ;
        RECT 161.675 -216.405 162.005 -216.075 ;
        RECT 161.675 -217.765 162.005 -217.435 ;
        RECT 161.675 -219.125 162.005 -218.795 ;
        RECT 161.675 -220.485 162.005 -220.155 ;
        RECT 161.675 -221.845 162.005 -221.515 ;
        RECT 161.675 -223.205 162.005 -222.875 ;
        RECT 161.675 -224.565 162.005 -224.235 ;
        RECT 161.675 -225.925 162.005 -225.595 ;
        RECT 161.675 -227.285 162.005 -226.955 ;
        RECT 161.675 -228.645 162.005 -228.315 ;
        RECT 161.675 -230.005 162.005 -229.675 ;
        RECT 161.675 -231.365 162.005 -231.035 ;
        RECT 161.675 -232.725 162.005 -232.395 ;
        RECT 161.675 -234.085 162.005 -233.755 ;
        RECT 161.675 -235.445 162.005 -235.115 ;
        RECT 161.675 -236.805 162.005 -236.475 ;
        RECT 161.675 -238.165 162.005 -237.835 ;
        RECT 161.675 -243.81 162.005 -242.68 ;
        RECT 161.68 -243.925 162 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 246.76 163.365 247.89 ;
        RECT 163.035 241.915 163.365 242.245 ;
        RECT 163.035 240.555 163.365 240.885 ;
        RECT 163.035 239.195 163.365 239.525 ;
        RECT 163.035 237.835 163.365 238.165 ;
        RECT 163.04 237.16 163.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 -1.525 163.365 -1.195 ;
        RECT 163.035 -2.885 163.365 -2.555 ;
        RECT 163.04 -3.56 163.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 -122.565 163.365 -122.235 ;
        RECT 163.035 -123.925 163.365 -123.595 ;
        RECT 163.035 -125.285 163.365 -124.955 ;
        RECT 163.035 -126.645 163.365 -126.315 ;
        RECT 163.035 -128.005 163.365 -127.675 ;
        RECT 163.035 -129.365 163.365 -129.035 ;
        RECT 163.035 -130.725 163.365 -130.395 ;
        RECT 163.035 -132.085 163.365 -131.755 ;
        RECT 163.035 -133.445 163.365 -133.115 ;
        RECT 163.035 -134.805 163.365 -134.475 ;
        RECT 163.035 -136.165 163.365 -135.835 ;
        RECT 163.035 -137.525 163.365 -137.195 ;
        RECT 163.035 -138.885 163.365 -138.555 ;
        RECT 163.035 -140.245 163.365 -139.915 ;
        RECT 163.035 -141.605 163.365 -141.275 ;
        RECT 163.035 -142.965 163.365 -142.635 ;
        RECT 163.035 -144.325 163.365 -143.995 ;
        RECT 163.035 -145.685 163.365 -145.355 ;
        RECT 163.035 -147.045 163.365 -146.715 ;
        RECT 163.035 -148.405 163.365 -148.075 ;
        RECT 163.035 -149.765 163.365 -149.435 ;
        RECT 163.035 -151.125 163.365 -150.795 ;
        RECT 163.035 -152.485 163.365 -152.155 ;
        RECT 163.035 -153.845 163.365 -153.515 ;
        RECT 163.035 -155.205 163.365 -154.875 ;
        RECT 163.035 -156.565 163.365 -156.235 ;
        RECT 163.035 -157.925 163.365 -157.595 ;
        RECT 163.035 -159.285 163.365 -158.955 ;
        RECT 163.035 -160.645 163.365 -160.315 ;
        RECT 163.035 -162.005 163.365 -161.675 ;
        RECT 163.035 -163.365 163.365 -163.035 ;
        RECT 163.035 -164.725 163.365 -164.395 ;
        RECT 163.035 -166.085 163.365 -165.755 ;
        RECT 163.035 -167.445 163.365 -167.115 ;
        RECT 163.035 -168.805 163.365 -168.475 ;
        RECT 163.035 -170.165 163.365 -169.835 ;
        RECT 163.035 -171.525 163.365 -171.195 ;
        RECT 163.035 -172.885 163.365 -172.555 ;
        RECT 163.035 -174.245 163.365 -173.915 ;
        RECT 163.035 -175.605 163.365 -175.275 ;
        RECT 163.035 -176.965 163.365 -176.635 ;
        RECT 163.035 -178.325 163.365 -177.995 ;
        RECT 163.035 -179.685 163.365 -179.355 ;
        RECT 163.035 -181.045 163.365 -180.715 ;
        RECT 163.035 -182.405 163.365 -182.075 ;
        RECT 163.035 -183.765 163.365 -183.435 ;
        RECT 163.035 -185.125 163.365 -184.795 ;
        RECT 163.035 -186.485 163.365 -186.155 ;
        RECT 163.035 -187.845 163.365 -187.515 ;
        RECT 163.035 -189.205 163.365 -188.875 ;
        RECT 163.035 -190.565 163.365 -190.235 ;
        RECT 163.035 -191.925 163.365 -191.595 ;
        RECT 163.035 -193.285 163.365 -192.955 ;
        RECT 163.035 -194.645 163.365 -194.315 ;
        RECT 163.035 -196.005 163.365 -195.675 ;
        RECT 163.035 -197.365 163.365 -197.035 ;
        RECT 163.035 -198.725 163.365 -198.395 ;
        RECT 163.035 -200.085 163.365 -199.755 ;
        RECT 163.035 -201.445 163.365 -201.115 ;
        RECT 163.035 -202.805 163.365 -202.475 ;
        RECT 163.035 -204.165 163.365 -203.835 ;
        RECT 163.035 -205.525 163.365 -205.195 ;
        RECT 163.035 -206.885 163.365 -206.555 ;
        RECT 163.035 -208.245 163.365 -207.915 ;
        RECT 163.035 -209.605 163.365 -209.275 ;
        RECT 163.035 -210.965 163.365 -210.635 ;
        RECT 163.035 -212.325 163.365 -211.995 ;
        RECT 163.035 -213.685 163.365 -213.355 ;
        RECT 163.035 -215.045 163.365 -214.715 ;
        RECT 163.035 -216.405 163.365 -216.075 ;
        RECT 163.035 -217.765 163.365 -217.435 ;
        RECT 163.035 -219.125 163.365 -218.795 ;
        RECT 163.035 -220.485 163.365 -220.155 ;
        RECT 163.035 -221.845 163.365 -221.515 ;
        RECT 163.035 -223.205 163.365 -222.875 ;
        RECT 163.035 -224.565 163.365 -224.235 ;
        RECT 163.035 -225.925 163.365 -225.595 ;
        RECT 163.035 -227.285 163.365 -226.955 ;
        RECT 163.035 -228.645 163.365 -228.315 ;
        RECT 163.035 -230.005 163.365 -229.675 ;
        RECT 163.035 -231.365 163.365 -231.035 ;
        RECT 163.035 -232.725 163.365 -232.395 ;
        RECT 163.035 -234.085 163.365 -233.755 ;
        RECT 163.035 -235.445 163.365 -235.115 ;
        RECT 163.035 -236.805 163.365 -236.475 ;
        RECT 163.035 -238.165 163.365 -237.835 ;
        RECT 163.035 -243.81 163.365 -242.68 ;
        RECT 163.04 -243.925 163.36 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 246.76 164.725 247.89 ;
        RECT 164.395 241.915 164.725 242.245 ;
        RECT 164.395 240.555 164.725 240.885 ;
        RECT 164.395 239.195 164.725 239.525 ;
        RECT 164.395 237.835 164.725 238.165 ;
        RECT 164.4 237.16 164.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 -1.525 164.725 -1.195 ;
        RECT 164.395 -2.885 164.725 -2.555 ;
        RECT 164.4 -3.56 164.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 -164.725 164.725 -164.395 ;
        RECT 164.395 -166.085 164.725 -165.755 ;
        RECT 164.395 -167.445 164.725 -167.115 ;
        RECT 164.395 -168.805 164.725 -168.475 ;
        RECT 164.395 -170.165 164.725 -169.835 ;
        RECT 164.395 -171.525 164.725 -171.195 ;
        RECT 164.395 -172.885 164.725 -172.555 ;
        RECT 164.395 -174.245 164.725 -173.915 ;
        RECT 164.395 -175.605 164.725 -175.275 ;
        RECT 164.395 -176.965 164.725 -176.635 ;
        RECT 164.395 -178.325 164.725 -177.995 ;
        RECT 164.395 -179.685 164.725 -179.355 ;
        RECT 164.395 -181.045 164.725 -180.715 ;
        RECT 164.395 -182.405 164.725 -182.075 ;
        RECT 164.395 -183.765 164.725 -183.435 ;
        RECT 164.395 -185.125 164.725 -184.795 ;
        RECT 164.395 -186.485 164.725 -186.155 ;
        RECT 164.395 -187.845 164.725 -187.515 ;
        RECT 164.395 -189.205 164.725 -188.875 ;
        RECT 164.395 -190.565 164.725 -190.235 ;
        RECT 164.395 -191.925 164.725 -191.595 ;
        RECT 164.395 -193.285 164.725 -192.955 ;
        RECT 164.395 -194.645 164.725 -194.315 ;
        RECT 164.395 -196.005 164.725 -195.675 ;
        RECT 164.395 -197.365 164.725 -197.035 ;
        RECT 164.395 -198.725 164.725 -198.395 ;
        RECT 164.395 -200.085 164.725 -199.755 ;
        RECT 164.395 -201.445 164.725 -201.115 ;
        RECT 164.395 -202.805 164.725 -202.475 ;
        RECT 164.395 -204.165 164.725 -203.835 ;
        RECT 164.395 -205.525 164.725 -205.195 ;
        RECT 164.395 -206.885 164.725 -206.555 ;
        RECT 164.395 -208.245 164.725 -207.915 ;
        RECT 164.395 -209.605 164.725 -209.275 ;
        RECT 164.395 -210.965 164.725 -210.635 ;
        RECT 164.395 -212.325 164.725 -211.995 ;
        RECT 164.395 -213.685 164.725 -213.355 ;
        RECT 164.395 -215.045 164.725 -214.715 ;
        RECT 164.395 -216.405 164.725 -216.075 ;
        RECT 164.395 -217.765 164.725 -217.435 ;
        RECT 164.395 -219.125 164.725 -218.795 ;
        RECT 164.395 -220.485 164.725 -220.155 ;
        RECT 164.395 -221.845 164.725 -221.515 ;
        RECT 164.395 -223.205 164.725 -222.875 ;
        RECT 164.395 -224.565 164.725 -224.235 ;
        RECT 164.395 -225.925 164.725 -225.595 ;
        RECT 164.395 -227.285 164.725 -226.955 ;
        RECT 164.395 -228.645 164.725 -228.315 ;
        RECT 164.395 -230.005 164.725 -229.675 ;
        RECT 164.395 -231.365 164.725 -231.035 ;
        RECT 164.395 -232.725 164.725 -232.395 ;
        RECT 164.395 -234.085 164.725 -233.755 ;
        RECT 164.395 -235.445 164.725 -235.115 ;
        RECT 164.395 -236.805 164.725 -236.475 ;
        RECT 164.395 -238.165 164.725 -237.835 ;
        RECT 164.395 -243.81 164.725 -242.68 ;
        RECT 164.4 -243.925 164.72 -122.235 ;
        RECT 164.395 -122.565 164.725 -122.235 ;
        RECT 164.395 -123.925 164.725 -123.595 ;
        RECT 164.395 -125.285 164.725 -124.955 ;
        RECT 164.395 -126.645 164.725 -126.315 ;
        RECT 164.395 -128.005 164.725 -127.675 ;
        RECT 164.395 -129.365 164.725 -129.035 ;
        RECT 164.395 -130.725 164.725 -130.395 ;
        RECT 164.395 -132.085 164.725 -131.755 ;
        RECT 164.395 -133.445 164.725 -133.115 ;
        RECT 164.395 -134.805 164.725 -134.475 ;
        RECT 164.395 -136.165 164.725 -135.835 ;
        RECT 164.395 -137.525 164.725 -137.195 ;
        RECT 164.395 -138.885 164.725 -138.555 ;
        RECT 164.395 -140.245 164.725 -139.915 ;
        RECT 164.395 -141.605 164.725 -141.275 ;
        RECT 164.395 -142.965 164.725 -142.635 ;
        RECT 164.395 -144.325 164.725 -143.995 ;
        RECT 164.395 -145.685 164.725 -145.355 ;
        RECT 164.395 -147.045 164.725 -146.715 ;
        RECT 164.395 -148.405 164.725 -148.075 ;
        RECT 164.395 -149.765 164.725 -149.435 ;
        RECT 164.395 -151.125 164.725 -150.795 ;
        RECT 164.395 -152.485 164.725 -152.155 ;
        RECT 164.395 -153.845 164.725 -153.515 ;
        RECT 164.395 -155.205 164.725 -154.875 ;
        RECT 164.395 -156.565 164.725 -156.235 ;
        RECT 164.395 -157.925 164.725 -157.595 ;
        RECT 164.395 -159.285 164.725 -158.955 ;
        RECT 164.395 -160.645 164.725 -160.315 ;
        RECT 164.395 -162.005 164.725 -161.675 ;
        RECT 164.395 -163.365 164.725 -163.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 246.76 130.725 247.89 ;
        RECT 130.395 241.915 130.725 242.245 ;
        RECT 130.395 240.555 130.725 240.885 ;
        RECT 130.395 239.195 130.725 239.525 ;
        RECT 130.395 237.835 130.725 238.165 ;
        RECT 130.4 237.16 130.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 -1.525 130.725 -1.195 ;
        RECT 130.395 -2.885 130.725 -2.555 ;
        RECT 130.4 -3.56 130.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 -122.565 130.725 -122.235 ;
        RECT 130.395 -123.925 130.725 -123.595 ;
        RECT 130.395 -125.285 130.725 -124.955 ;
        RECT 130.395 -126.645 130.725 -126.315 ;
        RECT 130.395 -128.005 130.725 -127.675 ;
        RECT 130.395 -129.365 130.725 -129.035 ;
        RECT 130.395 -130.725 130.725 -130.395 ;
        RECT 130.395 -132.085 130.725 -131.755 ;
        RECT 130.395 -133.445 130.725 -133.115 ;
        RECT 130.395 -134.805 130.725 -134.475 ;
        RECT 130.395 -136.165 130.725 -135.835 ;
        RECT 130.395 -137.525 130.725 -137.195 ;
        RECT 130.395 -138.885 130.725 -138.555 ;
        RECT 130.395 -140.245 130.725 -139.915 ;
        RECT 130.395 -141.605 130.725 -141.275 ;
        RECT 130.395 -142.965 130.725 -142.635 ;
        RECT 130.395 -144.325 130.725 -143.995 ;
        RECT 130.395 -145.685 130.725 -145.355 ;
        RECT 130.395 -147.045 130.725 -146.715 ;
        RECT 130.395 -148.405 130.725 -148.075 ;
        RECT 130.395 -149.765 130.725 -149.435 ;
        RECT 130.395 -151.125 130.725 -150.795 ;
        RECT 130.395 -152.485 130.725 -152.155 ;
        RECT 130.395 -153.845 130.725 -153.515 ;
        RECT 130.395 -155.205 130.725 -154.875 ;
        RECT 130.395 -156.565 130.725 -156.235 ;
        RECT 130.395 -157.925 130.725 -157.595 ;
        RECT 130.395 -159.285 130.725 -158.955 ;
        RECT 130.395 -160.645 130.725 -160.315 ;
        RECT 130.395 -162.005 130.725 -161.675 ;
        RECT 130.395 -163.365 130.725 -163.035 ;
        RECT 130.395 -164.725 130.725 -164.395 ;
        RECT 130.395 -166.085 130.725 -165.755 ;
        RECT 130.395 -167.445 130.725 -167.115 ;
        RECT 130.395 -168.805 130.725 -168.475 ;
        RECT 130.395 -170.165 130.725 -169.835 ;
        RECT 130.395 -171.525 130.725 -171.195 ;
        RECT 130.395 -172.885 130.725 -172.555 ;
        RECT 130.395 -174.245 130.725 -173.915 ;
        RECT 130.395 -175.605 130.725 -175.275 ;
        RECT 130.395 -176.965 130.725 -176.635 ;
        RECT 130.395 -178.325 130.725 -177.995 ;
        RECT 130.395 -179.685 130.725 -179.355 ;
        RECT 130.395 -181.045 130.725 -180.715 ;
        RECT 130.395 -182.405 130.725 -182.075 ;
        RECT 130.395 -183.765 130.725 -183.435 ;
        RECT 130.395 -185.125 130.725 -184.795 ;
        RECT 130.395 -186.485 130.725 -186.155 ;
        RECT 130.395 -187.845 130.725 -187.515 ;
        RECT 130.395 -189.205 130.725 -188.875 ;
        RECT 130.395 -190.565 130.725 -190.235 ;
        RECT 130.395 -191.925 130.725 -191.595 ;
        RECT 130.395 -193.285 130.725 -192.955 ;
        RECT 130.395 -194.645 130.725 -194.315 ;
        RECT 130.395 -196.005 130.725 -195.675 ;
        RECT 130.395 -197.365 130.725 -197.035 ;
        RECT 130.395 -198.725 130.725 -198.395 ;
        RECT 130.395 -200.085 130.725 -199.755 ;
        RECT 130.395 -201.445 130.725 -201.115 ;
        RECT 130.395 -202.805 130.725 -202.475 ;
        RECT 130.395 -204.165 130.725 -203.835 ;
        RECT 130.395 -205.525 130.725 -205.195 ;
        RECT 130.395 -206.885 130.725 -206.555 ;
        RECT 130.395 -208.245 130.725 -207.915 ;
        RECT 130.395 -209.605 130.725 -209.275 ;
        RECT 130.395 -210.965 130.725 -210.635 ;
        RECT 130.395 -212.325 130.725 -211.995 ;
        RECT 130.395 -213.685 130.725 -213.355 ;
        RECT 130.395 -215.045 130.725 -214.715 ;
        RECT 130.395 -216.405 130.725 -216.075 ;
        RECT 130.395 -217.765 130.725 -217.435 ;
        RECT 130.395 -219.125 130.725 -218.795 ;
        RECT 130.395 -220.485 130.725 -220.155 ;
        RECT 130.395 -221.845 130.725 -221.515 ;
        RECT 130.395 -223.205 130.725 -222.875 ;
        RECT 130.395 -224.565 130.725 -224.235 ;
        RECT 130.395 -225.925 130.725 -225.595 ;
        RECT 130.395 -227.285 130.725 -226.955 ;
        RECT 130.395 -228.645 130.725 -228.315 ;
        RECT 130.395 -230.005 130.725 -229.675 ;
        RECT 130.395 -231.365 130.725 -231.035 ;
        RECT 130.395 -232.725 130.725 -232.395 ;
        RECT 130.395 -234.085 130.725 -233.755 ;
        RECT 130.395 -235.445 130.725 -235.115 ;
        RECT 130.395 -236.805 130.725 -236.475 ;
        RECT 130.395 -238.165 130.725 -237.835 ;
        RECT 130.395 -243.81 130.725 -242.68 ;
        RECT 130.4 -243.925 130.72 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 246.76 132.085 247.89 ;
        RECT 131.755 241.915 132.085 242.245 ;
        RECT 131.755 240.555 132.085 240.885 ;
        RECT 131.755 239.195 132.085 239.525 ;
        RECT 131.755 237.835 132.085 238.165 ;
        RECT 131.76 237.16 132.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 -1.525 132.085 -1.195 ;
        RECT 131.755 -2.885 132.085 -2.555 ;
        RECT 131.76 -3.56 132.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 -122.565 132.085 -122.235 ;
        RECT 131.755 -123.925 132.085 -123.595 ;
        RECT 131.755 -125.285 132.085 -124.955 ;
        RECT 131.755 -126.645 132.085 -126.315 ;
        RECT 131.755 -128.005 132.085 -127.675 ;
        RECT 131.755 -129.365 132.085 -129.035 ;
        RECT 131.755 -130.725 132.085 -130.395 ;
        RECT 131.755 -132.085 132.085 -131.755 ;
        RECT 131.755 -133.445 132.085 -133.115 ;
        RECT 131.755 -134.805 132.085 -134.475 ;
        RECT 131.755 -136.165 132.085 -135.835 ;
        RECT 131.755 -137.525 132.085 -137.195 ;
        RECT 131.755 -138.885 132.085 -138.555 ;
        RECT 131.755 -140.245 132.085 -139.915 ;
        RECT 131.755 -141.605 132.085 -141.275 ;
        RECT 131.755 -142.965 132.085 -142.635 ;
        RECT 131.755 -144.325 132.085 -143.995 ;
        RECT 131.755 -145.685 132.085 -145.355 ;
        RECT 131.755 -147.045 132.085 -146.715 ;
        RECT 131.755 -148.405 132.085 -148.075 ;
        RECT 131.755 -149.765 132.085 -149.435 ;
        RECT 131.755 -151.125 132.085 -150.795 ;
        RECT 131.755 -152.485 132.085 -152.155 ;
        RECT 131.755 -153.845 132.085 -153.515 ;
        RECT 131.755 -155.205 132.085 -154.875 ;
        RECT 131.755 -156.565 132.085 -156.235 ;
        RECT 131.755 -157.925 132.085 -157.595 ;
        RECT 131.755 -159.285 132.085 -158.955 ;
        RECT 131.755 -160.645 132.085 -160.315 ;
        RECT 131.755 -162.005 132.085 -161.675 ;
        RECT 131.755 -163.365 132.085 -163.035 ;
        RECT 131.755 -164.725 132.085 -164.395 ;
        RECT 131.755 -166.085 132.085 -165.755 ;
        RECT 131.755 -167.445 132.085 -167.115 ;
        RECT 131.755 -168.805 132.085 -168.475 ;
        RECT 131.755 -170.165 132.085 -169.835 ;
        RECT 131.755 -171.525 132.085 -171.195 ;
        RECT 131.755 -172.885 132.085 -172.555 ;
        RECT 131.755 -174.245 132.085 -173.915 ;
        RECT 131.755 -175.605 132.085 -175.275 ;
        RECT 131.755 -176.965 132.085 -176.635 ;
        RECT 131.755 -178.325 132.085 -177.995 ;
        RECT 131.755 -179.685 132.085 -179.355 ;
        RECT 131.755 -181.045 132.085 -180.715 ;
        RECT 131.755 -182.405 132.085 -182.075 ;
        RECT 131.755 -183.765 132.085 -183.435 ;
        RECT 131.755 -185.125 132.085 -184.795 ;
        RECT 131.755 -186.485 132.085 -186.155 ;
        RECT 131.755 -187.845 132.085 -187.515 ;
        RECT 131.755 -189.205 132.085 -188.875 ;
        RECT 131.755 -190.565 132.085 -190.235 ;
        RECT 131.755 -191.925 132.085 -191.595 ;
        RECT 131.755 -193.285 132.085 -192.955 ;
        RECT 131.755 -194.645 132.085 -194.315 ;
        RECT 131.755 -196.005 132.085 -195.675 ;
        RECT 131.755 -197.365 132.085 -197.035 ;
        RECT 131.755 -198.725 132.085 -198.395 ;
        RECT 131.755 -200.085 132.085 -199.755 ;
        RECT 131.755 -201.445 132.085 -201.115 ;
        RECT 131.755 -202.805 132.085 -202.475 ;
        RECT 131.755 -204.165 132.085 -203.835 ;
        RECT 131.755 -205.525 132.085 -205.195 ;
        RECT 131.755 -206.885 132.085 -206.555 ;
        RECT 131.755 -208.245 132.085 -207.915 ;
        RECT 131.755 -209.605 132.085 -209.275 ;
        RECT 131.755 -210.965 132.085 -210.635 ;
        RECT 131.755 -212.325 132.085 -211.995 ;
        RECT 131.755 -213.685 132.085 -213.355 ;
        RECT 131.755 -215.045 132.085 -214.715 ;
        RECT 131.755 -216.405 132.085 -216.075 ;
        RECT 131.755 -217.765 132.085 -217.435 ;
        RECT 131.755 -219.125 132.085 -218.795 ;
        RECT 131.755 -220.485 132.085 -220.155 ;
        RECT 131.755 -221.845 132.085 -221.515 ;
        RECT 131.755 -223.205 132.085 -222.875 ;
        RECT 131.755 -224.565 132.085 -224.235 ;
        RECT 131.755 -225.925 132.085 -225.595 ;
        RECT 131.755 -227.285 132.085 -226.955 ;
        RECT 131.755 -228.645 132.085 -228.315 ;
        RECT 131.755 -230.005 132.085 -229.675 ;
        RECT 131.755 -231.365 132.085 -231.035 ;
        RECT 131.755 -232.725 132.085 -232.395 ;
        RECT 131.755 -234.085 132.085 -233.755 ;
        RECT 131.755 -235.445 132.085 -235.115 ;
        RECT 131.755 -236.805 132.085 -236.475 ;
        RECT 131.755 -238.165 132.085 -237.835 ;
        RECT 131.755 -243.81 132.085 -242.68 ;
        RECT 131.76 -243.925 132.08 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 246.76 133.445 247.89 ;
        RECT 133.115 241.915 133.445 242.245 ;
        RECT 133.115 240.555 133.445 240.885 ;
        RECT 133.115 239.195 133.445 239.525 ;
        RECT 133.115 237.835 133.445 238.165 ;
        RECT 133.12 237.16 133.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 -126.645 133.445 -126.315 ;
        RECT 133.115 -128.005 133.445 -127.675 ;
        RECT 133.115 -129.365 133.445 -129.035 ;
        RECT 133.115 -130.725 133.445 -130.395 ;
        RECT 133.115 -132.085 133.445 -131.755 ;
        RECT 133.115 -133.445 133.445 -133.115 ;
        RECT 133.115 -134.805 133.445 -134.475 ;
        RECT 133.115 -136.165 133.445 -135.835 ;
        RECT 133.115 -137.525 133.445 -137.195 ;
        RECT 133.115 -138.885 133.445 -138.555 ;
        RECT 133.115 -140.245 133.445 -139.915 ;
        RECT 133.115 -141.605 133.445 -141.275 ;
        RECT 133.115 -142.965 133.445 -142.635 ;
        RECT 133.115 -144.325 133.445 -143.995 ;
        RECT 133.115 -145.685 133.445 -145.355 ;
        RECT 133.115 -147.045 133.445 -146.715 ;
        RECT 133.115 -148.405 133.445 -148.075 ;
        RECT 133.115 -149.765 133.445 -149.435 ;
        RECT 133.115 -151.125 133.445 -150.795 ;
        RECT 133.115 -152.485 133.445 -152.155 ;
        RECT 133.115 -153.845 133.445 -153.515 ;
        RECT 133.115 -155.205 133.445 -154.875 ;
        RECT 133.115 -156.565 133.445 -156.235 ;
        RECT 133.115 -157.925 133.445 -157.595 ;
        RECT 133.115 -159.285 133.445 -158.955 ;
        RECT 133.115 -160.645 133.445 -160.315 ;
        RECT 133.115 -162.005 133.445 -161.675 ;
        RECT 133.115 -163.365 133.445 -163.035 ;
        RECT 133.115 -164.725 133.445 -164.395 ;
        RECT 133.115 -166.085 133.445 -165.755 ;
        RECT 133.115 -167.445 133.445 -167.115 ;
        RECT 133.115 -168.805 133.445 -168.475 ;
        RECT 133.115 -170.165 133.445 -169.835 ;
        RECT 133.115 -171.525 133.445 -171.195 ;
        RECT 133.115 -172.885 133.445 -172.555 ;
        RECT 133.115 -174.245 133.445 -173.915 ;
        RECT 133.115 -175.605 133.445 -175.275 ;
        RECT 133.115 -176.965 133.445 -176.635 ;
        RECT 133.115 -178.325 133.445 -177.995 ;
        RECT 133.115 -179.685 133.445 -179.355 ;
        RECT 133.115 -181.045 133.445 -180.715 ;
        RECT 133.115 -182.405 133.445 -182.075 ;
        RECT 133.115 -183.765 133.445 -183.435 ;
        RECT 133.115 -185.125 133.445 -184.795 ;
        RECT 133.115 -186.485 133.445 -186.155 ;
        RECT 133.115 -187.845 133.445 -187.515 ;
        RECT 133.115 -189.205 133.445 -188.875 ;
        RECT 133.115 -190.565 133.445 -190.235 ;
        RECT 133.115 -191.925 133.445 -191.595 ;
        RECT 133.115 -193.285 133.445 -192.955 ;
        RECT 133.115 -194.645 133.445 -194.315 ;
        RECT 133.115 -196.005 133.445 -195.675 ;
        RECT 133.115 -197.365 133.445 -197.035 ;
        RECT 133.115 -198.725 133.445 -198.395 ;
        RECT 133.115 -200.085 133.445 -199.755 ;
        RECT 133.115 -201.445 133.445 -201.115 ;
        RECT 133.115 -202.805 133.445 -202.475 ;
        RECT 133.115 -204.165 133.445 -203.835 ;
        RECT 133.115 -205.525 133.445 -205.195 ;
        RECT 133.115 -206.885 133.445 -206.555 ;
        RECT 133.115 -208.245 133.445 -207.915 ;
        RECT 133.115 -209.605 133.445 -209.275 ;
        RECT 133.115 -210.965 133.445 -210.635 ;
        RECT 133.115 -212.325 133.445 -211.995 ;
        RECT 133.115 -213.685 133.445 -213.355 ;
        RECT 133.115 -215.045 133.445 -214.715 ;
        RECT 133.115 -216.405 133.445 -216.075 ;
        RECT 133.115 -217.765 133.445 -217.435 ;
        RECT 133.115 -219.125 133.445 -218.795 ;
        RECT 133.115 -220.485 133.445 -220.155 ;
        RECT 133.115 -221.845 133.445 -221.515 ;
        RECT 133.115 -223.205 133.445 -222.875 ;
        RECT 133.115 -224.565 133.445 -224.235 ;
        RECT 133.115 -225.925 133.445 -225.595 ;
        RECT 133.115 -227.285 133.445 -226.955 ;
        RECT 133.115 -228.645 133.445 -228.315 ;
        RECT 133.115 -230.005 133.445 -229.675 ;
        RECT 133.115 -231.365 133.445 -231.035 ;
        RECT 133.115 -232.725 133.445 -232.395 ;
        RECT 133.115 -234.085 133.445 -233.755 ;
        RECT 133.115 -235.445 133.445 -235.115 ;
        RECT 133.115 -236.805 133.445 -236.475 ;
        RECT 133.115 -238.165 133.445 -237.835 ;
        RECT 133.115 -243.81 133.445 -242.68 ;
        RECT 133.12 -243.925 133.44 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.46 -125.535 133.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 246.76 134.805 247.89 ;
        RECT 134.475 241.915 134.805 242.245 ;
        RECT 134.475 240.555 134.805 240.885 ;
        RECT 134.475 239.195 134.805 239.525 ;
        RECT 134.475 237.835 134.805 238.165 ;
        RECT 134.48 237.16 134.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 246.76 136.165 247.89 ;
        RECT 135.835 241.915 136.165 242.245 ;
        RECT 135.835 240.555 136.165 240.885 ;
        RECT 135.835 239.195 136.165 239.525 ;
        RECT 135.835 237.835 136.165 238.165 ;
        RECT 135.84 237.16 136.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 -1.525 136.165 -1.195 ;
        RECT 135.835 -2.885 136.165 -2.555 ;
        RECT 135.84 -3.56 136.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 246.76 137.525 247.89 ;
        RECT 137.195 241.915 137.525 242.245 ;
        RECT 137.195 240.555 137.525 240.885 ;
        RECT 137.195 239.195 137.525 239.525 ;
        RECT 137.195 237.835 137.525 238.165 ;
        RECT 137.2 237.16 137.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 -1.525 137.525 -1.195 ;
        RECT 137.195 -2.885 137.525 -2.555 ;
        RECT 137.2 -3.56 137.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 -122.565 137.525 -122.235 ;
        RECT 137.195 -123.925 137.525 -123.595 ;
        RECT 137.195 -125.285 137.525 -124.955 ;
        RECT 137.195 -126.645 137.525 -126.315 ;
        RECT 137.195 -128.005 137.525 -127.675 ;
        RECT 137.195 -129.365 137.525 -129.035 ;
        RECT 137.195 -130.725 137.525 -130.395 ;
        RECT 137.195 -132.085 137.525 -131.755 ;
        RECT 137.195 -133.445 137.525 -133.115 ;
        RECT 137.195 -134.805 137.525 -134.475 ;
        RECT 137.195 -136.165 137.525 -135.835 ;
        RECT 137.195 -137.525 137.525 -137.195 ;
        RECT 137.195 -138.885 137.525 -138.555 ;
        RECT 137.195 -140.245 137.525 -139.915 ;
        RECT 137.195 -141.605 137.525 -141.275 ;
        RECT 137.195 -142.965 137.525 -142.635 ;
        RECT 137.195 -144.325 137.525 -143.995 ;
        RECT 137.195 -145.685 137.525 -145.355 ;
        RECT 137.195 -147.045 137.525 -146.715 ;
        RECT 137.195 -148.405 137.525 -148.075 ;
        RECT 137.195 -149.765 137.525 -149.435 ;
        RECT 137.195 -151.125 137.525 -150.795 ;
        RECT 137.195 -152.485 137.525 -152.155 ;
        RECT 137.195 -153.845 137.525 -153.515 ;
        RECT 137.195 -155.205 137.525 -154.875 ;
        RECT 137.195 -156.565 137.525 -156.235 ;
        RECT 137.195 -157.925 137.525 -157.595 ;
        RECT 137.195 -159.285 137.525 -158.955 ;
        RECT 137.195 -160.645 137.525 -160.315 ;
        RECT 137.195 -162.005 137.525 -161.675 ;
        RECT 137.195 -163.365 137.525 -163.035 ;
        RECT 137.195 -164.725 137.525 -164.395 ;
        RECT 137.195 -166.085 137.525 -165.755 ;
        RECT 137.195 -167.445 137.525 -167.115 ;
        RECT 137.195 -168.805 137.525 -168.475 ;
        RECT 137.195 -170.165 137.525 -169.835 ;
        RECT 137.195 -171.525 137.525 -171.195 ;
        RECT 137.195 -172.885 137.525 -172.555 ;
        RECT 137.195 -174.245 137.525 -173.915 ;
        RECT 137.195 -175.605 137.525 -175.275 ;
        RECT 137.195 -176.965 137.525 -176.635 ;
        RECT 137.195 -178.325 137.525 -177.995 ;
        RECT 137.195 -179.685 137.525 -179.355 ;
        RECT 137.195 -181.045 137.525 -180.715 ;
        RECT 137.195 -182.405 137.525 -182.075 ;
        RECT 137.195 -183.765 137.525 -183.435 ;
        RECT 137.195 -185.125 137.525 -184.795 ;
        RECT 137.195 -186.485 137.525 -186.155 ;
        RECT 137.195 -187.845 137.525 -187.515 ;
        RECT 137.195 -189.205 137.525 -188.875 ;
        RECT 137.195 -190.565 137.525 -190.235 ;
        RECT 137.195 -191.925 137.525 -191.595 ;
        RECT 137.195 -193.285 137.525 -192.955 ;
        RECT 137.195 -194.645 137.525 -194.315 ;
        RECT 137.195 -196.005 137.525 -195.675 ;
        RECT 137.195 -197.365 137.525 -197.035 ;
        RECT 137.195 -198.725 137.525 -198.395 ;
        RECT 137.195 -200.085 137.525 -199.755 ;
        RECT 137.195 -201.445 137.525 -201.115 ;
        RECT 137.195 -202.805 137.525 -202.475 ;
        RECT 137.195 -204.165 137.525 -203.835 ;
        RECT 137.195 -205.525 137.525 -205.195 ;
        RECT 137.195 -206.885 137.525 -206.555 ;
        RECT 137.195 -208.245 137.525 -207.915 ;
        RECT 137.195 -209.605 137.525 -209.275 ;
        RECT 137.195 -210.965 137.525 -210.635 ;
        RECT 137.195 -212.325 137.525 -211.995 ;
        RECT 137.195 -213.685 137.525 -213.355 ;
        RECT 137.195 -215.045 137.525 -214.715 ;
        RECT 137.195 -216.405 137.525 -216.075 ;
        RECT 137.195 -217.765 137.525 -217.435 ;
        RECT 137.195 -219.125 137.525 -218.795 ;
        RECT 137.195 -220.485 137.525 -220.155 ;
        RECT 137.195 -221.845 137.525 -221.515 ;
        RECT 137.195 -223.205 137.525 -222.875 ;
        RECT 137.195 -224.565 137.525 -224.235 ;
        RECT 137.195 -225.925 137.525 -225.595 ;
        RECT 137.195 -227.285 137.525 -226.955 ;
        RECT 137.195 -228.645 137.525 -228.315 ;
        RECT 137.195 -230.005 137.525 -229.675 ;
        RECT 137.195 -231.365 137.525 -231.035 ;
        RECT 137.195 -232.725 137.525 -232.395 ;
        RECT 137.195 -234.085 137.525 -233.755 ;
        RECT 137.195 -235.445 137.525 -235.115 ;
        RECT 137.195 -236.805 137.525 -236.475 ;
        RECT 137.195 -238.165 137.525 -237.835 ;
        RECT 137.195 -243.81 137.525 -242.68 ;
        RECT 137.2 -243.925 137.52 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 246.76 138.885 247.89 ;
        RECT 138.555 241.915 138.885 242.245 ;
        RECT 138.555 240.555 138.885 240.885 ;
        RECT 138.555 239.195 138.885 239.525 ;
        RECT 138.555 237.835 138.885 238.165 ;
        RECT 138.56 237.16 138.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 -1.525 138.885 -1.195 ;
        RECT 138.555 -2.885 138.885 -2.555 ;
        RECT 138.56 -3.56 138.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 -122.565 138.885 -122.235 ;
        RECT 138.555 -123.925 138.885 -123.595 ;
        RECT 138.555 -125.285 138.885 -124.955 ;
        RECT 138.555 -126.645 138.885 -126.315 ;
        RECT 138.555 -128.005 138.885 -127.675 ;
        RECT 138.555 -129.365 138.885 -129.035 ;
        RECT 138.555 -130.725 138.885 -130.395 ;
        RECT 138.555 -132.085 138.885 -131.755 ;
        RECT 138.555 -133.445 138.885 -133.115 ;
        RECT 138.555 -134.805 138.885 -134.475 ;
        RECT 138.555 -136.165 138.885 -135.835 ;
        RECT 138.555 -137.525 138.885 -137.195 ;
        RECT 138.555 -138.885 138.885 -138.555 ;
        RECT 138.555 -140.245 138.885 -139.915 ;
        RECT 138.555 -141.605 138.885 -141.275 ;
        RECT 138.555 -142.965 138.885 -142.635 ;
        RECT 138.555 -144.325 138.885 -143.995 ;
        RECT 138.555 -145.685 138.885 -145.355 ;
        RECT 138.555 -147.045 138.885 -146.715 ;
        RECT 138.555 -148.405 138.885 -148.075 ;
        RECT 138.555 -149.765 138.885 -149.435 ;
        RECT 138.555 -151.125 138.885 -150.795 ;
        RECT 138.555 -152.485 138.885 -152.155 ;
        RECT 138.555 -153.845 138.885 -153.515 ;
        RECT 138.555 -155.205 138.885 -154.875 ;
        RECT 138.555 -156.565 138.885 -156.235 ;
        RECT 138.555 -157.925 138.885 -157.595 ;
        RECT 138.555 -159.285 138.885 -158.955 ;
        RECT 138.555 -160.645 138.885 -160.315 ;
        RECT 138.555 -162.005 138.885 -161.675 ;
        RECT 138.555 -163.365 138.885 -163.035 ;
        RECT 138.555 -164.725 138.885 -164.395 ;
        RECT 138.555 -166.085 138.885 -165.755 ;
        RECT 138.555 -167.445 138.885 -167.115 ;
        RECT 138.555 -168.805 138.885 -168.475 ;
        RECT 138.555 -170.165 138.885 -169.835 ;
        RECT 138.555 -171.525 138.885 -171.195 ;
        RECT 138.555 -172.885 138.885 -172.555 ;
        RECT 138.555 -174.245 138.885 -173.915 ;
        RECT 138.555 -175.605 138.885 -175.275 ;
        RECT 138.555 -176.965 138.885 -176.635 ;
        RECT 138.555 -178.325 138.885 -177.995 ;
        RECT 138.555 -179.685 138.885 -179.355 ;
        RECT 138.555 -181.045 138.885 -180.715 ;
        RECT 138.555 -182.405 138.885 -182.075 ;
        RECT 138.555 -183.765 138.885 -183.435 ;
        RECT 138.555 -185.125 138.885 -184.795 ;
        RECT 138.555 -186.485 138.885 -186.155 ;
        RECT 138.555 -187.845 138.885 -187.515 ;
        RECT 138.555 -189.205 138.885 -188.875 ;
        RECT 138.555 -190.565 138.885 -190.235 ;
        RECT 138.555 -191.925 138.885 -191.595 ;
        RECT 138.555 -193.285 138.885 -192.955 ;
        RECT 138.555 -194.645 138.885 -194.315 ;
        RECT 138.555 -196.005 138.885 -195.675 ;
        RECT 138.555 -197.365 138.885 -197.035 ;
        RECT 138.555 -198.725 138.885 -198.395 ;
        RECT 138.555 -200.085 138.885 -199.755 ;
        RECT 138.555 -201.445 138.885 -201.115 ;
        RECT 138.555 -202.805 138.885 -202.475 ;
        RECT 138.555 -204.165 138.885 -203.835 ;
        RECT 138.555 -205.525 138.885 -205.195 ;
        RECT 138.555 -206.885 138.885 -206.555 ;
        RECT 138.555 -208.245 138.885 -207.915 ;
        RECT 138.555 -209.605 138.885 -209.275 ;
        RECT 138.555 -210.965 138.885 -210.635 ;
        RECT 138.555 -212.325 138.885 -211.995 ;
        RECT 138.555 -213.685 138.885 -213.355 ;
        RECT 138.555 -215.045 138.885 -214.715 ;
        RECT 138.555 -216.405 138.885 -216.075 ;
        RECT 138.555 -217.765 138.885 -217.435 ;
        RECT 138.555 -219.125 138.885 -218.795 ;
        RECT 138.555 -220.485 138.885 -220.155 ;
        RECT 138.555 -221.845 138.885 -221.515 ;
        RECT 138.555 -223.205 138.885 -222.875 ;
        RECT 138.555 -224.565 138.885 -224.235 ;
        RECT 138.555 -225.925 138.885 -225.595 ;
        RECT 138.555 -227.285 138.885 -226.955 ;
        RECT 138.555 -228.645 138.885 -228.315 ;
        RECT 138.555 -230.005 138.885 -229.675 ;
        RECT 138.555 -231.365 138.885 -231.035 ;
        RECT 138.555 -232.725 138.885 -232.395 ;
        RECT 138.555 -234.085 138.885 -233.755 ;
        RECT 138.555 -235.445 138.885 -235.115 ;
        RECT 138.555 -236.805 138.885 -236.475 ;
        RECT 138.555 -238.165 138.885 -237.835 ;
        RECT 138.555 -243.81 138.885 -242.68 ;
        RECT 138.56 -243.925 138.88 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 246.76 140.245 247.89 ;
        RECT 139.915 241.915 140.245 242.245 ;
        RECT 139.915 240.555 140.245 240.885 ;
        RECT 139.915 239.195 140.245 239.525 ;
        RECT 139.915 237.835 140.245 238.165 ;
        RECT 139.92 237.16 140.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 -1.525 140.245 -1.195 ;
        RECT 139.915 -2.885 140.245 -2.555 ;
        RECT 139.92 -3.56 140.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 -122.565 140.245 -122.235 ;
        RECT 139.915 -123.925 140.245 -123.595 ;
        RECT 139.915 -125.285 140.245 -124.955 ;
        RECT 139.915 -126.645 140.245 -126.315 ;
        RECT 139.915 -128.005 140.245 -127.675 ;
        RECT 139.915 -129.365 140.245 -129.035 ;
        RECT 139.915 -130.725 140.245 -130.395 ;
        RECT 139.915 -132.085 140.245 -131.755 ;
        RECT 139.915 -133.445 140.245 -133.115 ;
        RECT 139.915 -134.805 140.245 -134.475 ;
        RECT 139.915 -136.165 140.245 -135.835 ;
        RECT 139.915 -137.525 140.245 -137.195 ;
        RECT 139.915 -138.885 140.245 -138.555 ;
        RECT 139.915 -140.245 140.245 -139.915 ;
        RECT 139.915 -141.605 140.245 -141.275 ;
        RECT 139.915 -142.965 140.245 -142.635 ;
        RECT 139.915 -144.325 140.245 -143.995 ;
        RECT 139.915 -145.685 140.245 -145.355 ;
        RECT 139.915 -147.045 140.245 -146.715 ;
        RECT 139.915 -148.405 140.245 -148.075 ;
        RECT 139.915 -149.765 140.245 -149.435 ;
        RECT 139.915 -151.125 140.245 -150.795 ;
        RECT 139.915 -152.485 140.245 -152.155 ;
        RECT 139.915 -153.845 140.245 -153.515 ;
        RECT 139.915 -155.205 140.245 -154.875 ;
        RECT 139.915 -156.565 140.245 -156.235 ;
        RECT 139.915 -157.925 140.245 -157.595 ;
        RECT 139.915 -159.285 140.245 -158.955 ;
        RECT 139.915 -160.645 140.245 -160.315 ;
        RECT 139.915 -162.005 140.245 -161.675 ;
        RECT 139.915 -163.365 140.245 -163.035 ;
        RECT 139.915 -164.725 140.245 -164.395 ;
        RECT 139.915 -166.085 140.245 -165.755 ;
        RECT 139.915 -167.445 140.245 -167.115 ;
        RECT 139.915 -168.805 140.245 -168.475 ;
        RECT 139.915 -170.165 140.245 -169.835 ;
        RECT 139.915 -171.525 140.245 -171.195 ;
        RECT 139.915 -172.885 140.245 -172.555 ;
        RECT 139.915 -174.245 140.245 -173.915 ;
        RECT 139.915 -175.605 140.245 -175.275 ;
        RECT 139.915 -176.965 140.245 -176.635 ;
        RECT 139.915 -178.325 140.245 -177.995 ;
        RECT 139.915 -179.685 140.245 -179.355 ;
        RECT 139.915 -181.045 140.245 -180.715 ;
        RECT 139.915 -182.405 140.245 -182.075 ;
        RECT 139.915 -183.765 140.245 -183.435 ;
        RECT 139.915 -185.125 140.245 -184.795 ;
        RECT 139.915 -186.485 140.245 -186.155 ;
        RECT 139.915 -187.845 140.245 -187.515 ;
        RECT 139.915 -189.205 140.245 -188.875 ;
        RECT 139.915 -190.565 140.245 -190.235 ;
        RECT 139.915 -191.925 140.245 -191.595 ;
        RECT 139.915 -193.285 140.245 -192.955 ;
        RECT 139.915 -194.645 140.245 -194.315 ;
        RECT 139.915 -196.005 140.245 -195.675 ;
        RECT 139.915 -197.365 140.245 -197.035 ;
        RECT 139.915 -198.725 140.245 -198.395 ;
        RECT 139.915 -200.085 140.245 -199.755 ;
        RECT 139.915 -201.445 140.245 -201.115 ;
        RECT 139.915 -202.805 140.245 -202.475 ;
        RECT 139.915 -204.165 140.245 -203.835 ;
        RECT 139.915 -205.525 140.245 -205.195 ;
        RECT 139.915 -206.885 140.245 -206.555 ;
        RECT 139.915 -208.245 140.245 -207.915 ;
        RECT 139.915 -209.605 140.245 -209.275 ;
        RECT 139.915 -210.965 140.245 -210.635 ;
        RECT 139.915 -212.325 140.245 -211.995 ;
        RECT 139.915 -213.685 140.245 -213.355 ;
        RECT 139.915 -215.045 140.245 -214.715 ;
        RECT 139.915 -216.405 140.245 -216.075 ;
        RECT 139.915 -217.765 140.245 -217.435 ;
        RECT 139.915 -219.125 140.245 -218.795 ;
        RECT 139.915 -220.485 140.245 -220.155 ;
        RECT 139.915 -221.845 140.245 -221.515 ;
        RECT 139.915 -223.205 140.245 -222.875 ;
        RECT 139.915 -224.565 140.245 -224.235 ;
        RECT 139.915 -225.925 140.245 -225.595 ;
        RECT 139.915 -227.285 140.245 -226.955 ;
        RECT 139.915 -228.645 140.245 -228.315 ;
        RECT 139.915 -230.005 140.245 -229.675 ;
        RECT 139.915 -231.365 140.245 -231.035 ;
        RECT 139.915 -232.725 140.245 -232.395 ;
        RECT 139.915 -234.085 140.245 -233.755 ;
        RECT 139.915 -235.445 140.245 -235.115 ;
        RECT 139.915 -236.805 140.245 -236.475 ;
        RECT 139.915 -238.165 140.245 -237.835 ;
        RECT 139.915 -243.81 140.245 -242.68 ;
        RECT 139.92 -243.925 140.24 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 246.76 141.605 247.89 ;
        RECT 141.275 241.915 141.605 242.245 ;
        RECT 141.275 240.555 141.605 240.885 ;
        RECT 141.275 239.195 141.605 239.525 ;
        RECT 141.275 237.835 141.605 238.165 ;
        RECT 141.28 237.16 141.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -1.525 141.605 -1.195 ;
        RECT 141.275 -2.885 141.605 -2.555 ;
        RECT 141.28 -3.56 141.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -122.565 141.605 -122.235 ;
        RECT 141.275 -123.925 141.605 -123.595 ;
        RECT 141.275 -125.285 141.605 -124.955 ;
        RECT 141.275 -126.645 141.605 -126.315 ;
        RECT 141.275 -128.005 141.605 -127.675 ;
        RECT 141.275 -129.365 141.605 -129.035 ;
        RECT 141.275 -130.725 141.605 -130.395 ;
        RECT 141.275 -132.085 141.605 -131.755 ;
        RECT 141.275 -133.445 141.605 -133.115 ;
        RECT 141.275 -134.805 141.605 -134.475 ;
        RECT 141.275 -136.165 141.605 -135.835 ;
        RECT 141.275 -137.525 141.605 -137.195 ;
        RECT 141.275 -138.885 141.605 -138.555 ;
        RECT 141.275 -140.245 141.605 -139.915 ;
        RECT 141.275 -141.605 141.605 -141.275 ;
        RECT 141.275 -142.965 141.605 -142.635 ;
        RECT 141.275 -144.325 141.605 -143.995 ;
        RECT 141.275 -145.685 141.605 -145.355 ;
        RECT 141.275 -147.045 141.605 -146.715 ;
        RECT 141.275 -148.405 141.605 -148.075 ;
        RECT 141.275 -149.765 141.605 -149.435 ;
        RECT 141.275 -151.125 141.605 -150.795 ;
        RECT 141.275 -152.485 141.605 -152.155 ;
        RECT 141.275 -153.845 141.605 -153.515 ;
        RECT 141.275 -155.205 141.605 -154.875 ;
        RECT 141.275 -156.565 141.605 -156.235 ;
        RECT 141.275 -157.925 141.605 -157.595 ;
        RECT 141.275 -159.285 141.605 -158.955 ;
        RECT 141.275 -160.645 141.605 -160.315 ;
        RECT 141.275 -162.005 141.605 -161.675 ;
        RECT 141.275 -163.365 141.605 -163.035 ;
        RECT 141.275 -164.725 141.605 -164.395 ;
        RECT 141.275 -166.085 141.605 -165.755 ;
        RECT 141.275 -167.445 141.605 -167.115 ;
        RECT 141.275 -168.805 141.605 -168.475 ;
        RECT 141.275 -170.165 141.605 -169.835 ;
        RECT 141.275 -171.525 141.605 -171.195 ;
        RECT 141.275 -172.885 141.605 -172.555 ;
        RECT 141.275 -174.245 141.605 -173.915 ;
        RECT 141.275 -175.605 141.605 -175.275 ;
        RECT 141.275 -176.965 141.605 -176.635 ;
        RECT 141.275 -178.325 141.605 -177.995 ;
        RECT 141.275 -179.685 141.605 -179.355 ;
        RECT 141.275 -181.045 141.605 -180.715 ;
        RECT 141.275 -182.405 141.605 -182.075 ;
        RECT 141.275 -183.765 141.605 -183.435 ;
        RECT 141.275 -185.125 141.605 -184.795 ;
        RECT 141.275 -186.485 141.605 -186.155 ;
        RECT 141.275 -187.845 141.605 -187.515 ;
        RECT 141.275 -189.205 141.605 -188.875 ;
        RECT 141.275 -190.565 141.605 -190.235 ;
        RECT 141.275 -191.925 141.605 -191.595 ;
        RECT 141.275 -193.285 141.605 -192.955 ;
        RECT 141.275 -194.645 141.605 -194.315 ;
        RECT 141.275 -196.005 141.605 -195.675 ;
        RECT 141.275 -197.365 141.605 -197.035 ;
        RECT 141.275 -198.725 141.605 -198.395 ;
        RECT 141.275 -200.085 141.605 -199.755 ;
        RECT 141.275 -201.445 141.605 -201.115 ;
        RECT 141.275 -202.805 141.605 -202.475 ;
        RECT 141.275 -204.165 141.605 -203.835 ;
        RECT 141.275 -205.525 141.605 -205.195 ;
        RECT 141.275 -206.885 141.605 -206.555 ;
        RECT 141.275 -208.245 141.605 -207.915 ;
        RECT 141.275 -209.605 141.605 -209.275 ;
        RECT 141.275 -210.965 141.605 -210.635 ;
        RECT 141.275 -212.325 141.605 -211.995 ;
        RECT 141.275 -213.685 141.605 -213.355 ;
        RECT 141.275 -215.045 141.605 -214.715 ;
        RECT 141.275 -216.405 141.605 -216.075 ;
        RECT 141.275 -217.765 141.605 -217.435 ;
        RECT 141.275 -219.125 141.605 -218.795 ;
        RECT 141.275 -220.485 141.605 -220.155 ;
        RECT 141.275 -221.845 141.605 -221.515 ;
        RECT 141.275 -223.205 141.605 -222.875 ;
        RECT 141.275 -224.565 141.605 -224.235 ;
        RECT 141.275 -225.925 141.605 -225.595 ;
        RECT 141.275 -227.285 141.605 -226.955 ;
        RECT 141.275 -228.645 141.605 -228.315 ;
        RECT 141.275 -230.005 141.605 -229.675 ;
        RECT 141.275 -231.365 141.605 -231.035 ;
        RECT 141.275 -232.725 141.605 -232.395 ;
        RECT 141.275 -234.085 141.605 -233.755 ;
        RECT 141.275 -235.445 141.605 -235.115 ;
        RECT 141.275 -236.805 141.605 -236.475 ;
        RECT 141.275 -238.165 141.605 -237.835 ;
        RECT 141.275 -243.81 141.605 -242.68 ;
        RECT 141.28 -243.925 141.6 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 246.76 142.965 247.89 ;
        RECT 142.635 241.915 142.965 242.245 ;
        RECT 142.635 240.555 142.965 240.885 ;
        RECT 142.635 239.195 142.965 239.525 ;
        RECT 142.635 237.835 142.965 238.165 ;
        RECT 142.64 237.16 142.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 -1.525 142.965 -1.195 ;
        RECT 142.635 -2.885 142.965 -2.555 ;
        RECT 142.64 -3.56 142.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 -122.565 142.965 -122.235 ;
        RECT 142.635 -123.925 142.965 -123.595 ;
        RECT 142.635 -125.285 142.965 -124.955 ;
        RECT 142.635 -126.645 142.965 -126.315 ;
        RECT 142.635 -128.005 142.965 -127.675 ;
        RECT 142.635 -129.365 142.965 -129.035 ;
        RECT 142.635 -130.725 142.965 -130.395 ;
        RECT 142.635 -132.085 142.965 -131.755 ;
        RECT 142.635 -133.445 142.965 -133.115 ;
        RECT 142.635 -134.805 142.965 -134.475 ;
        RECT 142.635 -136.165 142.965 -135.835 ;
        RECT 142.635 -137.525 142.965 -137.195 ;
        RECT 142.635 -138.885 142.965 -138.555 ;
        RECT 142.635 -140.245 142.965 -139.915 ;
        RECT 142.635 -141.605 142.965 -141.275 ;
        RECT 142.635 -142.965 142.965 -142.635 ;
        RECT 142.635 -144.325 142.965 -143.995 ;
        RECT 142.635 -145.685 142.965 -145.355 ;
        RECT 142.635 -147.045 142.965 -146.715 ;
        RECT 142.635 -148.405 142.965 -148.075 ;
        RECT 142.635 -149.765 142.965 -149.435 ;
        RECT 142.635 -151.125 142.965 -150.795 ;
        RECT 142.635 -152.485 142.965 -152.155 ;
        RECT 142.635 -153.845 142.965 -153.515 ;
        RECT 142.635 -155.205 142.965 -154.875 ;
        RECT 142.635 -156.565 142.965 -156.235 ;
        RECT 142.635 -157.925 142.965 -157.595 ;
        RECT 142.635 -159.285 142.965 -158.955 ;
        RECT 142.635 -160.645 142.965 -160.315 ;
        RECT 142.635 -162.005 142.965 -161.675 ;
        RECT 142.635 -163.365 142.965 -163.035 ;
        RECT 142.635 -164.725 142.965 -164.395 ;
        RECT 142.635 -166.085 142.965 -165.755 ;
        RECT 142.635 -167.445 142.965 -167.115 ;
        RECT 142.635 -168.805 142.965 -168.475 ;
        RECT 142.635 -170.165 142.965 -169.835 ;
        RECT 142.635 -171.525 142.965 -171.195 ;
        RECT 142.635 -172.885 142.965 -172.555 ;
        RECT 142.635 -174.245 142.965 -173.915 ;
        RECT 142.635 -175.605 142.965 -175.275 ;
        RECT 142.635 -176.965 142.965 -176.635 ;
        RECT 142.635 -178.325 142.965 -177.995 ;
        RECT 142.635 -179.685 142.965 -179.355 ;
        RECT 142.635 -181.045 142.965 -180.715 ;
        RECT 142.635 -182.405 142.965 -182.075 ;
        RECT 142.635 -183.765 142.965 -183.435 ;
        RECT 142.635 -185.125 142.965 -184.795 ;
        RECT 142.635 -186.485 142.965 -186.155 ;
        RECT 142.635 -187.845 142.965 -187.515 ;
        RECT 142.635 -189.205 142.965 -188.875 ;
        RECT 142.635 -190.565 142.965 -190.235 ;
        RECT 142.635 -191.925 142.965 -191.595 ;
        RECT 142.635 -193.285 142.965 -192.955 ;
        RECT 142.635 -194.645 142.965 -194.315 ;
        RECT 142.635 -196.005 142.965 -195.675 ;
        RECT 142.635 -197.365 142.965 -197.035 ;
        RECT 142.635 -198.725 142.965 -198.395 ;
        RECT 142.635 -200.085 142.965 -199.755 ;
        RECT 142.635 -201.445 142.965 -201.115 ;
        RECT 142.635 -202.805 142.965 -202.475 ;
        RECT 142.635 -204.165 142.965 -203.835 ;
        RECT 142.635 -205.525 142.965 -205.195 ;
        RECT 142.635 -206.885 142.965 -206.555 ;
        RECT 142.635 -208.245 142.965 -207.915 ;
        RECT 142.635 -209.605 142.965 -209.275 ;
        RECT 142.635 -210.965 142.965 -210.635 ;
        RECT 142.635 -212.325 142.965 -211.995 ;
        RECT 142.635 -213.685 142.965 -213.355 ;
        RECT 142.635 -215.045 142.965 -214.715 ;
        RECT 142.635 -216.405 142.965 -216.075 ;
        RECT 142.635 -217.765 142.965 -217.435 ;
        RECT 142.635 -219.125 142.965 -218.795 ;
        RECT 142.635 -220.485 142.965 -220.155 ;
        RECT 142.635 -221.845 142.965 -221.515 ;
        RECT 142.635 -223.205 142.965 -222.875 ;
        RECT 142.635 -224.565 142.965 -224.235 ;
        RECT 142.635 -225.925 142.965 -225.595 ;
        RECT 142.635 -227.285 142.965 -226.955 ;
        RECT 142.635 -228.645 142.965 -228.315 ;
        RECT 142.635 -230.005 142.965 -229.675 ;
        RECT 142.635 -231.365 142.965 -231.035 ;
        RECT 142.635 -232.725 142.965 -232.395 ;
        RECT 142.635 -234.085 142.965 -233.755 ;
        RECT 142.635 -235.445 142.965 -235.115 ;
        RECT 142.635 -236.805 142.965 -236.475 ;
        RECT 142.635 -238.165 142.965 -237.835 ;
        RECT 142.635 -243.81 142.965 -242.68 ;
        RECT 142.64 -243.925 142.96 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 246.76 144.325 247.89 ;
        RECT 143.995 241.915 144.325 242.245 ;
        RECT 143.995 240.555 144.325 240.885 ;
        RECT 143.995 239.195 144.325 239.525 ;
        RECT 143.995 237.835 144.325 238.165 ;
        RECT 144 237.16 144.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 -126.645 144.325 -126.315 ;
        RECT 143.995 -128.005 144.325 -127.675 ;
        RECT 143.995 -129.365 144.325 -129.035 ;
        RECT 143.995 -130.725 144.325 -130.395 ;
        RECT 143.995 -132.085 144.325 -131.755 ;
        RECT 143.995 -133.445 144.325 -133.115 ;
        RECT 143.995 -134.805 144.325 -134.475 ;
        RECT 143.995 -136.165 144.325 -135.835 ;
        RECT 143.995 -137.525 144.325 -137.195 ;
        RECT 143.995 -138.885 144.325 -138.555 ;
        RECT 143.995 -140.245 144.325 -139.915 ;
        RECT 143.995 -141.605 144.325 -141.275 ;
        RECT 143.995 -142.965 144.325 -142.635 ;
        RECT 143.995 -144.325 144.325 -143.995 ;
        RECT 143.995 -145.685 144.325 -145.355 ;
        RECT 143.995 -147.045 144.325 -146.715 ;
        RECT 143.995 -148.405 144.325 -148.075 ;
        RECT 143.995 -149.765 144.325 -149.435 ;
        RECT 143.995 -151.125 144.325 -150.795 ;
        RECT 143.995 -152.485 144.325 -152.155 ;
        RECT 143.995 -153.845 144.325 -153.515 ;
        RECT 143.995 -155.205 144.325 -154.875 ;
        RECT 143.995 -156.565 144.325 -156.235 ;
        RECT 143.995 -157.925 144.325 -157.595 ;
        RECT 143.995 -159.285 144.325 -158.955 ;
        RECT 143.995 -160.645 144.325 -160.315 ;
        RECT 143.995 -162.005 144.325 -161.675 ;
        RECT 143.995 -163.365 144.325 -163.035 ;
        RECT 143.995 -164.725 144.325 -164.395 ;
        RECT 143.995 -166.085 144.325 -165.755 ;
        RECT 143.995 -167.445 144.325 -167.115 ;
        RECT 143.995 -168.805 144.325 -168.475 ;
        RECT 143.995 -170.165 144.325 -169.835 ;
        RECT 143.995 -171.525 144.325 -171.195 ;
        RECT 143.995 -172.885 144.325 -172.555 ;
        RECT 143.995 -174.245 144.325 -173.915 ;
        RECT 143.995 -175.605 144.325 -175.275 ;
        RECT 143.995 -176.965 144.325 -176.635 ;
        RECT 143.995 -178.325 144.325 -177.995 ;
        RECT 143.995 -179.685 144.325 -179.355 ;
        RECT 143.995 -181.045 144.325 -180.715 ;
        RECT 143.995 -182.405 144.325 -182.075 ;
        RECT 143.995 -183.765 144.325 -183.435 ;
        RECT 143.995 -185.125 144.325 -184.795 ;
        RECT 143.995 -186.485 144.325 -186.155 ;
        RECT 143.995 -187.845 144.325 -187.515 ;
        RECT 143.995 -189.205 144.325 -188.875 ;
        RECT 143.995 -190.565 144.325 -190.235 ;
        RECT 143.995 -191.925 144.325 -191.595 ;
        RECT 143.995 -193.285 144.325 -192.955 ;
        RECT 143.995 -194.645 144.325 -194.315 ;
        RECT 143.995 -196.005 144.325 -195.675 ;
        RECT 143.995 -197.365 144.325 -197.035 ;
        RECT 143.995 -198.725 144.325 -198.395 ;
        RECT 143.995 -200.085 144.325 -199.755 ;
        RECT 143.995 -201.445 144.325 -201.115 ;
        RECT 143.995 -202.805 144.325 -202.475 ;
        RECT 143.995 -204.165 144.325 -203.835 ;
        RECT 143.995 -205.525 144.325 -205.195 ;
        RECT 143.995 -206.885 144.325 -206.555 ;
        RECT 143.995 -208.245 144.325 -207.915 ;
        RECT 143.995 -209.605 144.325 -209.275 ;
        RECT 143.995 -210.965 144.325 -210.635 ;
        RECT 143.995 -212.325 144.325 -211.995 ;
        RECT 143.995 -213.685 144.325 -213.355 ;
        RECT 143.995 -215.045 144.325 -214.715 ;
        RECT 143.995 -216.405 144.325 -216.075 ;
        RECT 143.995 -217.765 144.325 -217.435 ;
        RECT 143.995 -219.125 144.325 -218.795 ;
        RECT 143.995 -220.485 144.325 -220.155 ;
        RECT 143.995 -221.845 144.325 -221.515 ;
        RECT 143.995 -223.205 144.325 -222.875 ;
        RECT 143.995 -224.565 144.325 -224.235 ;
        RECT 143.995 -225.925 144.325 -225.595 ;
        RECT 143.995 -227.285 144.325 -226.955 ;
        RECT 143.995 -228.645 144.325 -228.315 ;
        RECT 143.995 -230.005 144.325 -229.675 ;
        RECT 143.995 -231.365 144.325 -231.035 ;
        RECT 143.995 -232.725 144.325 -232.395 ;
        RECT 143.995 -234.085 144.325 -233.755 ;
        RECT 143.995 -235.445 144.325 -235.115 ;
        RECT 143.995 -236.805 144.325 -236.475 ;
        RECT 143.995 -238.165 144.325 -237.835 ;
        RECT 143.995 -243.81 144.325 -242.68 ;
        RECT 144 -243.925 144.32 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.36 -125.535 144.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 246.76 145.685 247.89 ;
        RECT 145.355 241.915 145.685 242.245 ;
        RECT 145.355 240.555 145.685 240.885 ;
        RECT 145.355 239.195 145.685 239.525 ;
        RECT 145.355 237.835 145.685 238.165 ;
        RECT 145.36 237.16 145.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 246.76 147.045 247.89 ;
        RECT 146.715 241.915 147.045 242.245 ;
        RECT 146.715 240.555 147.045 240.885 ;
        RECT 146.715 239.195 147.045 239.525 ;
        RECT 146.715 237.835 147.045 238.165 ;
        RECT 146.72 237.16 147.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 -1.525 147.045 -1.195 ;
        RECT 146.715 -2.885 147.045 -2.555 ;
        RECT 146.72 -3.56 147.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 246.76 148.405 247.89 ;
        RECT 148.075 241.915 148.405 242.245 ;
        RECT 148.075 240.555 148.405 240.885 ;
        RECT 148.075 239.195 148.405 239.525 ;
        RECT 148.075 237.835 148.405 238.165 ;
        RECT 148.08 237.16 148.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -1.525 148.405 -1.195 ;
        RECT 148.075 -2.885 148.405 -2.555 ;
        RECT 148.08 -3.56 148.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -191.925 148.405 -191.595 ;
        RECT 148.075 -193.285 148.405 -192.955 ;
        RECT 148.075 -194.645 148.405 -194.315 ;
        RECT 148.075 -196.005 148.405 -195.675 ;
        RECT 148.075 -197.365 148.405 -197.035 ;
        RECT 148.075 -198.725 148.405 -198.395 ;
        RECT 148.075 -200.085 148.405 -199.755 ;
        RECT 148.075 -201.445 148.405 -201.115 ;
        RECT 148.075 -202.805 148.405 -202.475 ;
        RECT 148.075 -204.165 148.405 -203.835 ;
        RECT 148.075 -205.525 148.405 -205.195 ;
        RECT 148.075 -206.885 148.405 -206.555 ;
        RECT 148.075 -208.245 148.405 -207.915 ;
        RECT 148.075 -209.605 148.405 -209.275 ;
        RECT 148.075 -210.965 148.405 -210.635 ;
        RECT 148.075 -212.325 148.405 -211.995 ;
        RECT 148.075 -213.685 148.405 -213.355 ;
        RECT 148.075 -215.045 148.405 -214.715 ;
        RECT 148.075 -216.405 148.405 -216.075 ;
        RECT 148.075 -217.765 148.405 -217.435 ;
        RECT 148.075 -219.125 148.405 -218.795 ;
        RECT 148.075 -220.485 148.405 -220.155 ;
        RECT 148.075 -221.845 148.405 -221.515 ;
        RECT 148.075 -223.205 148.405 -222.875 ;
        RECT 148.075 -224.565 148.405 -224.235 ;
        RECT 148.075 -225.925 148.405 -225.595 ;
        RECT 148.075 -227.285 148.405 -226.955 ;
        RECT 148.075 -228.645 148.405 -228.315 ;
        RECT 148.075 -230.005 148.405 -229.675 ;
        RECT 148.075 -231.365 148.405 -231.035 ;
        RECT 148.075 -232.725 148.405 -232.395 ;
        RECT 148.075 -234.085 148.405 -233.755 ;
        RECT 148.075 -235.445 148.405 -235.115 ;
        RECT 148.075 -236.805 148.405 -236.475 ;
        RECT 148.075 -238.165 148.405 -237.835 ;
        RECT 148.075 -243.81 148.405 -242.68 ;
        RECT 148.08 -243.925 148.4 -122.235 ;
        RECT 148.075 -122.565 148.405 -122.235 ;
        RECT 148.075 -123.925 148.405 -123.595 ;
        RECT 148.075 -125.285 148.405 -124.955 ;
        RECT 148.075 -126.645 148.405 -126.315 ;
        RECT 148.075 -128.005 148.405 -127.675 ;
        RECT 148.075 -129.365 148.405 -129.035 ;
        RECT 148.075 -130.725 148.405 -130.395 ;
        RECT 148.075 -132.085 148.405 -131.755 ;
        RECT 148.075 -133.445 148.405 -133.115 ;
        RECT 148.075 -134.805 148.405 -134.475 ;
        RECT 148.075 -136.165 148.405 -135.835 ;
        RECT 148.075 -137.525 148.405 -137.195 ;
        RECT 148.075 -138.885 148.405 -138.555 ;
        RECT 148.075 -140.245 148.405 -139.915 ;
        RECT 148.075 -141.605 148.405 -141.275 ;
        RECT 148.075 -142.965 148.405 -142.635 ;
        RECT 148.075 -144.325 148.405 -143.995 ;
        RECT 148.075 -145.685 148.405 -145.355 ;
        RECT 148.075 -147.045 148.405 -146.715 ;
        RECT 148.075 -148.405 148.405 -148.075 ;
        RECT 148.075 -149.765 148.405 -149.435 ;
        RECT 148.075 -151.125 148.405 -150.795 ;
        RECT 148.075 -152.485 148.405 -152.155 ;
        RECT 148.075 -153.845 148.405 -153.515 ;
        RECT 148.075 -155.205 148.405 -154.875 ;
        RECT 148.075 -156.565 148.405 -156.235 ;
        RECT 148.075 -157.925 148.405 -157.595 ;
        RECT 148.075 -159.285 148.405 -158.955 ;
        RECT 148.075 -160.645 148.405 -160.315 ;
        RECT 148.075 -162.005 148.405 -161.675 ;
        RECT 148.075 -163.365 148.405 -163.035 ;
        RECT 148.075 -164.725 148.405 -164.395 ;
        RECT 148.075 -166.085 148.405 -165.755 ;
        RECT 148.075 -167.445 148.405 -167.115 ;
        RECT 148.075 -168.805 148.405 -168.475 ;
        RECT 148.075 -170.165 148.405 -169.835 ;
        RECT 148.075 -171.525 148.405 -171.195 ;
        RECT 148.075 -172.885 148.405 -172.555 ;
        RECT 148.075 -174.245 148.405 -173.915 ;
        RECT 148.075 -175.605 148.405 -175.275 ;
        RECT 148.075 -176.965 148.405 -176.635 ;
        RECT 148.075 -178.325 148.405 -177.995 ;
        RECT 148.075 -179.685 148.405 -179.355 ;
        RECT 148.075 -181.045 148.405 -180.715 ;
        RECT 148.075 -182.405 148.405 -182.075 ;
        RECT 148.075 -183.765 148.405 -183.435 ;
        RECT 148.075 -185.125 148.405 -184.795 ;
        RECT 148.075 -186.485 148.405 -186.155 ;
        RECT 148.075 -187.845 148.405 -187.515 ;
        RECT 148.075 -189.205 148.405 -188.875 ;
        RECT 148.075 -190.565 148.405 -190.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 246.76 111.685 247.89 ;
        RECT 111.355 241.915 111.685 242.245 ;
        RECT 111.355 240.555 111.685 240.885 ;
        RECT 111.355 239.195 111.685 239.525 ;
        RECT 111.355 237.835 111.685 238.165 ;
        RECT 111.36 237.16 111.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 -126.645 111.685 -126.315 ;
        RECT 111.355 -128.005 111.685 -127.675 ;
        RECT 111.355 -129.365 111.685 -129.035 ;
        RECT 111.355 -130.725 111.685 -130.395 ;
        RECT 111.355 -132.085 111.685 -131.755 ;
        RECT 111.355 -133.445 111.685 -133.115 ;
        RECT 111.355 -134.805 111.685 -134.475 ;
        RECT 111.355 -136.165 111.685 -135.835 ;
        RECT 111.355 -137.525 111.685 -137.195 ;
        RECT 111.355 -138.885 111.685 -138.555 ;
        RECT 111.355 -140.245 111.685 -139.915 ;
        RECT 111.355 -141.605 111.685 -141.275 ;
        RECT 111.355 -142.965 111.685 -142.635 ;
        RECT 111.355 -144.325 111.685 -143.995 ;
        RECT 111.355 -145.685 111.685 -145.355 ;
        RECT 111.355 -147.045 111.685 -146.715 ;
        RECT 111.355 -148.405 111.685 -148.075 ;
        RECT 111.355 -149.765 111.685 -149.435 ;
        RECT 111.355 -151.125 111.685 -150.795 ;
        RECT 111.355 -152.485 111.685 -152.155 ;
        RECT 111.355 -153.845 111.685 -153.515 ;
        RECT 111.355 -155.205 111.685 -154.875 ;
        RECT 111.355 -156.565 111.685 -156.235 ;
        RECT 111.355 -157.925 111.685 -157.595 ;
        RECT 111.355 -159.285 111.685 -158.955 ;
        RECT 111.355 -160.645 111.685 -160.315 ;
        RECT 111.355 -162.005 111.685 -161.675 ;
        RECT 111.355 -163.365 111.685 -163.035 ;
        RECT 111.355 -164.725 111.685 -164.395 ;
        RECT 111.355 -166.085 111.685 -165.755 ;
        RECT 111.355 -167.445 111.685 -167.115 ;
        RECT 111.355 -168.805 111.685 -168.475 ;
        RECT 111.355 -170.165 111.685 -169.835 ;
        RECT 111.355 -171.525 111.685 -171.195 ;
        RECT 111.355 -172.885 111.685 -172.555 ;
        RECT 111.355 -174.245 111.685 -173.915 ;
        RECT 111.355 -175.605 111.685 -175.275 ;
        RECT 111.355 -176.965 111.685 -176.635 ;
        RECT 111.355 -178.325 111.685 -177.995 ;
        RECT 111.355 -179.685 111.685 -179.355 ;
        RECT 111.355 -181.045 111.685 -180.715 ;
        RECT 111.355 -182.405 111.685 -182.075 ;
        RECT 111.355 -183.765 111.685 -183.435 ;
        RECT 111.355 -185.125 111.685 -184.795 ;
        RECT 111.355 -186.485 111.685 -186.155 ;
        RECT 111.355 -187.845 111.685 -187.515 ;
        RECT 111.355 -189.205 111.685 -188.875 ;
        RECT 111.355 -190.565 111.685 -190.235 ;
        RECT 111.355 -191.925 111.685 -191.595 ;
        RECT 111.355 -193.285 111.685 -192.955 ;
        RECT 111.355 -194.645 111.685 -194.315 ;
        RECT 111.355 -196.005 111.685 -195.675 ;
        RECT 111.355 -197.365 111.685 -197.035 ;
        RECT 111.355 -198.725 111.685 -198.395 ;
        RECT 111.355 -200.085 111.685 -199.755 ;
        RECT 111.355 -201.445 111.685 -201.115 ;
        RECT 111.355 -202.805 111.685 -202.475 ;
        RECT 111.355 -204.165 111.685 -203.835 ;
        RECT 111.355 -205.525 111.685 -205.195 ;
        RECT 111.355 -206.885 111.685 -206.555 ;
        RECT 111.355 -208.245 111.685 -207.915 ;
        RECT 111.355 -209.605 111.685 -209.275 ;
        RECT 111.355 -210.965 111.685 -210.635 ;
        RECT 111.355 -212.325 111.685 -211.995 ;
        RECT 111.355 -213.685 111.685 -213.355 ;
        RECT 111.355 -215.045 111.685 -214.715 ;
        RECT 111.355 -216.405 111.685 -216.075 ;
        RECT 111.355 -217.765 111.685 -217.435 ;
        RECT 111.355 -219.125 111.685 -218.795 ;
        RECT 111.355 -220.485 111.685 -220.155 ;
        RECT 111.355 -221.845 111.685 -221.515 ;
        RECT 111.355 -223.205 111.685 -222.875 ;
        RECT 111.355 -224.565 111.685 -224.235 ;
        RECT 111.355 -225.925 111.685 -225.595 ;
        RECT 111.355 -227.285 111.685 -226.955 ;
        RECT 111.355 -228.645 111.685 -228.315 ;
        RECT 111.355 -230.005 111.685 -229.675 ;
        RECT 111.355 -231.365 111.685 -231.035 ;
        RECT 111.355 -232.725 111.685 -232.395 ;
        RECT 111.355 -234.085 111.685 -233.755 ;
        RECT 111.355 -235.445 111.685 -235.115 ;
        RECT 111.355 -236.805 111.685 -236.475 ;
        RECT 111.355 -238.165 111.685 -237.835 ;
        RECT 111.355 -243.81 111.685 -242.68 ;
        RECT 111.36 -243.925 111.68 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.66 -125.535 111.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 246.76 113.045 247.89 ;
        RECT 112.715 241.915 113.045 242.245 ;
        RECT 112.715 240.555 113.045 240.885 ;
        RECT 112.715 239.195 113.045 239.525 ;
        RECT 112.715 237.835 113.045 238.165 ;
        RECT 112.72 237.16 113.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 246.76 114.405 247.89 ;
        RECT 114.075 241.915 114.405 242.245 ;
        RECT 114.075 240.555 114.405 240.885 ;
        RECT 114.075 239.195 114.405 239.525 ;
        RECT 114.075 237.835 114.405 238.165 ;
        RECT 114.08 237.16 114.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 -1.525 114.405 -1.195 ;
        RECT 114.075 -2.885 114.405 -2.555 ;
        RECT 114.08 -3.56 114.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 246.76 115.765 247.89 ;
        RECT 115.435 241.915 115.765 242.245 ;
        RECT 115.435 240.555 115.765 240.885 ;
        RECT 115.435 239.195 115.765 239.525 ;
        RECT 115.435 237.835 115.765 238.165 ;
        RECT 115.44 237.16 115.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 -1.525 115.765 -1.195 ;
        RECT 115.435 -2.885 115.765 -2.555 ;
        RECT 115.44 -3.56 115.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 -122.565 115.765 -122.235 ;
        RECT 115.435 -123.925 115.765 -123.595 ;
        RECT 115.435 -125.285 115.765 -124.955 ;
        RECT 115.435 -126.645 115.765 -126.315 ;
        RECT 115.435 -128.005 115.765 -127.675 ;
        RECT 115.435 -129.365 115.765 -129.035 ;
        RECT 115.435 -130.725 115.765 -130.395 ;
        RECT 115.435 -132.085 115.765 -131.755 ;
        RECT 115.435 -133.445 115.765 -133.115 ;
        RECT 115.435 -134.805 115.765 -134.475 ;
        RECT 115.435 -136.165 115.765 -135.835 ;
        RECT 115.435 -137.525 115.765 -137.195 ;
        RECT 115.435 -138.885 115.765 -138.555 ;
        RECT 115.435 -140.245 115.765 -139.915 ;
        RECT 115.435 -141.605 115.765 -141.275 ;
        RECT 115.435 -142.965 115.765 -142.635 ;
        RECT 115.435 -144.325 115.765 -143.995 ;
        RECT 115.435 -145.685 115.765 -145.355 ;
        RECT 115.435 -147.045 115.765 -146.715 ;
        RECT 115.435 -148.405 115.765 -148.075 ;
        RECT 115.435 -149.765 115.765 -149.435 ;
        RECT 115.435 -151.125 115.765 -150.795 ;
        RECT 115.435 -152.485 115.765 -152.155 ;
        RECT 115.435 -153.845 115.765 -153.515 ;
        RECT 115.435 -155.205 115.765 -154.875 ;
        RECT 115.435 -156.565 115.765 -156.235 ;
        RECT 115.435 -157.925 115.765 -157.595 ;
        RECT 115.435 -159.285 115.765 -158.955 ;
        RECT 115.435 -160.645 115.765 -160.315 ;
        RECT 115.435 -162.005 115.765 -161.675 ;
        RECT 115.435 -163.365 115.765 -163.035 ;
        RECT 115.435 -164.725 115.765 -164.395 ;
        RECT 115.435 -166.085 115.765 -165.755 ;
        RECT 115.435 -167.445 115.765 -167.115 ;
        RECT 115.435 -168.805 115.765 -168.475 ;
        RECT 115.435 -170.165 115.765 -169.835 ;
        RECT 115.435 -171.525 115.765 -171.195 ;
        RECT 115.435 -172.885 115.765 -172.555 ;
        RECT 115.435 -174.245 115.765 -173.915 ;
        RECT 115.435 -175.605 115.765 -175.275 ;
        RECT 115.435 -176.965 115.765 -176.635 ;
        RECT 115.435 -178.325 115.765 -177.995 ;
        RECT 115.435 -179.685 115.765 -179.355 ;
        RECT 115.435 -181.045 115.765 -180.715 ;
        RECT 115.435 -182.405 115.765 -182.075 ;
        RECT 115.435 -183.765 115.765 -183.435 ;
        RECT 115.435 -185.125 115.765 -184.795 ;
        RECT 115.435 -186.485 115.765 -186.155 ;
        RECT 115.435 -187.845 115.765 -187.515 ;
        RECT 115.435 -189.205 115.765 -188.875 ;
        RECT 115.435 -190.565 115.765 -190.235 ;
        RECT 115.435 -191.925 115.765 -191.595 ;
        RECT 115.435 -193.285 115.765 -192.955 ;
        RECT 115.435 -194.645 115.765 -194.315 ;
        RECT 115.435 -196.005 115.765 -195.675 ;
        RECT 115.435 -197.365 115.765 -197.035 ;
        RECT 115.435 -198.725 115.765 -198.395 ;
        RECT 115.435 -200.085 115.765 -199.755 ;
        RECT 115.435 -201.445 115.765 -201.115 ;
        RECT 115.435 -202.805 115.765 -202.475 ;
        RECT 115.435 -204.165 115.765 -203.835 ;
        RECT 115.435 -205.525 115.765 -205.195 ;
        RECT 115.435 -206.885 115.765 -206.555 ;
        RECT 115.435 -208.245 115.765 -207.915 ;
        RECT 115.435 -209.605 115.765 -209.275 ;
        RECT 115.435 -210.965 115.765 -210.635 ;
        RECT 115.435 -212.325 115.765 -211.995 ;
        RECT 115.435 -213.685 115.765 -213.355 ;
        RECT 115.435 -215.045 115.765 -214.715 ;
        RECT 115.435 -216.405 115.765 -216.075 ;
        RECT 115.435 -217.765 115.765 -217.435 ;
        RECT 115.435 -219.125 115.765 -218.795 ;
        RECT 115.435 -220.485 115.765 -220.155 ;
        RECT 115.435 -221.845 115.765 -221.515 ;
        RECT 115.435 -223.205 115.765 -222.875 ;
        RECT 115.435 -224.565 115.765 -224.235 ;
        RECT 115.435 -225.925 115.765 -225.595 ;
        RECT 115.435 -227.285 115.765 -226.955 ;
        RECT 115.435 -228.645 115.765 -228.315 ;
        RECT 115.435 -230.005 115.765 -229.675 ;
        RECT 115.435 -231.365 115.765 -231.035 ;
        RECT 115.435 -232.725 115.765 -232.395 ;
        RECT 115.435 -234.085 115.765 -233.755 ;
        RECT 115.435 -235.445 115.765 -235.115 ;
        RECT 115.435 -236.805 115.765 -236.475 ;
        RECT 115.435 -238.165 115.765 -237.835 ;
        RECT 115.435 -243.81 115.765 -242.68 ;
        RECT 115.44 -243.925 115.76 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 246.76 117.125 247.89 ;
        RECT 116.795 241.915 117.125 242.245 ;
        RECT 116.795 240.555 117.125 240.885 ;
        RECT 116.795 239.195 117.125 239.525 ;
        RECT 116.795 237.835 117.125 238.165 ;
        RECT 116.8 237.16 117.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -1.525 117.125 -1.195 ;
        RECT 116.795 -2.885 117.125 -2.555 ;
        RECT 116.8 -3.56 117.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -122.565 117.125 -122.235 ;
        RECT 116.795 -123.925 117.125 -123.595 ;
        RECT 116.795 -125.285 117.125 -124.955 ;
        RECT 116.795 -126.645 117.125 -126.315 ;
        RECT 116.795 -128.005 117.125 -127.675 ;
        RECT 116.795 -129.365 117.125 -129.035 ;
        RECT 116.795 -130.725 117.125 -130.395 ;
        RECT 116.795 -132.085 117.125 -131.755 ;
        RECT 116.795 -133.445 117.125 -133.115 ;
        RECT 116.795 -134.805 117.125 -134.475 ;
        RECT 116.795 -136.165 117.125 -135.835 ;
        RECT 116.795 -137.525 117.125 -137.195 ;
        RECT 116.795 -138.885 117.125 -138.555 ;
        RECT 116.795 -140.245 117.125 -139.915 ;
        RECT 116.795 -141.605 117.125 -141.275 ;
        RECT 116.795 -142.965 117.125 -142.635 ;
        RECT 116.795 -144.325 117.125 -143.995 ;
        RECT 116.795 -145.685 117.125 -145.355 ;
        RECT 116.795 -147.045 117.125 -146.715 ;
        RECT 116.795 -148.405 117.125 -148.075 ;
        RECT 116.795 -149.765 117.125 -149.435 ;
        RECT 116.795 -151.125 117.125 -150.795 ;
        RECT 116.795 -152.485 117.125 -152.155 ;
        RECT 116.795 -153.845 117.125 -153.515 ;
        RECT 116.795 -155.205 117.125 -154.875 ;
        RECT 116.795 -156.565 117.125 -156.235 ;
        RECT 116.795 -157.925 117.125 -157.595 ;
        RECT 116.795 -159.285 117.125 -158.955 ;
        RECT 116.795 -160.645 117.125 -160.315 ;
        RECT 116.795 -162.005 117.125 -161.675 ;
        RECT 116.795 -163.365 117.125 -163.035 ;
        RECT 116.795 -164.725 117.125 -164.395 ;
        RECT 116.795 -166.085 117.125 -165.755 ;
        RECT 116.795 -167.445 117.125 -167.115 ;
        RECT 116.795 -168.805 117.125 -168.475 ;
        RECT 116.795 -170.165 117.125 -169.835 ;
        RECT 116.795 -171.525 117.125 -171.195 ;
        RECT 116.795 -172.885 117.125 -172.555 ;
        RECT 116.795 -174.245 117.125 -173.915 ;
        RECT 116.795 -175.605 117.125 -175.275 ;
        RECT 116.795 -176.965 117.125 -176.635 ;
        RECT 116.795 -178.325 117.125 -177.995 ;
        RECT 116.795 -179.685 117.125 -179.355 ;
        RECT 116.795 -181.045 117.125 -180.715 ;
        RECT 116.795 -182.405 117.125 -182.075 ;
        RECT 116.795 -183.765 117.125 -183.435 ;
        RECT 116.795 -185.125 117.125 -184.795 ;
        RECT 116.795 -186.485 117.125 -186.155 ;
        RECT 116.795 -187.845 117.125 -187.515 ;
        RECT 116.795 -189.205 117.125 -188.875 ;
        RECT 116.795 -190.565 117.125 -190.235 ;
        RECT 116.795 -191.925 117.125 -191.595 ;
        RECT 116.795 -193.285 117.125 -192.955 ;
        RECT 116.795 -194.645 117.125 -194.315 ;
        RECT 116.795 -196.005 117.125 -195.675 ;
        RECT 116.795 -197.365 117.125 -197.035 ;
        RECT 116.795 -198.725 117.125 -198.395 ;
        RECT 116.795 -200.085 117.125 -199.755 ;
        RECT 116.795 -201.445 117.125 -201.115 ;
        RECT 116.795 -202.805 117.125 -202.475 ;
        RECT 116.795 -204.165 117.125 -203.835 ;
        RECT 116.795 -205.525 117.125 -205.195 ;
        RECT 116.795 -206.885 117.125 -206.555 ;
        RECT 116.795 -208.245 117.125 -207.915 ;
        RECT 116.795 -209.605 117.125 -209.275 ;
        RECT 116.795 -210.965 117.125 -210.635 ;
        RECT 116.795 -212.325 117.125 -211.995 ;
        RECT 116.795 -213.685 117.125 -213.355 ;
        RECT 116.795 -215.045 117.125 -214.715 ;
        RECT 116.795 -216.405 117.125 -216.075 ;
        RECT 116.795 -217.765 117.125 -217.435 ;
        RECT 116.795 -219.125 117.125 -218.795 ;
        RECT 116.795 -220.485 117.125 -220.155 ;
        RECT 116.795 -221.845 117.125 -221.515 ;
        RECT 116.795 -223.205 117.125 -222.875 ;
        RECT 116.795 -224.565 117.125 -224.235 ;
        RECT 116.795 -225.925 117.125 -225.595 ;
        RECT 116.795 -227.285 117.125 -226.955 ;
        RECT 116.795 -228.645 117.125 -228.315 ;
        RECT 116.795 -230.005 117.125 -229.675 ;
        RECT 116.795 -231.365 117.125 -231.035 ;
        RECT 116.795 -232.725 117.125 -232.395 ;
        RECT 116.795 -234.085 117.125 -233.755 ;
        RECT 116.795 -235.445 117.125 -235.115 ;
        RECT 116.795 -236.805 117.125 -236.475 ;
        RECT 116.795 -238.165 117.125 -237.835 ;
        RECT 116.795 -243.81 117.125 -242.68 ;
        RECT 116.8 -243.925 117.12 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 246.76 118.485 247.89 ;
        RECT 118.155 241.915 118.485 242.245 ;
        RECT 118.155 240.555 118.485 240.885 ;
        RECT 118.155 239.195 118.485 239.525 ;
        RECT 118.155 237.835 118.485 238.165 ;
        RECT 118.16 237.16 118.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 -1.525 118.485 -1.195 ;
        RECT 118.155 -2.885 118.485 -2.555 ;
        RECT 118.16 -3.56 118.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 -122.565 118.485 -122.235 ;
        RECT 118.155 -123.925 118.485 -123.595 ;
        RECT 118.155 -125.285 118.485 -124.955 ;
        RECT 118.155 -126.645 118.485 -126.315 ;
        RECT 118.155 -128.005 118.485 -127.675 ;
        RECT 118.155 -129.365 118.485 -129.035 ;
        RECT 118.155 -130.725 118.485 -130.395 ;
        RECT 118.155 -132.085 118.485 -131.755 ;
        RECT 118.155 -133.445 118.485 -133.115 ;
        RECT 118.155 -134.805 118.485 -134.475 ;
        RECT 118.155 -136.165 118.485 -135.835 ;
        RECT 118.155 -137.525 118.485 -137.195 ;
        RECT 118.155 -138.885 118.485 -138.555 ;
        RECT 118.155 -140.245 118.485 -139.915 ;
        RECT 118.155 -141.605 118.485 -141.275 ;
        RECT 118.155 -142.965 118.485 -142.635 ;
        RECT 118.155 -144.325 118.485 -143.995 ;
        RECT 118.155 -145.685 118.485 -145.355 ;
        RECT 118.155 -147.045 118.485 -146.715 ;
        RECT 118.155 -148.405 118.485 -148.075 ;
        RECT 118.155 -149.765 118.485 -149.435 ;
        RECT 118.155 -151.125 118.485 -150.795 ;
        RECT 118.155 -152.485 118.485 -152.155 ;
        RECT 118.155 -153.845 118.485 -153.515 ;
        RECT 118.155 -155.205 118.485 -154.875 ;
        RECT 118.155 -156.565 118.485 -156.235 ;
        RECT 118.155 -157.925 118.485 -157.595 ;
        RECT 118.155 -159.285 118.485 -158.955 ;
        RECT 118.155 -160.645 118.485 -160.315 ;
        RECT 118.155 -162.005 118.485 -161.675 ;
        RECT 118.155 -163.365 118.485 -163.035 ;
        RECT 118.155 -164.725 118.485 -164.395 ;
        RECT 118.155 -166.085 118.485 -165.755 ;
        RECT 118.155 -167.445 118.485 -167.115 ;
        RECT 118.155 -168.805 118.485 -168.475 ;
        RECT 118.155 -170.165 118.485 -169.835 ;
        RECT 118.155 -171.525 118.485 -171.195 ;
        RECT 118.155 -172.885 118.485 -172.555 ;
        RECT 118.155 -174.245 118.485 -173.915 ;
        RECT 118.155 -175.605 118.485 -175.275 ;
        RECT 118.155 -176.965 118.485 -176.635 ;
        RECT 118.155 -178.325 118.485 -177.995 ;
        RECT 118.155 -179.685 118.485 -179.355 ;
        RECT 118.155 -181.045 118.485 -180.715 ;
        RECT 118.155 -182.405 118.485 -182.075 ;
        RECT 118.155 -183.765 118.485 -183.435 ;
        RECT 118.155 -185.125 118.485 -184.795 ;
        RECT 118.155 -186.485 118.485 -186.155 ;
        RECT 118.155 -187.845 118.485 -187.515 ;
        RECT 118.155 -189.205 118.485 -188.875 ;
        RECT 118.155 -190.565 118.485 -190.235 ;
        RECT 118.155 -191.925 118.485 -191.595 ;
        RECT 118.155 -193.285 118.485 -192.955 ;
        RECT 118.155 -194.645 118.485 -194.315 ;
        RECT 118.155 -196.005 118.485 -195.675 ;
        RECT 118.155 -197.365 118.485 -197.035 ;
        RECT 118.155 -198.725 118.485 -198.395 ;
        RECT 118.155 -200.085 118.485 -199.755 ;
        RECT 118.155 -201.445 118.485 -201.115 ;
        RECT 118.155 -202.805 118.485 -202.475 ;
        RECT 118.155 -204.165 118.485 -203.835 ;
        RECT 118.155 -205.525 118.485 -205.195 ;
        RECT 118.155 -206.885 118.485 -206.555 ;
        RECT 118.155 -208.245 118.485 -207.915 ;
        RECT 118.155 -209.605 118.485 -209.275 ;
        RECT 118.155 -210.965 118.485 -210.635 ;
        RECT 118.155 -212.325 118.485 -211.995 ;
        RECT 118.155 -213.685 118.485 -213.355 ;
        RECT 118.155 -215.045 118.485 -214.715 ;
        RECT 118.155 -216.405 118.485 -216.075 ;
        RECT 118.155 -217.765 118.485 -217.435 ;
        RECT 118.155 -219.125 118.485 -218.795 ;
        RECT 118.155 -220.485 118.485 -220.155 ;
        RECT 118.155 -221.845 118.485 -221.515 ;
        RECT 118.155 -223.205 118.485 -222.875 ;
        RECT 118.155 -224.565 118.485 -224.235 ;
        RECT 118.155 -225.925 118.485 -225.595 ;
        RECT 118.155 -227.285 118.485 -226.955 ;
        RECT 118.155 -228.645 118.485 -228.315 ;
        RECT 118.155 -230.005 118.485 -229.675 ;
        RECT 118.155 -231.365 118.485 -231.035 ;
        RECT 118.155 -232.725 118.485 -232.395 ;
        RECT 118.155 -234.085 118.485 -233.755 ;
        RECT 118.155 -235.445 118.485 -235.115 ;
        RECT 118.155 -236.805 118.485 -236.475 ;
        RECT 118.155 -238.165 118.485 -237.835 ;
        RECT 118.155 -243.81 118.485 -242.68 ;
        RECT 118.16 -243.925 118.48 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 246.76 119.845 247.89 ;
        RECT 119.515 241.915 119.845 242.245 ;
        RECT 119.515 240.555 119.845 240.885 ;
        RECT 119.515 239.195 119.845 239.525 ;
        RECT 119.515 237.835 119.845 238.165 ;
        RECT 119.52 237.16 119.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 -1.525 119.845 -1.195 ;
        RECT 119.515 -2.885 119.845 -2.555 ;
        RECT 119.52 -3.56 119.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 -122.565 119.845 -122.235 ;
        RECT 119.515 -123.925 119.845 -123.595 ;
        RECT 119.515 -125.285 119.845 -124.955 ;
        RECT 119.515 -126.645 119.845 -126.315 ;
        RECT 119.515 -128.005 119.845 -127.675 ;
        RECT 119.515 -129.365 119.845 -129.035 ;
        RECT 119.515 -130.725 119.845 -130.395 ;
        RECT 119.515 -132.085 119.845 -131.755 ;
        RECT 119.515 -133.445 119.845 -133.115 ;
        RECT 119.515 -134.805 119.845 -134.475 ;
        RECT 119.515 -136.165 119.845 -135.835 ;
        RECT 119.515 -137.525 119.845 -137.195 ;
        RECT 119.515 -138.885 119.845 -138.555 ;
        RECT 119.515 -140.245 119.845 -139.915 ;
        RECT 119.515 -141.605 119.845 -141.275 ;
        RECT 119.515 -142.965 119.845 -142.635 ;
        RECT 119.515 -144.325 119.845 -143.995 ;
        RECT 119.515 -145.685 119.845 -145.355 ;
        RECT 119.515 -147.045 119.845 -146.715 ;
        RECT 119.515 -148.405 119.845 -148.075 ;
        RECT 119.515 -149.765 119.845 -149.435 ;
        RECT 119.515 -151.125 119.845 -150.795 ;
        RECT 119.515 -152.485 119.845 -152.155 ;
        RECT 119.515 -153.845 119.845 -153.515 ;
        RECT 119.515 -155.205 119.845 -154.875 ;
        RECT 119.515 -156.565 119.845 -156.235 ;
        RECT 119.515 -157.925 119.845 -157.595 ;
        RECT 119.515 -159.285 119.845 -158.955 ;
        RECT 119.515 -160.645 119.845 -160.315 ;
        RECT 119.515 -162.005 119.845 -161.675 ;
        RECT 119.515 -163.365 119.845 -163.035 ;
        RECT 119.515 -164.725 119.845 -164.395 ;
        RECT 119.515 -166.085 119.845 -165.755 ;
        RECT 119.515 -167.445 119.845 -167.115 ;
        RECT 119.515 -168.805 119.845 -168.475 ;
        RECT 119.515 -170.165 119.845 -169.835 ;
        RECT 119.515 -171.525 119.845 -171.195 ;
        RECT 119.515 -172.885 119.845 -172.555 ;
        RECT 119.515 -174.245 119.845 -173.915 ;
        RECT 119.515 -175.605 119.845 -175.275 ;
        RECT 119.515 -176.965 119.845 -176.635 ;
        RECT 119.515 -178.325 119.845 -177.995 ;
        RECT 119.515 -179.685 119.845 -179.355 ;
        RECT 119.515 -181.045 119.845 -180.715 ;
        RECT 119.515 -182.405 119.845 -182.075 ;
        RECT 119.515 -183.765 119.845 -183.435 ;
        RECT 119.515 -185.125 119.845 -184.795 ;
        RECT 119.515 -186.485 119.845 -186.155 ;
        RECT 119.515 -187.845 119.845 -187.515 ;
        RECT 119.515 -189.205 119.845 -188.875 ;
        RECT 119.515 -190.565 119.845 -190.235 ;
        RECT 119.515 -191.925 119.845 -191.595 ;
        RECT 119.515 -193.285 119.845 -192.955 ;
        RECT 119.515 -194.645 119.845 -194.315 ;
        RECT 119.515 -196.005 119.845 -195.675 ;
        RECT 119.515 -197.365 119.845 -197.035 ;
        RECT 119.515 -198.725 119.845 -198.395 ;
        RECT 119.515 -200.085 119.845 -199.755 ;
        RECT 119.515 -201.445 119.845 -201.115 ;
        RECT 119.515 -202.805 119.845 -202.475 ;
        RECT 119.515 -204.165 119.845 -203.835 ;
        RECT 119.515 -205.525 119.845 -205.195 ;
        RECT 119.515 -206.885 119.845 -206.555 ;
        RECT 119.515 -208.245 119.845 -207.915 ;
        RECT 119.515 -209.605 119.845 -209.275 ;
        RECT 119.515 -210.965 119.845 -210.635 ;
        RECT 119.515 -212.325 119.845 -211.995 ;
        RECT 119.515 -213.685 119.845 -213.355 ;
        RECT 119.515 -215.045 119.845 -214.715 ;
        RECT 119.515 -216.405 119.845 -216.075 ;
        RECT 119.515 -217.765 119.845 -217.435 ;
        RECT 119.515 -219.125 119.845 -218.795 ;
        RECT 119.515 -220.485 119.845 -220.155 ;
        RECT 119.515 -221.845 119.845 -221.515 ;
        RECT 119.515 -223.205 119.845 -222.875 ;
        RECT 119.515 -224.565 119.845 -224.235 ;
        RECT 119.515 -225.925 119.845 -225.595 ;
        RECT 119.515 -227.285 119.845 -226.955 ;
        RECT 119.515 -228.645 119.845 -228.315 ;
        RECT 119.515 -230.005 119.845 -229.675 ;
        RECT 119.515 -231.365 119.845 -231.035 ;
        RECT 119.515 -232.725 119.845 -232.395 ;
        RECT 119.515 -234.085 119.845 -233.755 ;
        RECT 119.515 -235.445 119.845 -235.115 ;
        RECT 119.515 -236.805 119.845 -236.475 ;
        RECT 119.515 -238.165 119.845 -237.835 ;
        RECT 119.515 -243.81 119.845 -242.68 ;
        RECT 119.52 -243.925 119.84 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 246.76 121.205 247.89 ;
        RECT 120.875 241.915 121.205 242.245 ;
        RECT 120.875 240.555 121.205 240.885 ;
        RECT 120.875 239.195 121.205 239.525 ;
        RECT 120.875 237.835 121.205 238.165 ;
        RECT 120.88 237.16 121.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 -1.525 121.205 -1.195 ;
        RECT 120.875 -2.885 121.205 -2.555 ;
        RECT 120.88 -3.56 121.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 -122.565 121.205 -122.235 ;
        RECT 120.875 -123.925 121.205 -123.595 ;
        RECT 120.875 -125.285 121.205 -124.955 ;
        RECT 120.875 -126.645 121.205 -126.315 ;
        RECT 120.875 -128.005 121.205 -127.675 ;
        RECT 120.875 -129.365 121.205 -129.035 ;
        RECT 120.875 -130.725 121.205 -130.395 ;
        RECT 120.875 -132.085 121.205 -131.755 ;
        RECT 120.875 -133.445 121.205 -133.115 ;
        RECT 120.875 -134.805 121.205 -134.475 ;
        RECT 120.875 -136.165 121.205 -135.835 ;
        RECT 120.875 -137.525 121.205 -137.195 ;
        RECT 120.875 -138.885 121.205 -138.555 ;
        RECT 120.875 -140.245 121.205 -139.915 ;
        RECT 120.875 -141.605 121.205 -141.275 ;
        RECT 120.875 -142.965 121.205 -142.635 ;
        RECT 120.875 -144.325 121.205 -143.995 ;
        RECT 120.875 -145.685 121.205 -145.355 ;
        RECT 120.875 -147.045 121.205 -146.715 ;
        RECT 120.875 -148.405 121.205 -148.075 ;
        RECT 120.875 -149.765 121.205 -149.435 ;
        RECT 120.875 -151.125 121.205 -150.795 ;
        RECT 120.875 -152.485 121.205 -152.155 ;
        RECT 120.875 -153.845 121.205 -153.515 ;
        RECT 120.875 -155.205 121.205 -154.875 ;
        RECT 120.875 -156.565 121.205 -156.235 ;
        RECT 120.875 -157.925 121.205 -157.595 ;
        RECT 120.875 -159.285 121.205 -158.955 ;
        RECT 120.875 -160.645 121.205 -160.315 ;
        RECT 120.875 -162.005 121.205 -161.675 ;
        RECT 120.875 -163.365 121.205 -163.035 ;
        RECT 120.875 -164.725 121.205 -164.395 ;
        RECT 120.875 -166.085 121.205 -165.755 ;
        RECT 120.875 -167.445 121.205 -167.115 ;
        RECT 120.875 -168.805 121.205 -168.475 ;
        RECT 120.875 -170.165 121.205 -169.835 ;
        RECT 120.875 -171.525 121.205 -171.195 ;
        RECT 120.875 -172.885 121.205 -172.555 ;
        RECT 120.875 -174.245 121.205 -173.915 ;
        RECT 120.875 -175.605 121.205 -175.275 ;
        RECT 120.875 -176.965 121.205 -176.635 ;
        RECT 120.875 -178.325 121.205 -177.995 ;
        RECT 120.875 -179.685 121.205 -179.355 ;
        RECT 120.875 -181.045 121.205 -180.715 ;
        RECT 120.875 -182.405 121.205 -182.075 ;
        RECT 120.875 -183.765 121.205 -183.435 ;
        RECT 120.875 -185.125 121.205 -184.795 ;
        RECT 120.875 -186.485 121.205 -186.155 ;
        RECT 120.875 -187.845 121.205 -187.515 ;
        RECT 120.875 -189.205 121.205 -188.875 ;
        RECT 120.875 -190.565 121.205 -190.235 ;
        RECT 120.875 -191.925 121.205 -191.595 ;
        RECT 120.875 -193.285 121.205 -192.955 ;
        RECT 120.875 -194.645 121.205 -194.315 ;
        RECT 120.875 -196.005 121.205 -195.675 ;
        RECT 120.875 -197.365 121.205 -197.035 ;
        RECT 120.875 -198.725 121.205 -198.395 ;
        RECT 120.875 -200.085 121.205 -199.755 ;
        RECT 120.875 -201.445 121.205 -201.115 ;
        RECT 120.875 -202.805 121.205 -202.475 ;
        RECT 120.875 -204.165 121.205 -203.835 ;
        RECT 120.875 -205.525 121.205 -205.195 ;
        RECT 120.875 -206.885 121.205 -206.555 ;
        RECT 120.875 -208.245 121.205 -207.915 ;
        RECT 120.875 -209.605 121.205 -209.275 ;
        RECT 120.875 -210.965 121.205 -210.635 ;
        RECT 120.875 -212.325 121.205 -211.995 ;
        RECT 120.875 -213.685 121.205 -213.355 ;
        RECT 120.875 -215.045 121.205 -214.715 ;
        RECT 120.875 -216.405 121.205 -216.075 ;
        RECT 120.875 -217.765 121.205 -217.435 ;
        RECT 120.875 -219.125 121.205 -218.795 ;
        RECT 120.875 -220.485 121.205 -220.155 ;
        RECT 120.875 -221.845 121.205 -221.515 ;
        RECT 120.875 -223.205 121.205 -222.875 ;
        RECT 120.875 -224.565 121.205 -224.235 ;
        RECT 120.875 -225.925 121.205 -225.595 ;
        RECT 120.875 -227.285 121.205 -226.955 ;
        RECT 120.875 -228.645 121.205 -228.315 ;
        RECT 120.875 -230.005 121.205 -229.675 ;
        RECT 120.875 -231.365 121.205 -231.035 ;
        RECT 120.875 -232.725 121.205 -232.395 ;
        RECT 120.875 -234.085 121.205 -233.755 ;
        RECT 120.875 -235.445 121.205 -235.115 ;
        RECT 120.875 -236.805 121.205 -236.475 ;
        RECT 120.875 -238.165 121.205 -237.835 ;
        RECT 120.875 -243.81 121.205 -242.68 ;
        RECT 120.88 -243.925 121.2 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 246.76 122.565 247.89 ;
        RECT 122.235 241.915 122.565 242.245 ;
        RECT 122.235 240.555 122.565 240.885 ;
        RECT 122.235 239.195 122.565 239.525 ;
        RECT 122.235 237.835 122.565 238.165 ;
        RECT 122.24 237.16 122.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 -126.645 122.565 -126.315 ;
        RECT 122.235 -128.005 122.565 -127.675 ;
        RECT 122.235 -129.365 122.565 -129.035 ;
        RECT 122.235 -130.725 122.565 -130.395 ;
        RECT 122.235 -132.085 122.565 -131.755 ;
        RECT 122.235 -133.445 122.565 -133.115 ;
        RECT 122.235 -134.805 122.565 -134.475 ;
        RECT 122.235 -136.165 122.565 -135.835 ;
        RECT 122.235 -137.525 122.565 -137.195 ;
        RECT 122.235 -138.885 122.565 -138.555 ;
        RECT 122.235 -140.245 122.565 -139.915 ;
        RECT 122.235 -141.605 122.565 -141.275 ;
        RECT 122.235 -142.965 122.565 -142.635 ;
        RECT 122.235 -144.325 122.565 -143.995 ;
        RECT 122.235 -145.685 122.565 -145.355 ;
        RECT 122.235 -147.045 122.565 -146.715 ;
        RECT 122.235 -148.405 122.565 -148.075 ;
        RECT 122.235 -149.765 122.565 -149.435 ;
        RECT 122.235 -151.125 122.565 -150.795 ;
        RECT 122.235 -152.485 122.565 -152.155 ;
        RECT 122.235 -153.845 122.565 -153.515 ;
        RECT 122.235 -155.205 122.565 -154.875 ;
        RECT 122.235 -156.565 122.565 -156.235 ;
        RECT 122.235 -157.925 122.565 -157.595 ;
        RECT 122.235 -159.285 122.565 -158.955 ;
        RECT 122.235 -160.645 122.565 -160.315 ;
        RECT 122.235 -162.005 122.565 -161.675 ;
        RECT 122.235 -163.365 122.565 -163.035 ;
        RECT 122.235 -164.725 122.565 -164.395 ;
        RECT 122.235 -166.085 122.565 -165.755 ;
        RECT 122.235 -167.445 122.565 -167.115 ;
        RECT 122.235 -168.805 122.565 -168.475 ;
        RECT 122.235 -170.165 122.565 -169.835 ;
        RECT 122.235 -171.525 122.565 -171.195 ;
        RECT 122.235 -172.885 122.565 -172.555 ;
        RECT 122.235 -174.245 122.565 -173.915 ;
        RECT 122.235 -175.605 122.565 -175.275 ;
        RECT 122.235 -176.965 122.565 -176.635 ;
        RECT 122.235 -178.325 122.565 -177.995 ;
        RECT 122.235 -179.685 122.565 -179.355 ;
        RECT 122.235 -181.045 122.565 -180.715 ;
        RECT 122.235 -182.405 122.565 -182.075 ;
        RECT 122.235 -183.765 122.565 -183.435 ;
        RECT 122.235 -185.125 122.565 -184.795 ;
        RECT 122.235 -186.485 122.565 -186.155 ;
        RECT 122.235 -187.845 122.565 -187.515 ;
        RECT 122.235 -189.205 122.565 -188.875 ;
        RECT 122.235 -190.565 122.565 -190.235 ;
        RECT 122.235 -191.925 122.565 -191.595 ;
        RECT 122.235 -193.285 122.565 -192.955 ;
        RECT 122.235 -194.645 122.565 -194.315 ;
        RECT 122.235 -196.005 122.565 -195.675 ;
        RECT 122.235 -197.365 122.565 -197.035 ;
        RECT 122.235 -198.725 122.565 -198.395 ;
        RECT 122.235 -200.085 122.565 -199.755 ;
        RECT 122.235 -201.445 122.565 -201.115 ;
        RECT 122.235 -202.805 122.565 -202.475 ;
        RECT 122.235 -204.165 122.565 -203.835 ;
        RECT 122.235 -205.525 122.565 -205.195 ;
        RECT 122.235 -206.885 122.565 -206.555 ;
        RECT 122.235 -208.245 122.565 -207.915 ;
        RECT 122.235 -209.605 122.565 -209.275 ;
        RECT 122.235 -210.965 122.565 -210.635 ;
        RECT 122.235 -212.325 122.565 -211.995 ;
        RECT 122.235 -213.685 122.565 -213.355 ;
        RECT 122.235 -215.045 122.565 -214.715 ;
        RECT 122.235 -216.405 122.565 -216.075 ;
        RECT 122.235 -217.765 122.565 -217.435 ;
        RECT 122.235 -219.125 122.565 -218.795 ;
        RECT 122.235 -220.485 122.565 -220.155 ;
        RECT 122.235 -221.845 122.565 -221.515 ;
        RECT 122.235 -223.205 122.565 -222.875 ;
        RECT 122.235 -224.565 122.565 -224.235 ;
        RECT 122.235 -225.925 122.565 -225.595 ;
        RECT 122.235 -227.285 122.565 -226.955 ;
        RECT 122.235 -228.645 122.565 -228.315 ;
        RECT 122.235 -230.005 122.565 -229.675 ;
        RECT 122.235 -231.365 122.565 -231.035 ;
        RECT 122.235 -232.725 122.565 -232.395 ;
        RECT 122.235 -234.085 122.565 -233.755 ;
        RECT 122.235 -235.445 122.565 -235.115 ;
        RECT 122.235 -236.805 122.565 -236.475 ;
        RECT 122.235 -238.165 122.565 -237.835 ;
        RECT 122.235 -243.81 122.565 -242.68 ;
        RECT 122.24 -243.925 122.56 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.56 -125.535 122.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 246.76 123.925 247.89 ;
        RECT 123.595 241.915 123.925 242.245 ;
        RECT 123.595 240.555 123.925 240.885 ;
        RECT 123.595 239.195 123.925 239.525 ;
        RECT 123.595 237.835 123.925 238.165 ;
        RECT 123.6 237.16 123.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 246.76 125.285 247.89 ;
        RECT 124.955 241.915 125.285 242.245 ;
        RECT 124.955 240.555 125.285 240.885 ;
        RECT 124.955 239.195 125.285 239.525 ;
        RECT 124.955 237.835 125.285 238.165 ;
        RECT 124.96 237.16 125.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 -1.525 125.285 -1.195 ;
        RECT 124.955 -2.885 125.285 -2.555 ;
        RECT 124.96 -3.56 125.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 246.76 126.645 247.89 ;
        RECT 126.315 241.915 126.645 242.245 ;
        RECT 126.315 240.555 126.645 240.885 ;
        RECT 126.315 239.195 126.645 239.525 ;
        RECT 126.315 237.835 126.645 238.165 ;
        RECT 126.32 237.16 126.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 -1.525 126.645 -1.195 ;
        RECT 126.315 -2.885 126.645 -2.555 ;
        RECT 126.32 -3.56 126.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 -122.565 126.645 -122.235 ;
        RECT 126.315 -123.925 126.645 -123.595 ;
        RECT 126.315 -125.285 126.645 -124.955 ;
        RECT 126.315 -126.645 126.645 -126.315 ;
        RECT 126.315 -128.005 126.645 -127.675 ;
        RECT 126.315 -129.365 126.645 -129.035 ;
        RECT 126.315 -130.725 126.645 -130.395 ;
        RECT 126.315 -132.085 126.645 -131.755 ;
        RECT 126.315 -133.445 126.645 -133.115 ;
        RECT 126.315 -134.805 126.645 -134.475 ;
        RECT 126.315 -136.165 126.645 -135.835 ;
        RECT 126.315 -137.525 126.645 -137.195 ;
        RECT 126.315 -138.885 126.645 -138.555 ;
        RECT 126.315 -140.245 126.645 -139.915 ;
        RECT 126.315 -141.605 126.645 -141.275 ;
        RECT 126.315 -142.965 126.645 -142.635 ;
        RECT 126.315 -144.325 126.645 -143.995 ;
        RECT 126.315 -145.685 126.645 -145.355 ;
        RECT 126.315 -147.045 126.645 -146.715 ;
        RECT 126.315 -148.405 126.645 -148.075 ;
        RECT 126.315 -149.765 126.645 -149.435 ;
        RECT 126.315 -151.125 126.645 -150.795 ;
        RECT 126.315 -152.485 126.645 -152.155 ;
        RECT 126.315 -153.845 126.645 -153.515 ;
        RECT 126.315 -155.205 126.645 -154.875 ;
        RECT 126.315 -156.565 126.645 -156.235 ;
        RECT 126.315 -157.925 126.645 -157.595 ;
        RECT 126.315 -159.285 126.645 -158.955 ;
        RECT 126.315 -160.645 126.645 -160.315 ;
        RECT 126.315 -162.005 126.645 -161.675 ;
        RECT 126.315 -163.365 126.645 -163.035 ;
        RECT 126.315 -164.725 126.645 -164.395 ;
        RECT 126.315 -166.085 126.645 -165.755 ;
        RECT 126.315 -167.445 126.645 -167.115 ;
        RECT 126.315 -168.805 126.645 -168.475 ;
        RECT 126.315 -170.165 126.645 -169.835 ;
        RECT 126.315 -171.525 126.645 -171.195 ;
        RECT 126.315 -172.885 126.645 -172.555 ;
        RECT 126.315 -174.245 126.645 -173.915 ;
        RECT 126.315 -175.605 126.645 -175.275 ;
        RECT 126.315 -176.965 126.645 -176.635 ;
        RECT 126.315 -178.325 126.645 -177.995 ;
        RECT 126.315 -179.685 126.645 -179.355 ;
        RECT 126.315 -181.045 126.645 -180.715 ;
        RECT 126.315 -182.405 126.645 -182.075 ;
        RECT 126.315 -183.765 126.645 -183.435 ;
        RECT 126.315 -185.125 126.645 -184.795 ;
        RECT 126.315 -186.485 126.645 -186.155 ;
        RECT 126.315 -187.845 126.645 -187.515 ;
        RECT 126.315 -189.205 126.645 -188.875 ;
        RECT 126.315 -190.565 126.645 -190.235 ;
        RECT 126.315 -191.925 126.645 -191.595 ;
        RECT 126.315 -193.285 126.645 -192.955 ;
        RECT 126.315 -194.645 126.645 -194.315 ;
        RECT 126.315 -196.005 126.645 -195.675 ;
        RECT 126.315 -197.365 126.645 -197.035 ;
        RECT 126.315 -198.725 126.645 -198.395 ;
        RECT 126.315 -200.085 126.645 -199.755 ;
        RECT 126.315 -201.445 126.645 -201.115 ;
        RECT 126.315 -202.805 126.645 -202.475 ;
        RECT 126.315 -204.165 126.645 -203.835 ;
        RECT 126.315 -205.525 126.645 -205.195 ;
        RECT 126.315 -206.885 126.645 -206.555 ;
        RECT 126.315 -208.245 126.645 -207.915 ;
        RECT 126.315 -209.605 126.645 -209.275 ;
        RECT 126.315 -210.965 126.645 -210.635 ;
        RECT 126.315 -212.325 126.645 -211.995 ;
        RECT 126.315 -213.685 126.645 -213.355 ;
        RECT 126.315 -215.045 126.645 -214.715 ;
        RECT 126.315 -216.405 126.645 -216.075 ;
        RECT 126.315 -217.765 126.645 -217.435 ;
        RECT 126.315 -219.125 126.645 -218.795 ;
        RECT 126.315 -220.485 126.645 -220.155 ;
        RECT 126.315 -221.845 126.645 -221.515 ;
        RECT 126.315 -223.205 126.645 -222.875 ;
        RECT 126.315 -224.565 126.645 -224.235 ;
        RECT 126.315 -225.925 126.645 -225.595 ;
        RECT 126.315 -227.285 126.645 -226.955 ;
        RECT 126.315 -228.645 126.645 -228.315 ;
        RECT 126.315 -230.005 126.645 -229.675 ;
        RECT 126.315 -231.365 126.645 -231.035 ;
        RECT 126.315 -232.725 126.645 -232.395 ;
        RECT 126.315 -234.085 126.645 -233.755 ;
        RECT 126.315 -235.445 126.645 -235.115 ;
        RECT 126.315 -236.805 126.645 -236.475 ;
        RECT 126.315 -238.165 126.645 -237.835 ;
        RECT 126.315 -243.81 126.645 -242.68 ;
        RECT 126.32 -243.925 126.64 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 246.76 128.005 247.89 ;
        RECT 127.675 241.915 128.005 242.245 ;
        RECT 127.675 240.555 128.005 240.885 ;
        RECT 127.675 239.195 128.005 239.525 ;
        RECT 127.675 237.835 128.005 238.165 ;
        RECT 127.68 237.16 128 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 -1.525 128.005 -1.195 ;
        RECT 127.675 -2.885 128.005 -2.555 ;
        RECT 127.68 -3.56 128 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 -122.565 128.005 -122.235 ;
        RECT 127.675 -123.925 128.005 -123.595 ;
        RECT 127.675 -125.285 128.005 -124.955 ;
        RECT 127.675 -126.645 128.005 -126.315 ;
        RECT 127.675 -128.005 128.005 -127.675 ;
        RECT 127.675 -129.365 128.005 -129.035 ;
        RECT 127.675 -130.725 128.005 -130.395 ;
        RECT 127.675 -132.085 128.005 -131.755 ;
        RECT 127.675 -133.445 128.005 -133.115 ;
        RECT 127.675 -134.805 128.005 -134.475 ;
        RECT 127.675 -136.165 128.005 -135.835 ;
        RECT 127.675 -137.525 128.005 -137.195 ;
        RECT 127.675 -138.885 128.005 -138.555 ;
        RECT 127.675 -140.245 128.005 -139.915 ;
        RECT 127.675 -141.605 128.005 -141.275 ;
        RECT 127.675 -142.965 128.005 -142.635 ;
        RECT 127.675 -144.325 128.005 -143.995 ;
        RECT 127.675 -145.685 128.005 -145.355 ;
        RECT 127.675 -147.045 128.005 -146.715 ;
        RECT 127.675 -148.405 128.005 -148.075 ;
        RECT 127.675 -149.765 128.005 -149.435 ;
        RECT 127.675 -151.125 128.005 -150.795 ;
        RECT 127.675 -152.485 128.005 -152.155 ;
        RECT 127.675 -153.845 128.005 -153.515 ;
        RECT 127.675 -155.205 128.005 -154.875 ;
        RECT 127.675 -156.565 128.005 -156.235 ;
        RECT 127.675 -157.925 128.005 -157.595 ;
        RECT 127.675 -159.285 128.005 -158.955 ;
        RECT 127.675 -160.645 128.005 -160.315 ;
        RECT 127.675 -162.005 128.005 -161.675 ;
        RECT 127.675 -163.365 128.005 -163.035 ;
        RECT 127.675 -164.725 128.005 -164.395 ;
        RECT 127.675 -166.085 128.005 -165.755 ;
        RECT 127.675 -167.445 128.005 -167.115 ;
        RECT 127.675 -168.805 128.005 -168.475 ;
        RECT 127.675 -170.165 128.005 -169.835 ;
        RECT 127.675 -171.525 128.005 -171.195 ;
        RECT 127.675 -172.885 128.005 -172.555 ;
        RECT 127.675 -174.245 128.005 -173.915 ;
        RECT 127.675 -175.605 128.005 -175.275 ;
        RECT 127.675 -176.965 128.005 -176.635 ;
        RECT 127.675 -178.325 128.005 -177.995 ;
        RECT 127.675 -179.685 128.005 -179.355 ;
        RECT 127.675 -181.045 128.005 -180.715 ;
        RECT 127.675 -182.405 128.005 -182.075 ;
        RECT 127.675 -183.765 128.005 -183.435 ;
        RECT 127.675 -185.125 128.005 -184.795 ;
        RECT 127.675 -186.485 128.005 -186.155 ;
        RECT 127.675 -187.845 128.005 -187.515 ;
        RECT 127.675 -189.205 128.005 -188.875 ;
        RECT 127.675 -190.565 128.005 -190.235 ;
        RECT 127.675 -191.925 128.005 -191.595 ;
        RECT 127.675 -193.285 128.005 -192.955 ;
        RECT 127.675 -194.645 128.005 -194.315 ;
        RECT 127.675 -196.005 128.005 -195.675 ;
        RECT 127.675 -197.365 128.005 -197.035 ;
        RECT 127.675 -198.725 128.005 -198.395 ;
        RECT 127.675 -200.085 128.005 -199.755 ;
        RECT 127.675 -201.445 128.005 -201.115 ;
        RECT 127.675 -202.805 128.005 -202.475 ;
        RECT 127.675 -204.165 128.005 -203.835 ;
        RECT 127.675 -205.525 128.005 -205.195 ;
        RECT 127.675 -206.885 128.005 -206.555 ;
        RECT 127.675 -208.245 128.005 -207.915 ;
        RECT 127.675 -209.605 128.005 -209.275 ;
        RECT 127.675 -210.965 128.005 -210.635 ;
        RECT 127.675 -212.325 128.005 -211.995 ;
        RECT 127.675 -213.685 128.005 -213.355 ;
        RECT 127.675 -215.045 128.005 -214.715 ;
        RECT 127.675 -216.405 128.005 -216.075 ;
        RECT 127.675 -217.765 128.005 -217.435 ;
        RECT 127.675 -219.125 128.005 -218.795 ;
        RECT 127.675 -220.485 128.005 -220.155 ;
        RECT 127.675 -221.845 128.005 -221.515 ;
        RECT 127.675 -223.205 128.005 -222.875 ;
        RECT 127.675 -224.565 128.005 -224.235 ;
        RECT 127.675 -225.925 128.005 -225.595 ;
        RECT 127.675 -227.285 128.005 -226.955 ;
        RECT 127.675 -228.645 128.005 -228.315 ;
        RECT 127.675 -230.005 128.005 -229.675 ;
        RECT 127.675 -231.365 128.005 -231.035 ;
        RECT 127.675 -232.725 128.005 -232.395 ;
        RECT 127.675 -234.085 128.005 -233.755 ;
        RECT 127.675 -235.445 128.005 -235.115 ;
        RECT 127.675 -236.805 128.005 -236.475 ;
        RECT 127.675 -238.165 128.005 -237.835 ;
        RECT 127.675 -243.81 128.005 -242.68 ;
        RECT 127.68 -243.925 128 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 246.76 129.365 247.89 ;
        RECT 129.035 241.915 129.365 242.245 ;
        RECT 129.035 240.555 129.365 240.885 ;
        RECT 129.035 239.195 129.365 239.525 ;
        RECT 129.035 237.835 129.365 238.165 ;
        RECT 129.04 237.16 129.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -1.525 129.365 -1.195 ;
        RECT 129.035 -2.885 129.365 -2.555 ;
        RECT 129.04 -3.56 129.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -205.525 129.365 -205.195 ;
        RECT 129.035 -206.885 129.365 -206.555 ;
        RECT 129.035 -208.245 129.365 -207.915 ;
        RECT 129.035 -209.605 129.365 -209.275 ;
        RECT 129.035 -210.965 129.365 -210.635 ;
        RECT 129.035 -212.325 129.365 -211.995 ;
        RECT 129.035 -213.685 129.365 -213.355 ;
        RECT 129.035 -215.045 129.365 -214.715 ;
        RECT 129.035 -216.405 129.365 -216.075 ;
        RECT 129.035 -217.765 129.365 -217.435 ;
        RECT 129.035 -219.125 129.365 -218.795 ;
        RECT 129.035 -220.485 129.365 -220.155 ;
        RECT 129.035 -221.845 129.365 -221.515 ;
        RECT 129.035 -223.205 129.365 -222.875 ;
        RECT 129.035 -224.565 129.365 -224.235 ;
        RECT 129.035 -225.925 129.365 -225.595 ;
        RECT 129.035 -227.285 129.365 -226.955 ;
        RECT 129.035 -228.645 129.365 -228.315 ;
        RECT 129.035 -230.005 129.365 -229.675 ;
        RECT 129.035 -231.365 129.365 -231.035 ;
        RECT 129.035 -232.725 129.365 -232.395 ;
        RECT 129.035 -234.085 129.365 -233.755 ;
        RECT 129.035 -235.445 129.365 -235.115 ;
        RECT 129.035 -236.805 129.365 -236.475 ;
        RECT 129.035 -238.165 129.365 -237.835 ;
        RECT 129.035 -243.81 129.365 -242.68 ;
        RECT 129.04 -243.925 129.36 -122.235 ;
        RECT 129.035 -122.565 129.365 -122.235 ;
        RECT 129.035 -123.925 129.365 -123.595 ;
        RECT 129.035 -125.285 129.365 -124.955 ;
        RECT 129.035 -126.645 129.365 -126.315 ;
        RECT 129.035 -128.005 129.365 -127.675 ;
        RECT 129.035 -129.365 129.365 -129.035 ;
        RECT 129.035 -130.725 129.365 -130.395 ;
        RECT 129.035 -132.085 129.365 -131.755 ;
        RECT 129.035 -133.445 129.365 -133.115 ;
        RECT 129.035 -134.805 129.365 -134.475 ;
        RECT 129.035 -136.165 129.365 -135.835 ;
        RECT 129.035 -137.525 129.365 -137.195 ;
        RECT 129.035 -138.885 129.365 -138.555 ;
        RECT 129.035 -140.245 129.365 -139.915 ;
        RECT 129.035 -141.605 129.365 -141.275 ;
        RECT 129.035 -142.965 129.365 -142.635 ;
        RECT 129.035 -144.325 129.365 -143.995 ;
        RECT 129.035 -145.685 129.365 -145.355 ;
        RECT 129.035 -147.045 129.365 -146.715 ;
        RECT 129.035 -148.405 129.365 -148.075 ;
        RECT 129.035 -149.765 129.365 -149.435 ;
        RECT 129.035 -151.125 129.365 -150.795 ;
        RECT 129.035 -152.485 129.365 -152.155 ;
        RECT 129.035 -153.845 129.365 -153.515 ;
        RECT 129.035 -155.205 129.365 -154.875 ;
        RECT 129.035 -156.565 129.365 -156.235 ;
        RECT 129.035 -157.925 129.365 -157.595 ;
        RECT 129.035 -159.285 129.365 -158.955 ;
        RECT 129.035 -160.645 129.365 -160.315 ;
        RECT 129.035 -162.005 129.365 -161.675 ;
        RECT 129.035 -163.365 129.365 -163.035 ;
        RECT 129.035 -164.725 129.365 -164.395 ;
        RECT 129.035 -166.085 129.365 -165.755 ;
        RECT 129.035 -167.445 129.365 -167.115 ;
        RECT 129.035 -168.805 129.365 -168.475 ;
        RECT 129.035 -170.165 129.365 -169.835 ;
        RECT 129.035 -171.525 129.365 -171.195 ;
        RECT 129.035 -172.885 129.365 -172.555 ;
        RECT 129.035 -174.245 129.365 -173.915 ;
        RECT 129.035 -175.605 129.365 -175.275 ;
        RECT 129.035 -176.965 129.365 -176.635 ;
        RECT 129.035 -178.325 129.365 -177.995 ;
        RECT 129.035 -179.685 129.365 -179.355 ;
        RECT 129.035 -181.045 129.365 -180.715 ;
        RECT 129.035 -182.405 129.365 -182.075 ;
        RECT 129.035 -183.765 129.365 -183.435 ;
        RECT 129.035 -185.125 129.365 -184.795 ;
        RECT 129.035 -186.485 129.365 -186.155 ;
        RECT 129.035 -187.845 129.365 -187.515 ;
        RECT 129.035 -189.205 129.365 -188.875 ;
        RECT 129.035 -190.565 129.365 -190.235 ;
        RECT 129.035 -191.925 129.365 -191.595 ;
        RECT 129.035 -193.285 129.365 -192.955 ;
        RECT 129.035 -194.645 129.365 -194.315 ;
        RECT 129.035 -196.005 129.365 -195.675 ;
        RECT 129.035 -197.365 129.365 -197.035 ;
        RECT 129.035 -198.725 129.365 -198.395 ;
        RECT 129.035 -200.085 129.365 -199.755 ;
        RECT 129.035 -201.445 129.365 -201.115 ;
        RECT 129.035 -202.805 129.365 -202.475 ;
        RECT 129.035 -204.165 129.365 -203.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 -1.525 94.005 -1.195 ;
        RECT 93.675 -2.885 94.005 -2.555 ;
        RECT 93.68 -3.56 94 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 -122.565 94.005 -122.235 ;
        RECT 93.675 -123.925 94.005 -123.595 ;
        RECT 93.675 -125.285 94.005 -124.955 ;
        RECT 93.675 -126.645 94.005 -126.315 ;
        RECT 93.675 -128.005 94.005 -127.675 ;
        RECT 93.675 -129.365 94.005 -129.035 ;
        RECT 93.675 -130.725 94.005 -130.395 ;
        RECT 93.675 -132.085 94.005 -131.755 ;
        RECT 93.675 -133.445 94.005 -133.115 ;
        RECT 93.675 -134.805 94.005 -134.475 ;
        RECT 93.675 -136.165 94.005 -135.835 ;
        RECT 93.675 -137.525 94.005 -137.195 ;
        RECT 93.675 -138.885 94.005 -138.555 ;
        RECT 93.675 -140.245 94.005 -139.915 ;
        RECT 93.675 -141.605 94.005 -141.275 ;
        RECT 93.675 -142.965 94.005 -142.635 ;
        RECT 93.675 -144.325 94.005 -143.995 ;
        RECT 93.675 -145.685 94.005 -145.355 ;
        RECT 93.675 -147.045 94.005 -146.715 ;
        RECT 93.675 -148.405 94.005 -148.075 ;
        RECT 93.675 -149.765 94.005 -149.435 ;
        RECT 93.675 -151.125 94.005 -150.795 ;
        RECT 93.675 -152.485 94.005 -152.155 ;
        RECT 93.675 -153.845 94.005 -153.515 ;
        RECT 93.675 -155.205 94.005 -154.875 ;
        RECT 93.675 -156.565 94.005 -156.235 ;
        RECT 93.675 -157.925 94.005 -157.595 ;
        RECT 93.675 -159.285 94.005 -158.955 ;
        RECT 93.675 -160.645 94.005 -160.315 ;
        RECT 93.675 -162.005 94.005 -161.675 ;
        RECT 93.675 -163.365 94.005 -163.035 ;
        RECT 93.675 -164.725 94.005 -164.395 ;
        RECT 93.675 -166.085 94.005 -165.755 ;
        RECT 93.675 -167.445 94.005 -167.115 ;
        RECT 93.675 -168.805 94.005 -168.475 ;
        RECT 93.675 -170.165 94.005 -169.835 ;
        RECT 93.675 -171.525 94.005 -171.195 ;
        RECT 93.675 -172.885 94.005 -172.555 ;
        RECT 93.675 -174.245 94.005 -173.915 ;
        RECT 93.675 -175.605 94.005 -175.275 ;
        RECT 93.675 -176.965 94.005 -176.635 ;
        RECT 93.675 -178.325 94.005 -177.995 ;
        RECT 93.675 -179.685 94.005 -179.355 ;
        RECT 93.675 -181.045 94.005 -180.715 ;
        RECT 93.675 -182.405 94.005 -182.075 ;
        RECT 93.675 -183.765 94.005 -183.435 ;
        RECT 93.675 -185.125 94.005 -184.795 ;
        RECT 93.675 -186.485 94.005 -186.155 ;
        RECT 93.675 -187.845 94.005 -187.515 ;
        RECT 93.675 -189.205 94.005 -188.875 ;
        RECT 93.675 -190.565 94.005 -190.235 ;
        RECT 93.675 -191.925 94.005 -191.595 ;
        RECT 93.675 -193.285 94.005 -192.955 ;
        RECT 93.675 -194.645 94.005 -194.315 ;
        RECT 93.675 -196.005 94.005 -195.675 ;
        RECT 93.675 -197.365 94.005 -197.035 ;
        RECT 93.675 -198.725 94.005 -198.395 ;
        RECT 93.675 -200.085 94.005 -199.755 ;
        RECT 93.675 -201.445 94.005 -201.115 ;
        RECT 93.675 -202.805 94.005 -202.475 ;
        RECT 93.675 -204.165 94.005 -203.835 ;
        RECT 93.675 -205.525 94.005 -205.195 ;
        RECT 93.675 -206.885 94.005 -206.555 ;
        RECT 93.675 -208.245 94.005 -207.915 ;
        RECT 93.675 -209.605 94.005 -209.275 ;
        RECT 93.675 -210.965 94.005 -210.635 ;
        RECT 93.675 -212.325 94.005 -211.995 ;
        RECT 93.675 -213.685 94.005 -213.355 ;
        RECT 93.675 -215.045 94.005 -214.715 ;
        RECT 93.675 -216.405 94.005 -216.075 ;
        RECT 93.675 -217.765 94.005 -217.435 ;
        RECT 93.675 -219.125 94.005 -218.795 ;
        RECT 93.675 -220.485 94.005 -220.155 ;
        RECT 93.675 -221.845 94.005 -221.515 ;
        RECT 93.675 -223.205 94.005 -222.875 ;
        RECT 93.675 -224.565 94.005 -224.235 ;
        RECT 93.675 -225.925 94.005 -225.595 ;
        RECT 93.675 -227.285 94.005 -226.955 ;
        RECT 93.675 -228.645 94.005 -228.315 ;
        RECT 93.675 -230.005 94.005 -229.675 ;
        RECT 93.675 -231.365 94.005 -231.035 ;
        RECT 93.675 -232.725 94.005 -232.395 ;
        RECT 93.675 -234.085 94.005 -233.755 ;
        RECT 93.675 -235.445 94.005 -235.115 ;
        RECT 93.675 -236.805 94.005 -236.475 ;
        RECT 93.675 -238.165 94.005 -237.835 ;
        RECT 93.675 -243.81 94.005 -242.68 ;
        RECT 93.68 -243.925 94 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 246.76 95.365 247.89 ;
        RECT 95.035 241.915 95.365 242.245 ;
        RECT 95.035 240.555 95.365 240.885 ;
        RECT 95.035 239.195 95.365 239.525 ;
        RECT 95.035 237.835 95.365 238.165 ;
        RECT 95.04 237.16 95.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 -1.525 95.365 -1.195 ;
        RECT 95.035 -2.885 95.365 -2.555 ;
        RECT 95.04 -3.56 95.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 -122.565 95.365 -122.235 ;
        RECT 95.035 -123.925 95.365 -123.595 ;
        RECT 95.035 -125.285 95.365 -124.955 ;
        RECT 95.035 -126.645 95.365 -126.315 ;
        RECT 95.035 -128.005 95.365 -127.675 ;
        RECT 95.035 -129.365 95.365 -129.035 ;
        RECT 95.035 -130.725 95.365 -130.395 ;
        RECT 95.035 -132.085 95.365 -131.755 ;
        RECT 95.035 -133.445 95.365 -133.115 ;
        RECT 95.035 -134.805 95.365 -134.475 ;
        RECT 95.035 -136.165 95.365 -135.835 ;
        RECT 95.035 -137.525 95.365 -137.195 ;
        RECT 95.035 -138.885 95.365 -138.555 ;
        RECT 95.035 -140.245 95.365 -139.915 ;
        RECT 95.035 -141.605 95.365 -141.275 ;
        RECT 95.035 -142.965 95.365 -142.635 ;
        RECT 95.035 -144.325 95.365 -143.995 ;
        RECT 95.035 -145.685 95.365 -145.355 ;
        RECT 95.035 -147.045 95.365 -146.715 ;
        RECT 95.035 -148.405 95.365 -148.075 ;
        RECT 95.035 -149.765 95.365 -149.435 ;
        RECT 95.035 -151.125 95.365 -150.795 ;
        RECT 95.035 -152.485 95.365 -152.155 ;
        RECT 95.035 -153.845 95.365 -153.515 ;
        RECT 95.035 -155.205 95.365 -154.875 ;
        RECT 95.035 -156.565 95.365 -156.235 ;
        RECT 95.035 -157.925 95.365 -157.595 ;
        RECT 95.035 -159.285 95.365 -158.955 ;
        RECT 95.035 -160.645 95.365 -160.315 ;
        RECT 95.035 -162.005 95.365 -161.675 ;
        RECT 95.035 -163.365 95.365 -163.035 ;
        RECT 95.035 -164.725 95.365 -164.395 ;
        RECT 95.035 -166.085 95.365 -165.755 ;
        RECT 95.035 -167.445 95.365 -167.115 ;
        RECT 95.035 -168.805 95.365 -168.475 ;
        RECT 95.035 -170.165 95.365 -169.835 ;
        RECT 95.035 -171.525 95.365 -171.195 ;
        RECT 95.035 -172.885 95.365 -172.555 ;
        RECT 95.035 -174.245 95.365 -173.915 ;
        RECT 95.035 -175.605 95.365 -175.275 ;
        RECT 95.035 -176.965 95.365 -176.635 ;
        RECT 95.035 -178.325 95.365 -177.995 ;
        RECT 95.035 -179.685 95.365 -179.355 ;
        RECT 95.035 -181.045 95.365 -180.715 ;
        RECT 95.035 -182.405 95.365 -182.075 ;
        RECT 95.035 -183.765 95.365 -183.435 ;
        RECT 95.035 -185.125 95.365 -184.795 ;
        RECT 95.035 -186.485 95.365 -186.155 ;
        RECT 95.035 -187.845 95.365 -187.515 ;
        RECT 95.035 -189.205 95.365 -188.875 ;
        RECT 95.035 -190.565 95.365 -190.235 ;
        RECT 95.035 -191.925 95.365 -191.595 ;
        RECT 95.035 -193.285 95.365 -192.955 ;
        RECT 95.035 -194.645 95.365 -194.315 ;
        RECT 95.035 -196.005 95.365 -195.675 ;
        RECT 95.035 -197.365 95.365 -197.035 ;
        RECT 95.035 -198.725 95.365 -198.395 ;
        RECT 95.035 -200.085 95.365 -199.755 ;
        RECT 95.035 -201.445 95.365 -201.115 ;
        RECT 95.035 -202.805 95.365 -202.475 ;
        RECT 95.035 -204.165 95.365 -203.835 ;
        RECT 95.035 -205.525 95.365 -205.195 ;
        RECT 95.035 -206.885 95.365 -206.555 ;
        RECT 95.035 -208.245 95.365 -207.915 ;
        RECT 95.035 -209.605 95.365 -209.275 ;
        RECT 95.035 -210.965 95.365 -210.635 ;
        RECT 95.035 -212.325 95.365 -211.995 ;
        RECT 95.035 -213.685 95.365 -213.355 ;
        RECT 95.035 -215.045 95.365 -214.715 ;
        RECT 95.035 -216.405 95.365 -216.075 ;
        RECT 95.035 -217.765 95.365 -217.435 ;
        RECT 95.035 -219.125 95.365 -218.795 ;
        RECT 95.035 -220.485 95.365 -220.155 ;
        RECT 95.035 -221.845 95.365 -221.515 ;
        RECT 95.035 -223.205 95.365 -222.875 ;
        RECT 95.035 -224.565 95.365 -224.235 ;
        RECT 95.035 -225.925 95.365 -225.595 ;
        RECT 95.035 -227.285 95.365 -226.955 ;
        RECT 95.035 -228.645 95.365 -228.315 ;
        RECT 95.035 -230.005 95.365 -229.675 ;
        RECT 95.035 -231.365 95.365 -231.035 ;
        RECT 95.035 -232.725 95.365 -232.395 ;
        RECT 95.035 -234.085 95.365 -233.755 ;
        RECT 95.035 -235.445 95.365 -235.115 ;
        RECT 95.035 -236.805 95.365 -236.475 ;
        RECT 95.035 -238.165 95.365 -237.835 ;
        RECT 95.035 -243.81 95.365 -242.68 ;
        RECT 95.04 -243.925 95.36 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 246.76 96.725 247.89 ;
        RECT 96.395 241.915 96.725 242.245 ;
        RECT 96.395 240.555 96.725 240.885 ;
        RECT 96.395 239.195 96.725 239.525 ;
        RECT 96.395 237.835 96.725 238.165 ;
        RECT 96.4 237.16 96.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -1.525 96.725 -1.195 ;
        RECT 96.395 -2.885 96.725 -2.555 ;
        RECT 96.4 -3.56 96.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -122.565 96.725 -122.235 ;
        RECT 96.395 -123.925 96.725 -123.595 ;
        RECT 96.395 -125.285 96.725 -124.955 ;
        RECT 96.395 -126.645 96.725 -126.315 ;
        RECT 96.395 -128.005 96.725 -127.675 ;
        RECT 96.395 -129.365 96.725 -129.035 ;
        RECT 96.395 -130.725 96.725 -130.395 ;
        RECT 96.395 -132.085 96.725 -131.755 ;
        RECT 96.395 -133.445 96.725 -133.115 ;
        RECT 96.395 -134.805 96.725 -134.475 ;
        RECT 96.395 -136.165 96.725 -135.835 ;
        RECT 96.395 -137.525 96.725 -137.195 ;
        RECT 96.395 -138.885 96.725 -138.555 ;
        RECT 96.395 -140.245 96.725 -139.915 ;
        RECT 96.395 -141.605 96.725 -141.275 ;
        RECT 96.395 -142.965 96.725 -142.635 ;
        RECT 96.395 -144.325 96.725 -143.995 ;
        RECT 96.395 -145.685 96.725 -145.355 ;
        RECT 96.395 -147.045 96.725 -146.715 ;
        RECT 96.395 -148.405 96.725 -148.075 ;
        RECT 96.395 -149.765 96.725 -149.435 ;
        RECT 96.395 -151.125 96.725 -150.795 ;
        RECT 96.395 -152.485 96.725 -152.155 ;
        RECT 96.395 -153.845 96.725 -153.515 ;
        RECT 96.395 -155.205 96.725 -154.875 ;
        RECT 96.395 -156.565 96.725 -156.235 ;
        RECT 96.395 -157.925 96.725 -157.595 ;
        RECT 96.395 -159.285 96.725 -158.955 ;
        RECT 96.395 -160.645 96.725 -160.315 ;
        RECT 96.395 -162.005 96.725 -161.675 ;
        RECT 96.395 -163.365 96.725 -163.035 ;
        RECT 96.395 -164.725 96.725 -164.395 ;
        RECT 96.395 -166.085 96.725 -165.755 ;
        RECT 96.395 -167.445 96.725 -167.115 ;
        RECT 96.395 -168.805 96.725 -168.475 ;
        RECT 96.395 -170.165 96.725 -169.835 ;
        RECT 96.395 -171.525 96.725 -171.195 ;
        RECT 96.395 -172.885 96.725 -172.555 ;
        RECT 96.395 -174.245 96.725 -173.915 ;
        RECT 96.395 -175.605 96.725 -175.275 ;
        RECT 96.395 -176.965 96.725 -176.635 ;
        RECT 96.395 -178.325 96.725 -177.995 ;
        RECT 96.395 -179.685 96.725 -179.355 ;
        RECT 96.395 -181.045 96.725 -180.715 ;
        RECT 96.395 -182.405 96.725 -182.075 ;
        RECT 96.395 -183.765 96.725 -183.435 ;
        RECT 96.395 -185.125 96.725 -184.795 ;
        RECT 96.395 -186.485 96.725 -186.155 ;
        RECT 96.395 -187.845 96.725 -187.515 ;
        RECT 96.395 -189.205 96.725 -188.875 ;
        RECT 96.395 -190.565 96.725 -190.235 ;
        RECT 96.395 -191.925 96.725 -191.595 ;
        RECT 96.395 -193.285 96.725 -192.955 ;
        RECT 96.395 -194.645 96.725 -194.315 ;
        RECT 96.395 -196.005 96.725 -195.675 ;
        RECT 96.395 -197.365 96.725 -197.035 ;
        RECT 96.395 -198.725 96.725 -198.395 ;
        RECT 96.395 -200.085 96.725 -199.755 ;
        RECT 96.395 -201.445 96.725 -201.115 ;
        RECT 96.395 -202.805 96.725 -202.475 ;
        RECT 96.395 -204.165 96.725 -203.835 ;
        RECT 96.395 -205.525 96.725 -205.195 ;
        RECT 96.395 -206.885 96.725 -206.555 ;
        RECT 96.395 -208.245 96.725 -207.915 ;
        RECT 96.395 -209.605 96.725 -209.275 ;
        RECT 96.395 -210.965 96.725 -210.635 ;
        RECT 96.395 -212.325 96.725 -211.995 ;
        RECT 96.395 -213.685 96.725 -213.355 ;
        RECT 96.395 -215.045 96.725 -214.715 ;
        RECT 96.395 -216.405 96.725 -216.075 ;
        RECT 96.395 -217.765 96.725 -217.435 ;
        RECT 96.395 -219.125 96.725 -218.795 ;
        RECT 96.395 -220.485 96.725 -220.155 ;
        RECT 96.395 -221.845 96.725 -221.515 ;
        RECT 96.395 -223.205 96.725 -222.875 ;
        RECT 96.395 -224.565 96.725 -224.235 ;
        RECT 96.395 -225.925 96.725 -225.595 ;
        RECT 96.395 -227.285 96.725 -226.955 ;
        RECT 96.395 -228.645 96.725 -228.315 ;
        RECT 96.395 -230.005 96.725 -229.675 ;
        RECT 96.395 -231.365 96.725 -231.035 ;
        RECT 96.395 -232.725 96.725 -232.395 ;
        RECT 96.395 -234.085 96.725 -233.755 ;
        RECT 96.395 -235.445 96.725 -235.115 ;
        RECT 96.395 -236.805 96.725 -236.475 ;
        RECT 96.395 -238.165 96.725 -237.835 ;
        RECT 96.395 -243.81 96.725 -242.68 ;
        RECT 96.4 -243.925 96.72 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 246.76 98.085 247.89 ;
        RECT 97.755 241.915 98.085 242.245 ;
        RECT 97.755 240.555 98.085 240.885 ;
        RECT 97.755 239.195 98.085 239.525 ;
        RECT 97.755 237.835 98.085 238.165 ;
        RECT 97.76 237.16 98.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 -1.525 98.085 -1.195 ;
        RECT 97.755 -2.885 98.085 -2.555 ;
        RECT 97.76 -3.56 98.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 -122.565 98.085 -122.235 ;
        RECT 97.755 -123.925 98.085 -123.595 ;
        RECT 97.755 -125.285 98.085 -124.955 ;
        RECT 97.755 -126.645 98.085 -126.315 ;
        RECT 97.755 -128.005 98.085 -127.675 ;
        RECT 97.755 -129.365 98.085 -129.035 ;
        RECT 97.755 -130.725 98.085 -130.395 ;
        RECT 97.755 -132.085 98.085 -131.755 ;
        RECT 97.755 -133.445 98.085 -133.115 ;
        RECT 97.755 -134.805 98.085 -134.475 ;
        RECT 97.755 -136.165 98.085 -135.835 ;
        RECT 97.755 -137.525 98.085 -137.195 ;
        RECT 97.755 -138.885 98.085 -138.555 ;
        RECT 97.755 -140.245 98.085 -139.915 ;
        RECT 97.755 -141.605 98.085 -141.275 ;
        RECT 97.755 -142.965 98.085 -142.635 ;
        RECT 97.755 -144.325 98.085 -143.995 ;
        RECT 97.755 -145.685 98.085 -145.355 ;
        RECT 97.755 -147.045 98.085 -146.715 ;
        RECT 97.755 -148.405 98.085 -148.075 ;
        RECT 97.755 -149.765 98.085 -149.435 ;
        RECT 97.755 -151.125 98.085 -150.795 ;
        RECT 97.755 -152.485 98.085 -152.155 ;
        RECT 97.755 -153.845 98.085 -153.515 ;
        RECT 97.755 -155.205 98.085 -154.875 ;
        RECT 97.755 -156.565 98.085 -156.235 ;
        RECT 97.755 -157.925 98.085 -157.595 ;
        RECT 97.755 -159.285 98.085 -158.955 ;
        RECT 97.755 -160.645 98.085 -160.315 ;
        RECT 97.755 -162.005 98.085 -161.675 ;
        RECT 97.755 -163.365 98.085 -163.035 ;
        RECT 97.755 -164.725 98.085 -164.395 ;
        RECT 97.755 -166.085 98.085 -165.755 ;
        RECT 97.755 -167.445 98.085 -167.115 ;
        RECT 97.755 -168.805 98.085 -168.475 ;
        RECT 97.755 -170.165 98.085 -169.835 ;
        RECT 97.755 -171.525 98.085 -171.195 ;
        RECT 97.755 -172.885 98.085 -172.555 ;
        RECT 97.755 -174.245 98.085 -173.915 ;
        RECT 97.755 -175.605 98.085 -175.275 ;
        RECT 97.755 -176.965 98.085 -176.635 ;
        RECT 97.755 -178.325 98.085 -177.995 ;
        RECT 97.755 -179.685 98.085 -179.355 ;
        RECT 97.755 -181.045 98.085 -180.715 ;
        RECT 97.755 -182.405 98.085 -182.075 ;
        RECT 97.755 -183.765 98.085 -183.435 ;
        RECT 97.755 -185.125 98.085 -184.795 ;
        RECT 97.755 -186.485 98.085 -186.155 ;
        RECT 97.755 -187.845 98.085 -187.515 ;
        RECT 97.755 -189.205 98.085 -188.875 ;
        RECT 97.755 -190.565 98.085 -190.235 ;
        RECT 97.755 -191.925 98.085 -191.595 ;
        RECT 97.755 -193.285 98.085 -192.955 ;
        RECT 97.755 -194.645 98.085 -194.315 ;
        RECT 97.755 -196.005 98.085 -195.675 ;
        RECT 97.755 -197.365 98.085 -197.035 ;
        RECT 97.755 -198.725 98.085 -198.395 ;
        RECT 97.755 -200.085 98.085 -199.755 ;
        RECT 97.755 -201.445 98.085 -201.115 ;
        RECT 97.755 -202.805 98.085 -202.475 ;
        RECT 97.755 -204.165 98.085 -203.835 ;
        RECT 97.755 -205.525 98.085 -205.195 ;
        RECT 97.755 -206.885 98.085 -206.555 ;
        RECT 97.755 -208.245 98.085 -207.915 ;
        RECT 97.755 -209.605 98.085 -209.275 ;
        RECT 97.755 -210.965 98.085 -210.635 ;
        RECT 97.755 -212.325 98.085 -211.995 ;
        RECT 97.755 -213.685 98.085 -213.355 ;
        RECT 97.755 -215.045 98.085 -214.715 ;
        RECT 97.755 -216.405 98.085 -216.075 ;
        RECT 97.755 -217.765 98.085 -217.435 ;
        RECT 97.755 -219.125 98.085 -218.795 ;
        RECT 97.755 -220.485 98.085 -220.155 ;
        RECT 97.755 -221.845 98.085 -221.515 ;
        RECT 97.755 -223.205 98.085 -222.875 ;
        RECT 97.755 -224.565 98.085 -224.235 ;
        RECT 97.755 -225.925 98.085 -225.595 ;
        RECT 97.755 -227.285 98.085 -226.955 ;
        RECT 97.755 -228.645 98.085 -228.315 ;
        RECT 97.755 -230.005 98.085 -229.675 ;
        RECT 97.755 -231.365 98.085 -231.035 ;
        RECT 97.755 -232.725 98.085 -232.395 ;
        RECT 97.755 -234.085 98.085 -233.755 ;
        RECT 97.755 -235.445 98.085 -235.115 ;
        RECT 97.755 -236.805 98.085 -236.475 ;
        RECT 97.755 -238.165 98.085 -237.835 ;
        RECT 97.755 -243.81 98.085 -242.68 ;
        RECT 97.76 -243.925 98.08 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 246.76 99.445 247.89 ;
        RECT 99.115 241.915 99.445 242.245 ;
        RECT 99.115 240.555 99.445 240.885 ;
        RECT 99.115 239.195 99.445 239.525 ;
        RECT 99.115 237.835 99.445 238.165 ;
        RECT 99.12 237.16 99.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -1.525 99.445 -1.195 ;
        RECT 99.115 -2.885 99.445 -2.555 ;
        RECT 99.12 -3.56 99.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -122.565 99.445 -122.235 ;
        RECT 99.115 -123.925 99.445 -123.595 ;
        RECT 99.115 -125.285 99.445 -124.955 ;
        RECT 99.115 -126.645 99.445 -126.315 ;
        RECT 99.115 -128.005 99.445 -127.675 ;
        RECT 99.115 -129.365 99.445 -129.035 ;
        RECT 99.115 -130.725 99.445 -130.395 ;
        RECT 99.115 -132.085 99.445 -131.755 ;
        RECT 99.115 -133.445 99.445 -133.115 ;
        RECT 99.115 -134.805 99.445 -134.475 ;
        RECT 99.115 -136.165 99.445 -135.835 ;
        RECT 99.115 -137.525 99.445 -137.195 ;
        RECT 99.115 -138.885 99.445 -138.555 ;
        RECT 99.115 -140.245 99.445 -139.915 ;
        RECT 99.115 -141.605 99.445 -141.275 ;
        RECT 99.115 -142.965 99.445 -142.635 ;
        RECT 99.115 -144.325 99.445 -143.995 ;
        RECT 99.115 -145.685 99.445 -145.355 ;
        RECT 99.115 -147.045 99.445 -146.715 ;
        RECT 99.115 -148.405 99.445 -148.075 ;
        RECT 99.115 -149.765 99.445 -149.435 ;
        RECT 99.115 -151.125 99.445 -150.795 ;
        RECT 99.115 -152.485 99.445 -152.155 ;
        RECT 99.115 -153.845 99.445 -153.515 ;
        RECT 99.115 -155.205 99.445 -154.875 ;
        RECT 99.115 -156.565 99.445 -156.235 ;
        RECT 99.115 -157.925 99.445 -157.595 ;
        RECT 99.115 -159.285 99.445 -158.955 ;
        RECT 99.115 -160.645 99.445 -160.315 ;
        RECT 99.115 -162.005 99.445 -161.675 ;
        RECT 99.115 -163.365 99.445 -163.035 ;
        RECT 99.115 -164.725 99.445 -164.395 ;
        RECT 99.115 -166.085 99.445 -165.755 ;
        RECT 99.115 -167.445 99.445 -167.115 ;
        RECT 99.115 -168.805 99.445 -168.475 ;
        RECT 99.115 -170.165 99.445 -169.835 ;
        RECT 99.115 -171.525 99.445 -171.195 ;
        RECT 99.115 -172.885 99.445 -172.555 ;
        RECT 99.115 -174.245 99.445 -173.915 ;
        RECT 99.115 -175.605 99.445 -175.275 ;
        RECT 99.115 -176.965 99.445 -176.635 ;
        RECT 99.115 -178.325 99.445 -177.995 ;
        RECT 99.115 -179.685 99.445 -179.355 ;
        RECT 99.115 -181.045 99.445 -180.715 ;
        RECT 99.115 -182.405 99.445 -182.075 ;
        RECT 99.115 -183.765 99.445 -183.435 ;
        RECT 99.115 -185.125 99.445 -184.795 ;
        RECT 99.115 -186.485 99.445 -186.155 ;
        RECT 99.115 -187.845 99.445 -187.515 ;
        RECT 99.115 -189.205 99.445 -188.875 ;
        RECT 99.115 -190.565 99.445 -190.235 ;
        RECT 99.115 -191.925 99.445 -191.595 ;
        RECT 99.115 -193.285 99.445 -192.955 ;
        RECT 99.115 -194.645 99.445 -194.315 ;
        RECT 99.115 -196.005 99.445 -195.675 ;
        RECT 99.115 -197.365 99.445 -197.035 ;
        RECT 99.115 -198.725 99.445 -198.395 ;
        RECT 99.115 -200.085 99.445 -199.755 ;
        RECT 99.115 -201.445 99.445 -201.115 ;
        RECT 99.115 -202.805 99.445 -202.475 ;
        RECT 99.115 -204.165 99.445 -203.835 ;
        RECT 99.115 -205.525 99.445 -205.195 ;
        RECT 99.115 -206.885 99.445 -206.555 ;
        RECT 99.115 -208.245 99.445 -207.915 ;
        RECT 99.115 -209.605 99.445 -209.275 ;
        RECT 99.115 -210.965 99.445 -210.635 ;
        RECT 99.115 -212.325 99.445 -211.995 ;
        RECT 99.115 -213.685 99.445 -213.355 ;
        RECT 99.115 -215.045 99.445 -214.715 ;
        RECT 99.115 -216.405 99.445 -216.075 ;
        RECT 99.115 -217.765 99.445 -217.435 ;
        RECT 99.115 -219.125 99.445 -218.795 ;
        RECT 99.115 -220.485 99.445 -220.155 ;
        RECT 99.115 -221.845 99.445 -221.515 ;
        RECT 99.115 -223.205 99.445 -222.875 ;
        RECT 99.115 -224.565 99.445 -224.235 ;
        RECT 99.115 -225.925 99.445 -225.595 ;
        RECT 99.115 -227.285 99.445 -226.955 ;
        RECT 99.115 -228.645 99.445 -228.315 ;
        RECT 99.115 -230.005 99.445 -229.675 ;
        RECT 99.115 -231.365 99.445 -231.035 ;
        RECT 99.115 -232.725 99.445 -232.395 ;
        RECT 99.115 -234.085 99.445 -233.755 ;
        RECT 99.115 -235.445 99.445 -235.115 ;
        RECT 99.115 -236.805 99.445 -236.475 ;
        RECT 99.115 -238.165 99.445 -237.835 ;
        RECT 99.115 -243.81 99.445 -242.68 ;
        RECT 99.12 -243.925 99.44 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 246.76 100.805 247.89 ;
        RECT 100.475 241.915 100.805 242.245 ;
        RECT 100.475 240.555 100.805 240.885 ;
        RECT 100.475 239.195 100.805 239.525 ;
        RECT 100.475 237.835 100.805 238.165 ;
        RECT 100.48 237.16 100.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 -126.645 100.805 -126.315 ;
        RECT 100.475 -128.005 100.805 -127.675 ;
        RECT 100.475 -129.365 100.805 -129.035 ;
        RECT 100.475 -130.725 100.805 -130.395 ;
        RECT 100.475 -132.085 100.805 -131.755 ;
        RECT 100.475 -133.445 100.805 -133.115 ;
        RECT 100.475 -134.805 100.805 -134.475 ;
        RECT 100.475 -136.165 100.805 -135.835 ;
        RECT 100.475 -137.525 100.805 -137.195 ;
        RECT 100.475 -138.885 100.805 -138.555 ;
        RECT 100.475 -140.245 100.805 -139.915 ;
        RECT 100.475 -141.605 100.805 -141.275 ;
        RECT 100.475 -142.965 100.805 -142.635 ;
        RECT 100.475 -144.325 100.805 -143.995 ;
        RECT 100.475 -145.685 100.805 -145.355 ;
        RECT 100.475 -147.045 100.805 -146.715 ;
        RECT 100.475 -148.405 100.805 -148.075 ;
        RECT 100.475 -149.765 100.805 -149.435 ;
        RECT 100.475 -151.125 100.805 -150.795 ;
        RECT 100.475 -152.485 100.805 -152.155 ;
        RECT 100.475 -153.845 100.805 -153.515 ;
        RECT 100.475 -155.205 100.805 -154.875 ;
        RECT 100.475 -156.565 100.805 -156.235 ;
        RECT 100.475 -157.925 100.805 -157.595 ;
        RECT 100.475 -159.285 100.805 -158.955 ;
        RECT 100.475 -160.645 100.805 -160.315 ;
        RECT 100.475 -162.005 100.805 -161.675 ;
        RECT 100.475 -163.365 100.805 -163.035 ;
        RECT 100.475 -164.725 100.805 -164.395 ;
        RECT 100.475 -166.085 100.805 -165.755 ;
        RECT 100.475 -167.445 100.805 -167.115 ;
        RECT 100.475 -168.805 100.805 -168.475 ;
        RECT 100.475 -170.165 100.805 -169.835 ;
        RECT 100.475 -171.525 100.805 -171.195 ;
        RECT 100.475 -172.885 100.805 -172.555 ;
        RECT 100.475 -174.245 100.805 -173.915 ;
        RECT 100.475 -175.605 100.805 -175.275 ;
        RECT 100.475 -176.965 100.805 -176.635 ;
        RECT 100.475 -178.325 100.805 -177.995 ;
        RECT 100.475 -179.685 100.805 -179.355 ;
        RECT 100.475 -181.045 100.805 -180.715 ;
        RECT 100.475 -182.405 100.805 -182.075 ;
        RECT 100.475 -183.765 100.805 -183.435 ;
        RECT 100.475 -185.125 100.805 -184.795 ;
        RECT 100.475 -186.485 100.805 -186.155 ;
        RECT 100.475 -187.845 100.805 -187.515 ;
        RECT 100.475 -189.205 100.805 -188.875 ;
        RECT 100.475 -190.565 100.805 -190.235 ;
        RECT 100.475 -191.925 100.805 -191.595 ;
        RECT 100.475 -193.285 100.805 -192.955 ;
        RECT 100.475 -194.645 100.805 -194.315 ;
        RECT 100.475 -196.005 100.805 -195.675 ;
        RECT 100.475 -197.365 100.805 -197.035 ;
        RECT 100.475 -198.725 100.805 -198.395 ;
        RECT 100.475 -200.085 100.805 -199.755 ;
        RECT 100.475 -201.445 100.805 -201.115 ;
        RECT 100.475 -202.805 100.805 -202.475 ;
        RECT 100.475 -204.165 100.805 -203.835 ;
        RECT 100.475 -205.525 100.805 -205.195 ;
        RECT 100.475 -206.885 100.805 -206.555 ;
        RECT 100.475 -208.245 100.805 -207.915 ;
        RECT 100.475 -209.605 100.805 -209.275 ;
        RECT 100.475 -210.965 100.805 -210.635 ;
        RECT 100.475 -212.325 100.805 -211.995 ;
        RECT 100.475 -213.685 100.805 -213.355 ;
        RECT 100.475 -215.045 100.805 -214.715 ;
        RECT 100.475 -216.405 100.805 -216.075 ;
        RECT 100.475 -217.765 100.805 -217.435 ;
        RECT 100.475 -219.125 100.805 -218.795 ;
        RECT 100.475 -220.485 100.805 -220.155 ;
        RECT 100.475 -221.845 100.805 -221.515 ;
        RECT 100.475 -223.205 100.805 -222.875 ;
        RECT 100.475 -224.565 100.805 -224.235 ;
        RECT 100.475 -225.925 100.805 -225.595 ;
        RECT 100.475 -227.285 100.805 -226.955 ;
        RECT 100.475 -228.645 100.805 -228.315 ;
        RECT 100.475 -230.005 100.805 -229.675 ;
        RECT 100.475 -231.365 100.805 -231.035 ;
        RECT 100.475 -232.725 100.805 -232.395 ;
        RECT 100.475 -234.085 100.805 -233.755 ;
        RECT 100.475 -235.445 100.805 -235.115 ;
        RECT 100.475 -236.805 100.805 -236.475 ;
        RECT 100.475 -238.165 100.805 -237.835 ;
        RECT 100.475 -243.81 100.805 -242.68 ;
        RECT 100.48 -243.925 100.8 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.76 -125.535 101.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 246.76 102.165 247.89 ;
        RECT 101.835 241.915 102.165 242.245 ;
        RECT 101.835 240.555 102.165 240.885 ;
        RECT 101.835 239.195 102.165 239.525 ;
        RECT 101.835 237.835 102.165 238.165 ;
        RECT 101.84 237.16 102.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 246.76 103.525 247.89 ;
        RECT 103.195 241.915 103.525 242.245 ;
        RECT 103.195 240.555 103.525 240.885 ;
        RECT 103.195 239.195 103.525 239.525 ;
        RECT 103.195 237.835 103.525 238.165 ;
        RECT 103.2 237.16 103.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 -1.525 103.525 -1.195 ;
        RECT 103.195 -2.885 103.525 -2.555 ;
        RECT 103.2 -3.56 103.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 246.76 104.885 247.89 ;
        RECT 104.555 241.915 104.885 242.245 ;
        RECT 104.555 240.555 104.885 240.885 ;
        RECT 104.555 239.195 104.885 239.525 ;
        RECT 104.555 237.835 104.885 238.165 ;
        RECT 104.56 237.16 104.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 -1.525 104.885 -1.195 ;
        RECT 104.555 -2.885 104.885 -2.555 ;
        RECT 104.56 -3.56 104.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 -122.565 104.885 -122.235 ;
        RECT 104.555 -123.925 104.885 -123.595 ;
        RECT 104.555 -125.285 104.885 -124.955 ;
        RECT 104.555 -126.645 104.885 -126.315 ;
        RECT 104.555 -128.005 104.885 -127.675 ;
        RECT 104.555 -129.365 104.885 -129.035 ;
        RECT 104.555 -130.725 104.885 -130.395 ;
        RECT 104.555 -132.085 104.885 -131.755 ;
        RECT 104.555 -133.445 104.885 -133.115 ;
        RECT 104.555 -134.805 104.885 -134.475 ;
        RECT 104.555 -136.165 104.885 -135.835 ;
        RECT 104.555 -137.525 104.885 -137.195 ;
        RECT 104.555 -138.885 104.885 -138.555 ;
        RECT 104.555 -140.245 104.885 -139.915 ;
        RECT 104.555 -141.605 104.885 -141.275 ;
        RECT 104.555 -142.965 104.885 -142.635 ;
        RECT 104.555 -144.325 104.885 -143.995 ;
        RECT 104.555 -145.685 104.885 -145.355 ;
        RECT 104.555 -147.045 104.885 -146.715 ;
        RECT 104.555 -148.405 104.885 -148.075 ;
        RECT 104.555 -149.765 104.885 -149.435 ;
        RECT 104.555 -151.125 104.885 -150.795 ;
        RECT 104.555 -152.485 104.885 -152.155 ;
        RECT 104.555 -153.845 104.885 -153.515 ;
        RECT 104.555 -155.205 104.885 -154.875 ;
        RECT 104.555 -156.565 104.885 -156.235 ;
        RECT 104.555 -157.925 104.885 -157.595 ;
        RECT 104.555 -159.285 104.885 -158.955 ;
        RECT 104.555 -160.645 104.885 -160.315 ;
        RECT 104.555 -162.005 104.885 -161.675 ;
        RECT 104.555 -163.365 104.885 -163.035 ;
        RECT 104.555 -164.725 104.885 -164.395 ;
        RECT 104.555 -166.085 104.885 -165.755 ;
        RECT 104.555 -167.445 104.885 -167.115 ;
        RECT 104.555 -168.805 104.885 -168.475 ;
        RECT 104.555 -170.165 104.885 -169.835 ;
        RECT 104.555 -171.525 104.885 -171.195 ;
        RECT 104.555 -172.885 104.885 -172.555 ;
        RECT 104.555 -174.245 104.885 -173.915 ;
        RECT 104.555 -175.605 104.885 -175.275 ;
        RECT 104.555 -176.965 104.885 -176.635 ;
        RECT 104.555 -178.325 104.885 -177.995 ;
        RECT 104.555 -179.685 104.885 -179.355 ;
        RECT 104.555 -181.045 104.885 -180.715 ;
        RECT 104.555 -182.405 104.885 -182.075 ;
        RECT 104.555 -183.765 104.885 -183.435 ;
        RECT 104.555 -185.125 104.885 -184.795 ;
        RECT 104.555 -186.485 104.885 -186.155 ;
        RECT 104.555 -187.845 104.885 -187.515 ;
        RECT 104.555 -189.205 104.885 -188.875 ;
        RECT 104.555 -190.565 104.885 -190.235 ;
        RECT 104.555 -191.925 104.885 -191.595 ;
        RECT 104.555 -193.285 104.885 -192.955 ;
        RECT 104.555 -194.645 104.885 -194.315 ;
        RECT 104.555 -196.005 104.885 -195.675 ;
        RECT 104.555 -197.365 104.885 -197.035 ;
        RECT 104.555 -198.725 104.885 -198.395 ;
        RECT 104.555 -200.085 104.885 -199.755 ;
        RECT 104.555 -201.445 104.885 -201.115 ;
        RECT 104.555 -202.805 104.885 -202.475 ;
        RECT 104.555 -204.165 104.885 -203.835 ;
        RECT 104.555 -205.525 104.885 -205.195 ;
        RECT 104.555 -206.885 104.885 -206.555 ;
        RECT 104.555 -208.245 104.885 -207.915 ;
        RECT 104.555 -209.605 104.885 -209.275 ;
        RECT 104.555 -210.965 104.885 -210.635 ;
        RECT 104.555 -212.325 104.885 -211.995 ;
        RECT 104.555 -213.685 104.885 -213.355 ;
        RECT 104.555 -215.045 104.885 -214.715 ;
        RECT 104.555 -216.405 104.885 -216.075 ;
        RECT 104.555 -217.765 104.885 -217.435 ;
        RECT 104.555 -219.125 104.885 -218.795 ;
        RECT 104.555 -220.485 104.885 -220.155 ;
        RECT 104.555 -221.845 104.885 -221.515 ;
        RECT 104.555 -223.205 104.885 -222.875 ;
        RECT 104.555 -224.565 104.885 -224.235 ;
        RECT 104.555 -225.925 104.885 -225.595 ;
        RECT 104.555 -227.285 104.885 -226.955 ;
        RECT 104.555 -228.645 104.885 -228.315 ;
        RECT 104.555 -230.005 104.885 -229.675 ;
        RECT 104.555 -231.365 104.885 -231.035 ;
        RECT 104.555 -232.725 104.885 -232.395 ;
        RECT 104.555 -234.085 104.885 -233.755 ;
        RECT 104.555 -235.445 104.885 -235.115 ;
        RECT 104.555 -236.805 104.885 -236.475 ;
        RECT 104.555 -238.165 104.885 -237.835 ;
        RECT 104.555 -243.81 104.885 -242.68 ;
        RECT 104.56 -243.925 104.88 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 246.76 106.245 247.89 ;
        RECT 105.915 241.915 106.245 242.245 ;
        RECT 105.915 240.555 106.245 240.885 ;
        RECT 105.915 239.195 106.245 239.525 ;
        RECT 105.915 237.835 106.245 238.165 ;
        RECT 105.92 237.16 106.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 -1.525 106.245 -1.195 ;
        RECT 105.915 -2.885 106.245 -2.555 ;
        RECT 105.92 -3.56 106.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 -122.565 106.245 -122.235 ;
        RECT 105.915 -123.925 106.245 -123.595 ;
        RECT 105.915 -125.285 106.245 -124.955 ;
        RECT 105.915 -126.645 106.245 -126.315 ;
        RECT 105.915 -128.005 106.245 -127.675 ;
        RECT 105.915 -129.365 106.245 -129.035 ;
        RECT 105.915 -130.725 106.245 -130.395 ;
        RECT 105.915 -132.085 106.245 -131.755 ;
        RECT 105.915 -133.445 106.245 -133.115 ;
        RECT 105.915 -134.805 106.245 -134.475 ;
        RECT 105.915 -136.165 106.245 -135.835 ;
        RECT 105.915 -137.525 106.245 -137.195 ;
        RECT 105.915 -138.885 106.245 -138.555 ;
        RECT 105.915 -140.245 106.245 -139.915 ;
        RECT 105.915 -141.605 106.245 -141.275 ;
        RECT 105.915 -142.965 106.245 -142.635 ;
        RECT 105.915 -144.325 106.245 -143.995 ;
        RECT 105.915 -145.685 106.245 -145.355 ;
        RECT 105.915 -147.045 106.245 -146.715 ;
        RECT 105.915 -148.405 106.245 -148.075 ;
        RECT 105.915 -149.765 106.245 -149.435 ;
        RECT 105.915 -151.125 106.245 -150.795 ;
        RECT 105.915 -152.485 106.245 -152.155 ;
        RECT 105.915 -153.845 106.245 -153.515 ;
        RECT 105.915 -155.205 106.245 -154.875 ;
        RECT 105.915 -156.565 106.245 -156.235 ;
        RECT 105.915 -157.925 106.245 -157.595 ;
        RECT 105.915 -159.285 106.245 -158.955 ;
        RECT 105.915 -160.645 106.245 -160.315 ;
        RECT 105.915 -162.005 106.245 -161.675 ;
        RECT 105.915 -163.365 106.245 -163.035 ;
        RECT 105.915 -164.725 106.245 -164.395 ;
        RECT 105.915 -166.085 106.245 -165.755 ;
        RECT 105.915 -167.445 106.245 -167.115 ;
        RECT 105.915 -168.805 106.245 -168.475 ;
        RECT 105.915 -170.165 106.245 -169.835 ;
        RECT 105.915 -171.525 106.245 -171.195 ;
        RECT 105.915 -172.885 106.245 -172.555 ;
        RECT 105.915 -174.245 106.245 -173.915 ;
        RECT 105.915 -175.605 106.245 -175.275 ;
        RECT 105.915 -176.965 106.245 -176.635 ;
        RECT 105.915 -178.325 106.245 -177.995 ;
        RECT 105.915 -179.685 106.245 -179.355 ;
        RECT 105.915 -181.045 106.245 -180.715 ;
        RECT 105.915 -182.405 106.245 -182.075 ;
        RECT 105.915 -183.765 106.245 -183.435 ;
        RECT 105.915 -185.125 106.245 -184.795 ;
        RECT 105.915 -186.485 106.245 -186.155 ;
        RECT 105.915 -187.845 106.245 -187.515 ;
        RECT 105.915 -189.205 106.245 -188.875 ;
        RECT 105.915 -190.565 106.245 -190.235 ;
        RECT 105.915 -191.925 106.245 -191.595 ;
        RECT 105.915 -193.285 106.245 -192.955 ;
        RECT 105.915 -194.645 106.245 -194.315 ;
        RECT 105.915 -196.005 106.245 -195.675 ;
        RECT 105.915 -197.365 106.245 -197.035 ;
        RECT 105.915 -198.725 106.245 -198.395 ;
        RECT 105.915 -200.085 106.245 -199.755 ;
        RECT 105.915 -201.445 106.245 -201.115 ;
        RECT 105.915 -202.805 106.245 -202.475 ;
        RECT 105.915 -204.165 106.245 -203.835 ;
        RECT 105.915 -205.525 106.245 -205.195 ;
        RECT 105.915 -206.885 106.245 -206.555 ;
        RECT 105.915 -208.245 106.245 -207.915 ;
        RECT 105.915 -209.605 106.245 -209.275 ;
        RECT 105.915 -210.965 106.245 -210.635 ;
        RECT 105.915 -212.325 106.245 -211.995 ;
        RECT 105.915 -213.685 106.245 -213.355 ;
        RECT 105.915 -215.045 106.245 -214.715 ;
        RECT 105.915 -216.405 106.245 -216.075 ;
        RECT 105.915 -217.765 106.245 -217.435 ;
        RECT 105.915 -219.125 106.245 -218.795 ;
        RECT 105.915 -220.485 106.245 -220.155 ;
        RECT 105.915 -221.845 106.245 -221.515 ;
        RECT 105.915 -223.205 106.245 -222.875 ;
        RECT 105.915 -224.565 106.245 -224.235 ;
        RECT 105.915 -225.925 106.245 -225.595 ;
        RECT 105.915 -227.285 106.245 -226.955 ;
        RECT 105.915 -228.645 106.245 -228.315 ;
        RECT 105.915 -230.005 106.245 -229.675 ;
        RECT 105.915 -231.365 106.245 -231.035 ;
        RECT 105.915 -232.725 106.245 -232.395 ;
        RECT 105.915 -234.085 106.245 -233.755 ;
        RECT 105.915 -235.445 106.245 -235.115 ;
        RECT 105.915 -236.805 106.245 -236.475 ;
        RECT 105.915 -238.165 106.245 -237.835 ;
        RECT 105.915 -243.81 106.245 -242.68 ;
        RECT 105.92 -243.925 106.24 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 246.76 107.605 247.89 ;
        RECT 107.275 241.915 107.605 242.245 ;
        RECT 107.275 240.555 107.605 240.885 ;
        RECT 107.275 239.195 107.605 239.525 ;
        RECT 107.275 237.835 107.605 238.165 ;
        RECT 107.28 237.16 107.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 -1.525 107.605 -1.195 ;
        RECT 107.275 -2.885 107.605 -2.555 ;
        RECT 107.28 -3.56 107.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 -122.565 107.605 -122.235 ;
        RECT 107.275 -123.925 107.605 -123.595 ;
        RECT 107.275 -125.285 107.605 -124.955 ;
        RECT 107.275 -126.645 107.605 -126.315 ;
        RECT 107.275 -128.005 107.605 -127.675 ;
        RECT 107.275 -129.365 107.605 -129.035 ;
        RECT 107.275 -130.725 107.605 -130.395 ;
        RECT 107.275 -132.085 107.605 -131.755 ;
        RECT 107.275 -133.445 107.605 -133.115 ;
        RECT 107.275 -134.805 107.605 -134.475 ;
        RECT 107.275 -136.165 107.605 -135.835 ;
        RECT 107.275 -137.525 107.605 -137.195 ;
        RECT 107.275 -138.885 107.605 -138.555 ;
        RECT 107.275 -140.245 107.605 -139.915 ;
        RECT 107.275 -141.605 107.605 -141.275 ;
        RECT 107.275 -142.965 107.605 -142.635 ;
        RECT 107.275 -144.325 107.605 -143.995 ;
        RECT 107.275 -145.685 107.605 -145.355 ;
        RECT 107.275 -147.045 107.605 -146.715 ;
        RECT 107.275 -148.405 107.605 -148.075 ;
        RECT 107.275 -149.765 107.605 -149.435 ;
        RECT 107.275 -151.125 107.605 -150.795 ;
        RECT 107.275 -152.485 107.605 -152.155 ;
        RECT 107.275 -153.845 107.605 -153.515 ;
        RECT 107.275 -155.205 107.605 -154.875 ;
        RECT 107.275 -156.565 107.605 -156.235 ;
        RECT 107.275 -157.925 107.605 -157.595 ;
        RECT 107.275 -159.285 107.605 -158.955 ;
        RECT 107.275 -160.645 107.605 -160.315 ;
        RECT 107.275 -162.005 107.605 -161.675 ;
        RECT 107.275 -163.365 107.605 -163.035 ;
        RECT 107.275 -164.725 107.605 -164.395 ;
        RECT 107.275 -166.085 107.605 -165.755 ;
        RECT 107.275 -167.445 107.605 -167.115 ;
        RECT 107.275 -168.805 107.605 -168.475 ;
        RECT 107.275 -170.165 107.605 -169.835 ;
        RECT 107.275 -171.525 107.605 -171.195 ;
        RECT 107.275 -172.885 107.605 -172.555 ;
        RECT 107.275 -174.245 107.605 -173.915 ;
        RECT 107.275 -175.605 107.605 -175.275 ;
        RECT 107.275 -176.965 107.605 -176.635 ;
        RECT 107.275 -178.325 107.605 -177.995 ;
        RECT 107.275 -179.685 107.605 -179.355 ;
        RECT 107.275 -181.045 107.605 -180.715 ;
        RECT 107.275 -182.405 107.605 -182.075 ;
        RECT 107.275 -183.765 107.605 -183.435 ;
        RECT 107.275 -185.125 107.605 -184.795 ;
        RECT 107.275 -186.485 107.605 -186.155 ;
        RECT 107.275 -187.845 107.605 -187.515 ;
        RECT 107.275 -189.205 107.605 -188.875 ;
        RECT 107.275 -190.565 107.605 -190.235 ;
        RECT 107.275 -191.925 107.605 -191.595 ;
        RECT 107.275 -193.285 107.605 -192.955 ;
        RECT 107.275 -194.645 107.605 -194.315 ;
        RECT 107.275 -196.005 107.605 -195.675 ;
        RECT 107.275 -197.365 107.605 -197.035 ;
        RECT 107.275 -198.725 107.605 -198.395 ;
        RECT 107.275 -200.085 107.605 -199.755 ;
        RECT 107.275 -201.445 107.605 -201.115 ;
        RECT 107.275 -202.805 107.605 -202.475 ;
        RECT 107.275 -204.165 107.605 -203.835 ;
        RECT 107.275 -205.525 107.605 -205.195 ;
        RECT 107.275 -206.885 107.605 -206.555 ;
        RECT 107.275 -208.245 107.605 -207.915 ;
        RECT 107.275 -209.605 107.605 -209.275 ;
        RECT 107.275 -210.965 107.605 -210.635 ;
        RECT 107.275 -212.325 107.605 -211.995 ;
        RECT 107.275 -213.685 107.605 -213.355 ;
        RECT 107.275 -215.045 107.605 -214.715 ;
        RECT 107.275 -216.405 107.605 -216.075 ;
        RECT 107.275 -217.765 107.605 -217.435 ;
        RECT 107.275 -219.125 107.605 -218.795 ;
        RECT 107.275 -220.485 107.605 -220.155 ;
        RECT 107.275 -221.845 107.605 -221.515 ;
        RECT 107.275 -223.205 107.605 -222.875 ;
        RECT 107.275 -224.565 107.605 -224.235 ;
        RECT 107.275 -225.925 107.605 -225.595 ;
        RECT 107.275 -227.285 107.605 -226.955 ;
        RECT 107.275 -228.645 107.605 -228.315 ;
        RECT 107.275 -230.005 107.605 -229.675 ;
        RECT 107.275 -231.365 107.605 -231.035 ;
        RECT 107.275 -232.725 107.605 -232.395 ;
        RECT 107.275 -234.085 107.605 -233.755 ;
        RECT 107.275 -235.445 107.605 -235.115 ;
        RECT 107.275 -236.805 107.605 -236.475 ;
        RECT 107.275 -238.165 107.605 -237.835 ;
        RECT 107.275 -243.81 107.605 -242.68 ;
        RECT 107.28 -243.925 107.6 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 246.76 108.965 247.89 ;
        RECT 108.635 241.915 108.965 242.245 ;
        RECT 108.635 240.555 108.965 240.885 ;
        RECT 108.635 239.195 108.965 239.525 ;
        RECT 108.635 237.835 108.965 238.165 ;
        RECT 108.64 237.16 108.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 -1.525 108.965 -1.195 ;
        RECT 108.635 -2.885 108.965 -2.555 ;
        RECT 108.64 -3.56 108.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 -122.565 108.965 -122.235 ;
        RECT 108.635 -123.925 108.965 -123.595 ;
        RECT 108.635 -125.285 108.965 -124.955 ;
        RECT 108.635 -126.645 108.965 -126.315 ;
        RECT 108.635 -128.005 108.965 -127.675 ;
        RECT 108.635 -129.365 108.965 -129.035 ;
        RECT 108.635 -130.725 108.965 -130.395 ;
        RECT 108.635 -132.085 108.965 -131.755 ;
        RECT 108.635 -133.445 108.965 -133.115 ;
        RECT 108.635 -134.805 108.965 -134.475 ;
        RECT 108.635 -136.165 108.965 -135.835 ;
        RECT 108.635 -137.525 108.965 -137.195 ;
        RECT 108.635 -138.885 108.965 -138.555 ;
        RECT 108.635 -140.245 108.965 -139.915 ;
        RECT 108.635 -141.605 108.965 -141.275 ;
        RECT 108.635 -142.965 108.965 -142.635 ;
        RECT 108.635 -144.325 108.965 -143.995 ;
        RECT 108.635 -145.685 108.965 -145.355 ;
        RECT 108.635 -147.045 108.965 -146.715 ;
        RECT 108.635 -148.405 108.965 -148.075 ;
        RECT 108.635 -149.765 108.965 -149.435 ;
        RECT 108.635 -151.125 108.965 -150.795 ;
        RECT 108.635 -152.485 108.965 -152.155 ;
        RECT 108.635 -153.845 108.965 -153.515 ;
        RECT 108.635 -155.205 108.965 -154.875 ;
        RECT 108.635 -156.565 108.965 -156.235 ;
        RECT 108.635 -157.925 108.965 -157.595 ;
        RECT 108.635 -159.285 108.965 -158.955 ;
        RECT 108.635 -160.645 108.965 -160.315 ;
        RECT 108.635 -162.005 108.965 -161.675 ;
        RECT 108.635 -163.365 108.965 -163.035 ;
        RECT 108.635 -164.725 108.965 -164.395 ;
        RECT 108.635 -166.085 108.965 -165.755 ;
        RECT 108.635 -167.445 108.965 -167.115 ;
        RECT 108.635 -168.805 108.965 -168.475 ;
        RECT 108.635 -170.165 108.965 -169.835 ;
        RECT 108.635 -171.525 108.965 -171.195 ;
        RECT 108.635 -172.885 108.965 -172.555 ;
        RECT 108.635 -174.245 108.965 -173.915 ;
        RECT 108.635 -175.605 108.965 -175.275 ;
        RECT 108.635 -176.965 108.965 -176.635 ;
        RECT 108.635 -178.325 108.965 -177.995 ;
        RECT 108.635 -179.685 108.965 -179.355 ;
        RECT 108.635 -181.045 108.965 -180.715 ;
        RECT 108.635 -182.405 108.965 -182.075 ;
        RECT 108.635 -183.765 108.965 -183.435 ;
        RECT 108.635 -185.125 108.965 -184.795 ;
        RECT 108.635 -186.485 108.965 -186.155 ;
        RECT 108.635 -187.845 108.965 -187.515 ;
        RECT 108.635 -189.205 108.965 -188.875 ;
        RECT 108.635 -190.565 108.965 -190.235 ;
        RECT 108.635 -191.925 108.965 -191.595 ;
        RECT 108.635 -193.285 108.965 -192.955 ;
        RECT 108.635 -194.645 108.965 -194.315 ;
        RECT 108.635 -196.005 108.965 -195.675 ;
        RECT 108.635 -197.365 108.965 -197.035 ;
        RECT 108.635 -198.725 108.965 -198.395 ;
        RECT 108.635 -200.085 108.965 -199.755 ;
        RECT 108.635 -201.445 108.965 -201.115 ;
        RECT 108.635 -202.805 108.965 -202.475 ;
        RECT 108.635 -204.165 108.965 -203.835 ;
        RECT 108.635 -205.525 108.965 -205.195 ;
        RECT 108.635 -206.885 108.965 -206.555 ;
        RECT 108.635 -208.245 108.965 -207.915 ;
        RECT 108.635 -209.605 108.965 -209.275 ;
        RECT 108.635 -210.965 108.965 -210.635 ;
        RECT 108.635 -212.325 108.965 -211.995 ;
        RECT 108.635 -213.685 108.965 -213.355 ;
        RECT 108.635 -215.045 108.965 -214.715 ;
        RECT 108.635 -216.405 108.965 -216.075 ;
        RECT 108.635 -217.765 108.965 -217.435 ;
        RECT 108.635 -219.125 108.965 -218.795 ;
        RECT 108.635 -220.485 108.965 -220.155 ;
        RECT 108.635 -221.845 108.965 -221.515 ;
        RECT 108.635 -223.205 108.965 -222.875 ;
        RECT 108.635 -224.565 108.965 -224.235 ;
        RECT 108.635 -225.925 108.965 -225.595 ;
        RECT 108.635 -227.285 108.965 -226.955 ;
        RECT 108.635 -228.645 108.965 -228.315 ;
        RECT 108.635 -230.005 108.965 -229.675 ;
        RECT 108.635 -231.365 108.965 -231.035 ;
        RECT 108.635 -232.725 108.965 -232.395 ;
        RECT 108.635 -234.085 108.965 -233.755 ;
        RECT 108.635 -235.445 108.965 -235.115 ;
        RECT 108.635 -236.805 108.965 -236.475 ;
        RECT 108.635 -238.165 108.965 -237.835 ;
        RECT 108.635 -243.81 108.965 -242.68 ;
        RECT 108.64 -243.925 108.96 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 246.76 110.325 247.89 ;
        RECT 109.995 241.915 110.325 242.245 ;
        RECT 109.995 240.555 110.325 240.885 ;
        RECT 109.995 239.195 110.325 239.525 ;
        RECT 109.995 237.835 110.325 238.165 ;
        RECT 110 237.16 110.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 -1.525 110.325 -1.195 ;
        RECT 109.995 -2.885 110.325 -2.555 ;
        RECT 110 -3.56 110.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 -219.125 110.325 -218.795 ;
        RECT 109.995 -220.485 110.325 -220.155 ;
        RECT 109.995 -221.845 110.325 -221.515 ;
        RECT 109.995 -223.205 110.325 -222.875 ;
        RECT 109.995 -224.565 110.325 -224.235 ;
        RECT 109.995 -225.925 110.325 -225.595 ;
        RECT 109.995 -227.285 110.325 -226.955 ;
        RECT 109.995 -228.645 110.325 -228.315 ;
        RECT 109.995 -230.005 110.325 -229.675 ;
        RECT 109.995 -231.365 110.325 -231.035 ;
        RECT 109.995 -232.725 110.325 -232.395 ;
        RECT 109.995 -234.085 110.325 -233.755 ;
        RECT 109.995 -235.445 110.325 -235.115 ;
        RECT 109.995 -236.805 110.325 -236.475 ;
        RECT 109.995 -238.165 110.325 -237.835 ;
        RECT 109.995 -243.81 110.325 -242.68 ;
        RECT 110 -243.925 110.32 -122.235 ;
        RECT 109.995 -122.565 110.325 -122.235 ;
        RECT 109.995 -123.925 110.325 -123.595 ;
        RECT 109.995 -125.285 110.325 -124.955 ;
        RECT 109.995 -126.645 110.325 -126.315 ;
        RECT 109.995 -128.005 110.325 -127.675 ;
        RECT 109.995 -129.365 110.325 -129.035 ;
        RECT 109.995 -130.725 110.325 -130.395 ;
        RECT 109.995 -132.085 110.325 -131.755 ;
        RECT 109.995 -133.445 110.325 -133.115 ;
        RECT 109.995 -134.805 110.325 -134.475 ;
        RECT 109.995 -136.165 110.325 -135.835 ;
        RECT 109.995 -137.525 110.325 -137.195 ;
        RECT 109.995 -138.885 110.325 -138.555 ;
        RECT 109.995 -140.245 110.325 -139.915 ;
        RECT 109.995 -141.605 110.325 -141.275 ;
        RECT 109.995 -142.965 110.325 -142.635 ;
        RECT 109.995 -144.325 110.325 -143.995 ;
        RECT 109.995 -145.685 110.325 -145.355 ;
        RECT 109.995 -147.045 110.325 -146.715 ;
        RECT 109.995 -148.405 110.325 -148.075 ;
        RECT 109.995 -149.765 110.325 -149.435 ;
        RECT 109.995 -151.125 110.325 -150.795 ;
        RECT 109.995 -152.485 110.325 -152.155 ;
        RECT 109.995 -153.845 110.325 -153.515 ;
        RECT 109.995 -155.205 110.325 -154.875 ;
        RECT 109.995 -156.565 110.325 -156.235 ;
        RECT 109.995 -157.925 110.325 -157.595 ;
        RECT 109.995 -159.285 110.325 -158.955 ;
        RECT 109.995 -160.645 110.325 -160.315 ;
        RECT 109.995 -162.005 110.325 -161.675 ;
        RECT 109.995 -163.365 110.325 -163.035 ;
        RECT 109.995 -164.725 110.325 -164.395 ;
        RECT 109.995 -166.085 110.325 -165.755 ;
        RECT 109.995 -167.445 110.325 -167.115 ;
        RECT 109.995 -168.805 110.325 -168.475 ;
        RECT 109.995 -170.165 110.325 -169.835 ;
        RECT 109.995 -171.525 110.325 -171.195 ;
        RECT 109.995 -172.885 110.325 -172.555 ;
        RECT 109.995 -174.245 110.325 -173.915 ;
        RECT 109.995 -175.605 110.325 -175.275 ;
        RECT 109.995 -176.965 110.325 -176.635 ;
        RECT 109.995 -178.325 110.325 -177.995 ;
        RECT 109.995 -179.685 110.325 -179.355 ;
        RECT 109.995 -181.045 110.325 -180.715 ;
        RECT 109.995 -182.405 110.325 -182.075 ;
        RECT 109.995 -183.765 110.325 -183.435 ;
        RECT 109.995 -185.125 110.325 -184.795 ;
        RECT 109.995 -186.485 110.325 -186.155 ;
        RECT 109.995 -187.845 110.325 -187.515 ;
        RECT 109.995 -189.205 110.325 -188.875 ;
        RECT 109.995 -190.565 110.325 -190.235 ;
        RECT 109.995 -191.925 110.325 -191.595 ;
        RECT 109.995 -193.285 110.325 -192.955 ;
        RECT 109.995 -194.645 110.325 -194.315 ;
        RECT 109.995 -196.005 110.325 -195.675 ;
        RECT 109.995 -197.365 110.325 -197.035 ;
        RECT 109.995 -198.725 110.325 -198.395 ;
        RECT 109.995 -200.085 110.325 -199.755 ;
        RECT 109.995 -201.445 110.325 -201.115 ;
        RECT 109.995 -202.805 110.325 -202.475 ;
        RECT 109.995 -204.165 110.325 -203.835 ;
        RECT 109.995 -205.525 110.325 -205.195 ;
        RECT 109.995 -206.885 110.325 -206.555 ;
        RECT 109.995 -208.245 110.325 -207.915 ;
        RECT 109.995 -209.605 110.325 -209.275 ;
        RECT 109.995 -210.965 110.325 -210.635 ;
        RECT 109.995 -212.325 110.325 -211.995 ;
        RECT 109.995 -213.685 110.325 -213.355 ;
        RECT 109.995 -215.045 110.325 -214.715 ;
        RECT 109.995 -216.405 110.325 -216.075 ;
        RECT 109.995 -217.765 110.325 -217.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 246.76 74.965 247.89 ;
        RECT 74.635 241.915 74.965 242.245 ;
        RECT 74.635 240.555 74.965 240.885 ;
        RECT 74.635 239.195 74.965 239.525 ;
        RECT 74.635 237.835 74.965 238.165 ;
        RECT 74.64 237.16 74.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -1.525 74.965 -1.195 ;
        RECT 74.635 -2.885 74.965 -2.555 ;
        RECT 74.64 -3.56 74.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -122.565 74.965 -122.235 ;
        RECT 74.635 -123.925 74.965 -123.595 ;
        RECT 74.635 -125.285 74.965 -124.955 ;
        RECT 74.635 -126.645 74.965 -126.315 ;
        RECT 74.635 -128.005 74.965 -127.675 ;
        RECT 74.635 -129.365 74.965 -129.035 ;
        RECT 74.635 -130.725 74.965 -130.395 ;
        RECT 74.635 -132.085 74.965 -131.755 ;
        RECT 74.635 -133.445 74.965 -133.115 ;
        RECT 74.635 -134.805 74.965 -134.475 ;
        RECT 74.635 -136.165 74.965 -135.835 ;
        RECT 74.635 -137.525 74.965 -137.195 ;
        RECT 74.635 -138.885 74.965 -138.555 ;
        RECT 74.635 -140.245 74.965 -139.915 ;
        RECT 74.635 -141.605 74.965 -141.275 ;
        RECT 74.635 -142.965 74.965 -142.635 ;
        RECT 74.635 -144.325 74.965 -143.995 ;
        RECT 74.635 -145.685 74.965 -145.355 ;
        RECT 74.635 -147.045 74.965 -146.715 ;
        RECT 74.635 -148.405 74.965 -148.075 ;
        RECT 74.635 -149.765 74.965 -149.435 ;
        RECT 74.635 -151.125 74.965 -150.795 ;
        RECT 74.635 -152.485 74.965 -152.155 ;
        RECT 74.635 -153.845 74.965 -153.515 ;
        RECT 74.635 -155.205 74.965 -154.875 ;
        RECT 74.635 -156.565 74.965 -156.235 ;
        RECT 74.635 -157.925 74.965 -157.595 ;
        RECT 74.635 -159.285 74.965 -158.955 ;
        RECT 74.635 -160.645 74.965 -160.315 ;
        RECT 74.635 -162.005 74.965 -161.675 ;
        RECT 74.635 -163.365 74.965 -163.035 ;
        RECT 74.635 -164.725 74.965 -164.395 ;
        RECT 74.635 -166.085 74.965 -165.755 ;
        RECT 74.635 -167.445 74.965 -167.115 ;
        RECT 74.635 -168.805 74.965 -168.475 ;
        RECT 74.635 -170.165 74.965 -169.835 ;
        RECT 74.635 -171.525 74.965 -171.195 ;
        RECT 74.635 -172.885 74.965 -172.555 ;
        RECT 74.635 -174.245 74.965 -173.915 ;
        RECT 74.635 -175.605 74.965 -175.275 ;
        RECT 74.635 -176.965 74.965 -176.635 ;
        RECT 74.635 -178.325 74.965 -177.995 ;
        RECT 74.635 -179.685 74.965 -179.355 ;
        RECT 74.635 -181.045 74.965 -180.715 ;
        RECT 74.635 -182.405 74.965 -182.075 ;
        RECT 74.635 -183.765 74.965 -183.435 ;
        RECT 74.635 -185.125 74.965 -184.795 ;
        RECT 74.635 -186.485 74.965 -186.155 ;
        RECT 74.635 -187.845 74.965 -187.515 ;
        RECT 74.635 -189.205 74.965 -188.875 ;
        RECT 74.635 -190.565 74.965 -190.235 ;
        RECT 74.635 -191.925 74.965 -191.595 ;
        RECT 74.635 -193.285 74.965 -192.955 ;
        RECT 74.635 -194.645 74.965 -194.315 ;
        RECT 74.635 -196.005 74.965 -195.675 ;
        RECT 74.635 -197.365 74.965 -197.035 ;
        RECT 74.635 -198.725 74.965 -198.395 ;
        RECT 74.635 -200.085 74.965 -199.755 ;
        RECT 74.635 -201.445 74.965 -201.115 ;
        RECT 74.635 -202.805 74.965 -202.475 ;
        RECT 74.635 -204.165 74.965 -203.835 ;
        RECT 74.635 -205.525 74.965 -205.195 ;
        RECT 74.635 -206.885 74.965 -206.555 ;
        RECT 74.635 -208.245 74.965 -207.915 ;
        RECT 74.635 -209.605 74.965 -209.275 ;
        RECT 74.635 -210.965 74.965 -210.635 ;
        RECT 74.635 -212.325 74.965 -211.995 ;
        RECT 74.635 -213.685 74.965 -213.355 ;
        RECT 74.635 -215.045 74.965 -214.715 ;
        RECT 74.635 -216.405 74.965 -216.075 ;
        RECT 74.635 -217.765 74.965 -217.435 ;
        RECT 74.635 -219.125 74.965 -218.795 ;
        RECT 74.635 -220.485 74.965 -220.155 ;
        RECT 74.635 -221.845 74.965 -221.515 ;
        RECT 74.635 -223.205 74.965 -222.875 ;
        RECT 74.635 -224.565 74.965 -224.235 ;
        RECT 74.635 -225.925 74.965 -225.595 ;
        RECT 74.635 -227.285 74.965 -226.955 ;
        RECT 74.635 -228.645 74.965 -228.315 ;
        RECT 74.635 -230.005 74.965 -229.675 ;
        RECT 74.635 -231.365 74.965 -231.035 ;
        RECT 74.635 -232.725 74.965 -232.395 ;
        RECT 74.635 -234.085 74.965 -233.755 ;
        RECT 74.635 -235.445 74.965 -235.115 ;
        RECT 74.635 -236.805 74.965 -236.475 ;
        RECT 74.635 -238.165 74.965 -237.835 ;
        RECT 74.635 -243.81 74.965 -242.68 ;
        RECT 74.64 -243.925 74.96 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 246.76 76.325 247.89 ;
        RECT 75.995 241.915 76.325 242.245 ;
        RECT 75.995 240.555 76.325 240.885 ;
        RECT 75.995 239.195 76.325 239.525 ;
        RECT 75.995 237.835 76.325 238.165 ;
        RECT 76 237.16 76.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 -1.525 76.325 -1.195 ;
        RECT 75.995 -2.885 76.325 -2.555 ;
        RECT 76 -3.56 76.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 -122.565 76.325 -122.235 ;
        RECT 75.995 -123.925 76.325 -123.595 ;
        RECT 75.995 -125.285 76.325 -124.955 ;
        RECT 75.995 -126.645 76.325 -126.315 ;
        RECT 75.995 -128.005 76.325 -127.675 ;
        RECT 75.995 -129.365 76.325 -129.035 ;
        RECT 75.995 -130.725 76.325 -130.395 ;
        RECT 75.995 -132.085 76.325 -131.755 ;
        RECT 75.995 -133.445 76.325 -133.115 ;
        RECT 75.995 -134.805 76.325 -134.475 ;
        RECT 75.995 -136.165 76.325 -135.835 ;
        RECT 75.995 -137.525 76.325 -137.195 ;
        RECT 75.995 -138.885 76.325 -138.555 ;
        RECT 75.995 -140.245 76.325 -139.915 ;
        RECT 75.995 -141.605 76.325 -141.275 ;
        RECT 75.995 -142.965 76.325 -142.635 ;
        RECT 75.995 -144.325 76.325 -143.995 ;
        RECT 75.995 -145.685 76.325 -145.355 ;
        RECT 75.995 -147.045 76.325 -146.715 ;
        RECT 75.995 -148.405 76.325 -148.075 ;
        RECT 75.995 -149.765 76.325 -149.435 ;
        RECT 75.995 -151.125 76.325 -150.795 ;
        RECT 75.995 -152.485 76.325 -152.155 ;
        RECT 75.995 -153.845 76.325 -153.515 ;
        RECT 75.995 -155.205 76.325 -154.875 ;
        RECT 75.995 -156.565 76.325 -156.235 ;
        RECT 75.995 -157.925 76.325 -157.595 ;
        RECT 75.995 -159.285 76.325 -158.955 ;
        RECT 75.995 -160.645 76.325 -160.315 ;
        RECT 75.995 -162.005 76.325 -161.675 ;
        RECT 75.995 -163.365 76.325 -163.035 ;
        RECT 75.995 -164.725 76.325 -164.395 ;
        RECT 75.995 -166.085 76.325 -165.755 ;
        RECT 75.995 -167.445 76.325 -167.115 ;
        RECT 75.995 -168.805 76.325 -168.475 ;
        RECT 75.995 -170.165 76.325 -169.835 ;
        RECT 75.995 -171.525 76.325 -171.195 ;
        RECT 75.995 -172.885 76.325 -172.555 ;
        RECT 75.995 -174.245 76.325 -173.915 ;
        RECT 75.995 -175.605 76.325 -175.275 ;
        RECT 75.995 -176.965 76.325 -176.635 ;
        RECT 75.995 -178.325 76.325 -177.995 ;
        RECT 75.995 -179.685 76.325 -179.355 ;
        RECT 75.995 -181.045 76.325 -180.715 ;
        RECT 75.995 -182.405 76.325 -182.075 ;
        RECT 75.995 -183.765 76.325 -183.435 ;
        RECT 75.995 -185.125 76.325 -184.795 ;
        RECT 75.995 -186.485 76.325 -186.155 ;
        RECT 75.995 -187.845 76.325 -187.515 ;
        RECT 75.995 -189.205 76.325 -188.875 ;
        RECT 75.995 -190.565 76.325 -190.235 ;
        RECT 75.995 -191.925 76.325 -191.595 ;
        RECT 75.995 -193.285 76.325 -192.955 ;
        RECT 75.995 -194.645 76.325 -194.315 ;
        RECT 75.995 -196.005 76.325 -195.675 ;
        RECT 75.995 -197.365 76.325 -197.035 ;
        RECT 75.995 -198.725 76.325 -198.395 ;
        RECT 75.995 -200.085 76.325 -199.755 ;
        RECT 75.995 -201.445 76.325 -201.115 ;
        RECT 75.995 -202.805 76.325 -202.475 ;
        RECT 75.995 -204.165 76.325 -203.835 ;
        RECT 75.995 -205.525 76.325 -205.195 ;
        RECT 75.995 -206.885 76.325 -206.555 ;
        RECT 75.995 -208.245 76.325 -207.915 ;
        RECT 75.995 -209.605 76.325 -209.275 ;
        RECT 75.995 -210.965 76.325 -210.635 ;
        RECT 75.995 -212.325 76.325 -211.995 ;
        RECT 75.995 -213.685 76.325 -213.355 ;
        RECT 75.995 -215.045 76.325 -214.715 ;
        RECT 75.995 -216.405 76.325 -216.075 ;
        RECT 75.995 -217.765 76.325 -217.435 ;
        RECT 75.995 -219.125 76.325 -218.795 ;
        RECT 75.995 -220.485 76.325 -220.155 ;
        RECT 75.995 -221.845 76.325 -221.515 ;
        RECT 75.995 -223.205 76.325 -222.875 ;
        RECT 75.995 -224.565 76.325 -224.235 ;
        RECT 75.995 -225.925 76.325 -225.595 ;
        RECT 75.995 -227.285 76.325 -226.955 ;
        RECT 75.995 -228.645 76.325 -228.315 ;
        RECT 75.995 -230.005 76.325 -229.675 ;
        RECT 75.995 -231.365 76.325 -231.035 ;
        RECT 75.995 -232.725 76.325 -232.395 ;
        RECT 75.995 -234.085 76.325 -233.755 ;
        RECT 75.995 -235.445 76.325 -235.115 ;
        RECT 75.995 -236.805 76.325 -236.475 ;
        RECT 75.995 -238.165 76.325 -237.835 ;
        RECT 75.995 -243.81 76.325 -242.68 ;
        RECT 76 -243.925 76.32 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 246.76 77.685 247.89 ;
        RECT 77.355 241.915 77.685 242.245 ;
        RECT 77.355 240.555 77.685 240.885 ;
        RECT 77.355 239.195 77.685 239.525 ;
        RECT 77.355 237.835 77.685 238.165 ;
        RECT 77.36 237.16 77.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 -1.525 77.685 -1.195 ;
        RECT 77.355 -2.885 77.685 -2.555 ;
        RECT 77.36 -3.56 77.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 -122.565 77.685 -122.235 ;
        RECT 77.355 -123.925 77.685 -123.595 ;
        RECT 77.355 -125.285 77.685 -124.955 ;
        RECT 77.355 -126.645 77.685 -126.315 ;
        RECT 77.355 -128.005 77.685 -127.675 ;
        RECT 77.355 -129.365 77.685 -129.035 ;
        RECT 77.355 -130.725 77.685 -130.395 ;
        RECT 77.355 -132.085 77.685 -131.755 ;
        RECT 77.355 -133.445 77.685 -133.115 ;
        RECT 77.355 -134.805 77.685 -134.475 ;
        RECT 77.355 -136.165 77.685 -135.835 ;
        RECT 77.355 -137.525 77.685 -137.195 ;
        RECT 77.355 -138.885 77.685 -138.555 ;
        RECT 77.355 -140.245 77.685 -139.915 ;
        RECT 77.355 -141.605 77.685 -141.275 ;
        RECT 77.355 -142.965 77.685 -142.635 ;
        RECT 77.355 -144.325 77.685 -143.995 ;
        RECT 77.355 -145.685 77.685 -145.355 ;
        RECT 77.355 -147.045 77.685 -146.715 ;
        RECT 77.355 -148.405 77.685 -148.075 ;
        RECT 77.355 -149.765 77.685 -149.435 ;
        RECT 77.355 -151.125 77.685 -150.795 ;
        RECT 77.355 -152.485 77.685 -152.155 ;
        RECT 77.355 -153.845 77.685 -153.515 ;
        RECT 77.355 -155.205 77.685 -154.875 ;
        RECT 77.355 -156.565 77.685 -156.235 ;
        RECT 77.355 -157.925 77.685 -157.595 ;
        RECT 77.355 -159.285 77.685 -158.955 ;
        RECT 77.355 -160.645 77.685 -160.315 ;
        RECT 77.355 -162.005 77.685 -161.675 ;
        RECT 77.355 -163.365 77.685 -163.035 ;
        RECT 77.355 -164.725 77.685 -164.395 ;
        RECT 77.355 -166.085 77.685 -165.755 ;
        RECT 77.355 -167.445 77.685 -167.115 ;
        RECT 77.355 -168.805 77.685 -168.475 ;
        RECT 77.355 -170.165 77.685 -169.835 ;
        RECT 77.355 -171.525 77.685 -171.195 ;
        RECT 77.355 -172.885 77.685 -172.555 ;
        RECT 77.355 -174.245 77.685 -173.915 ;
        RECT 77.355 -175.605 77.685 -175.275 ;
        RECT 77.355 -176.965 77.685 -176.635 ;
        RECT 77.355 -178.325 77.685 -177.995 ;
        RECT 77.355 -179.685 77.685 -179.355 ;
        RECT 77.355 -181.045 77.685 -180.715 ;
        RECT 77.355 -182.405 77.685 -182.075 ;
        RECT 77.355 -183.765 77.685 -183.435 ;
        RECT 77.355 -185.125 77.685 -184.795 ;
        RECT 77.355 -186.485 77.685 -186.155 ;
        RECT 77.355 -187.845 77.685 -187.515 ;
        RECT 77.355 -189.205 77.685 -188.875 ;
        RECT 77.355 -190.565 77.685 -190.235 ;
        RECT 77.355 -191.925 77.685 -191.595 ;
        RECT 77.355 -193.285 77.685 -192.955 ;
        RECT 77.355 -194.645 77.685 -194.315 ;
        RECT 77.355 -196.005 77.685 -195.675 ;
        RECT 77.355 -197.365 77.685 -197.035 ;
        RECT 77.355 -198.725 77.685 -198.395 ;
        RECT 77.355 -200.085 77.685 -199.755 ;
        RECT 77.355 -201.445 77.685 -201.115 ;
        RECT 77.355 -202.805 77.685 -202.475 ;
        RECT 77.355 -204.165 77.685 -203.835 ;
        RECT 77.355 -205.525 77.685 -205.195 ;
        RECT 77.355 -206.885 77.685 -206.555 ;
        RECT 77.355 -208.245 77.685 -207.915 ;
        RECT 77.355 -209.605 77.685 -209.275 ;
        RECT 77.355 -210.965 77.685 -210.635 ;
        RECT 77.355 -212.325 77.685 -211.995 ;
        RECT 77.355 -213.685 77.685 -213.355 ;
        RECT 77.355 -215.045 77.685 -214.715 ;
        RECT 77.355 -216.405 77.685 -216.075 ;
        RECT 77.355 -217.765 77.685 -217.435 ;
        RECT 77.355 -219.125 77.685 -218.795 ;
        RECT 77.355 -220.485 77.685 -220.155 ;
        RECT 77.355 -221.845 77.685 -221.515 ;
        RECT 77.355 -223.205 77.685 -222.875 ;
        RECT 77.355 -224.565 77.685 -224.235 ;
        RECT 77.355 -225.925 77.685 -225.595 ;
        RECT 77.355 -227.285 77.685 -226.955 ;
        RECT 77.355 -228.645 77.685 -228.315 ;
        RECT 77.355 -230.005 77.685 -229.675 ;
        RECT 77.355 -231.365 77.685 -231.035 ;
        RECT 77.355 -232.725 77.685 -232.395 ;
        RECT 77.355 -234.085 77.685 -233.755 ;
        RECT 77.355 -235.445 77.685 -235.115 ;
        RECT 77.355 -236.805 77.685 -236.475 ;
        RECT 77.355 -238.165 77.685 -237.835 ;
        RECT 77.355 -243.81 77.685 -242.68 ;
        RECT 77.36 -243.925 77.68 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 246.76 79.045 247.89 ;
        RECT 78.715 241.915 79.045 242.245 ;
        RECT 78.715 240.555 79.045 240.885 ;
        RECT 78.715 239.195 79.045 239.525 ;
        RECT 78.715 237.835 79.045 238.165 ;
        RECT 78.72 237.16 79.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 -126.645 79.045 -126.315 ;
        RECT 78.715 -128.005 79.045 -127.675 ;
        RECT 78.715 -129.365 79.045 -129.035 ;
        RECT 78.715 -130.725 79.045 -130.395 ;
        RECT 78.715 -132.085 79.045 -131.755 ;
        RECT 78.715 -133.445 79.045 -133.115 ;
        RECT 78.715 -134.805 79.045 -134.475 ;
        RECT 78.715 -136.165 79.045 -135.835 ;
        RECT 78.715 -137.525 79.045 -137.195 ;
        RECT 78.715 -138.885 79.045 -138.555 ;
        RECT 78.715 -140.245 79.045 -139.915 ;
        RECT 78.715 -141.605 79.045 -141.275 ;
        RECT 78.715 -142.965 79.045 -142.635 ;
        RECT 78.715 -144.325 79.045 -143.995 ;
        RECT 78.715 -145.685 79.045 -145.355 ;
        RECT 78.715 -147.045 79.045 -146.715 ;
        RECT 78.715 -148.405 79.045 -148.075 ;
        RECT 78.715 -149.765 79.045 -149.435 ;
        RECT 78.715 -151.125 79.045 -150.795 ;
        RECT 78.715 -152.485 79.045 -152.155 ;
        RECT 78.715 -153.845 79.045 -153.515 ;
        RECT 78.715 -155.205 79.045 -154.875 ;
        RECT 78.715 -156.565 79.045 -156.235 ;
        RECT 78.715 -157.925 79.045 -157.595 ;
        RECT 78.715 -159.285 79.045 -158.955 ;
        RECT 78.715 -160.645 79.045 -160.315 ;
        RECT 78.715 -162.005 79.045 -161.675 ;
        RECT 78.715 -163.365 79.045 -163.035 ;
        RECT 78.715 -164.725 79.045 -164.395 ;
        RECT 78.715 -166.085 79.045 -165.755 ;
        RECT 78.715 -167.445 79.045 -167.115 ;
        RECT 78.715 -168.805 79.045 -168.475 ;
        RECT 78.715 -170.165 79.045 -169.835 ;
        RECT 78.715 -171.525 79.045 -171.195 ;
        RECT 78.715 -172.885 79.045 -172.555 ;
        RECT 78.715 -174.245 79.045 -173.915 ;
        RECT 78.715 -175.605 79.045 -175.275 ;
        RECT 78.715 -176.965 79.045 -176.635 ;
        RECT 78.715 -178.325 79.045 -177.995 ;
        RECT 78.715 -179.685 79.045 -179.355 ;
        RECT 78.715 -181.045 79.045 -180.715 ;
        RECT 78.715 -182.405 79.045 -182.075 ;
        RECT 78.715 -183.765 79.045 -183.435 ;
        RECT 78.715 -185.125 79.045 -184.795 ;
        RECT 78.715 -186.485 79.045 -186.155 ;
        RECT 78.715 -187.845 79.045 -187.515 ;
        RECT 78.715 -189.205 79.045 -188.875 ;
        RECT 78.715 -190.565 79.045 -190.235 ;
        RECT 78.715 -191.925 79.045 -191.595 ;
        RECT 78.715 -193.285 79.045 -192.955 ;
        RECT 78.715 -194.645 79.045 -194.315 ;
        RECT 78.715 -196.005 79.045 -195.675 ;
        RECT 78.715 -197.365 79.045 -197.035 ;
        RECT 78.715 -198.725 79.045 -198.395 ;
        RECT 78.715 -200.085 79.045 -199.755 ;
        RECT 78.715 -201.445 79.045 -201.115 ;
        RECT 78.715 -202.805 79.045 -202.475 ;
        RECT 78.715 -204.165 79.045 -203.835 ;
        RECT 78.715 -205.525 79.045 -205.195 ;
        RECT 78.715 -206.885 79.045 -206.555 ;
        RECT 78.715 -208.245 79.045 -207.915 ;
        RECT 78.715 -209.605 79.045 -209.275 ;
        RECT 78.715 -210.965 79.045 -210.635 ;
        RECT 78.715 -212.325 79.045 -211.995 ;
        RECT 78.715 -213.685 79.045 -213.355 ;
        RECT 78.715 -215.045 79.045 -214.715 ;
        RECT 78.715 -216.405 79.045 -216.075 ;
        RECT 78.715 -217.765 79.045 -217.435 ;
        RECT 78.715 -219.125 79.045 -218.795 ;
        RECT 78.715 -220.485 79.045 -220.155 ;
        RECT 78.715 -221.845 79.045 -221.515 ;
        RECT 78.715 -223.205 79.045 -222.875 ;
        RECT 78.715 -224.565 79.045 -224.235 ;
        RECT 78.715 -225.925 79.045 -225.595 ;
        RECT 78.715 -227.285 79.045 -226.955 ;
        RECT 78.715 -228.645 79.045 -228.315 ;
        RECT 78.715 -230.005 79.045 -229.675 ;
        RECT 78.715 -231.365 79.045 -231.035 ;
        RECT 78.715 -232.725 79.045 -232.395 ;
        RECT 78.715 -234.085 79.045 -233.755 ;
        RECT 78.715 -235.445 79.045 -235.115 ;
        RECT 78.715 -236.805 79.045 -236.475 ;
        RECT 78.715 -238.165 79.045 -237.835 ;
        RECT 78.715 -243.81 79.045 -242.68 ;
        RECT 78.72 -243.925 79.04 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.96 -125.535 79.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 246.76 80.405 247.89 ;
        RECT 80.075 241.915 80.405 242.245 ;
        RECT 80.075 240.555 80.405 240.885 ;
        RECT 80.075 239.195 80.405 239.525 ;
        RECT 80.075 237.835 80.405 238.165 ;
        RECT 80.08 237.16 80.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 246.76 81.765 247.89 ;
        RECT 81.435 241.915 81.765 242.245 ;
        RECT 81.435 240.555 81.765 240.885 ;
        RECT 81.435 239.195 81.765 239.525 ;
        RECT 81.435 237.835 81.765 238.165 ;
        RECT 81.44 237.16 81.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 -1.525 81.765 -1.195 ;
        RECT 81.435 -2.885 81.765 -2.555 ;
        RECT 81.44 -3.56 81.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 246.76 83.125 247.89 ;
        RECT 82.795 241.915 83.125 242.245 ;
        RECT 82.795 240.555 83.125 240.885 ;
        RECT 82.795 239.195 83.125 239.525 ;
        RECT 82.795 237.835 83.125 238.165 ;
        RECT 82.8 237.16 83.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 -1.525 83.125 -1.195 ;
        RECT 82.795 -2.885 83.125 -2.555 ;
        RECT 82.8 -3.56 83.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 -122.565 83.125 -122.235 ;
        RECT 82.795 -123.925 83.125 -123.595 ;
        RECT 82.795 -125.285 83.125 -124.955 ;
        RECT 82.795 -126.645 83.125 -126.315 ;
        RECT 82.795 -128.005 83.125 -127.675 ;
        RECT 82.795 -129.365 83.125 -129.035 ;
        RECT 82.795 -130.725 83.125 -130.395 ;
        RECT 82.795 -132.085 83.125 -131.755 ;
        RECT 82.795 -133.445 83.125 -133.115 ;
        RECT 82.795 -134.805 83.125 -134.475 ;
        RECT 82.795 -136.165 83.125 -135.835 ;
        RECT 82.795 -137.525 83.125 -137.195 ;
        RECT 82.795 -138.885 83.125 -138.555 ;
        RECT 82.795 -140.245 83.125 -139.915 ;
        RECT 82.795 -141.605 83.125 -141.275 ;
        RECT 82.795 -142.965 83.125 -142.635 ;
        RECT 82.795 -144.325 83.125 -143.995 ;
        RECT 82.795 -145.685 83.125 -145.355 ;
        RECT 82.795 -147.045 83.125 -146.715 ;
        RECT 82.795 -148.405 83.125 -148.075 ;
        RECT 82.795 -149.765 83.125 -149.435 ;
        RECT 82.795 -151.125 83.125 -150.795 ;
        RECT 82.795 -152.485 83.125 -152.155 ;
        RECT 82.795 -153.845 83.125 -153.515 ;
        RECT 82.795 -155.205 83.125 -154.875 ;
        RECT 82.795 -156.565 83.125 -156.235 ;
        RECT 82.795 -157.925 83.125 -157.595 ;
        RECT 82.795 -159.285 83.125 -158.955 ;
        RECT 82.795 -160.645 83.125 -160.315 ;
        RECT 82.795 -162.005 83.125 -161.675 ;
        RECT 82.795 -163.365 83.125 -163.035 ;
        RECT 82.795 -164.725 83.125 -164.395 ;
        RECT 82.795 -166.085 83.125 -165.755 ;
        RECT 82.795 -167.445 83.125 -167.115 ;
        RECT 82.795 -168.805 83.125 -168.475 ;
        RECT 82.795 -170.165 83.125 -169.835 ;
        RECT 82.795 -171.525 83.125 -171.195 ;
        RECT 82.795 -172.885 83.125 -172.555 ;
        RECT 82.795 -174.245 83.125 -173.915 ;
        RECT 82.795 -175.605 83.125 -175.275 ;
        RECT 82.795 -176.965 83.125 -176.635 ;
        RECT 82.795 -178.325 83.125 -177.995 ;
        RECT 82.795 -179.685 83.125 -179.355 ;
        RECT 82.795 -181.045 83.125 -180.715 ;
        RECT 82.795 -182.405 83.125 -182.075 ;
        RECT 82.795 -183.765 83.125 -183.435 ;
        RECT 82.795 -185.125 83.125 -184.795 ;
        RECT 82.795 -186.485 83.125 -186.155 ;
        RECT 82.795 -187.845 83.125 -187.515 ;
        RECT 82.795 -189.205 83.125 -188.875 ;
        RECT 82.795 -190.565 83.125 -190.235 ;
        RECT 82.795 -191.925 83.125 -191.595 ;
        RECT 82.795 -193.285 83.125 -192.955 ;
        RECT 82.795 -194.645 83.125 -194.315 ;
        RECT 82.795 -196.005 83.125 -195.675 ;
        RECT 82.795 -197.365 83.125 -197.035 ;
        RECT 82.795 -198.725 83.125 -198.395 ;
        RECT 82.795 -200.085 83.125 -199.755 ;
        RECT 82.795 -201.445 83.125 -201.115 ;
        RECT 82.795 -202.805 83.125 -202.475 ;
        RECT 82.795 -204.165 83.125 -203.835 ;
        RECT 82.795 -205.525 83.125 -205.195 ;
        RECT 82.795 -206.885 83.125 -206.555 ;
        RECT 82.795 -208.245 83.125 -207.915 ;
        RECT 82.795 -209.605 83.125 -209.275 ;
        RECT 82.795 -210.965 83.125 -210.635 ;
        RECT 82.795 -212.325 83.125 -211.995 ;
        RECT 82.795 -213.685 83.125 -213.355 ;
        RECT 82.795 -215.045 83.125 -214.715 ;
        RECT 82.795 -216.405 83.125 -216.075 ;
        RECT 82.795 -217.765 83.125 -217.435 ;
        RECT 82.795 -219.125 83.125 -218.795 ;
        RECT 82.795 -220.485 83.125 -220.155 ;
        RECT 82.795 -221.845 83.125 -221.515 ;
        RECT 82.795 -223.205 83.125 -222.875 ;
        RECT 82.795 -224.565 83.125 -224.235 ;
        RECT 82.795 -225.925 83.125 -225.595 ;
        RECT 82.795 -227.285 83.125 -226.955 ;
        RECT 82.795 -228.645 83.125 -228.315 ;
        RECT 82.795 -230.005 83.125 -229.675 ;
        RECT 82.795 -231.365 83.125 -231.035 ;
        RECT 82.795 -232.725 83.125 -232.395 ;
        RECT 82.795 -234.085 83.125 -233.755 ;
        RECT 82.795 -235.445 83.125 -235.115 ;
        RECT 82.795 -236.805 83.125 -236.475 ;
        RECT 82.795 -238.165 83.125 -237.835 ;
        RECT 82.795 -243.81 83.125 -242.68 ;
        RECT 82.8 -243.925 83.12 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 246.76 84.485 247.89 ;
        RECT 84.155 241.915 84.485 242.245 ;
        RECT 84.155 240.555 84.485 240.885 ;
        RECT 84.155 239.195 84.485 239.525 ;
        RECT 84.155 237.835 84.485 238.165 ;
        RECT 84.16 237.16 84.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -1.525 84.485 -1.195 ;
        RECT 84.155 -2.885 84.485 -2.555 ;
        RECT 84.16 -3.56 84.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -122.565 84.485 -122.235 ;
        RECT 84.155 -123.925 84.485 -123.595 ;
        RECT 84.155 -125.285 84.485 -124.955 ;
        RECT 84.155 -126.645 84.485 -126.315 ;
        RECT 84.155 -128.005 84.485 -127.675 ;
        RECT 84.155 -129.365 84.485 -129.035 ;
        RECT 84.155 -130.725 84.485 -130.395 ;
        RECT 84.155 -132.085 84.485 -131.755 ;
        RECT 84.155 -133.445 84.485 -133.115 ;
        RECT 84.155 -134.805 84.485 -134.475 ;
        RECT 84.155 -136.165 84.485 -135.835 ;
        RECT 84.155 -137.525 84.485 -137.195 ;
        RECT 84.155 -138.885 84.485 -138.555 ;
        RECT 84.155 -140.245 84.485 -139.915 ;
        RECT 84.155 -141.605 84.485 -141.275 ;
        RECT 84.155 -142.965 84.485 -142.635 ;
        RECT 84.155 -144.325 84.485 -143.995 ;
        RECT 84.155 -145.685 84.485 -145.355 ;
        RECT 84.155 -147.045 84.485 -146.715 ;
        RECT 84.155 -148.405 84.485 -148.075 ;
        RECT 84.155 -149.765 84.485 -149.435 ;
        RECT 84.155 -151.125 84.485 -150.795 ;
        RECT 84.155 -152.485 84.485 -152.155 ;
        RECT 84.155 -153.845 84.485 -153.515 ;
        RECT 84.155 -155.205 84.485 -154.875 ;
        RECT 84.155 -156.565 84.485 -156.235 ;
        RECT 84.155 -157.925 84.485 -157.595 ;
        RECT 84.155 -159.285 84.485 -158.955 ;
        RECT 84.155 -160.645 84.485 -160.315 ;
        RECT 84.155 -162.005 84.485 -161.675 ;
        RECT 84.155 -163.365 84.485 -163.035 ;
        RECT 84.155 -164.725 84.485 -164.395 ;
        RECT 84.155 -166.085 84.485 -165.755 ;
        RECT 84.155 -167.445 84.485 -167.115 ;
        RECT 84.155 -168.805 84.485 -168.475 ;
        RECT 84.155 -170.165 84.485 -169.835 ;
        RECT 84.155 -171.525 84.485 -171.195 ;
        RECT 84.155 -172.885 84.485 -172.555 ;
        RECT 84.155 -174.245 84.485 -173.915 ;
        RECT 84.155 -175.605 84.485 -175.275 ;
        RECT 84.155 -176.965 84.485 -176.635 ;
        RECT 84.155 -178.325 84.485 -177.995 ;
        RECT 84.155 -179.685 84.485 -179.355 ;
        RECT 84.155 -181.045 84.485 -180.715 ;
        RECT 84.155 -182.405 84.485 -182.075 ;
        RECT 84.155 -183.765 84.485 -183.435 ;
        RECT 84.155 -185.125 84.485 -184.795 ;
        RECT 84.155 -186.485 84.485 -186.155 ;
        RECT 84.155 -187.845 84.485 -187.515 ;
        RECT 84.155 -189.205 84.485 -188.875 ;
        RECT 84.155 -190.565 84.485 -190.235 ;
        RECT 84.155 -191.925 84.485 -191.595 ;
        RECT 84.155 -193.285 84.485 -192.955 ;
        RECT 84.155 -194.645 84.485 -194.315 ;
        RECT 84.155 -196.005 84.485 -195.675 ;
        RECT 84.155 -197.365 84.485 -197.035 ;
        RECT 84.155 -198.725 84.485 -198.395 ;
        RECT 84.155 -200.085 84.485 -199.755 ;
        RECT 84.155 -201.445 84.485 -201.115 ;
        RECT 84.155 -202.805 84.485 -202.475 ;
        RECT 84.155 -204.165 84.485 -203.835 ;
        RECT 84.155 -205.525 84.485 -205.195 ;
        RECT 84.155 -206.885 84.485 -206.555 ;
        RECT 84.155 -208.245 84.485 -207.915 ;
        RECT 84.155 -209.605 84.485 -209.275 ;
        RECT 84.155 -210.965 84.485 -210.635 ;
        RECT 84.155 -212.325 84.485 -211.995 ;
        RECT 84.155 -213.685 84.485 -213.355 ;
        RECT 84.155 -215.045 84.485 -214.715 ;
        RECT 84.155 -216.405 84.485 -216.075 ;
        RECT 84.155 -217.765 84.485 -217.435 ;
        RECT 84.155 -219.125 84.485 -218.795 ;
        RECT 84.155 -220.485 84.485 -220.155 ;
        RECT 84.155 -221.845 84.485 -221.515 ;
        RECT 84.155 -223.205 84.485 -222.875 ;
        RECT 84.155 -224.565 84.485 -224.235 ;
        RECT 84.155 -225.925 84.485 -225.595 ;
        RECT 84.155 -227.285 84.485 -226.955 ;
        RECT 84.155 -228.645 84.485 -228.315 ;
        RECT 84.155 -230.005 84.485 -229.675 ;
        RECT 84.155 -231.365 84.485 -231.035 ;
        RECT 84.155 -232.725 84.485 -232.395 ;
        RECT 84.155 -234.085 84.485 -233.755 ;
        RECT 84.155 -235.445 84.485 -235.115 ;
        RECT 84.155 -236.805 84.485 -236.475 ;
        RECT 84.155 -238.165 84.485 -237.835 ;
        RECT 84.155 -243.81 84.485 -242.68 ;
        RECT 84.16 -243.925 84.48 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 246.76 85.845 247.89 ;
        RECT 85.515 241.915 85.845 242.245 ;
        RECT 85.515 240.555 85.845 240.885 ;
        RECT 85.515 239.195 85.845 239.525 ;
        RECT 85.515 237.835 85.845 238.165 ;
        RECT 85.52 237.16 85.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 -1.525 85.845 -1.195 ;
        RECT 85.515 -2.885 85.845 -2.555 ;
        RECT 85.52 -3.56 85.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 -122.565 85.845 -122.235 ;
        RECT 85.515 -123.925 85.845 -123.595 ;
        RECT 85.515 -125.285 85.845 -124.955 ;
        RECT 85.515 -126.645 85.845 -126.315 ;
        RECT 85.515 -128.005 85.845 -127.675 ;
        RECT 85.515 -129.365 85.845 -129.035 ;
        RECT 85.515 -130.725 85.845 -130.395 ;
        RECT 85.515 -132.085 85.845 -131.755 ;
        RECT 85.515 -133.445 85.845 -133.115 ;
        RECT 85.515 -134.805 85.845 -134.475 ;
        RECT 85.515 -136.165 85.845 -135.835 ;
        RECT 85.515 -137.525 85.845 -137.195 ;
        RECT 85.515 -138.885 85.845 -138.555 ;
        RECT 85.515 -140.245 85.845 -139.915 ;
        RECT 85.515 -141.605 85.845 -141.275 ;
        RECT 85.515 -142.965 85.845 -142.635 ;
        RECT 85.515 -144.325 85.845 -143.995 ;
        RECT 85.515 -145.685 85.845 -145.355 ;
        RECT 85.515 -147.045 85.845 -146.715 ;
        RECT 85.515 -148.405 85.845 -148.075 ;
        RECT 85.515 -149.765 85.845 -149.435 ;
        RECT 85.515 -151.125 85.845 -150.795 ;
        RECT 85.515 -152.485 85.845 -152.155 ;
        RECT 85.515 -153.845 85.845 -153.515 ;
        RECT 85.515 -155.205 85.845 -154.875 ;
        RECT 85.515 -156.565 85.845 -156.235 ;
        RECT 85.515 -157.925 85.845 -157.595 ;
        RECT 85.515 -159.285 85.845 -158.955 ;
        RECT 85.515 -160.645 85.845 -160.315 ;
        RECT 85.515 -162.005 85.845 -161.675 ;
        RECT 85.515 -163.365 85.845 -163.035 ;
        RECT 85.515 -164.725 85.845 -164.395 ;
        RECT 85.515 -166.085 85.845 -165.755 ;
        RECT 85.515 -167.445 85.845 -167.115 ;
        RECT 85.515 -168.805 85.845 -168.475 ;
        RECT 85.515 -170.165 85.845 -169.835 ;
        RECT 85.515 -171.525 85.845 -171.195 ;
        RECT 85.515 -172.885 85.845 -172.555 ;
        RECT 85.515 -174.245 85.845 -173.915 ;
        RECT 85.515 -175.605 85.845 -175.275 ;
        RECT 85.515 -176.965 85.845 -176.635 ;
        RECT 85.515 -178.325 85.845 -177.995 ;
        RECT 85.515 -179.685 85.845 -179.355 ;
        RECT 85.515 -181.045 85.845 -180.715 ;
        RECT 85.515 -182.405 85.845 -182.075 ;
        RECT 85.515 -183.765 85.845 -183.435 ;
        RECT 85.515 -185.125 85.845 -184.795 ;
        RECT 85.515 -186.485 85.845 -186.155 ;
        RECT 85.515 -187.845 85.845 -187.515 ;
        RECT 85.515 -189.205 85.845 -188.875 ;
        RECT 85.515 -190.565 85.845 -190.235 ;
        RECT 85.515 -191.925 85.845 -191.595 ;
        RECT 85.515 -193.285 85.845 -192.955 ;
        RECT 85.515 -194.645 85.845 -194.315 ;
        RECT 85.515 -196.005 85.845 -195.675 ;
        RECT 85.515 -197.365 85.845 -197.035 ;
        RECT 85.515 -198.725 85.845 -198.395 ;
        RECT 85.515 -200.085 85.845 -199.755 ;
        RECT 85.515 -201.445 85.845 -201.115 ;
        RECT 85.515 -202.805 85.845 -202.475 ;
        RECT 85.515 -204.165 85.845 -203.835 ;
        RECT 85.515 -205.525 85.845 -205.195 ;
        RECT 85.515 -206.885 85.845 -206.555 ;
        RECT 85.515 -208.245 85.845 -207.915 ;
        RECT 85.515 -209.605 85.845 -209.275 ;
        RECT 85.515 -210.965 85.845 -210.635 ;
        RECT 85.515 -212.325 85.845 -211.995 ;
        RECT 85.515 -213.685 85.845 -213.355 ;
        RECT 85.515 -215.045 85.845 -214.715 ;
        RECT 85.515 -216.405 85.845 -216.075 ;
        RECT 85.515 -217.765 85.845 -217.435 ;
        RECT 85.515 -219.125 85.845 -218.795 ;
        RECT 85.515 -220.485 85.845 -220.155 ;
        RECT 85.515 -221.845 85.845 -221.515 ;
        RECT 85.515 -223.205 85.845 -222.875 ;
        RECT 85.515 -224.565 85.845 -224.235 ;
        RECT 85.515 -225.925 85.845 -225.595 ;
        RECT 85.515 -227.285 85.845 -226.955 ;
        RECT 85.515 -228.645 85.845 -228.315 ;
        RECT 85.515 -230.005 85.845 -229.675 ;
        RECT 85.515 -231.365 85.845 -231.035 ;
        RECT 85.515 -232.725 85.845 -232.395 ;
        RECT 85.515 -234.085 85.845 -233.755 ;
        RECT 85.515 -235.445 85.845 -235.115 ;
        RECT 85.515 -236.805 85.845 -236.475 ;
        RECT 85.515 -238.165 85.845 -237.835 ;
        RECT 85.515 -243.81 85.845 -242.68 ;
        RECT 85.52 -243.925 85.84 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 246.76 87.205 247.89 ;
        RECT 86.875 241.915 87.205 242.245 ;
        RECT 86.875 240.555 87.205 240.885 ;
        RECT 86.875 239.195 87.205 239.525 ;
        RECT 86.875 237.835 87.205 238.165 ;
        RECT 86.88 237.16 87.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -1.525 87.205 -1.195 ;
        RECT 86.875 -2.885 87.205 -2.555 ;
        RECT 86.88 -3.56 87.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -122.565 87.205 -122.235 ;
        RECT 86.875 -123.925 87.205 -123.595 ;
        RECT 86.875 -125.285 87.205 -124.955 ;
        RECT 86.875 -126.645 87.205 -126.315 ;
        RECT 86.875 -128.005 87.205 -127.675 ;
        RECT 86.875 -129.365 87.205 -129.035 ;
        RECT 86.875 -130.725 87.205 -130.395 ;
        RECT 86.875 -132.085 87.205 -131.755 ;
        RECT 86.875 -133.445 87.205 -133.115 ;
        RECT 86.875 -134.805 87.205 -134.475 ;
        RECT 86.875 -136.165 87.205 -135.835 ;
        RECT 86.875 -137.525 87.205 -137.195 ;
        RECT 86.875 -138.885 87.205 -138.555 ;
        RECT 86.875 -140.245 87.205 -139.915 ;
        RECT 86.875 -141.605 87.205 -141.275 ;
        RECT 86.875 -142.965 87.205 -142.635 ;
        RECT 86.875 -144.325 87.205 -143.995 ;
        RECT 86.875 -145.685 87.205 -145.355 ;
        RECT 86.875 -147.045 87.205 -146.715 ;
        RECT 86.875 -148.405 87.205 -148.075 ;
        RECT 86.875 -149.765 87.205 -149.435 ;
        RECT 86.875 -151.125 87.205 -150.795 ;
        RECT 86.875 -152.485 87.205 -152.155 ;
        RECT 86.875 -153.845 87.205 -153.515 ;
        RECT 86.875 -155.205 87.205 -154.875 ;
        RECT 86.875 -156.565 87.205 -156.235 ;
        RECT 86.875 -157.925 87.205 -157.595 ;
        RECT 86.875 -159.285 87.205 -158.955 ;
        RECT 86.875 -160.645 87.205 -160.315 ;
        RECT 86.875 -162.005 87.205 -161.675 ;
        RECT 86.875 -163.365 87.205 -163.035 ;
        RECT 86.875 -164.725 87.205 -164.395 ;
        RECT 86.875 -166.085 87.205 -165.755 ;
        RECT 86.875 -167.445 87.205 -167.115 ;
        RECT 86.875 -168.805 87.205 -168.475 ;
        RECT 86.875 -170.165 87.205 -169.835 ;
        RECT 86.875 -171.525 87.205 -171.195 ;
        RECT 86.875 -172.885 87.205 -172.555 ;
        RECT 86.875 -174.245 87.205 -173.915 ;
        RECT 86.875 -175.605 87.205 -175.275 ;
        RECT 86.875 -176.965 87.205 -176.635 ;
        RECT 86.875 -178.325 87.205 -177.995 ;
        RECT 86.875 -179.685 87.205 -179.355 ;
        RECT 86.875 -181.045 87.205 -180.715 ;
        RECT 86.875 -182.405 87.205 -182.075 ;
        RECT 86.875 -183.765 87.205 -183.435 ;
        RECT 86.875 -185.125 87.205 -184.795 ;
        RECT 86.875 -186.485 87.205 -186.155 ;
        RECT 86.875 -187.845 87.205 -187.515 ;
        RECT 86.875 -189.205 87.205 -188.875 ;
        RECT 86.875 -190.565 87.205 -190.235 ;
        RECT 86.875 -191.925 87.205 -191.595 ;
        RECT 86.875 -193.285 87.205 -192.955 ;
        RECT 86.875 -194.645 87.205 -194.315 ;
        RECT 86.875 -196.005 87.205 -195.675 ;
        RECT 86.875 -197.365 87.205 -197.035 ;
        RECT 86.875 -198.725 87.205 -198.395 ;
        RECT 86.875 -200.085 87.205 -199.755 ;
        RECT 86.875 -201.445 87.205 -201.115 ;
        RECT 86.875 -202.805 87.205 -202.475 ;
        RECT 86.875 -204.165 87.205 -203.835 ;
        RECT 86.875 -205.525 87.205 -205.195 ;
        RECT 86.875 -206.885 87.205 -206.555 ;
        RECT 86.875 -208.245 87.205 -207.915 ;
        RECT 86.875 -209.605 87.205 -209.275 ;
        RECT 86.875 -210.965 87.205 -210.635 ;
        RECT 86.875 -212.325 87.205 -211.995 ;
        RECT 86.875 -213.685 87.205 -213.355 ;
        RECT 86.875 -215.045 87.205 -214.715 ;
        RECT 86.875 -216.405 87.205 -216.075 ;
        RECT 86.875 -217.765 87.205 -217.435 ;
        RECT 86.875 -219.125 87.205 -218.795 ;
        RECT 86.875 -220.485 87.205 -220.155 ;
        RECT 86.875 -221.845 87.205 -221.515 ;
        RECT 86.875 -223.205 87.205 -222.875 ;
        RECT 86.875 -224.565 87.205 -224.235 ;
        RECT 86.875 -225.925 87.205 -225.595 ;
        RECT 86.875 -227.285 87.205 -226.955 ;
        RECT 86.875 -228.645 87.205 -228.315 ;
        RECT 86.875 -230.005 87.205 -229.675 ;
        RECT 86.875 -231.365 87.205 -231.035 ;
        RECT 86.875 -232.725 87.205 -232.395 ;
        RECT 86.875 -234.085 87.205 -233.755 ;
        RECT 86.875 -235.445 87.205 -235.115 ;
        RECT 86.875 -236.805 87.205 -236.475 ;
        RECT 86.875 -238.165 87.205 -237.835 ;
        RECT 86.875 -243.81 87.205 -242.68 ;
        RECT 86.88 -243.925 87.2 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 246.76 88.565 247.89 ;
        RECT 88.235 241.915 88.565 242.245 ;
        RECT 88.235 240.555 88.565 240.885 ;
        RECT 88.235 239.195 88.565 239.525 ;
        RECT 88.235 237.835 88.565 238.165 ;
        RECT 88.24 237.16 88.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 -1.525 88.565 -1.195 ;
        RECT 88.235 -2.885 88.565 -2.555 ;
        RECT 88.24 -3.56 88.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 -122.565 88.565 -122.235 ;
        RECT 88.235 -123.925 88.565 -123.595 ;
        RECT 88.235 -125.285 88.565 -124.955 ;
        RECT 88.235 -126.645 88.565 -126.315 ;
        RECT 88.235 -128.005 88.565 -127.675 ;
        RECT 88.235 -129.365 88.565 -129.035 ;
        RECT 88.235 -130.725 88.565 -130.395 ;
        RECT 88.235 -132.085 88.565 -131.755 ;
        RECT 88.235 -133.445 88.565 -133.115 ;
        RECT 88.235 -134.805 88.565 -134.475 ;
        RECT 88.235 -136.165 88.565 -135.835 ;
        RECT 88.235 -137.525 88.565 -137.195 ;
        RECT 88.235 -138.885 88.565 -138.555 ;
        RECT 88.235 -140.245 88.565 -139.915 ;
        RECT 88.235 -141.605 88.565 -141.275 ;
        RECT 88.235 -142.965 88.565 -142.635 ;
        RECT 88.235 -144.325 88.565 -143.995 ;
        RECT 88.235 -145.685 88.565 -145.355 ;
        RECT 88.235 -147.045 88.565 -146.715 ;
        RECT 88.235 -148.405 88.565 -148.075 ;
        RECT 88.235 -149.765 88.565 -149.435 ;
        RECT 88.235 -151.125 88.565 -150.795 ;
        RECT 88.235 -152.485 88.565 -152.155 ;
        RECT 88.235 -153.845 88.565 -153.515 ;
        RECT 88.235 -155.205 88.565 -154.875 ;
        RECT 88.235 -156.565 88.565 -156.235 ;
        RECT 88.235 -157.925 88.565 -157.595 ;
        RECT 88.235 -159.285 88.565 -158.955 ;
        RECT 88.235 -160.645 88.565 -160.315 ;
        RECT 88.235 -162.005 88.565 -161.675 ;
        RECT 88.235 -163.365 88.565 -163.035 ;
        RECT 88.235 -164.725 88.565 -164.395 ;
        RECT 88.235 -166.085 88.565 -165.755 ;
        RECT 88.235 -167.445 88.565 -167.115 ;
        RECT 88.235 -168.805 88.565 -168.475 ;
        RECT 88.235 -170.165 88.565 -169.835 ;
        RECT 88.235 -171.525 88.565 -171.195 ;
        RECT 88.235 -172.885 88.565 -172.555 ;
        RECT 88.235 -174.245 88.565 -173.915 ;
        RECT 88.235 -175.605 88.565 -175.275 ;
        RECT 88.235 -176.965 88.565 -176.635 ;
        RECT 88.235 -178.325 88.565 -177.995 ;
        RECT 88.235 -179.685 88.565 -179.355 ;
        RECT 88.235 -181.045 88.565 -180.715 ;
        RECT 88.235 -182.405 88.565 -182.075 ;
        RECT 88.235 -183.765 88.565 -183.435 ;
        RECT 88.235 -185.125 88.565 -184.795 ;
        RECT 88.235 -186.485 88.565 -186.155 ;
        RECT 88.235 -187.845 88.565 -187.515 ;
        RECT 88.235 -189.205 88.565 -188.875 ;
        RECT 88.235 -190.565 88.565 -190.235 ;
        RECT 88.235 -191.925 88.565 -191.595 ;
        RECT 88.235 -193.285 88.565 -192.955 ;
        RECT 88.235 -194.645 88.565 -194.315 ;
        RECT 88.235 -196.005 88.565 -195.675 ;
        RECT 88.235 -197.365 88.565 -197.035 ;
        RECT 88.235 -198.725 88.565 -198.395 ;
        RECT 88.235 -200.085 88.565 -199.755 ;
        RECT 88.235 -201.445 88.565 -201.115 ;
        RECT 88.235 -202.805 88.565 -202.475 ;
        RECT 88.235 -204.165 88.565 -203.835 ;
        RECT 88.235 -205.525 88.565 -205.195 ;
        RECT 88.235 -206.885 88.565 -206.555 ;
        RECT 88.235 -208.245 88.565 -207.915 ;
        RECT 88.235 -209.605 88.565 -209.275 ;
        RECT 88.235 -210.965 88.565 -210.635 ;
        RECT 88.235 -212.325 88.565 -211.995 ;
        RECT 88.235 -213.685 88.565 -213.355 ;
        RECT 88.235 -215.045 88.565 -214.715 ;
        RECT 88.235 -216.405 88.565 -216.075 ;
        RECT 88.235 -217.765 88.565 -217.435 ;
        RECT 88.235 -219.125 88.565 -218.795 ;
        RECT 88.235 -220.485 88.565 -220.155 ;
        RECT 88.235 -221.845 88.565 -221.515 ;
        RECT 88.235 -223.205 88.565 -222.875 ;
        RECT 88.235 -224.565 88.565 -224.235 ;
        RECT 88.235 -225.925 88.565 -225.595 ;
        RECT 88.235 -227.285 88.565 -226.955 ;
        RECT 88.235 -228.645 88.565 -228.315 ;
        RECT 88.235 -230.005 88.565 -229.675 ;
        RECT 88.235 -231.365 88.565 -231.035 ;
        RECT 88.235 -232.725 88.565 -232.395 ;
        RECT 88.235 -234.085 88.565 -233.755 ;
        RECT 88.235 -235.445 88.565 -235.115 ;
        RECT 88.235 -236.805 88.565 -236.475 ;
        RECT 88.235 -238.165 88.565 -237.835 ;
        RECT 88.235 -243.81 88.565 -242.68 ;
        RECT 88.24 -243.925 88.56 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 246.76 89.925 247.89 ;
        RECT 89.595 241.915 89.925 242.245 ;
        RECT 89.595 240.555 89.925 240.885 ;
        RECT 89.595 239.195 89.925 239.525 ;
        RECT 89.595 237.835 89.925 238.165 ;
        RECT 89.6 237.16 89.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 -126.645 89.925 -126.315 ;
        RECT 89.595 -128.005 89.925 -127.675 ;
        RECT 89.595 -129.365 89.925 -129.035 ;
        RECT 89.595 -130.725 89.925 -130.395 ;
        RECT 89.595 -132.085 89.925 -131.755 ;
        RECT 89.595 -133.445 89.925 -133.115 ;
        RECT 89.595 -134.805 89.925 -134.475 ;
        RECT 89.595 -136.165 89.925 -135.835 ;
        RECT 89.595 -137.525 89.925 -137.195 ;
        RECT 89.595 -138.885 89.925 -138.555 ;
        RECT 89.595 -140.245 89.925 -139.915 ;
        RECT 89.595 -141.605 89.925 -141.275 ;
        RECT 89.595 -142.965 89.925 -142.635 ;
        RECT 89.595 -144.325 89.925 -143.995 ;
        RECT 89.595 -145.685 89.925 -145.355 ;
        RECT 89.595 -147.045 89.925 -146.715 ;
        RECT 89.595 -148.405 89.925 -148.075 ;
        RECT 89.595 -149.765 89.925 -149.435 ;
        RECT 89.595 -151.125 89.925 -150.795 ;
        RECT 89.595 -152.485 89.925 -152.155 ;
        RECT 89.595 -153.845 89.925 -153.515 ;
        RECT 89.595 -155.205 89.925 -154.875 ;
        RECT 89.595 -156.565 89.925 -156.235 ;
        RECT 89.595 -157.925 89.925 -157.595 ;
        RECT 89.595 -159.285 89.925 -158.955 ;
        RECT 89.595 -160.645 89.925 -160.315 ;
        RECT 89.595 -162.005 89.925 -161.675 ;
        RECT 89.595 -163.365 89.925 -163.035 ;
        RECT 89.595 -164.725 89.925 -164.395 ;
        RECT 89.595 -166.085 89.925 -165.755 ;
        RECT 89.595 -167.445 89.925 -167.115 ;
        RECT 89.595 -168.805 89.925 -168.475 ;
        RECT 89.595 -170.165 89.925 -169.835 ;
        RECT 89.595 -171.525 89.925 -171.195 ;
        RECT 89.595 -172.885 89.925 -172.555 ;
        RECT 89.595 -174.245 89.925 -173.915 ;
        RECT 89.595 -175.605 89.925 -175.275 ;
        RECT 89.595 -176.965 89.925 -176.635 ;
        RECT 89.595 -178.325 89.925 -177.995 ;
        RECT 89.595 -179.685 89.925 -179.355 ;
        RECT 89.595 -181.045 89.925 -180.715 ;
        RECT 89.595 -182.405 89.925 -182.075 ;
        RECT 89.595 -183.765 89.925 -183.435 ;
        RECT 89.595 -185.125 89.925 -184.795 ;
        RECT 89.595 -186.485 89.925 -186.155 ;
        RECT 89.595 -187.845 89.925 -187.515 ;
        RECT 89.595 -189.205 89.925 -188.875 ;
        RECT 89.595 -190.565 89.925 -190.235 ;
        RECT 89.595 -191.925 89.925 -191.595 ;
        RECT 89.595 -193.285 89.925 -192.955 ;
        RECT 89.595 -194.645 89.925 -194.315 ;
        RECT 89.595 -196.005 89.925 -195.675 ;
        RECT 89.595 -197.365 89.925 -197.035 ;
        RECT 89.595 -198.725 89.925 -198.395 ;
        RECT 89.595 -200.085 89.925 -199.755 ;
        RECT 89.595 -201.445 89.925 -201.115 ;
        RECT 89.595 -202.805 89.925 -202.475 ;
        RECT 89.595 -204.165 89.925 -203.835 ;
        RECT 89.595 -205.525 89.925 -205.195 ;
        RECT 89.595 -206.885 89.925 -206.555 ;
        RECT 89.595 -208.245 89.925 -207.915 ;
        RECT 89.595 -209.605 89.925 -209.275 ;
        RECT 89.595 -210.965 89.925 -210.635 ;
        RECT 89.595 -212.325 89.925 -211.995 ;
        RECT 89.595 -213.685 89.925 -213.355 ;
        RECT 89.595 -215.045 89.925 -214.715 ;
        RECT 89.595 -216.405 89.925 -216.075 ;
        RECT 89.595 -217.765 89.925 -217.435 ;
        RECT 89.595 -219.125 89.925 -218.795 ;
        RECT 89.595 -220.485 89.925 -220.155 ;
        RECT 89.595 -221.845 89.925 -221.515 ;
        RECT 89.595 -223.205 89.925 -222.875 ;
        RECT 89.595 -224.565 89.925 -224.235 ;
        RECT 89.595 -225.925 89.925 -225.595 ;
        RECT 89.595 -227.285 89.925 -226.955 ;
        RECT 89.595 -228.645 89.925 -228.315 ;
        RECT 89.595 -230.005 89.925 -229.675 ;
        RECT 89.595 -231.365 89.925 -231.035 ;
        RECT 89.595 -232.725 89.925 -232.395 ;
        RECT 89.595 -234.085 89.925 -233.755 ;
        RECT 89.595 -235.445 89.925 -235.115 ;
        RECT 89.595 -236.805 89.925 -236.475 ;
        RECT 89.595 -238.165 89.925 -237.835 ;
        RECT 89.595 -243.81 89.925 -242.68 ;
        RECT 89.6 -243.925 89.92 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.86 -125.535 90.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 246.76 91.285 247.89 ;
        RECT 90.955 241.915 91.285 242.245 ;
        RECT 90.955 240.555 91.285 240.885 ;
        RECT 90.955 239.195 91.285 239.525 ;
        RECT 90.955 237.835 91.285 238.165 ;
        RECT 90.96 237.16 91.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 246.76 92.645 247.89 ;
        RECT 92.315 241.915 92.645 242.245 ;
        RECT 92.315 240.555 92.645 240.885 ;
        RECT 92.315 239.195 92.645 239.525 ;
        RECT 92.315 237.835 92.645 238.165 ;
        RECT 92.32 237.16 92.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -1.525 92.645 -1.195 ;
        RECT 92.315 -2.885 92.645 -2.555 ;
        RECT 92.32 -3.56 92.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 246.76 94.005 247.89 ;
        RECT 93.675 241.915 94.005 242.245 ;
        RECT 93.675 240.555 94.005 240.885 ;
        RECT 93.675 239.195 94.005 239.525 ;
        RECT 93.675 237.835 94.005 238.165 ;
        RECT 93.68 237.16 94 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 246.76 55.925 247.89 ;
        RECT 55.595 241.915 55.925 242.245 ;
        RECT 55.595 240.555 55.925 240.885 ;
        RECT 55.595 239.195 55.925 239.525 ;
        RECT 55.595 237.835 55.925 238.165 ;
        RECT 55.6 237.16 55.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 -1.525 55.925 -1.195 ;
        RECT 55.595 -2.885 55.925 -2.555 ;
        RECT 55.6 -3.56 55.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 -122.565 55.925 -122.235 ;
        RECT 55.595 -123.925 55.925 -123.595 ;
        RECT 55.595 -125.285 55.925 -124.955 ;
        RECT 55.595 -126.645 55.925 -126.315 ;
        RECT 55.595 -128.005 55.925 -127.675 ;
        RECT 55.595 -129.365 55.925 -129.035 ;
        RECT 55.595 -130.725 55.925 -130.395 ;
        RECT 55.595 -132.085 55.925 -131.755 ;
        RECT 55.595 -133.445 55.925 -133.115 ;
        RECT 55.595 -134.805 55.925 -134.475 ;
        RECT 55.595 -136.165 55.925 -135.835 ;
        RECT 55.595 -137.525 55.925 -137.195 ;
        RECT 55.595 -138.885 55.925 -138.555 ;
        RECT 55.595 -140.245 55.925 -139.915 ;
        RECT 55.595 -141.605 55.925 -141.275 ;
        RECT 55.595 -142.965 55.925 -142.635 ;
        RECT 55.595 -144.325 55.925 -143.995 ;
        RECT 55.595 -145.685 55.925 -145.355 ;
        RECT 55.595 -147.045 55.925 -146.715 ;
        RECT 55.595 -148.405 55.925 -148.075 ;
        RECT 55.595 -149.765 55.925 -149.435 ;
        RECT 55.595 -151.125 55.925 -150.795 ;
        RECT 55.595 -152.485 55.925 -152.155 ;
        RECT 55.595 -153.845 55.925 -153.515 ;
        RECT 55.595 -155.205 55.925 -154.875 ;
        RECT 55.595 -156.565 55.925 -156.235 ;
        RECT 55.595 -157.925 55.925 -157.595 ;
        RECT 55.595 -159.285 55.925 -158.955 ;
        RECT 55.595 -160.645 55.925 -160.315 ;
        RECT 55.595 -162.005 55.925 -161.675 ;
        RECT 55.595 -163.365 55.925 -163.035 ;
        RECT 55.595 -164.725 55.925 -164.395 ;
        RECT 55.595 -166.085 55.925 -165.755 ;
        RECT 55.595 -167.445 55.925 -167.115 ;
        RECT 55.595 -168.805 55.925 -168.475 ;
        RECT 55.595 -170.165 55.925 -169.835 ;
        RECT 55.595 -171.525 55.925 -171.195 ;
        RECT 55.595 -172.885 55.925 -172.555 ;
        RECT 55.595 -174.245 55.925 -173.915 ;
        RECT 55.595 -175.605 55.925 -175.275 ;
        RECT 55.595 -176.965 55.925 -176.635 ;
        RECT 55.595 -178.325 55.925 -177.995 ;
        RECT 55.595 -179.685 55.925 -179.355 ;
        RECT 55.595 -181.045 55.925 -180.715 ;
        RECT 55.595 -182.405 55.925 -182.075 ;
        RECT 55.595 -183.765 55.925 -183.435 ;
        RECT 55.595 -185.125 55.925 -184.795 ;
        RECT 55.595 -186.485 55.925 -186.155 ;
        RECT 55.595 -187.845 55.925 -187.515 ;
        RECT 55.595 -189.205 55.925 -188.875 ;
        RECT 55.595 -190.565 55.925 -190.235 ;
        RECT 55.595 -191.925 55.925 -191.595 ;
        RECT 55.595 -193.285 55.925 -192.955 ;
        RECT 55.595 -194.645 55.925 -194.315 ;
        RECT 55.595 -196.005 55.925 -195.675 ;
        RECT 55.595 -197.365 55.925 -197.035 ;
        RECT 55.595 -198.725 55.925 -198.395 ;
        RECT 55.595 -200.085 55.925 -199.755 ;
        RECT 55.595 -201.445 55.925 -201.115 ;
        RECT 55.595 -202.805 55.925 -202.475 ;
        RECT 55.595 -204.165 55.925 -203.835 ;
        RECT 55.595 -205.525 55.925 -205.195 ;
        RECT 55.595 -206.885 55.925 -206.555 ;
        RECT 55.595 -208.245 55.925 -207.915 ;
        RECT 55.595 -209.605 55.925 -209.275 ;
        RECT 55.595 -210.965 55.925 -210.635 ;
        RECT 55.595 -212.325 55.925 -211.995 ;
        RECT 55.595 -213.685 55.925 -213.355 ;
        RECT 55.595 -215.045 55.925 -214.715 ;
        RECT 55.595 -216.405 55.925 -216.075 ;
        RECT 55.595 -217.765 55.925 -217.435 ;
        RECT 55.595 -219.125 55.925 -218.795 ;
        RECT 55.595 -220.485 55.925 -220.155 ;
        RECT 55.595 -221.845 55.925 -221.515 ;
        RECT 55.595 -223.205 55.925 -222.875 ;
        RECT 55.595 -224.565 55.925 -224.235 ;
        RECT 55.595 -225.925 55.925 -225.595 ;
        RECT 55.595 -227.285 55.925 -226.955 ;
        RECT 55.595 -228.645 55.925 -228.315 ;
        RECT 55.595 -230.005 55.925 -229.675 ;
        RECT 55.595 -231.365 55.925 -231.035 ;
        RECT 55.595 -232.725 55.925 -232.395 ;
        RECT 55.595 -234.085 55.925 -233.755 ;
        RECT 55.595 -235.445 55.925 -235.115 ;
        RECT 55.595 -236.805 55.925 -236.475 ;
        RECT 55.595 -238.165 55.925 -237.835 ;
        RECT 55.595 -243.81 55.925 -242.68 ;
        RECT 55.6 -243.925 55.92 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 246.76 57.285 247.89 ;
        RECT 56.955 241.915 57.285 242.245 ;
        RECT 56.955 240.555 57.285 240.885 ;
        RECT 56.955 239.195 57.285 239.525 ;
        RECT 56.955 237.835 57.285 238.165 ;
        RECT 56.96 237.16 57.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 -126.645 57.285 -126.315 ;
        RECT 56.955 -128.005 57.285 -127.675 ;
        RECT 56.955 -129.365 57.285 -129.035 ;
        RECT 56.955 -130.725 57.285 -130.395 ;
        RECT 56.955 -132.085 57.285 -131.755 ;
        RECT 56.955 -133.445 57.285 -133.115 ;
        RECT 56.955 -134.805 57.285 -134.475 ;
        RECT 56.955 -136.165 57.285 -135.835 ;
        RECT 56.955 -137.525 57.285 -137.195 ;
        RECT 56.955 -138.885 57.285 -138.555 ;
        RECT 56.955 -140.245 57.285 -139.915 ;
        RECT 56.955 -141.605 57.285 -141.275 ;
        RECT 56.955 -142.965 57.285 -142.635 ;
        RECT 56.955 -144.325 57.285 -143.995 ;
        RECT 56.955 -145.685 57.285 -145.355 ;
        RECT 56.955 -147.045 57.285 -146.715 ;
        RECT 56.955 -148.405 57.285 -148.075 ;
        RECT 56.955 -149.765 57.285 -149.435 ;
        RECT 56.955 -151.125 57.285 -150.795 ;
        RECT 56.955 -152.485 57.285 -152.155 ;
        RECT 56.955 -153.845 57.285 -153.515 ;
        RECT 56.955 -155.205 57.285 -154.875 ;
        RECT 56.955 -156.565 57.285 -156.235 ;
        RECT 56.955 -157.925 57.285 -157.595 ;
        RECT 56.955 -159.285 57.285 -158.955 ;
        RECT 56.955 -160.645 57.285 -160.315 ;
        RECT 56.955 -162.005 57.285 -161.675 ;
        RECT 56.955 -163.365 57.285 -163.035 ;
        RECT 56.955 -164.725 57.285 -164.395 ;
        RECT 56.955 -166.085 57.285 -165.755 ;
        RECT 56.955 -167.445 57.285 -167.115 ;
        RECT 56.955 -168.805 57.285 -168.475 ;
        RECT 56.955 -170.165 57.285 -169.835 ;
        RECT 56.955 -171.525 57.285 -171.195 ;
        RECT 56.955 -172.885 57.285 -172.555 ;
        RECT 56.955 -174.245 57.285 -173.915 ;
        RECT 56.955 -175.605 57.285 -175.275 ;
        RECT 56.955 -176.965 57.285 -176.635 ;
        RECT 56.955 -178.325 57.285 -177.995 ;
        RECT 56.955 -179.685 57.285 -179.355 ;
        RECT 56.955 -181.045 57.285 -180.715 ;
        RECT 56.955 -182.405 57.285 -182.075 ;
        RECT 56.955 -183.765 57.285 -183.435 ;
        RECT 56.955 -185.125 57.285 -184.795 ;
        RECT 56.955 -186.485 57.285 -186.155 ;
        RECT 56.955 -187.845 57.285 -187.515 ;
        RECT 56.955 -189.205 57.285 -188.875 ;
        RECT 56.955 -190.565 57.285 -190.235 ;
        RECT 56.955 -191.925 57.285 -191.595 ;
        RECT 56.955 -193.285 57.285 -192.955 ;
        RECT 56.955 -194.645 57.285 -194.315 ;
        RECT 56.955 -196.005 57.285 -195.675 ;
        RECT 56.955 -197.365 57.285 -197.035 ;
        RECT 56.955 -198.725 57.285 -198.395 ;
        RECT 56.955 -200.085 57.285 -199.755 ;
        RECT 56.955 -201.445 57.285 -201.115 ;
        RECT 56.955 -202.805 57.285 -202.475 ;
        RECT 56.955 -204.165 57.285 -203.835 ;
        RECT 56.955 -205.525 57.285 -205.195 ;
        RECT 56.955 -206.885 57.285 -206.555 ;
        RECT 56.955 -208.245 57.285 -207.915 ;
        RECT 56.955 -209.605 57.285 -209.275 ;
        RECT 56.955 -210.965 57.285 -210.635 ;
        RECT 56.955 -212.325 57.285 -211.995 ;
        RECT 56.955 -213.685 57.285 -213.355 ;
        RECT 56.955 -215.045 57.285 -214.715 ;
        RECT 56.955 -216.405 57.285 -216.075 ;
        RECT 56.955 -217.765 57.285 -217.435 ;
        RECT 56.955 -219.125 57.285 -218.795 ;
        RECT 56.955 -220.485 57.285 -220.155 ;
        RECT 56.955 -221.845 57.285 -221.515 ;
        RECT 56.955 -223.205 57.285 -222.875 ;
        RECT 56.955 -224.565 57.285 -224.235 ;
        RECT 56.955 -225.925 57.285 -225.595 ;
        RECT 56.955 -227.285 57.285 -226.955 ;
        RECT 56.955 -228.645 57.285 -228.315 ;
        RECT 56.955 -230.005 57.285 -229.675 ;
        RECT 56.955 -231.365 57.285 -231.035 ;
        RECT 56.955 -232.725 57.285 -232.395 ;
        RECT 56.955 -234.085 57.285 -233.755 ;
        RECT 56.955 -235.445 57.285 -235.115 ;
        RECT 56.955 -236.805 57.285 -236.475 ;
        RECT 56.955 -238.165 57.285 -237.835 ;
        RECT 56.955 -243.81 57.285 -242.68 ;
        RECT 56.96 -243.925 57.28 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.16 -125.535 57.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.315 246.76 58.645 247.89 ;
        RECT 58.315 241.915 58.645 242.245 ;
        RECT 58.315 240.555 58.645 240.885 ;
        RECT 58.315 239.195 58.645 239.525 ;
        RECT 58.315 237.835 58.645 238.165 ;
        RECT 58.32 237.16 58.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 246.76 60.005 247.89 ;
        RECT 59.675 241.915 60.005 242.245 ;
        RECT 59.675 240.555 60.005 240.885 ;
        RECT 59.675 239.195 60.005 239.525 ;
        RECT 59.675 237.835 60.005 238.165 ;
        RECT 59.68 237.16 60 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 -1.525 60.005 -1.195 ;
        RECT 59.675 -2.885 60.005 -2.555 ;
        RECT 59.68 -3.56 60 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 246.76 61.365 247.89 ;
        RECT 61.035 241.915 61.365 242.245 ;
        RECT 61.035 240.555 61.365 240.885 ;
        RECT 61.035 239.195 61.365 239.525 ;
        RECT 61.035 237.835 61.365 238.165 ;
        RECT 61.04 237.16 61.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 -1.525 61.365 -1.195 ;
        RECT 61.035 -2.885 61.365 -2.555 ;
        RECT 61.04 -3.56 61.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 -122.565 61.365 -122.235 ;
        RECT 61.035 -123.925 61.365 -123.595 ;
        RECT 61.035 -125.285 61.365 -124.955 ;
        RECT 61.035 -126.645 61.365 -126.315 ;
        RECT 61.035 -128.005 61.365 -127.675 ;
        RECT 61.035 -129.365 61.365 -129.035 ;
        RECT 61.035 -130.725 61.365 -130.395 ;
        RECT 61.035 -132.085 61.365 -131.755 ;
        RECT 61.035 -133.445 61.365 -133.115 ;
        RECT 61.035 -134.805 61.365 -134.475 ;
        RECT 61.035 -136.165 61.365 -135.835 ;
        RECT 61.035 -137.525 61.365 -137.195 ;
        RECT 61.035 -138.885 61.365 -138.555 ;
        RECT 61.035 -140.245 61.365 -139.915 ;
        RECT 61.035 -141.605 61.365 -141.275 ;
        RECT 61.035 -142.965 61.365 -142.635 ;
        RECT 61.035 -144.325 61.365 -143.995 ;
        RECT 61.035 -145.685 61.365 -145.355 ;
        RECT 61.035 -147.045 61.365 -146.715 ;
        RECT 61.035 -148.405 61.365 -148.075 ;
        RECT 61.035 -149.765 61.365 -149.435 ;
        RECT 61.035 -151.125 61.365 -150.795 ;
        RECT 61.035 -152.485 61.365 -152.155 ;
        RECT 61.035 -153.845 61.365 -153.515 ;
        RECT 61.035 -155.205 61.365 -154.875 ;
        RECT 61.035 -156.565 61.365 -156.235 ;
        RECT 61.035 -157.925 61.365 -157.595 ;
        RECT 61.035 -159.285 61.365 -158.955 ;
        RECT 61.035 -160.645 61.365 -160.315 ;
        RECT 61.035 -162.005 61.365 -161.675 ;
        RECT 61.035 -163.365 61.365 -163.035 ;
        RECT 61.035 -164.725 61.365 -164.395 ;
        RECT 61.035 -166.085 61.365 -165.755 ;
        RECT 61.035 -167.445 61.365 -167.115 ;
        RECT 61.035 -168.805 61.365 -168.475 ;
        RECT 61.035 -170.165 61.365 -169.835 ;
        RECT 61.035 -171.525 61.365 -171.195 ;
        RECT 61.035 -172.885 61.365 -172.555 ;
        RECT 61.035 -174.245 61.365 -173.915 ;
        RECT 61.035 -175.605 61.365 -175.275 ;
        RECT 61.035 -176.965 61.365 -176.635 ;
        RECT 61.035 -178.325 61.365 -177.995 ;
        RECT 61.035 -179.685 61.365 -179.355 ;
        RECT 61.035 -181.045 61.365 -180.715 ;
        RECT 61.035 -182.405 61.365 -182.075 ;
        RECT 61.035 -183.765 61.365 -183.435 ;
        RECT 61.035 -185.125 61.365 -184.795 ;
        RECT 61.035 -186.485 61.365 -186.155 ;
        RECT 61.035 -187.845 61.365 -187.515 ;
        RECT 61.035 -189.205 61.365 -188.875 ;
        RECT 61.035 -190.565 61.365 -190.235 ;
        RECT 61.035 -191.925 61.365 -191.595 ;
        RECT 61.035 -193.285 61.365 -192.955 ;
        RECT 61.035 -194.645 61.365 -194.315 ;
        RECT 61.035 -196.005 61.365 -195.675 ;
        RECT 61.035 -197.365 61.365 -197.035 ;
        RECT 61.035 -198.725 61.365 -198.395 ;
        RECT 61.035 -200.085 61.365 -199.755 ;
        RECT 61.035 -201.445 61.365 -201.115 ;
        RECT 61.035 -202.805 61.365 -202.475 ;
        RECT 61.035 -204.165 61.365 -203.835 ;
        RECT 61.035 -205.525 61.365 -205.195 ;
        RECT 61.035 -206.885 61.365 -206.555 ;
        RECT 61.035 -208.245 61.365 -207.915 ;
        RECT 61.035 -209.605 61.365 -209.275 ;
        RECT 61.035 -210.965 61.365 -210.635 ;
        RECT 61.035 -212.325 61.365 -211.995 ;
        RECT 61.035 -213.685 61.365 -213.355 ;
        RECT 61.035 -215.045 61.365 -214.715 ;
        RECT 61.035 -216.405 61.365 -216.075 ;
        RECT 61.035 -217.765 61.365 -217.435 ;
        RECT 61.035 -219.125 61.365 -218.795 ;
        RECT 61.035 -220.485 61.365 -220.155 ;
        RECT 61.035 -221.845 61.365 -221.515 ;
        RECT 61.035 -223.205 61.365 -222.875 ;
        RECT 61.035 -224.565 61.365 -224.235 ;
        RECT 61.035 -225.925 61.365 -225.595 ;
        RECT 61.035 -227.285 61.365 -226.955 ;
        RECT 61.035 -228.645 61.365 -228.315 ;
        RECT 61.035 -230.005 61.365 -229.675 ;
        RECT 61.035 -231.365 61.365 -231.035 ;
        RECT 61.035 -232.725 61.365 -232.395 ;
        RECT 61.035 -234.085 61.365 -233.755 ;
        RECT 61.035 -235.445 61.365 -235.115 ;
        RECT 61.035 -236.805 61.365 -236.475 ;
        RECT 61.035 -238.165 61.365 -237.835 ;
        RECT 61.035 -243.81 61.365 -242.68 ;
        RECT 61.04 -243.925 61.36 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 246.76 62.725 247.89 ;
        RECT 62.395 241.915 62.725 242.245 ;
        RECT 62.395 240.555 62.725 240.885 ;
        RECT 62.395 239.195 62.725 239.525 ;
        RECT 62.395 237.835 62.725 238.165 ;
        RECT 62.4 237.16 62.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -1.525 62.725 -1.195 ;
        RECT 62.395 -2.885 62.725 -2.555 ;
        RECT 62.4 -3.56 62.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -122.565 62.725 -122.235 ;
        RECT 62.395 -123.925 62.725 -123.595 ;
        RECT 62.395 -125.285 62.725 -124.955 ;
        RECT 62.395 -126.645 62.725 -126.315 ;
        RECT 62.395 -128.005 62.725 -127.675 ;
        RECT 62.395 -129.365 62.725 -129.035 ;
        RECT 62.395 -130.725 62.725 -130.395 ;
        RECT 62.395 -132.085 62.725 -131.755 ;
        RECT 62.395 -133.445 62.725 -133.115 ;
        RECT 62.395 -134.805 62.725 -134.475 ;
        RECT 62.395 -136.165 62.725 -135.835 ;
        RECT 62.395 -137.525 62.725 -137.195 ;
        RECT 62.395 -138.885 62.725 -138.555 ;
        RECT 62.395 -140.245 62.725 -139.915 ;
        RECT 62.395 -141.605 62.725 -141.275 ;
        RECT 62.395 -142.965 62.725 -142.635 ;
        RECT 62.395 -144.325 62.725 -143.995 ;
        RECT 62.395 -145.685 62.725 -145.355 ;
        RECT 62.395 -147.045 62.725 -146.715 ;
        RECT 62.395 -148.405 62.725 -148.075 ;
        RECT 62.395 -149.765 62.725 -149.435 ;
        RECT 62.395 -151.125 62.725 -150.795 ;
        RECT 62.395 -152.485 62.725 -152.155 ;
        RECT 62.395 -153.845 62.725 -153.515 ;
        RECT 62.395 -155.205 62.725 -154.875 ;
        RECT 62.395 -156.565 62.725 -156.235 ;
        RECT 62.395 -157.925 62.725 -157.595 ;
        RECT 62.395 -159.285 62.725 -158.955 ;
        RECT 62.395 -160.645 62.725 -160.315 ;
        RECT 62.395 -162.005 62.725 -161.675 ;
        RECT 62.395 -163.365 62.725 -163.035 ;
        RECT 62.395 -164.725 62.725 -164.395 ;
        RECT 62.395 -166.085 62.725 -165.755 ;
        RECT 62.395 -167.445 62.725 -167.115 ;
        RECT 62.395 -168.805 62.725 -168.475 ;
        RECT 62.395 -170.165 62.725 -169.835 ;
        RECT 62.395 -171.525 62.725 -171.195 ;
        RECT 62.395 -172.885 62.725 -172.555 ;
        RECT 62.395 -174.245 62.725 -173.915 ;
        RECT 62.395 -175.605 62.725 -175.275 ;
        RECT 62.395 -176.965 62.725 -176.635 ;
        RECT 62.395 -178.325 62.725 -177.995 ;
        RECT 62.395 -179.685 62.725 -179.355 ;
        RECT 62.395 -181.045 62.725 -180.715 ;
        RECT 62.395 -182.405 62.725 -182.075 ;
        RECT 62.395 -183.765 62.725 -183.435 ;
        RECT 62.395 -185.125 62.725 -184.795 ;
        RECT 62.395 -186.485 62.725 -186.155 ;
        RECT 62.395 -187.845 62.725 -187.515 ;
        RECT 62.395 -189.205 62.725 -188.875 ;
        RECT 62.395 -190.565 62.725 -190.235 ;
        RECT 62.395 -191.925 62.725 -191.595 ;
        RECT 62.395 -193.285 62.725 -192.955 ;
        RECT 62.395 -194.645 62.725 -194.315 ;
        RECT 62.395 -196.005 62.725 -195.675 ;
        RECT 62.395 -197.365 62.725 -197.035 ;
        RECT 62.395 -198.725 62.725 -198.395 ;
        RECT 62.395 -200.085 62.725 -199.755 ;
        RECT 62.395 -201.445 62.725 -201.115 ;
        RECT 62.395 -202.805 62.725 -202.475 ;
        RECT 62.395 -204.165 62.725 -203.835 ;
        RECT 62.395 -205.525 62.725 -205.195 ;
        RECT 62.395 -206.885 62.725 -206.555 ;
        RECT 62.395 -208.245 62.725 -207.915 ;
        RECT 62.395 -209.605 62.725 -209.275 ;
        RECT 62.395 -210.965 62.725 -210.635 ;
        RECT 62.395 -212.325 62.725 -211.995 ;
        RECT 62.395 -213.685 62.725 -213.355 ;
        RECT 62.395 -215.045 62.725 -214.715 ;
        RECT 62.395 -216.405 62.725 -216.075 ;
        RECT 62.395 -217.765 62.725 -217.435 ;
        RECT 62.395 -219.125 62.725 -218.795 ;
        RECT 62.395 -220.485 62.725 -220.155 ;
        RECT 62.395 -221.845 62.725 -221.515 ;
        RECT 62.395 -223.205 62.725 -222.875 ;
        RECT 62.395 -224.565 62.725 -224.235 ;
        RECT 62.395 -225.925 62.725 -225.595 ;
        RECT 62.395 -227.285 62.725 -226.955 ;
        RECT 62.395 -228.645 62.725 -228.315 ;
        RECT 62.395 -230.005 62.725 -229.675 ;
        RECT 62.395 -231.365 62.725 -231.035 ;
        RECT 62.395 -232.725 62.725 -232.395 ;
        RECT 62.395 -234.085 62.725 -233.755 ;
        RECT 62.395 -235.445 62.725 -235.115 ;
        RECT 62.395 -236.805 62.725 -236.475 ;
        RECT 62.395 -238.165 62.725 -237.835 ;
        RECT 62.395 -243.81 62.725 -242.68 ;
        RECT 62.4 -243.925 62.72 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 246.76 64.085 247.89 ;
        RECT 63.755 241.915 64.085 242.245 ;
        RECT 63.755 240.555 64.085 240.885 ;
        RECT 63.755 239.195 64.085 239.525 ;
        RECT 63.755 237.835 64.085 238.165 ;
        RECT 63.76 237.16 64.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 -1.525 64.085 -1.195 ;
        RECT 63.755 -2.885 64.085 -2.555 ;
        RECT 63.76 -3.56 64.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 -122.565 64.085 -122.235 ;
        RECT 63.755 -123.925 64.085 -123.595 ;
        RECT 63.755 -125.285 64.085 -124.955 ;
        RECT 63.755 -126.645 64.085 -126.315 ;
        RECT 63.755 -128.005 64.085 -127.675 ;
        RECT 63.755 -129.365 64.085 -129.035 ;
        RECT 63.755 -130.725 64.085 -130.395 ;
        RECT 63.755 -132.085 64.085 -131.755 ;
        RECT 63.755 -133.445 64.085 -133.115 ;
        RECT 63.755 -134.805 64.085 -134.475 ;
        RECT 63.755 -136.165 64.085 -135.835 ;
        RECT 63.755 -137.525 64.085 -137.195 ;
        RECT 63.755 -138.885 64.085 -138.555 ;
        RECT 63.755 -140.245 64.085 -139.915 ;
        RECT 63.755 -141.605 64.085 -141.275 ;
        RECT 63.755 -142.965 64.085 -142.635 ;
        RECT 63.755 -144.325 64.085 -143.995 ;
        RECT 63.755 -145.685 64.085 -145.355 ;
        RECT 63.755 -147.045 64.085 -146.715 ;
        RECT 63.755 -148.405 64.085 -148.075 ;
        RECT 63.755 -149.765 64.085 -149.435 ;
        RECT 63.755 -151.125 64.085 -150.795 ;
        RECT 63.755 -152.485 64.085 -152.155 ;
        RECT 63.755 -153.845 64.085 -153.515 ;
        RECT 63.755 -155.205 64.085 -154.875 ;
        RECT 63.755 -156.565 64.085 -156.235 ;
        RECT 63.755 -157.925 64.085 -157.595 ;
        RECT 63.755 -159.285 64.085 -158.955 ;
        RECT 63.755 -160.645 64.085 -160.315 ;
        RECT 63.755 -162.005 64.085 -161.675 ;
        RECT 63.755 -163.365 64.085 -163.035 ;
        RECT 63.755 -164.725 64.085 -164.395 ;
        RECT 63.755 -166.085 64.085 -165.755 ;
        RECT 63.755 -167.445 64.085 -167.115 ;
        RECT 63.755 -168.805 64.085 -168.475 ;
        RECT 63.755 -170.165 64.085 -169.835 ;
        RECT 63.755 -171.525 64.085 -171.195 ;
        RECT 63.755 -172.885 64.085 -172.555 ;
        RECT 63.755 -174.245 64.085 -173.915 ;
        RECT 63.755 -175.605 64.085 -175.275 ;
        RECT 63.755 -176.965 64.085 -176.635 ;
        RECT 63.755 -178.325 64.085 -177.995 ;
        RECT 63.755 -179.685 64.085 -179.355 ;
        RECT 63.755 -181.045 64.085 -180.715 ;
        RECT 63.755 -182.405 64.085 -182.075 ;
        RECT 63.755 -183.765 64.085 -183.435 ;
        RECT 63.755 -185.125 64.085 -184.795 ;
        RECT 63.755 -186.485 64.085 -186.155 ;
        RECT 63.755 -187.845 64.085 -187.515 ;
        RECT 63.755 -189.205 64.085 -188.875 ;
        RECT 63.755 -190.565 64.085 -190.235 ;
        RECT 63.755 -191.925 64.085 -191.595 ;
        RECT 63.755 -193.285 64.085 -192.955 ;
        RECT 63.755 -194.645 64.085 -194.315 ;
        RECT 63.755 -196.005 64.085 -195.675 ;
        RECT 63.755 -197.365 64.085 -197.035 ;
        RECT 63.755 -198.725 64.085 -198.395 ;
        RECT 63.755 -200.085 64.085 -199.755 ;
        RECT 63.755 -201.445 64.085 -201.115 ;
        RECT 63.755 -202.805 64.085 -202.475 ;
        RECT 63.755 -204.165 64.085 -203.835 ;
        RECT 63.755 -205.525 64.085 -205.195 ;
        RECT 63.755 -206.885 64.085 -206.555 ;
        RECT 63.755 -208.245 64.085 -207.915 ;
        RECT 63.755 -209.605 64.085 -209.275 ;
        RECT 63.755 -210.965 64.085 -210.635 ;
        RECT 63.755 -212.325 64.085 -211.995 ;
        RECT 63.755 -213.685 64.085 -213.355 ;
        RECT 63.755 -215.045 64.085 -214.715 ;
        RECT 63.755 -216.405 64.085 -216.075 ;
        RECT 63.755 -217.765 64.085 -217.435 ;
        RECT 63.755 -219.125 64.085 -218.795 ;
        RECT 63.755 -220.485 64.085 -220.155 ;
        RECT 63.755 -221.845 64.085 -221.515 ;
        RECT 63.755 -223.205 64.085 -222.875 ;
        RECT 63.755 -224.565 64.085 -224.235 ;
        RECT 63.755 -225.925 64.085 -225.595 ;
        RECT 63.755 -227.285 64.085 -226.955 ;
        RECT 63.755 -228.645 64.085 -228.315 ;
        RECT 63.755 -230.005 64.085 -229.675 ;
        RECT 63.755 -231.365 64.085 -231.035 ;
        RECT 63.755 -232.725 64.085 -232.395 ;
        RECT 63.755 -234.085 64.085 -233.755 ;
        RECT 63.755 -235.445 64.085 -235.115 ;
        RECT 63.755 -236.805 64.085 -236.475 ;
        RECT 63.755 -238.165 64.085 -237.835 ;
        RECT 63.755 -243.81 64.085 -242.68 ;
        RECT 63.76 -243.925 64.08 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 246.76 65.445 247.89 ;
        RECT 65.115 241.915 65.445 242.245 ;
        RECT 65.115 240.555 65.445 240.885 ;
        RECT 65.115 239.195 65.445 239.525 ;
        RECT 65.115 237.835 65.445 238.165 ;
        RECT 65.12 237.16 65.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 -1.525 65.445 -1.195 ;
        RECT 65.115 -2.885 65.445 -2.555 ;
        RECT 65.12 -3.56 65.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 -122.565 65.445 -122.235 ;
        RECT 65.115 -123.925 65.445 -123.595 ;
        RECT 65.115 -125.285 65.445 -124.955 ;
        RECT 65.115 -126.645 65.445 -126.315 ;
        RECT 65.115 -128.005 65.445 -127.675 ;
        RECT 65.115 -129.365 65.445 -129.035 ;
        RECT 65.115 -130.725 65.445 -130.395 ;
        RECT 65.115 -132.085 65.445 -131.755 ;
        RECT 65.115 -133.445 65.445 -133.115 ;
        RECT 65.115 -134.805 65.445 -134.475 ;
        RECT 65.115 -136.165 65.445 -135.835 ;
        RECT 65.115 -137.525 65.445 -137.195 ;
        RECT 65.115 -138.885 65.445 -138.555 ;
        RECT 65.115 -140.245 65.445 -139.915 ;
        RECT 65.115 -141.605 65.445 -141.275 ;
        RECT 65.115 -142.965 65.445 -142.635 ;
        RECT 65.115 -144.325 65.445 -143.995 ;
        RECT 65.115 -145.685 65.445 -145.355 ;
        RECT 65.115 -147.045 65.445 -146.715 ;
        RECT 65.115 -148.405 65.445 -148.075 ;
        RECT 65.115 -149.765 65.445 -149.435 ;
        RECT 65.115 -151.125 65.445 -150.795 ;
        RECT 65.115 -152.485 65.445 -152.155 ;
        RECT 65.115 -153.845 65.445 -153.515 ;
        RECT 65.115 -155.205 65.445 -154.875 ;
        RECT 65.115 -156.565 65.445 -156.235 ;
        RECT 65.115 -157.925 65.445 -157.595 ;
        RECT 65.115 -159.285 65.445 -158.955 ;
        RECT 65.115 -160.645 65.445 -160.315 ;
        RECT 65.115 -162.005 65.445 -161.675 ;
        RECT 65.115 -163.365 65.445 -163.035 ;
        RECT 65.115 -164.725 65.445 -164.395 ;
        RECT 65.115 -166.085 65.445 -165.755 ;
        RECT 65.115 -167.445 65.445 -167.115 ;
        RECT 65.115 -168.805 65.445 -168.475 ;
        RECT 65.115 -170.165 65.445 -169.835 ;
        RECT 65.115 -171.525 65.445 -171.195 ;
        RECT 65.115 -172.885 65.445 -172.555 ;
        RECT 65.115 -174.245 65.445 -173.915 ;
        RECT 65.115 -175.605 65.445 -175.275 ;
        RECT 65.115 -176.965 65.445 -176.635 ;
        RECT 65.115 -178.325 65.445 -177.995 ;
        RECT 65.115 -179.685 65.445 -179.355 ;
        RECT 65.115 -181.045 65.445 -180.715 ;
        RECT 65.115 -182.405 65.445 -182.075 ;
        RECT 65.115 -183.765 65.445 -183.435 ;
        RECT 65.115 -185.125 65.445 -184.795 ;
        RECT 65.115 -186.485 65.445 -186.155 ;
        RECT 65.115 -187.845 65.445 -187.515 ;
        RECT 65.115 -189.205 65.445 -188.875 ;
        RECT 65.115 -190.565 65.445 -190.235 ;
        RECT 65.115 -191.925 65.445 -191.595 ;
        RECT 65.115 -193.285 65.445 -192.955 ;
        RECT 65.115 -194.645 65.445 -194.315 ;
        RECT 65.115 -196.005 65.445 -195.675 ;
        RECT 65.115 -197.365 65.445 -197.035 ;
        RECT 65.115 -198.725 65.445 -198.395 ;
        RECT 65.115 -200.085 65.445 -199.755 ;
        RECT 65.115 -201.445 65.445 -201.115 ;
        RECT 65.115 -202.805 65.445 -202.475 ;
        RECT 65.115 -204.165 65.445 -203.835 ;
        RECT 65.115 -205.525 65.445 -205.195 ;
        RECT 65.115 -206.885 65.445 -206.555 ;
        RECT 65.115 -208.245 65.445 -207.915 ;
        RECT 65.115 -209.605 65.445 -209.275 ;
        RECT 65.115 -210.965 65.445 -210.635 ;
        RECT 65.115 -212.325 65.445 -211.995 ;
        RECT 65.115 -213.685 65.445 -213.355 ;
        RECT 65.115 -215.045 65.445 -214.715 ;
        RECT 65.115 -216.405 65.445 -216.075 ;
        RECT 65.115 -217.765 65.445 -217.435 ;
        RECT 65.115 -219.125 65.445 -218.795 ;
        RECT 65.115 -220.485 65.445 -220.155 ;
        RECT 65.115 -221.845 65.445 -221.515 ;
        RECT 65.115 -223.205 65.445 -222.875 ;
        RECT 65.115 -224.565 65.445 -224.235 ;
        RECT 65.115 -225.925 65.445 -225.595 ;
        RECT 65.115 -227.285 65.445 -226.955 ;
        RECT 65.115 -228.645 65.445 -228.315 ;
        RECT 65.115 -230.005 65.445 -229.675 ;
        RECT 65.115 -231.365 65.445 -231.035 ;
        RECT 65.115 -232.725 65.445 -232.395 ;
        RECT 65.115 -234.085 65.445 -233.755 ;
        RECT 65.115 -235.445 65.445 -235.115 ;
        RECT 65.115 -236.805 65.445 -236.475 ;
        RECT 65.115 -238.165 65.445 -237.835 ;
        RECT 65.115 -243.81 65.445 -242.68 ;
        RECT 65.12 -243.925 65.44 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 246.76 66.805 247.89 ;
        RECT 66.475 241.915 66.805 242.245 ;
        RECT 66.475 240.555 66.805 240.885 ;
        RECT 66.475 239.195 66.805 239.525 ;
        RECT 66.475 237.835 66.805 238.165 ;
        RECT 66.48 237.16 66.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 -1.525 66.805 -1.195 ;
        RECT 66.475 -2.885 66.805 -2.555 ;
        RECT 66.48 -3.56 66.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 -122.565 66.805 -122.235 ;
        RECT 66.475 -123.925 66.805 -123.595 ;
        RECT 66.475 -125.285 66.805 -124.955 ;
        RECT 66.475 -126.645 66.805 -126.315 ;
        RECT 66.475 -128.005 66.805 -127.675 ;
        RECT 66.475 -129.365 66.805 -129.035 ;
        RECT 66.475 -130.725 66.805 -130.395 ;
        RECT 66.475 -132.085 66.805 -131.755 ;
        RECT 66.475 -133.445 66.805 -133.115 ;
        RECT 66.475 -134.805 66.805 -134.475 ;
        RECT 66.475 -136.165 66.805 -135.835 ;
        RECT 66.475 -137.525 66.805 -137.195 ;
        RECT 66.475 -138.885 66.805 -138.555 ;
        RECT 66.475 -140.245 66.805 -139.915 ;
        RECT 66.475 -141.605 66.805 -141.275 ;
        RECT 66.475 -142.965 66.805 -142.635 ;
        RECT 66.475 -144.325 66.805 -143.995 ;
        RECT 66.475 -145.685 66.805 -145.355 ;
        RECT 66.475 -147.045 66.805 -146.715 ;
        RECT 66.475 -148.405 66.805 -148.075 ;
        RECT 66.475 -149.765 66.805 -149.435 ;
        RECT 66.475 -151.125 66.805 -150.795 ;
        RECT 66.475 -152.485 66.805 -152.155 ;
        RECT 66.475 -153.845 66.805 -153.515 ;
        RECT 66.475 -155.205 66.805 -154.875 ;
        RECT 66.475 -156.565 66.805 -156.235 ;
        RECT 66.475 -157.925 66.805 -157.595 ;
        RECT 66.475 -159.285 66.805 -158.955 ;
        RECT 66.475 -160.645 66.805 -160.315 ;
        RECT 66.475 -162.005 66.805 -161.675 ;
        RECT 66.475 -163.365 66.805 -163.035 ;
        RECT 66.475 -164.725 66.805 -164.395 ;
        RECT 66.475 -166.085 66.805 -165.755 ;
        RECT 66.475 -167.445 66.805 -167.115 ;
        RECT 66.475 -168.805 66.805 -168.475 ;
        RECT 66.475 -170.165 66.805 -169.835 ;
        RECT 66.475 -171.525 66.805 -171.195 ;
        RECT 66.475 -172.885 66.805 -172.555 ;
        RECT 66.475 -174.245 66.805 -173.915 ;
        RECT 66.475 -175.605 66.805 -175.275 ;
        RECT 66.475 -176.965 66.805 -176.635 ;
        RECT 66.475 -178.325 66.805 -177.995 ;
        RECT 66.475 -179.685 66.805 -179.355 ;
        RECT 66.475 -181.045 66.805 -180.715 ;
        RECT 66.475 -182.405 66.805 -182.075 ;
        RECT 66.475 -183.765 66.805 -183.435 ;
        RECT 66.475 -185.125 66.805 -184.795 ;
        RECT 66.475 -186.485 66.805 -186.155 ;
        RECT 66.475 -187.845 66.805 -187.515 ;
        RECT 66.475 -189.205 66.805 -188.875 ;
        RECT 66.475 -190.565 66.805 -190.235 ;
        RECT 66.475 -191.925 66.805 -191.595 ;
        RECT 66.475 -193.285 66.805 -192.955 ;
        RECT 66.475 -194.645 66.805 -194.315 ;
        RECT 66.475 -196.005 66.805 -195.675 ;
        RECT 66.475 -197.365 66.805 -197.035 ;
        RECT 66.475 -198.725 66.805 -198.395 ;
        RECT 66.475 -200.085 66.805 -199.755 ;
        RECT 66.475 -201.445 66.805 -201.115 ;
        RECT 66.475 -202.805 66.805 -202.475 ;
        RECT 66.475 -204.165 66.805 -203.835 ;
        RECT 66.475 -205.525 66.805 -205.195 ;
        RECT 66.475 -206.885 66.805 -206.555 ;
        RECT 66.475 -208.245 66.805 -207.915 ;
        RECT 66.475 -209.605 66.805 -209.275 ;
        RECT 66.475 -210.965 66.805 -210.635 ;
        RECT 66.475 -212.325 66.805 -211.995 ;
        RECT 66.475 -213.685 66.805 -213.355 ;
        RECT 66.475 -215.045 66.805 -214.715 ;
        RECT 66.475 -216.405 66.805 -216.075 ;
        RECT 66.475 -217.765 66.805 -217.435 ;
        RECT 66.475 -219.125 66.805 -218.795 ;
        RECT 66.475 -220.485 66.805 -220.155 ;
        RECT 66.475 -221.845 66.805 -221.515 ;
        RECT 66.475 -223.205 66.805 -222.875 ;
        RECT 66.475 -224.565 66.805 -224.235 ;
        RECT 66.475 -225.925 66.805 -225.595 ;
        RECT 66.475 -227.285 66.805 -226.955 ;
        RECT 66.475 -228.645 66.805 -228.315 ;
        RECT 66.475 -230.005 66.805 -229.675 ;
        RECT 66.475 -231.365 66.805 -231.035 ;
        RECT 66.475 -232.725 66.805 -232.395 ;
        RECT 66.475 -234.085 66.805 -233.755 ;
        RECT 66.475 -235.445 66.805 -235.115 ;
        RECT 66.475 -236.805 66.805 -236.475 ;
        RECT 66.475 -238.165 66.805 -237.835 ;
        RECT 66.475 -243.81 66.805 -242.68 ;
        RECT 66.48 -243.925 66.8 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 246.76 68.165 247.89 ;
        RECT 67.835 241.915 68.165 242.245 ;
        RECT 67.835 240.555 68.165 240.885 ;
        RECT 67.835 239.195 68.165 239.525 ;
        RECT 67.835 237.835 68.165 238.165 ;
        RECT 67.84 237.16 68.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 -126.645 68.165 -126.315 ;
        RECT 67.835 -128.005 68.165 -127.675 ;
        RECT 67.835 -129.365 68.165 -129.035 ;
        RECT 67.835 -130.725 68.165 -130.395 ;
        RECT 67.835 -132.085 68.165 -131.755 ;
        RECT 67.835 -133.445 68.165 -133.115 ;
        RECT 67.835 -134.805 68.165 -134.475 ;
        RECT 67.835 -136.165 68.165 -135.835 ;
        RECT 67.835 -137.525 68.165 -137.195 ;
        RECT 67.835 -138.885 68.165 -138.555 ;
        RECT 67.835 -140.245 68.165 -139.915 ;
        RECT 67.835 -141.605 68.165 -141.275 ;
        RECT 67.835 -142.965 68.165 -142.635 ;
        RECT 67.835 -144.325 68.165 -143.995 ;
        RECT 67.835 -145.685 68.165 -145.355 ;
        RECT 67.835 -147.045 68.165 -146.715 ;
        RECT 67.835 -148.405 68.165 -148.075 ;
        RECT 67.835 -149.765 68.165 -149.435 ;
        RECT 67.835 -151.125 68.165 -150.795 ;
        RECT 67.835 -152.485 68.165 -152.155 ;
        RECT 67.835 -153.845 68.165 -153.515 ;
        RECT 67.835 -155.205 68.165 -154.875 ;
        RECT 67.835 -156.565 68.165 -156.235 ;
        RECT 67.835 -157.925 68.165 -157.595 ;
        RECT 67.835 -159.285 68.165 -158.955 ;
        RECT 67.835 -160.645 68.165 -160.315 ;
        RECT 67.835 -162.005 68.165 -161.675 ;
        RECT 67.835 -163.365 68.165 -163.035 ;
        RECT 67.835 -164.725 68.165 -164.395 ;
        RECT 67.835 -166.085 68.165 -165.755 ;
        RECT 67.835 -167.445 68.165 -167.115 ;
        RECT 67.835 -168.805 68.165 -168.475 ;
        RECT 67.835 -170.165 68.165 -169.835 ;
        RECT 67.835 -171.525 68.165 -171.195 ;
        RECT 67.835 -172.885 68.165 -172.555 ;
        RECT 67.835 -174.245 68.165 -173.915 ;
        RECT 67.835 -175.605 68.165 -175.275 ;
        RECT 67.835 -176.965 68.165 -176.635 ;
        RECT 67.835 -178.325 68.165 -177.995 ;
        RECT 67.835 -179.685 68.165 -179.355 ;
        RECT 67.835 -181.045 68.165 -180.715 ;
        RECT 67.835 -182.405 68.165 -182.075 ;
        RECT 67.835 -183.765 68.165 -183.435 ;
        RECT 67.835 -185.125 68.165 -184.795 ;
        RECT 67.835 -186.485 68.165 -186.155 ;
        RECT 67.835 -187.845 68.165 -187.515 ;
        RECT 67.835 -189.205 68.165 -188.875 ;
        RECT 67.835 -190.565 68.165 -190.235 ;
        RECT 67.835 -191.925 68.165 -191.595 ;
        RECT 67.835 -193.285 68.165 -192.955 ;
        RECT 67.835 -194.645 68.165 -194.315 ;
        RECT 67.835 -196.005 68.165 -195.675 ;
        RECT 67.835 -197.365 68.165 -197.035 ;
        RECT 67.835 -198.725 68.165 -198.395 ;
        RECT 67.835 -200.085 68.165 -199.755 ;
        RECT 67.835 -201.445 68.165 -201.115 ;
        RECT 67.835 -202.805 68.165 -202.475 ;
        RECT 67.835 -204.165 68.165 -203.835 ;
        RECT 67.835 -205.525 68.165 -205.195 ;
        RECT 67.835 -206.885 68.165 -206.555 ;
        RECT 67.835 -208.245 68.165 -207.915 ;
        RECT 67.835 -209.605 68.165 -209.275 ;
        RECT 67.835 -210.965 68.165 -210.635 ;
        RECT 67.835 -212.325 68.165 -211.995 ;
        RECT 67.835 -213.685 68.165 -213.355 ;
        RECT 67.835 -215.045 68.165 -214.715 ;
        RECT 67.835 -216.405 68.165 -216.075 ;
        RECT 67.835 -217.765 68.165 -217.435 ;
        RECT 67.835 -219.125 68.165 -218.795 ;
        RECT 67.835 -220.485 68.165 -220.155 ;
        RECT 67.835 -221.845 68.165 -221.515 ;
        RECT 67.835 -223.205 68.165 -222.875 ;
        RECT 67.835 -224.565 68.165 -224.235 ;
        RECT 67.835 -225.925 68.165 -225.595 ;
        RECT 67.835 -227.285 68.165 -226.955 ;
        RECT 67.835 -228.645 68.165 -228.315 ;
        RECT 67.835 -230.005 68.165 -229.675 ;
        RECT 67.835 -231.365 68.165 -231.035 ;
        RECT 67.835 -232.725 68.165 -232.395 ;
        RECT 67.835 -234.085 68.165 -233.755 ;
        RECT 67.835 -235.445 68.165 -235.115 ;
        RECT 67.835 -236.805 68.165 -236.475 ;
        RECT 67.835 -238.165 68.165 -237.835 ;
        RECT 67.835 -243.81 68.165 -242.68 ;
        RECT 67.84 -243.925 68.16 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.06 -125.535 68.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 246.76 69.525 247.89 ;
        RECT 69.195 241.915 69.525 242.245 ;
        RECT 69.195 240.555 69.525 240.885 ;
        RECT 69.195 239.195 69.525 239.525 ;
        RECT 69.195 237.835 69.525 238.165 ;
        RECT 69.2 237.16 69.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 246.76 70.885 247.89 ;
        RECT 70.555 241.915 70.885 242.245 ;
        RECT 70.555 240.555 70.885 240.885 ;
        RECT 70.555 239.195 70.885 239.525 ;
        RECT 70.555 237.835 70.885 238.165 ;
        RECT 70.56 237.16 70.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 -1.525 70.885 -1.195 ;
        RECT 70.555 -2.885 70.885 -2.555 ;
        RECT 70.56 -3.56 70.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 246.76 72.245 247.89 ;
        RECT 71.915 241.915 72.245 242.245 ;
        RECT 71.915 240.555 72.245 240.885 ;
        RECT 71.915 239.195 72.245 239.525 ;
        RECT 71.915 237.835 72.245 238.165 ;
        RECT 71.92 237.16 72.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -1.525 72.245 -1.195 ;
        RECT 71.915 -2.885 72.245 -2.555 ;
        RECT 71.92 -3.56 72.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -122.565 72.245 -122.235 ;
        RECT 71.915 -123.925 72.245 -123.595 ;
        RECT 71.915 -125.285 72.245 -124.955 ;
        RECT 71.915 -126.645 72.245 -126.315 ;
        RECT 71.915 -128.005 72.245 -127.675 ;
        RECT 71.915 -129.365 72.245 -129.035 ;
        RECT 71.915 -130.725 72.245 -130.395 ;
        RECT 71.915 -132.085 72.245 -131.755 ;
        RECT 71.915 -133.445 72.245 -133.115 ;
        RECT 71.915 -134.805 72.245 -134.475 ;
        RECT 71.915 -136.165 72.245 -135.835 ;
        RECT 71.915 -137.525 72.245 -137.195 ;
        RECT 71.915 -138.885 72.245 -138.555 ;
        RECT 71.915 -140.245 72.245 -139.915 ;
        RECT 71.915 -141.605 72.245 -141.275 ;
        RECT 71.915 -142.965 72.245 -142.635 ;
        RECT 71.915 -144.325 72.245 -143.995 ;
        RECT 71.915 -145.685 72.245 -145.355 ;
        RECT 71.915 -147.045 72.245 -146.715 ;
        RECT 71.915 -148.405 72.245 -148.075 ;
        RECT 71.915 -149.765 72.245 -149.435 ;
        RECT 71.915 -151.125 72.245 -150.795 ;
        RECT 71.915 -152.485 72.245 -152.155 ;
        RECT 71.915 -153.845 72.245 -153.515 ;
        RECT 71.915 -155.205 72.245 -154.875 ;
        RECT 71.915 -156.565 72.245 -156.235 ;
        RECT 71.915 -157.925 72.245 -157.595 ;
        RECT 71.915 -159.285 72.245 -158.955 ;
        RECT 71.915 -160.645 72.245 -160.315 ;
        RECT 71.915 -162.005 72.245 -161.675 ;
        RECT 71.915 -163.365 72.245 -163.035 ;
        RECT 71.915 -164.725 72.245 -164.395 ;
        RECT 71.915 -166.085 72.245 -165.755 ;
        RECT 71.915 -167.445 72.245 -167.115 ;
        RECT 71.915 -168.805 72.245 -168.475 ;
        RECT 71.915 -170.165 72.245 -169.835 ;
        RECT 71.915 -171.525 72.245 -171.195 ;
        RECT 71.915 -172.885 72.245 -172.555 ;
        RECT 71.915 -174.245 72.245 -173.915 ;
        RECT 71.915 -175.605 72.245 -175.275 ;
        RECT 71.915 -176.965 72.245 -176.635 ;
        RECT 71.915 -178.325 72.245 -177.995 ;
        RECT 71.915 -179.685 72.245 -179.355 ;
        RECT 71.915 -181.045 72.245 -180.715 ;
        RECT 71.915 -182.405 72.245 -182.075 ;
        RECT 71.915 -183.765 72.245 -183.435 ;
        RECT 71.915 -185.125 72.245 -184.795 ;
        RECT 71.915 -186.485 72.245 -186.155 ;
        RECT 71.915 -187.845 72.245 -187.515 ;
        RECT 71.915 -189.205 72.245 -188.875 ;
        RECT 71.915 -190.565 72.245 -190.235 ;
        RECT 71.915 -191.925 72.245 -191.595 ;
        RECT 71.915 -193.285 72.245 -192.955 ;
        RECT 71.915 -194.645 72.245 -194.315 ;
        RECT 71.915 -196.005 72.245 -195.675 ;
        RECT 71.915 -197.365 72.245 -197.035 ;
        RECT 71.915 -198.725 72.245 -198.395 ;
        RECT 71.915 -200.085 72.245 -199.755 ;
        RECT 71.915 -201.445 72.245 -201.115 ;
        RECT 71.915 -202.805 72.245 -202.475 ;
        RECT 71.915 -204.165 72.245 -203.835 ;
        RECT 71.915 -205.525 72.245 -205.195 ;
        RECT 71.915 -206.885 72.245 -206.555 ;
        RECT 71.915 -208.245 72.245 -207.915 ;
        RECT 71.915 -209.605 72.245 -209.275 ;
        RECT 71.915 -210.965 72.245 -210.635 ;
        RECT 71.915 -212.325 72.245 -211.995 ;
        RECT 71.915 -213.685 72.245 -213.355 ;
        RECT 71.915 -215.045 72.245 -214.715 ;
        RECT 71.915 -216.405 72.245 -216.075 ;
        RECT 71.915 -217.765 72.245 -217.435 ;
        RECT 71.915 -219.125 72.245 -218.795 ;
        RECT 71.915 -220.485 72.245 -220.155 ;
        RECT 71.915 -221.845 72.245 -221.515 ;
        RECT 71.915 -223.205 72.245 -222.875 ;
        RECT 71.915 -224.565 72.245 -224.235 ;
        RECT 71.915 -225.925 72.245 -225.595 ;
        RECT 71.915 -227.285 72.245 -226.955 ;
        RECT 71.915 -228.645 72.245 -228.315 ;
        RECT 71.915 -230.005 72.245 -229.675 ;
        RECT 71.915 -231.365 72.245 -231.035 ;
        RECT 71.915 -232.725 72.245 -232.395 ;
        RECT 71.915 -234.085 72.245 -233.755 ;
        RECT 71.915 -235.445 72.245 -235.115 ;
        RECT 71.915 -236.805 72.245 -236.475 ;
        RECT 71.915 -238.165 72.245 -237.835 ;
        RECT 71.915 -243.81 72.245 -242.68 ;
        RECT 71.92 -243.925 72.24 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 246.76 73.605 247.89 ;
        RECT 73.275 241.915 73.605 242.245 ;
        RECT 73.275 240.555 73.605 240.885 ;
        RECT 73.275 239.195 73.605 239.525 ;
        RECT 73.275 237.835 73.605 238.165 ;
        RECT 73.28 237.16 73.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 -1.525 73.605 -1.195 ;
        RECT 73.275 -2.885 73.605 -2.555 ;
        RECT 73.28 -3.56 73.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 -128.005 73.605 -127.675 ;
        RECT 73.275 -129.365 73.605 -129.035 ;
        RECT 73.275 -130.725 73.605 -130.395 ;
        RECT 73.275 -132.085 73.605 -131.755 ;
        RECT 73.275 -133.445 73.605 -133.115 ;
        RECT 73.275 -134.805 73.605 -134.475 ;
        RECT 73.275 -136.165 73.605 -135.835 ;
        RECT 73.275 -137.525 73.605 -137.195 ;
        RECT 73.275 -138.885 73.605 -138.555 ;
        RECT 73.275 -140.245 73.605 -139.915 ;
        RECT 73.275 -141.605 73.605 -141.275 ;
        RECT 73.275 -142.965 73.605 -142.635 ;
        RECT 73.275 -144.325 73.605 -143.995 ;
        RECT 73.275 -145.685 73.605 -145.355 ;
        RECT 73.275 -147.045 73.605 -146.715 ;
        RECT 73.275 -148.405 73.605 -148.075 ;
        RECT 73.275 -149.765 73.605 -149.435 ;
        RECT 73.275 -151.125 73.605 -150.795 ;
        RECT 73.275 -152.485 73.605 -152.155 ;
        RECT 73.275 -153.845 73.605 -153.515 ;
        RECT 73.275 -155.205 73.605 -154.875 ;
        RECT 73.275 -156.565 73.605 -156.235 ;
        RECT 73.275 -157.925 73.605 -157.595 ;
        RECT 73.275 -159.285 73.605 -158.955 ;
        RECT 73.275 -160.645 73.605 -160.315 ;
        RECT 73.275 -162.005 73.605 -161.675 ;
        RECT 73.275 -163.365 73.605 -163.035 ;
        RECT 73.275 -164.725 73.605 -164.395 ;
        RECT 73.275 -166.085 73.605 -165.755 ;
        RECT 73.275 -167.445 73.605 -167.115 ;
        RECT 73.275 -168.805 73.605 -168.475 ;
        RECT 73.275 -170.165 73.605 -169.835 ;
        RECT 73.275 -171.525 73.605 -171.195 ;
        RECT 73.275 -172.885 73.605 -172.555 ;
        RECT 73.275 -174.245 73.605 -173.915 ;
        RECT 73.275 -175.605 73.605 -175.275 ;
        RECT 73.275 -176.965 73.605 -176.635 ;
        RECT 73.275 -178.325 73.605 -177.995 ;
        RECT 73.275 -179.685 73.605 -179.355 ;
        RECT 73.275 -181.045 73.605 -180.715 ;
        RECT 73.275 -182.405 73.605 -182.075 ;
        RECT 73.275 -183.765 73.605 -183.435 ;
        RECT 73.275 -185.125 73.605 -184.795 ;
        RECT 73.275 -186.485 73.605 -186.155 ;
        RECT 73.275 -187.845 73.605 -187.515 ;
        RECT 73.275 -189.205 73.605 -188.875 ;
        RECT 73.275 -190.565 73.605 -190.235 ;
        RECT 73.275 -191.925 73.605 -191.595 ;
        RECT 73.275 -193.285 73.605 -192.955 ;
        RECT 73.275 -194.645 73.605 -194.315 ;
        RECT 73.275 -196.005 73.605 -195.675 ;
        RECT 73.275 -197.365 73.605 -197.035 ;
        RECT 73.275 -198.725 73.605 -198.395 ;
        RECT 73.275 -200.085 73.605 -199.755 ;
        RECT 73.275 -201.445 73.605 -201.115 ;
        RECT 73.275 -202.805 73.605 -202.475 ;
        RECT 73.275 -204.165 73.605 -203.835 ;
        RECT 73.275 -205.525 73.605 -205.195 ;
        RECT 73.275 -206.885 73.605 -206.555 ;
        RECT 73.275 -208.245 73.605 -207.915 ;
        RECT 73.275 -209.605 73.605 -209.275 ;
        RECT 73.275 -210.965 73.605 -210.635 ;
        RECT 73.275 -212.325 73.605 -211.995 ;
        RECT 73.275 -213.685 73.605 -213.355 ;
        RECT 73.275 -215.045 73.605 -214.715 ;
        RECT 73.275 -216.405 73.605 -216.075 ;
        RECT 73.275 -217.765 73.605 -217.435 ;
        RECT 73.275 -219.125 73.605 -218.795 ;
        RECT 73.275 -220.485 73.605 -220.155 ;
        RECT 73.275 -221.845 73.605 -221.515 ;
        RECT 73.275 -223.205 73.605 -222.875 ;
        RECT 73.275 -224.565 73.605 -224.235 ;
        RECT 73.275 -225.925 73.605 -225.595 ;
        RECT 73.275 -227.285 73.605 -226.955 ;
        RECT 73.275 -228.645 73.605 -228.315 ;
        RECT 73.275 -230.005 73.605 -229.675 ;
        RECT 73.275 -231.365 73.605 -231.035 ;
        RECT 73.275 -232.725 73.605 -232.395 ;
        RECT 73.275 -234.085 73.605 -233.755 ;
        RECT 73.275 -235.445 73.605 -235.115 ;
        RECT 73.275 -236.805 73.605 -236.475 ;
        RECT 73.275 -238.165 73.605 -237.835 ;
        RECT 73.275 -243.81 73.605 -242.68 ;
        RECT 73.28 -243.925 73.6 -122.235 ;
        RECT 73.275 -122.565 73.605 -122.235 ;
        RECT 73.275 -123.925 73.605 -123.595 ;
        RECT 73.275 -125.285 73.605 -124.955 ;
        RECT 73.275 -126.645 73.605 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.36 -125.535 35.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 246.76 36.885 247.89 ;
        RECT 36.555 241.915 36.885 242.245 ;
        RECT 36.555 240.555 36.885 240.885 ;
        RECT 36.555 239.195 36.885 239.525 ;
        RECT 36.555 237.835 36.885 238.165 ;
        RECT 36.56 237.16 36.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 246.76 38.245 247.89 ;
        RECT 37.915 241.915 38.245 242.245 ;
        RECT 37.915 240.555 38.245 240.885 ;
        RECT 37.915 239.195 38.245 239.525 ;
        RECT 37.915 237.835 38.245 238.165 ;
        RECT 37.92 237.16 38.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 -1.525 38.245 -1.195 ;
        RECT 37.915 -2.885 38.245 -2.555 ;
        RECT 37.92 -3.56 38.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 246.76 39.605 247.89 ;
        RECT 39.275 241.915 39.605 242.245 ;
        RECT 39.275 240.555 39.605 240.885 ;
        RECT 39.275 239.195 39.605 239.525 ;
        RECT 39.275 237.835 39.605 238.165 ;
        RECT 39.28 237.16 39.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 -1.525 39.605 -1.195 ;
        RECT 39.275 -2.885 39.605 -2.555 ;
        RECT 39.28 -3.56 39.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 -122.565 39.605 -122.235 ;
        RECT 39.275 -123.925 39.605 -123.595 ;
        RECT 39.275 -125.285 39.605 -124.955 ;
        RECT 39.275 -126.645 39.605 -126.315 ;
        RECT 39.275 -128.005 39.605 -127.675 ;
        RECT 39.275 -129.365 39.605 -129.035 ;
        RECT 39.275 -130.725 39.605 -130.395 ;
        RECT 39.275 -132.085 39.605 -131.755 ;
        RECT 39.275 -133.445 39.605 -133.115 ;
        RECT 39.275 -134.805 39.605 -134.475 ;
        RECT 39.275 -136.165 39.605 -135.835 ;
        RECT 39.275 -137.525 39.605 -137.195 ;
        RECT 39.275 -138.885 39.605 -138.555 ;
        RECT 39.275 -140.245 39.605 -139.915 ;
        RECT 39.275 -141.605 39.605 -141.275 ;
        RECT 39.275 -142.965 39.605 -142.635 ;
        RECT 39.275 -144.325 39.605 -143.995 ;
        RECT 39.275 -145.685 39.605 -145.355 ;
        RECT 39.275 -147.045 39.605 -146.715 ;
        RECT 39.275 -148.405 39.605 -148.075 ;
        RECT 39.275 -149.765 39.605 -149.435 ;
        RECT 39.275 -151.125 39.605 -150.795 ;
        RECT 39.275 -152.485 39.605 -152.155 ;
        RECT 39.275 -153.845 39.605 -153.515 ;
        RECT 39.275 -155.205 39.605 -154.875 ;
        RECT 39.275 -156.565 39.605 -156.235 ;
        RECT 39.275 -157.925 39.605 -157.595 ;
        RECT 39.275 -159.285 39.605 -158.955 ;
        RECT 39.275 -160.645 39.605 -160.315 ;
        RECT 39.275 -162.005 39.605 -161.675 ;
        RECT 39.275 -163.365 39.605 -163.035 ;
        RECT 39.275 -164.725 39.605 -164.395 ;
        RECT 39.275 -166.085 39.605 -165.755 ;
        RECT 39.275 -167.445 39.605 -167.115 ;
        RECT 39.275 -168.805 39.605 -168.475 ;
        RECT 39.275 -170.165 39.605 -169.835 ;
        RECT 39.275 -171.525 39.605 -171.195 ;
        RECT 39.275 -172.885 39.605 -172.555 ;
        RECT 39.275 -174.245 39.605 -173.915 ;
        RECT 39.275 -175.605 39.605 -175.275 ;
        RECT 39.275 -176.965 39.605 -176.635 ;
        RECT 39.275 -178.325 39.605 -177.995 ;
        RECT 39.275 -179.685 39.605 -179.355 ;
        RECT 39.275 -181.045 39.605 -180.715 ;
        RECT 39.275 -182.405 39.605 -182.075 ;
        RECT 39.275 -183.765 39.605 -183.435 ;
        RECT 39.275 -185.125 39.605 -184.795 ;
        RECT 39.275 -186.485 39.605 -186.155 ;
        RECT 39.275 -187.845 39.605 -187.515 ;
        RECT 39.275 -189.205 39.605 -188.875 ;
        RECT 39.275 -190.565 39.605 -190.235 ;
        RECT 39.275 -191.925 39.605 -191.595 ;
        RECT 39.275 -193.285 39.605 -192.955 ;
        RECT 39.275 -194.645 39.605 -194.315 ;
        RECT 39.275 -196.005 39.605 -195.675 ;
        RECT 39.275 -197.365 39.605 -197.035 ;
        RECT 39.275 -198.725 39.605 -198.395 ;
        RECT 39.275 -200.085 39.605 -199.755 ;
        RECT 39.275 -201.445 39.605 -201.115 ;
        RECT 39.275 -202.805 39.605 -202.475 ;
        RECT 39.275 -204.165 39.605 -203.835 ;
        RECT 39.275 -205.525 39.605 -205.195 ;
        RECT 39.275 -206.885 39.605 -206.555 ;
        RECT 39.275 -208.245 39.605 -207.915 ;
        RECT 39.275 -209.605 39.605 -209.275 ;
        RECT 39.275 -210.965 39.605 -210.635 ;
        RECT 39.275 -212.325 39.605 -211.995 ;
        RECT 39.275 -213.685 39.605 -213.355 ;
        RECT 39.275 -215.045 39.605 -214.715 ;
        RECT 39.275 -216.405 39.605 -216.075 ;
        RECT 39.275 -217.765 39.605 -217.435 ;
        RECT 39.275 -219.125 39.605 -218.795 ;
        RECT 39.275 -220.485 39.605 -220.155 ;
        RECT 39.275 -221.845 39.605 -221.515 ;
        RECT 39.275 -223.205 39.605 -222.875 ;
        RECT 39.275 -224.565 39.605 -224.235 ;
        RECT 39.275 -225.925 39.605 -225.595 ;
        RECT 39.275 -227.285 39.605 -226.955 ;
        RECT 39.275 -228.645 39.605 -228.315 ;
        RECT 39.275 -230.005 39.605 -229.675 ;
        RECT 39.275 -231.365 39.605 -231.035 ;
        RECT 39.275 -232.725 39.605 -232.395 ;
        RECT 39.275 -234.085 39.605 -233.755 ;
        RECT 39.275 -235.445 39.605 -235.115 ;
        RECT 39.275 -236.805 39.605 -236.475 ;
        RECT 39.275 -238.165 39.605 -237.835 ;
        RECT 39.275 -243.81 39.605 -242.68 ;
        RECT 39.28 -243.925 39.6 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 246.76 40.965 247.89 ;
        RECT 40.635 241.915 40.965 242.245 ;
        RECT 40.635 240.555 40.965 240.885 ;
        RECT 40.635 239.195 40.965 239.525 ;
        RECT 40.635 237.835 40.965 238.165 ;
        RECT 40.64 237.16 40.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 -1.525 40.965 -1.195 ;
        RECT 40.635 -2.885 40.965 -2.555 ;
        RECT 40.64 -3.56 40.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 -122.565 40.965 -122.235 ;
        RECT 40.635 -123.925 40.965 -123.595 ;
        RECT 40.635 -125.285 40.965 -124.955 ;
        RECT 40.635 -126.645 40.965 -126.315 ;
        RECT 40.635 -128.005 40.965 -127.675 ;
        RECT 40.635 -129.365 40.965 -129.035 ;
        RECT 40.635 -130.725 40.965 -130.395 ;
        RECT 40.635 -132.085 40.965 -131.755 ;
        RECT 40.635 -133.445 40.965 -133.115 ;
        RECT 40.635 -134.805 40.965 -134.475 ;
        RECT 40.635 -136.165 40.965 -135.835 ;
        RECT 40.635 -137.525 40.965 -137.195 ;
        RECT 40.635 -138.885 40.965 -138.555 ;
        RECT 40.635 -140.245 40.965 -139.915 ;
        RECT 40.635 -141.605 40.965 -141.275 ;
        RECT 40.635 -142.965 40.965 -142.635 ;
        RECT 40.635 -144.325 40.965 -143.995 ;
        RECT 40.635 -145.685 40.965 -145.355 ;
        RECT 40.635 -147.045 40.965 -146.715 ;
        RECT 40.635 -148.405 40.965 -148.075 ;
        RECT 40.635 -149.765 40.965 -149.435 ;
        RECT 40.635 -151.125 40.965 -150.795 ;
        RECT 40.635 -152.485 40.965 -152.155 ;
        RECT 40.635 -153.845 40.965 -153.515 ;
        RECT 40.635 -155.205 40.965 -154.875 ;
        RECT 40.635 -156.565 40.965 -156.235 ;
        RECT 40.635 -157.925 40.965 -157.595 ;
        RECT 40.635 -159.285 40.965 -158.955 ;
        RECT 40.635 -160.645 40.965 -160.315 ;
        RECT 40.635 -162.005 40.965 -161.675 ;
        RECT 40.635 -163.365 40.965 -163.035 ;
        RECT 40.635 -164.725 40.965 -164.395 ;
        RECT 40.635 -166.085 40.965 -165.755 ;
        RECT 40.635 -167.445 40.965 -167.115 ;
        RECT 40.635 -168.805 40.965 -168.475 ;
        RECT 40.635 -170.165 40.965 -169.835 ;
        RECT 40.635 -171.525 40.965 -171.195 ;
        RECT 40.635 -172.885 40.965 -172.555 ;
        RECT 40.635 -174.245 40.965 -173.915 ;
        RECT 40.635 -175.605 40.965 -175.275 ;
        RECT 40.635 -176.965 40.965 -176.635 ;
        RECT 40.635 -178.325 40.965 -177.995 ;
        RECT 40.635 -179.685 40.965 -179.355 ;
        RECT 40.635 -181.045 40.965 -180.715 ;
        RECT 40.635 -182.405 40.965 -182.075 ;
        RECT 40.635 -183.765 40.965 -183.435 ;
        RECT 40.635 -185.125 40.965 -184.795 ;
        RECT 40.635 -186.485 40.965 -186.155 ;
        RECT 40.635 -187.845 40.965 -187.515 ;
        RECT 40.635 -189.205 40.965 -188.875 ;
        RECT 40.635 -190.565 40.965 -190.235 ;
        RECT 40.635 -191.925 40.965 -191.595 ;
        RECT 40.635 -193.285 40.965 -192.955 ;
        RECT 40.635 -194.645 40.965 -194.315 ;
        RECT 40.635 -196.005 40.965 -195.675 ;
        RECT 40.635 -197.365 40.965 -197.035 ;
        RECT 40.635 -198.725 40.965 -198.395 ;
        RECT 40.635 -200.085 40.965 -199.755 ;
        RECT 40.635 -201.445 40.965 -201.115 ;
        RECT 40.635 -202.805 40.965 -202.475 ;
        RECT 40.635 -204.165 40.965 -203.835 ;
        RECT 40.635 -205.525 40.965 -205.195 ;
        RECT 40.635 -206.885 40.965 -206.555 ;
        RECT 40.635 -208.245 40.965 -207.915 ;
        RECT 40.635 -209.605 40.965 -209.275 ;
        RECT 40.635 -210.965 40.965 -210.635 ;
        RECT 40.635 -212.325 40.965 -211.995 ;
        RECT 40.635 -213.685 40.965 -213.355 ;
        RECT 40.635 -215.045 40.965 -214.715 ;
        RECT 40.635 -216.405 40.965 -216.075 ;
        RECT 40.635 -217.765 40.965 -217.435 ;
        RECT 40.635 -219.125 40.965 -218.795 ;
        RECT 40.635 -220.485 40.965 -220.155 ;
        RECT 40.635 -221.845 40.965 -221.515 ;
        RECT 40.635 -223.205 40.965 -222.875 ;
        RECT 40.635 -224.565 40.965 -224.235 ;
        RECT 40.635 -225.925 40.965 -225.595 ;
        RECT 40.635 -227.285 40.965 -226.955 ;
        RECT 40.635 -228.645 40.965 -228.315 ;
        RECT 40.635 -230.005 40.965 -229.675 ;
        RECT 40.635 -231.365 40.965 -231.035 ;
        RECT 40.635 -232.725 40.965 -232.395 ;
        RECT 40.635 -234.085 40.965 -233.755 ;
        RECT 40.635 -235.445 40.965 -235.115 ;
        RECT 40.635 -236.805 40.965 -236.475 ;
        RECT 40.635 -238.165 40.965 -237.835 ;
        RECT 40.635 -243.81 40.965 -242.68 ;
        RECT 40.64 -243.925 40.96 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 246.76 42.325 247.89 ;
        RECT 41.995 241.915 42.325 242.245 ;
        RECT 41.995 240.555 42.325 240.885 ;
        RECT 41.995 239.195 42.325 239.525 ;
        RECT 41.995 237.835 42.325 238.165 ;
        RECT 42 237.16 42.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 -1.525 42.325 -1.195 ;
        RECT 41.995 -2.885 42.325 -2.555 ;
        RECT 42 -3.56 42.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 -122.565 42.325 -122.235 ;
        RECT 41.995 -123.925 42.325 -123.595 ;
        RECT 41.995 -125.285 42.325 -124.955 ;
        RECT 41.995 -126.645 42.325 -126.315 ;
        RECT 41.995 -128.005 42.325 -127.675 ;
        RECT 41.995 -129.365 42.325 -129.035 ;
        RECT 41.995 -130.725 42.325 -130.395 ;
        RECT 41.995 -132.085 42.325 -131.755 ;
        RECT 41.995 -133.445 42.325 -133.115 ;
        RECT 41.995 -134.805 42.325 -134.475 ;
        RECT 41.995 -136.165 42.325 -135.835 ;
        RECT 41.995 -137.525 42.325 -137.195 ;
        RECT 41.995 -138.885 42.325 -138.555 ;
        RECT 41.995 -140.245 42.325 -139.915 ;
        RECT 41.995 -141.605 42.325 -141.275 ;
        RECT 41.995 -142.965 42.325 -142.635 ;
        RECT 41.995 -144.325 42.325 -143.995 ;
        RECT 41.995 -145.685 42.325 -145.355 ;
        RECT 41.995 -147.045 42.325 -146.715 ;
        RECT 41.995 -148.405 42.325 -148.075 ;
        RECT 41.995 -149.765 42.325 -149.435 ;
        RECT 41.995 -151.125 42.325 -150.795 ;
        RECT 41.995 -152.485 42.325 -152.155 ;
        RECT 41.995 -153.845 42.325 -153.515 ;
        RECT 41.995 -155.205 42.325 -154.875 ;
        RECT 41.995 -156.565 42.325 -156.235 ;
        RECT 41.995 -157.925 42.325 -157.595 ;
        RECT 41.995 -159.285 42.325 -158.955 ;
        RECT 41.995 -160.645 42.325 -160.315 ;
        RECT 41.995 -162.005 42.325 -161.675 ;
        RECT 41.995 -163.365 42.325 -163.035 ;
        RECT 41.995 -164.725 42.325 -164.395 ;
        RECT 41.995 -166.085 42.325 -165.755 ;
        RECT 41.995 -167.445 42.325 -167.115 ;
        RECT 41.995 -168.805 42.325 -168.475 ;
        RECT 41.995 -170.165 42.325 -169.835 ;
        RECT 41.995 -171.525 42.325 -171.195 ;
        RECT 41.995 -172.885 42.325 -172.555 ;
        RECT 41.995 -174.245 42.325 -173.915 ;
        RECT 41.995 -175.605 42.325 -175.275 ;
        RECT 41.995 -176.965 42.325 -176.635 ;
        RECT 41.995 -178.325 42.325 -177.995 ;
        RECT 41.995 -179.685 42.325 -179.355 ;
        RECT 41.995 -181.045 42.325 -180.715 ;
        RECT 41.995 -182.405 42.325 -182.075 ;
        RECT 41.995 -183.765 42.325 -183.435 ;
        RECT 41.995 -185.125 42.325 -184.795 ;
        RECT 41.995 -186.485 42.325 -186.155 ;
        RECT 41.995 -187.845 42.325 -187.515 ;
        RECT 41.995 -189.205 42.325 -188.875 ;
        RECT 41.995 -190.565 42.325 -190.235 ;
        RECT 41.995 -191.925 42.325 -191.595 ;
        RECT 41.995 -193.285 42.325 -192.955 ;
        RECT 41.995 -194.645 42.325 -194.315 ;
        RECT 41.995 -196.005 42.325 -195.675 ;
        RECT 41.995 -197.365 42.325 -197.035 ;
        RECT 41.995 -198.725 42.325 -198.395 ;
        RECT 41.995 -200.085 42.325 -199.755 ;
        RECT 41.995 -201.445 42.325 -201.115 ;
        RECT 41.995 -202.805 42.325 -202.475 ;
        RECT 41.995 -204.165 42.325 -203.835 ;
        RECT 41.995 -205.525 42.325 -205.195 ;
        RECT 41.995 -206.885 42.325 -206.555 ;
        RECT 41.995 -208.245 42.325 -207.915 ;
        RECT 41.995 -209.605 42.325 -209.275 ;
        RECT 41.995 -210.965 42.325 -210.635 ;
        RECT 41.995 -212.325 42.325 -211.995 ;
        RECT 41.995 -213.685 42.325 -213.355 ;
        RECT 41.995 -215.045 42.325 -214.715 ;
        RECT 41.995 -216.405 42.325 -216.075 ;
        RECT 41.995 -217.765 42.325 -217.435 ;
        RECT 41.995 -219.125 42.325 -218.795 ;
        RECT 41.995 -220.485 42.325 -220.155 ;
        RECT 41.995 -221.845 42.325 -221.515 ;
        RECT 41.995 -223.205 42.325 -222.875 ;
        RECT 41.995 -224.565 42.325 -224.235 ;
        RECT 41.995 -225.925 42.325 -225.595 ;
        RECT 41.995 -227.285 42.325 -226.955 ;
        RECT 41.995 -228.645 42.325 -228.315 ;
        RECT 41.995 -230.005 42.325 -229.675 ;
        RECT 41.995 -231.365 42.325 -231.035 ;
        RECT 41.995 -232.725 42.325 -232.395 ;
        RECT 41.995 -234.085 42.325 -233.755 ;
        RECT 41.995 -235.445 42.325 -235.115 ;
        RECT 41.995 -236.805 42.325 -236.475 ;
        RECT 41.995 -238.165 42.325 -237.835 ;
        RECT 41.995 -243.81 42.325 -242.68 ;
        RECT 42 -243.925 42.32 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 246.76 43.685 247.89 ;
        RECT 43.355 241.915 43.685 242.245 ;
        RECT 43.355 240.555 43.685 240.885 ;
        RECT 43.355 239.195 43.685 239.525 ;
        RECT 43.355 237.835 43.685 238.165 ;
        RECT 43.36 237.16 43.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -1.525 43.685 -1.195 ;
        RECT 43.355 -2.885 43.685 -2.555 ;
        RECT 43.36 -3.56 43.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -122.565 43.685 -122.235 ;
        RECT 43.355 -123.925 43.685 -123.595 ;
        RECT 43.355 -125.285 43.685 -124.955 ;
        RECT 43.355 -126.645 43.685 -126.315 ;
        RECT 43.355 -128.005 43.685 -127.675 ;
        RECT 43.355 -129.365 43.685 -129.035 ;
        RECT 43.355 -130.725 43.685 -130.395 ;
        RECT 43.355 -132.085 43.685 -131.755 ;
        RECT 43.355 -133.445 43.685 -133.115 ;
        RECT 43.355 -134.805 43.685 -134.475 ;
        RECT 43.355 -136.165 43.685 -135.835 ;
        RECT 43.355 -137.525 43.685 -137.195 ;
        RECT 43.355 -138.885 43.685 -138.555 ;
        RECT 43.355 -140.245 43.685 -139.915 ;
        RECT 43.355 -141.605 43.685 -141.275 ;
        RECT 43.355 -142.965 43.685 -142.635 ;
        RECT 43.355 -144.325 43.685 -143.995 ;
        RECT 43.355 -145.685 43.685 -145.355 ;
        RECT 43.355 -147.045 43.685 -146.715 ;
        RECT 43.355 -148.405 43.685 -148.075 ;
        RECT 43.355 -149.765 43.685 -149.435 ;
        RECT 43.355 -151.125 43.685 -150.795 ;
        RECT 43.355 -152.485 43.685 -152.155 ;
        RECT 43.355 -153.845 43.685 -153.515 ;
        RECT 43.355 -155.205 43.685 -154.875 ;
        RECT 43.355 -156.565 43.685 -156.235 ;
        RECT 43.355 -157.925 43.685 -157.595 ;
        RECT 43.355 -159.285 43.685 -158.955 ;
        RECT 43.355 -160.645 43.685 -160.315 ;
        RECT 43.355 -162.005 43.685 -161.675 ;
        RECT 43.355 -163.365 43.685 -163.035 ;
        RECT 43.355 -164.725 43.685 -164.395 ;
        RECT 43.355 -166.085 43.685 -165.755 ;
        RECT 43.355 -167.445 43.685 -167.115 ;
        RECT 43.355 -168.805 43.685 -168.475 ;
        RECT 43.355 -170.165 43.685 -169.835 ;
        RECT 43.355 -171.525 43.685 -171.195 ;
        RECT 43.355 -172.885 43.685 -172.555 ;
        RECT 43.355 -174.245 43.685 -173.915 ;
        RECT 43.355 -175.605 43.685 -175.275 ;
        RECT 43.355 -176.965 43.685 -176.635 ;
        RECT 43.355 -178.325 43.685 -177.995 ;
        RECT 43.355 -179.685 43.685 -179.355 ;
        RECT 43.355 -181.045 43.685 -180.715 ;
        RECT 43.355 -182.405 43.685 -182.075 ;
        RECT 43.355 -183.765 43.685 -183.435 ;
        RECT 43.355 -185.125 43.685 -184.795 ;
        RECT 43.355 -186.485 43.685 -186.155 ;
        RECT 43.355 -187.845 43.685 -187.515 ;
        RECT 43.355 -189.205 43.685 -188.875 ;
        RECT 43.355 -190.565 43.685 -190.235 ;
        RECT 43.355 -191.925 43.685 -191.595 ;
        RECT 43.355 -193.285 43.685 -192.955 ;
        RECT 43.355 -194.645 43.685 -194.315 ;
        RECT 43.355 -196.005 43.685 -195.675 ;
        RECT 43.355 -197.365 43.685 -197.035 ;
        RECT 43.355 -198.725 43.685 -198.395 ;
        RECT 43.355 -200.085 43.685 -199.755 ;
        RECT 43.355 -201.445 43.685 -201.115 ;
        RECT 43.355 -202.805 43.685 -202.475 ;
        RECT 43.355 -204.165 43.685 -203.835 ;
        RECT 43.355 -205.525 43.685 -205.195 ;
        RECT 43.355 -206.885 43.685 -206.555 ;
        RECT 43.355 -208.245 43.685 -207.915 ;
        RECT 43.355 -209.605 43.685 -209.275 ;
        RECT 43.355 -210.965 43.685 -210.635 ;
        RECT 43.355 -212.325 43.685 -211.995 ;
        RECT 43.355 -213.685 43.685 -213.355 ;
        RECT 43.355 -215.045 43.685 -214.715 ;
        RECT 43.355 -216.405 43.685 -216.075 ;
        RECT 43.355 -217.765 43.685 -217.435 ;
        RECT 43.355 -219.125 43.685 -218.795 ;
        RECT 43.355 -220.485 43.685 -220.155 ;
        RECT 43.355 -221.845 43.685 -221.515 ;
        RECT 43.355 -223.205 43.685 -222.875 ;
        RECT 43.355 -224.565 43.685 -224.235 ;
        RECT 43.355 -225.925 43.685 -225.595 ;
        RECT 43.355 -227.285 43.685 -226.955 ;
        RECT 43.355 -228.645 43.685 -228.315 ;
        RECT 43.355 -230.005 43.685 -229.675 ;
        RECT 43.355 -231.365 43.685 -231.035 ;
        RECT 43.355 -232.725 43.685 -232.395 ;
        RECT 43.355 -234.085 43.685 -233.755 ;
        RECT 43.355 -235.445 43.685 -235.115 ;
        RECT 43.355 -236.805 43.685 -236.475 ;
        RECT 43.355 -238.165 43.685 -237.835 ;
        RECT 43.355 -243.81 43.685 -242.68 ;
        RECT 43.36 -243.925 43.68 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 246.76 45.045 247.89 ;
        RECT 44.715 241.915 45.045 242.245 ;
        RECT 44.715 240.555 45.045 240.885 ;
        RECT 44.715 239.195 45.045 239.525 ;
        RECT 44.715 237.835 45.045 238.165 ;
        RECT 44.72 237.16 45.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 -1.525 45.045 -1.195 ;
        RECT 44.715 -2.885 45.045 -2.555 ;
        RECT 44.72 -3.56 45.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 -122.565 45.045 -122.235 ;
        RECT 44.715 -123.925 45.045 -123.595 ;
        RECT 44.715 -125.285 45.045 -124.955 ;
        RECT 44.715 -126.645 45.045 -126.315 ;
        RECT 44.715 -128.005 45.045 -127.675 ;
        RECT 44.715 -129.365 45.045 -129.035 ;
        RECT 44.715 -130.725 45.045 -130.395 ;
        RECT 44.715 -132.085 45.045 -131.755 ;
        RECT 44.715 -133.445 45.045 -133.115 ;
        RECT 44.715 -134.805 45.045 -134.475 ;
        RECT 44.715 -136.165 45.045 -135.835 ;
        RECT 44.715 -137.525 45.045 -137.195 ;
        RECT 44.715 -138.885 45.045 -138.555 ;
        RECT 44.715 -140.245 45.045 -139.915 ;
        RECT 44.715 -141.605 45.045 -141.275 ;
        RECT 44.715 -142.965 45.045 -142.635 ;
        RECT 44.715 -144.325 45.045 -143.995 ;
        RECT 44.715 -145.685 45.045 -145.355 ;
        RECT 44.715 -147.045 45.045 -146.715 ;
        RECT 44.715 -148.405 45.045 -148.075 ;
        RECT 44.715 -149.765 45.045 -149.435 ;
        RECT 44.715 -151.125 45.045 -150.795 ;
        RECT 44.715 -152.485 45.045 -152.155 ;
        RECT 44.715 -153.845 45.045 -153.515 ;
        RECT 44.715 -155.205 45.045 -154.875 ;
        RECT 44.715 -156.565 45.045 -156.235 ;
        RECT 44.715 -157.925 45.045 -157.595 ;
        RECT 44.715 -159.285 45.045 -158.955 ;
        RECT 44.715 -160.645 45.045 -160.315 ;
        RECT 44.715 -162.005 45.045 -161.675 ;
        RECT 44.715 -163.365 45.045 -163.035 ;
        RECT 44.715 -164.725 45.045 -164.395 ;
        RECT 44.715 -166.085 45.045 -165.755 ;
        RECT 44.715 -167.445 45.045 -167.115 ;
        RECT 44.715 -168.805 45.045 -168.475 ;
        RECT 44.715 -170.165 45.045 -169.835 ;
        RECT 44.715 -171.525 45.045 -171.195 ;
        RECT 44.715 -172.885 45.045 -172.555 ;
        RECT 44.715 -174.245 45.045 -173.915 ;
        RECT 44.715 -175.605 45.045 -175.275 ;
        RECT 44.715 -176.965 45.045 -176.635 ;
        RECT 44.715 -178.325 45.045 -177.995 ;
        RECT 44.715 -179.685 45.045 -179.355 ;
        RECT 44.715 -181.045 45.045 -180.715 ;
        RECT 44.715 -182.405 45.045 -182.075 ;
        RECT 44.715 -183.765 45.045 -183.435 ;
        RECT 44.715 -185.125 45.045 -184.795 ;
        RECT 44.715 -186.485 45.045 -186.155 ;
        RECT 44.715 -187.845 45.045 -187.515 ;
        RECT 44.715 -189.205 45.045 -188.875 ;
        RECT 44.715 -190.565 45.045 -190.235 ;
        RECT 44.715 -191.925 45.045 -191.595 ;
        RECT 44.715 -193.285 45.045 -192.955 ;
        RECT 44.715 -194.645 45.045 -194.315 ;
        RECT 44.715 -196.005 45.045 -195.675 ;
        RECT 44.715 -197.365 45.045 -197.035 ;
        RECT 44.715 -198.725 45.045 -198.395 ;
        RECT 44.715 -200.085 45.045 -199.755 ;
        RECT 44.715 -201.445 45.045 -201.115 ;
        RECT 44.715 -202.805 45.045 -202.475 ;
        RECT 44.715 -204.165 45.045 -203.835 ;
        RECT 44.715 -205.525 45.045 -205.195 ;
        RECT 44.715 -206.885 45.045 -206.555 ;
        RECT 44.715 -208.245 45.045 -207.915 ;
        RECT 44.715 -209.605 45.045 -209.275 ;
        RECT 44.715 -210.965 45.045 -210.635 ;
        RECT 44.715 -212.325 45.045 -211.995 ;
        RECT 44.715 -213.685 45.045 -213.355 ;
        RECT 44.715 -215.045 45.045 -214.715 ;
        RECT 44.715 -216.405 45.045 -216.075 ;
        RECT 44.715 -217.765 45.045 -217.435 ;
        RECT 44.715 -219.125 45.045 -218.795 ;
        RECT 44.715 -220.485 45.045 -220.155 ;
        RECT 44.715 -221.845 45.045 -221.515 ;
        RECT 44.715 -223.205 45.045 -222.875 ;
        RECT 44.715 -224.565 45.045 -224.235 ;
        RECT 44.715 -225.925 45.045 -225.595 ;
        RECT 44.715 -227.285 45.045 -226.955 ;
        RECT 44.715 -228.645 45.045 -228.315 ;
        RECT 44.715 -230.005 45.045 -229.675 ;
        RECT 44.715 -231.365 45.045 -231.035 ;
        RECT 44.715 -232.725 45.045 -232.395 ;
        RECT 44.715 -234.085 45.045 -233.755 ;
        RECT 44.715 -235.445 45.045 -235.115 ;
        RECT 44.715 -236.805 45.045 -236.475 ;
        RECT 44.715 -238.165 45.045 -237.835 ;
        RECT 44.715 -243.81 45.045 -242.68 ;
        RECT 44.72 -243.925 45.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 246.76 46.405 247.89 ;
        RECT 46.075 241.915 46.405 242.245 ;
        RECT 46.075 240.555 46.405 240.885 ;
        RECT 46.075 239.195 46.405 239.525 ;
        RECT 46.075 237.835 46.405 238.165 ;
        RECT 46.08 237.16 46.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 -126.645 46.405 -126.315 ;
        RECT 46.075 -128.005 46.405 -127.675 ;
        RECT 46.075 -129.365 46.405 -129.035 ;
        RECT 46.075 -130.725 46.405 -130.395 ;
        RECT 46.075 -132.085 46.405 -131.755 ;
        RECT 46.075 -133.445 46.405 -133.115 ;
        RECT 46.075 -134.805 46.405 -134.475 ;
        RECT 46.075 -136.165 46.405 -135.835 ;
        RECT 46.075 -137.525 46.405 -137.195 ;
        RECT 46.075 -138.885 46.405 -138.555 ;
        RECT 46.075 -140.245 46.405 -139.915 ;
        RECT 46.075 -141.605 46.405 -141.275 ;
        RECT 46.075 -142.965 46.405 -142.635 ;
        RECT 46.075 -144.325 46.405 -143.995 ;
        RECT 46.075 -145.685 46.405 -145.355 ;
        RECT 46.075 -147.045 46.405 -146.715 ;
        RECT 46.075 -148.405 46.405 -148.075 ;
        RECT 46.075 -149.765 46.405 -149.435 ;
        RECT 46.075 -151.125 46.405 -150.795 ;
        RECT 46.075 -152.485 46.405 -152.155 ;
        RECT 46.075 -153.845 46.405 -153.515 ;
        RECT 46.075 -155.205 46.405 -154.875 ;
        RECT 46.075 -156.565 46.405 -156.235 ;
        RECT 46.075 -157.925 46.405 -157.595 ;
        RECT 46.075 -159.285 46.405 -158.955 ;
        RECT 46.075 -160.645 46.405 -160.315 ;
        RECT 46.075 -162.005 46.405 -161.675 ;
        RECT 46.075 -163.365 46.405 -163.035 ;
        RECT 46.075 -164.725 46.405 -164.395 ;
        RECT 46.075 -166.085 46.405 -165.755 ;
        RECT 46.075 -167.445 46.405 -167.115 ;
        RECT 46.075 -168.805 46.405 -168.475 ;
        RECT 46.075 -170.165 46.405 -169.835 ;
        RECT 46.075 -171.525 46.405 -171.195 ;
        RECT 46.075 -172.885 46.405 -172.555 ;
        RECT 46.075 -174.245 46.405 -173.915 ;
        RECT 46.075 -175.605 46.405 -175.275 ;
        RECT 46.075 -176.965 46.405 -176.635 ;
        RECT 46.075 -178.325 46.405 -177.995 ;
        RECT 46.075 -179.685 46.405 -179.355 ;
        RECT 46.075 -181.045 46.405 -180.715 ;
        RECT 46.075 -182.405 46.405 -182.075 ;
        RECT 46.075 -183.765 46.405 -183.435 ;
        RECT 46.075 -185.125 46.405 -184.795 ;
        RECT 46.075 -186.485 46.405 -186.155 ;
        RECT 46.075 -187.845 46.405 -187.515 ;
        RECT 46.075 -189.205 46.405 -188.875 ;
        RECT 46.075 -190.565 46.405 -190.235 ;
        RECT 46.075 -191.925 46.405 -191.595 ;
        RECT 46.075 -193.285 46.405 -192.955 ;
        RECT 46.075 -194.645 46.405 -194.315 ;
        RECT 46.075 -196.005 46.405 -195.675 ;
        RECT 46.075 -197.365 46.405 -197.035 ;
        RECT 46.075 -198.725 46.405 -198.395 ;
        RECT 46.075 -200.085 46.405 -199.755 ;
        RECT 46.075 -201.445 46.405 -201.115 ;
        RECT 46.075 -202.805 46.405 -202.475 ;
        RECT 46.075 -204.165 46.405 -203.835 ;
        RECT 46.075 -205.525 46.405 -205.195 ;
        RECT 46.075 -206.885 46.405 -206.555 ;
        RECT 46.075 -208.245 46.405 -207.915 ;
        RECT 46.075 -209.605 46.405 -209.275 ;
        RECT 46.075 -210.965 46.405 -210.635 ;
        RECT 46.075 -212.325 46.405 -211.995 ;
        RECT 46.075 -213.685 46.405 -213.355 ;
        RECT 46.075 -215.045 46.405 -214.715 ;
        RECT 46.075 -216.405 46.405 -216.075 ;
        RECT 46.075 -217.765 46.405 -217.435 ;
        RECT 46.075 -219.125 46.405 -218.795 ;
        RECT 46.075 -220.485 46.405 -220.155 ;
        RECT 46.075 -221.845 46.405 -221.515 ;
        RECT 46.075 -223.205 46.405 -222.875 ;
        RECT 46.075 -224.565 46.405 -224.235 ;
        RECT 46.075 -225.925 46.405 -225.595 ;
        RECT 46.075 -227.285 46.405 -226.955 ;
        RECT 46.075 -228.645 46.405 -228.315 ;
        RECT 46.075 -230.005 46.405 -229.675 ;
        RECT 46.075 -231.365 46.405 -231.035 ;
        RECT 46.075 -232.725 46.405 -232.395 ;
        RECT 46.075 -234.085 46.405 -233.755 ;
        RECT 46.075 -235.445 46.405 -235.115 ;
        RECT 46.075 -236.805 46.405 -236.475 ;
        RECT 46.075 -238.165 46.405 -237.835 ;
        RECT 46.075 -243.81 46.405 -242.68 ;
        RECT 46.08 -243.925 46.4 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.26 -125.535 46.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 246.76 47.765 247.89 ;
        RECT 47.435 241.915 47.765 242.245 ;
        RECT 47.435 240.555 47.765 240.885 ;
        RECT 47.435 239.195 47.765 239.525 ;
        RECT 47.435 237.835 47.765 238.165 ;
        RECT 47.44 237.16 47.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 246.76 49.125 247.89 ;
        RECT 48.795 241.915 49.125 242.245 ;
        RECT 48.795 240.555 49.125 240.885 ;
        RECT 48.795 239.195 49.125 239.525 ;
        RECT 48.795 237.835 49.125 238.165 ;
        RECT 48.8 237.16 49.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 -1.525 49.125 -1.195 ;
        RECT 48.795 -2.885 49.125 -2.555 ;
        RECT 48.8 -3.56 49.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 246.76 50.485 247.89 ;
        RECT 50.155 241.915 50.485 242.245 ;
        RECT 50.155 240.555 50.485 240.885 ;
        RECT 50.155 239.195 50.485 239.525 ;
        RECT 50.155 237.835 50.485 238.165 ;
        RECT 50.16 237.16 50.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -1.525 50.485 -1.195 ;
        RECT 50.155 -2.885 50.485 -2.555 ;
        RECT 50.16 -3.56 50.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -122.565 50.485 -122.235 ;
        RECT 50.155 -123.925 50.485 -123.595 ;
        RECT 50.155 -125.285 50.485 -124.955 ;
        RECT 50.155 -126.645 50.485 -126.315 ;
        RECT 50.155 -128.005 50.485 -127.675 ;
        RECT 50.155 -129.365 50.485 -129.035 ;
        RECT 50.155 -130.725 50.485 -130.395 ;
        RECT 50.155 -132.085 50.485 -131.755 ;
        RECT 50.155 -133.445 50.485 -133.115 ;
        RECT 50.155 -134.805 50.485 -134.475 ;
        RECT 50.155 -136.165 50.485 -135.835 ;
        RECT 50.155 -137.525 50.485 -137.195 ;
        RECT 50.155 -138.885 50.485 -138.555 ;
        RECT 50.155 -140.245 50.485 -139.915 ;
        RECT 50.155 -141.605 50.485 -141.275 ;
        RECT 50.155 -142.965 50.485 -142.635 ;
        RECT 50.155 -144.325 50.485 -143.995 ;
        RECT 50.155 -145.685 50.485 -145.355 ;
        RECT 50.155 -147.045 50.485 -146.715 ;
        RECT 50.155 -148.405 50.485 -148.075 ;
        RECT 50.155 -149.765 50.485 -149.435 ;
        RECT 50.155 -151.125 50.485 -150.795 ;
        RECT 50.155 -152.485 50.485 -152.155 ;
        RECT 50.155 -153.845 50.485 -153.515 ;
        RECT 50.155 -155.205 50.485 -154.875 ;
        RECT 50.155 -156.565 50.485 -156.235 ;
        RECT 50.155 -157.925 50.485 -157.595 ;
        RECT 50.155 -159.285 50.485 -158.955 ;
        RECT 50.155 -160.645 50.485 -160.315 ;
        RECT 50.155 -162.005 50.485 -161.675 ;
        RECT 50.155 -163.365 50.485 -163.035 ;
        RECT 50.155 -164.725 50.485 -164.395 ;
        RECT 50.155 -166.085 50.485 -165.755 ;
        RECT 50.155 -167.445 50.485 -167.115 ;
        RECT 50.155 -168.805 50.485 -168.475 ;
        RECT 50.155 -170.165 50.485 -169.835 ;
        RECT 50.155 -171.525 50.485 -171.195 ;
        RECT 50.155 -172.885 50.485 -172.555 ;
        RECT 50.155 -174.245 50.485 -173.915 ;
        RECT 50.155 -175.605 50.485 -175.275 ;
        RECT 50.155 -176.965 50.485 -176.635 ;
        RECT 50.155 -178.325 50.485 -177.995 ;
        RECT 50.155 -179.685 50.485 -179.355 ;
        RECT 50.155 -181.045 50.485 -180.715 ;
        RECT 50.155 -182.405 50.485 -182.075 ;
        RECT 50.155 -183.765 50.485 -183.435 ;
        RECT 50.155 -185.125 50.485 -184.795 ;
        RECT 50.155 -186.485 50.485 -186.155 ;
        RECT 50.155 -187.845 50.485 -187.515 ;
        RECT 50.155 -189.205 50.485 -188.875 ;
        RECT 50.155 -190.565 50.485 -190.235 ;
        RECT 50.155 -191.925 50.485 -191.595 ;
        RECT 50.155 -193.285 50.485 -192.955 ;
        RECT 50.155 -194.645 50.485 -194.315 ;
        RECT 50.155 -196.005 50.485 -195.675 ;
        RECT 50.155 -197.365 50.485 -197.035 ;
        RECT 50.155 -198.725 50.485 -198.395 ;
        RECT 50.155 -200.085 50.485 -199.755 ;
        RECT 50.155 -201.445 50.485 -201.115 ;
        RECT 50.155 -202.805 50.485 -202.475 ;
        RECT 50.155 -204.165 50.485 -203.835 ;
        RECT 50.155 -205.525 50.485 -205.195 ;
        RECT 50.155 -206.885 50.485 -206.555 ;
        RECT 50.155 -208.245 50.485 -207.915 ;
        RECT 50.155 -209.605 50.485 -209.275 ;
        RECT 50.155 -210.965 50.485 -210.635 ;
        RECT 50.155 -212.325 50.485 -211.995 ;
        RECT 50.155 -213.685 50.485 -213.355 ;
        RECT 50.155 -215.045 50.485 -214.715 ;
        RECT 50.155 -216.405 50.485 -216.075 ;
        RECT 50.155 -217.765 50.485 -217.435 ;
        RECT 50.155 -219.125 50.485 -218.795 ;
        RECT 50.155 -220.485 50.485 -220.155 ;
        RECT 50.155 -221.845 50.485 -221.515 ;
        RECT 50.155 -223.205 50.485 -222.875 ;
        RECT 50.155 -224.565 50.485 -224.235 ;
        RECT 50.155 -225.925 50.485 -225.595 ;
        RECT 50.155 -227.285 50.485 -226.955 ;
        RECT 50.155 -228.645 50.485 -228.315 ;
        RECT 50.155 -230.005 50.485 -229.675 ;
        RECT 50.155 -231.365 50.485 -231.035 ;
        RECT 50.155 -232.725 50.485 -232.395 ;
        RECT 50.155 -234.085 50.485 -233.755 ;
        RECT 50.155 -235.445 50.485 -235.115 ;
        RECT 50.155 -236.805 50.485 -236.475 ;
        RECT 50.155 -238.165 50.485 -237.835 ;
        RECT 50.155 -243.81 50.485 -242.68 ;
        RECT 50.16 -243.925 50.48 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 246.76 51.845 247.89 ;
        RECT 51.515 241.915 51.845 242.245 ;
        RECT 51.515 240.555 51.845 240.885 ;
        RECT 51.515 239.195 51.845 239.525 ;
        RECT 51.515 237.835 51.845 238.165 ;
        RECT 51.52 237.16 51.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 -1.525 51.845 -1.195 ;
        RECT 51.515 -2.885 51.845 -2.555 ;
        RECT 51.52 -3.56 51.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 -122.565 51.845 -122.235 ;
        RECT 51.515 -123.925 51.845 -123.595 ;
        RECT 51.515 -125.285 51.845 -124.955 ;
        RECT 51.515 -126.645 51.845 -126.315 ;
        RECT 51.515 -128.005 51.845 -127.675 ;
        RECT 51.515 -129.365 51.845 -129.035 ;
        RECT 51.515 -130.725 51.845 -130.395 ;
        RECT 51.515 -132.085 51.845 -131.755 ;
        RECT 51.515 -133.445 51.845 -133.115 ;
        RECT 51.515 -134.805 51.845 -134.475 ;
        RECT 51.515 -136.165 51.845 -135.835 ;
        RECT 51.515 -137.525 51.845 -137.195 ;
        RECT 51.515 -138.885 51.845 -138.555 ;
        RECT 51.515 -140.245 51.845 -139.915 ;
        RECT 51.515 -141.605 51.845 -141.275 ;
        RECT 51.515 -142.965 51.845 -142.635 ;
        RECT 51.515 -144.325 51.845 -143.995 ;
        RECT 51.515 -145.685 51.845 -145.355 ;
        RECT 51.515 -147.045 51.845 -146.715 ;
        RECT 51.515 -148.405 51.845 -148.075 ;
        RECT 51.515 -149.765 51.845 -149.435 ;
        RECT 51.515 -151.125 51.845 -150.795 ;
        RECT 51.515 -152.485 51.845 -152.155 ;
        RECT 51.515 -153.845 51.845 -153.515 ;
        RECT 51.515 -155.205 51.845 -154.875 ;
        RECT 51.515 -156.565 51.845 -156.235 ;
        RECT 51.515 -157.925 51.845 -157.595 ;
        RECT 51.515 -159.285 51.845 -158.955 ;
        RECT 51.515 -160.645 51.845 -160.315 ;
        RECT 51.515 -162.005 51.845 -161.675 ;
        RECT 51.515 -163.365 51.845 -163.035 ;
        RECT 51.515 -164.725 51.845 -164.395 ;
        RECT 51.515 -166.085 51.845 -165.755 ;
        RECT 51.515 -167.445 51.845 -167.115 ;
        RECT 51.515 -168.805 51.845 -168.475 ;
        RECT 51.515 -170.165 51.845 -169.835 ;
        RECT 51.515 -171.525 51.845 -171.195 ;
        RECT 51.515 -172.885 51.845 -172.555 ;
        RECT 51.515 -174.245 51.845 -173.915 ;
        RECT 51.515 -175.605 51.845 -175.275 ;
        RECT 51.515 -176.965 51.845 -176.635 ;
        RECT 51.515 -178.325 51.845 -177.995 ;
        RECT 51.515 -179.685 51.845 -179.355 ;
        RECT 51.515 -181.045 51.845 -180.715 ;
        RECT 51.515 -182.405 51.845 -182.075 ;
        RECT 51.515 -183.765 51.845 -183.435 ;
        RECT 51.515 -185.125 51.845 -184.795 ;
        RECT 51.515 -186.485 51.845 -186.155 ;
        RECT 51.515 -187.845 51.845 -187.515 ;
        RECT 51.515 -189.205 51.845 -188.875 ;
        RECT 51.515 -190.565 51.845 -190.235 ;
        RECT 51.515 -191.925 51.845 -191.595 ;
        RECT 51.515 -193.285 51.845 -192.955 ;
        RECT 51.515 -194.645 51.845 -194.315 ;
        RECT 51.515 -196.005 51.845 -195.675 ;
        RECT 51.515 -197.365 51.845 -197.035 ;
        RECT 51.515 -198.725 51.845 -198.395 ;
        RECT 51.515 -200.085 51.845 -199.755 ;
        RECT 51.515 -201.445 51.845 -201.115 ;
        RECT 51.515 -202.805 51.845 -202.475 ;
        RECT 51.515 -204.165 51.845 -203.835 ;
        RECT 51.515 -205.525 51.845 -205.195 ;
        RECT 51.515 -206.885 51.845 -206.555 ;
        RECT 51.515 -208.245 51.845 -207.915 ;
        RECT 51.515 -209.605 51.845 -209.275 ;
        RECT 51.515 -210.965 51.845 -210.635 ;
        RECT 51.515 -212.325 51.845 -211.995 ;
        RECT 51.515 -213.685 51.845 -213.355 ;
        RECT 51.515 -215.045 51.845 -214.715 ;
        RECT 51.515 -216.405 51.845 -216.075 ;
        RECT 51.515 -217.765 51.845 -217.435 ;
        RECT 51.515 -219.125 51.845 -218.795 ;
        RECT 51.515 -220.485 51.845 -220.155 ;
        RECT 51.515 -221.845 51.845 -221.515 ;
        RECT 51.515 -223.205 51.845 -222.875 ;
        RECT 51.515 -224.565 51.845 -224.235 ;
        RECT 51.515 -225.925 51.845 -225.595 ;
        RECT 51.515 -227.285 51.845 -226.955 ;
        RECT 51.515 -228.645 51.845 -228.315 ;
        RECT 51.515 -230.005 51.845 -229.675 ;
        RECT 51.515 -231.365 51.845 -231.035 ;
        RECT 51.515 -232.725 51.845 -232.395 ;
        RECT 51.515 -234.085 51.845 -233.755 ;
        RECT 51.515 -235.445 51.845 -235.115 ;
        RECT 51.515 -236.805 51.845 -236.475 ;
        RECT 51.515 -238.165 51.845 -237.835 ;
        RECT 51.515 -243.81 51.845 -242.68 ;
        RECT 51.52 -243.925 51.84 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 246.76 53.205 247.89 ;
        RECT 52.875 241.915 53.205 242.245 ;
        RECT 52.875 240.555 53.205 240.885 ;
        RECT 52.875 239.195 53.205 239.525 ;
        RECT 52.875 237.835 53.205 238.165 ;
        RECT 52.88 237.16 53.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 -1.525 53.205 -1.195 ;
        RECT 52.875 -2.885 53.205 -2.555 ;
        RECT 52.88 -3.56 53.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 -122.565 53.205 -122.235 ;
        RECT 52.875 -123.925 53.205 -123.595 ;
        RECT 52.875 -125.285 53.205 -124.955 ;
        RECT 52.875 -126.645 53.205 -126.315 ;
        RECT 52.875 -128.005 53.205 -127.675 ;
        RECT 52.875 -129.365 53.205 -129.035 ;
        RECT 52.875 -130.725 53.205 -130.395 ;
        RECT 52.875 -132.085 53.205 -131.755 ;
        RECT 52.875 -133.445 53.205 -133.115 ;
        RECT 52.875 -134.805 53.205 -134.475 ;
        RECT 52.875 -136.165 53.205 -135.835 ;
        RECT 52.875 -137.525 53.205 -137.195 ;
        RECT 52.875 -138.885 53.205 -138.555 ;
        RECT 52.875 -140.245 53.205 -139.915 ;
        RECT 52.875 -141.605 53.205 -141.275 ;
        RECT 52.875 -142.965 53.205 -142.635 ;
        RECT 52.875 -144.325 53.205 -143.995 ;
        RECT 52.875 -145.685 53.205 -145.355 ;
        RECT 52.875 -147.045 53.205 -146.715 ;
        RECT 52.875 -148.405 53.205 -148.075 ;
        RECT 52.875 -149.765 53.205 -149.435 ;
        RECT 52.875 -151.125 53.205 -150.795 ;
        RECT 52.875 -152.485 53.205 -152.155 ;
        RECT 52.875 -153.845 53.205 -153.515 ;
        RECT 52.875 -155.205 53.205 -154.875 ;
        RECT 52.875 -156.565 53.205 -156.235 ;
        RECT 52.875 -157.925 53.205 -157.595 ;
        RECT 52.875 -159.285 53.205 -158.955 ;
        RECT 52.875 -160.645 53.205 -160.315 ;
        RECT 52.875 -162.005 53.205 -161.675 ;
        RECT 52.875 -163.365 53.205 -163.035 ;
        RECT 52.875 -164.725 53.205 -164.395 ;
        RECT 52.875 -166.085 53.205 -165.755 ;
        RECT 52.875 -167.445 53.205 -167.115 ;
        RECT 52.875 -168.805 53.205 -168.475 ;
        RECT 52.875 -170.165 53.205 -169.835 ;
        RECT 52.875 -171.525 53.205 -171.195 ;
        RECT 52.875 -172.885 53.205 -172.555 ;
        RECT 52.875 -174.245 53.205 -173.915 ;
        RECT 52.875 -175.605 53.205 -175.275 ;
        RECT 52.875 -176.965 53.205 -176.635 ;
        RECT 52.875 -178.325 53.205 -177.995 ;
        RECT 52.875 -179.685 53.205 -179.355 ;
        RECT 52.875 -181.045 53.205 -180.715 ;
        RECT 52.875 -182.405 53.205 -182.075 ;
        RECT 52.875 -183.765 53.205 -183.435 ;
        RECT 52.875 -185.125 53.205 -184.795 ;
        RECT 52.875 -186.485 53.205 -186.155 ;
        RECT 52.875 -187.845 53.205 -187.515 ;
        RECT 52.875 -189.205 53.205 -188.875 ;
        RECT 52.875 -190.565 53.205 -190.235 ;
        RECT 52.875 -191.925 53.205 -191.595 ;
        RECT 52.875 -193.285 53.205 -192.955 ;
        RECT 52.875 -194.645 53.205 -194.315 ;
        RECT 52.875 -196.005 53.205 -195.675 ;
        RECT 52.875 -197.365 53.205 -197.035 ;
        RECT 52.875 -198.725 53.205 -198.395 ;
        RECT 52.875 -200.085 53.205 -199.755 ;
        RECT 52.875 -201.445 53.205 -201.115 ;
        RECT 52.875 -202.805 53.205 -202.475 ;
        RECT 52.875 -204.165 53.205 -203.835 ;
        RECT 52.875 -205.525 53.205 -205.195 ;
        RECT 52.875 -206.885 53.205 -206.555 ;
        RECT 52.875 -208.245 53.205 -207.915 ;
        RECT 52.875 -209.605 53.205 -209.275 ;
        RECT 52.875 -210.965 53.205 -210.635 ;
        RECT 52.875 -212.325 53.205 -211.995 ;
        RECT 52.875 -213.685 53.205 -213.355 ;
        RECT 52.875 -215.045 53.205 -214.715 ;
        RECT 52.875 -216.405 53.205 -216.075 ;
        RECT 52.875 -217.765 53.205 -217.435 ;
        RECT 52.875 -219.125 53.205 -218.795 ;
        RECT 52.875 -220.485 53.205 -220.155 ;
        RECT 52.875 -221.845 53.205 -221.515 ;
        RECT 52.875 -223.205 53.205 -222.875 ;
        RECT 52.875 -224.565 53.205 -224.235 ;
        RECT 52.875 -225.925 53.205 -225.595 ;
        RECT 52.875 -227.285 53.205 -226.955 ;
        RECT 52.875 -228.645 53.205 -228.315 ;
        RECT 52.875 -230.005 53.205 -229.675 ;
        RECT 52.875 -231.365 53.205 -231.035 ;
        RECT 52.875 -232.725 53.205 -232.395 ;
        RECT 52.875 -234.085 53.205 -233.755 ;
        RECT 52.875 -235.445 53.205 -235.115 ;
        RECT 52.875 -236.805 53.205 -236.475 ;
        RECT 52.875 -238.165 53.205 -237.835 ;
        RECT 52.875 -243.81 53.205 -242.68 ;
        RECT 52.88 -243.925 53.2 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 246.76 54.565 247.89 ;
        RECT 54.235 241.915 54.565 242.245 ;
        RECT 54.235 240.555 54.565 240.885 ;
        RECT 54.235 239.195 54.565 239.525 ;
        RECT 54.235 237.835 54.565 238.165 ;
        RECT 54.24 237.16 54.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 -1.525 54.565 -1.195 ;
        RECT 54.235 -2.885 54.565 -2.555 ;
        RECT 54.24 -3.56 54.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 -141.605 54.565 -141.275 ;
        RECT 54.235 -142.965 54.565 -142.635 ;
        RECT 54.235 -144.325 54.565 -143.995 ;
        RECT 54.235 -145.685 54.565 -145.355 ;
        RECT 54.235 -147.045 54.565 -146.715 ;
        RECT 54.235 -148.405 54.565 -148.075 ;
        RECT 54.235 -149.765 54.565 -149.435 ;
        RECT 54.235 -151.125 54.565 -150.795 ;
        RECT 54.235 -152.485 54.565 -152.155 ;
        RECT 54.235 -153.845 54.565 -153.515 ;
        RECT 54.235 -155.205 54.565 -154.875 ;
        RECT 54.235 -156.565 54.565 -156.235 ;
        RECT 54.235 -157.925 54.565 -157.595 ;
        RECT 54.235 -159.285 54.565 -158.955 ;
        RECT 54.235 -160.645 54.565 -160.315 ;
        RECT 54.235 -162.005 54.565 -161.675 ;
        RECT 54.235 -163.365 54.565 -163.035 ;
        RECT 54.235 -164.725 54.565 -164.395 ;
        RECT 54.235 -166.085 54.565 -165.755 ;
        RECT 54.235 -167.445 54.565 -167.115 ;
        RECT 54.235 -168.805 54.565 -168.475 ;
        RECT 54.235 -170.165 54.565 -169.835 ;
        RECT 54.235 -171.525 54.565 -171.195 ;
        RECT 54.235 -172.885 54.565 -172.555 ;
        RECT 54.235 -174.245 54.565 -173.915 ;
        RECT 54.235 -175.605 54.565 -175.275 ;
        RECT 54.235 -176.965 54.565 -176.635 ;
        RECT 54.235 -178.325 54.565 -177.995 ;
        RECT 54.235 -179.685 54.565 -179.355 ;
        RECT 54.235 -181.045 54.565 -180.715 ;
        RECT 54.235 -182.405 54.565 -182.075 ;
        RECT 54.235 -183.765 54.565 -183.435 ;
        RECT 54.235 -185.125 54.565 -184.795 ;
        RECT 54.235 -186.485 54.565 -186.155 ;
        RECT 54.235 -187.845 54.565 -187.515 ;
        RECT 54.235 -189.205 54.565 -188.875 ;
        RECT 54.235 -190.565 54.565 -190.235 ;
        RECT 54.235 -191.925 54.565 -191.595 ;
        RECT 54.235 -193.285 54.565 -192.955 ;
        RECT 54.235 -194.645 54.565 -194.315 ;
        RECT 54.235 -196.005 54.565 -195.675 ;
        RECT 54.235 -197.365 54.565 -197.035 ;
        RECT 54.235 -198.725 54.565 -198.395 ;
        RECT 54.235 -200.085 54.565 -199.755 ;
        RECT 54.235 -201.445 54.565 -201.115 ;
        RECT 54.235 -202.805 54.565 -202.475 ;
        RECT 54.235 -204.165 54.565 -203.835 ;
        RECT 54.235 -205.525 54.565 -205.195 ;
        RECT 54.235 -206.885 54.565 -206.555 ;
        RECT 54.235 -208.245 54.565 -207.915 ;
        RECT 54.235 -209.605 54.565 -209.275 ;
        RECT 54.235 -210.965 54.565 -210.635 ;
        RECT 54.235 -212.325 54.565 -211.995 ;
        RECT 54.235 -213.685 54.565 -213.355 ;
        RECT 54.235 -215.045 54.565 -214.715 ;
        RECT 54.235 -216.405 54.565 -216.075 ;
        RECT 54.235 -217.765 54.565 -217.435 ;
        RECT 54.235 -219.125 54.565 -218.795 ;
        RECT 54.235 -220.485 54.565 -220.155 ;
        RECT 54.235 -221.845 54.565 -221.515 ;
        RECT 54.235 -223.205 54.565 -222.875 ;
        RECT 54.235 -224.565 54.565 -224.235 ;
        RECT 54.235 -225.925 54.565 -225.595 ;
        RECT 54.235 -227.285 54.565 -226.955 ;
        RECT 54.235 -228.645 54.565 -228.315 ;
        RECT 54.235 -230.005 54.565 -229.675 ;
        RECT 54.235 -231.365 54.565 -231.035 ;
        RECT 54.235 -232.725 54.565 -232.395 ;
        RECT 54.235 -234.085 54.565 -233.755 ;
        RECT 54.235 -235.445 54.565 -235.115 ;
        RECT 54.235 -236.805 54.565 -236.475 ;
        RECT 54.235 -238.165 54.565 -237.835 ;
        RECT 54.235 -243.81 54.565 -242.68 ;
        RECT 54.24 -243.925 54.56 -122.235 ;
        RECT 54.235 -122.565 54.565 -122.235 ;
        RECT 54.235 -123.925 54.565 -123.595 ;
        RECT 54.235 -125.285 54.565 -124.955 ;
        RECT 54.235 -126.645 54.565 -126.315 ;
        RECT 54.235 -128.005 54.565 -127.675 ;
        RECT 54.235 -129.365 54.565 -129.035 ;
        RECT 54.235 -130.725 54.565 -130.395 ;
        RECT 54.235 -132.085 54.565 -131.755 ;
        RECT 54.235 -133.445 54.565 -133.115 ;
        RECT 54.235 -134.805 54.565 -134.475 ;
        RECT 54.235 -136.165 54.565 -135.835 ;
        RECT 54.235 -137.525 54.565 -137.195 ;
        RECT 54.235 -138.885 54.565 -138.555 ;
        RECT 54.235 -140.245 54.565 -139.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 246.76 20.565 247.89 ;
        RECT 20.235 241.915 20.565 242.245 ;
        RECT 20.235 240.555 20.565 240.885 ;
        RECT 20.235 239.195 20.565 239.525 ;
        RECT 20.235 237.835 20.565 238.165 ;
        RECT 20.24 237.16 20.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -1.525 20.565 -1.195 ;
        RECT 20.235 -2.885 20.565 -2.555 ;
        RECT 20.24 -3.56 20.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -122.565 20.565 -122.235 ;
        RECT 20.235 -123.925 20.565 -123.595 ;
        RECT 20.235 -125.285 20.565 -124.955 ;
        RECT 20.235 -126.645 20.565 -126.315 ;
        RECT 20.235 -128.005 20.565 -127.675 ;
        RECT 20.235 -129.365 20.565 -129.035 ;
        RECT 20.235 -130.725 20.565 -130.395 ;
        RECT 20.235 -132.085 20.565 -131.755 ;
        RECT 20.235 -133.445 20.565 -133.115 ;
        RECT 20.235 -134.805 20.565 -134.475 ;
        RECT 20.235 -136.165 20.565 -135.835 ;
        RECT 20.235 -137.525 20.565 -137.195 ;
        RECT 20.235 -138.885 20.565 -138.555 ;
        RECT 20.235 -140.245 20.565 -139.915 ;
        RECT 20.235 -141.605 20.565 -141.275 ;
        RECT 20.235 -142.965 20.565 -142.635 ;
        RECT 20.235 -144.325 20.565 -143.995 ;
        RECT 20.235 -145.685 20.565 -145.355 ;
        RECT 20.235 -147.045 20.565 -146.715 ;
        RECT 20.235 -148.405 20.565 -148.075 ;
        RECT 20.235 -149.765 20.565 -149.435 ;
        RECT 20.235 -151.125 20.565 -150.795 ;
        RECT 20.235 -152.485 20.565 -152.155 ;
        RECT 20.235 -153.845 20.565 -153.515 ;
        RECT 20.235 -155.205 20.565 -154.875 ;
        RECT 20.235 -156.565 20.565 -156.235 ;
        RECT 20.235 -157.925 20.565 -157.595 ;
        RECT 20.235 -159.285 20.565 -158.955 ;
        RECT 20.235 -160.645 20.565 -160.315 ;
        RECT 20.235 -162.005 20.565 -161.675 ;
        RECT 20.235 -163.365 20.565 -163.035 ;
        RECT 20.235 -164.725 20.565 -164.395 ;
        RECT 20.235 -166.085 20.565 -165.755 ;
        RECT 20.235 -167.445 20.565 -167.115 ;
        RECT 20.235 -168.805 20.565 -168.475 ;
        RECT 20.235 -170.165 20.565 -169.835 ;
        RECT 20.235 -171.525 20.565 -171.195 ;
        RECT 20.235 -172.885 20.565 -172.555 ;
        RECT 20.235 -174.245 20.565 -173.915 ;
        RECT 20.235 -175.605 20.565 -175.275 ;
        RECT 20.235 -176.965 20.565 -176.635 ;
        RECT 20.235 -178.325 20.565 -177.995 ;
        RECT 20.235 -179.685 20.565 -179.355 ;
        RECT 20.235 -181.045 20.565 -180.715 ;
        RECT 20.235 -182.405 20.565 -182.075 ;
        RECT 20.235 -183.765 20.565 -183.435 ;
        RECT 20.235 -185.125 20.565 -184.795 ;
        RECT 20.235 -186.485 20.565 -186.155 ;
        RECT 20.235 -187.845 20.565 -187.515 ;
        RECT 20.235 -189.205 20.565 -188.875 ;
        RECT 20.235 -190.565 20.565 -190.235 ;
        RECT 20.235 -191.925 20.565 -191.595 ;
        RECT 20.235 -193.285 20.565 -192.955 ;
        RECT 20.235 -194.645 20.565 -194.315 ;
        RECT 20.235 -196.005 20.565 -195.675 ;
        RECT 20.235 -197.365 20.565 -197.035 ;
        RECT 20.235 -198.725 20.565 -198.395 ;
        RECT 20.235 -200.085 20.565 -199.755 ;
        RECT 20.235 -201.445 20.565 -201.115 ;
        RECT 20.235 -202.805 20.565 -202.475 ;
        RECT 20.235 -204.165 20.565 -203.835 ;
        RECT 20.235 -205.525 20.565 -205.195 ;
        RECT 20.235 -206.885 20.565 -206.555 ;
        RECT 20.235 -208.245 20.565 -207.915 ;
        RECT 20.235 -209.605 20.565 -209.275 ;
        RECT 20.235 -210.965 20.565 -210.635 ;
        RECT 20.235 -212.325 20.565 -211.995 ;
        RECT 20.235 -213.685 20.565 -213.355 ;
        RECT 20.235 -215.045 20.565 -214.715 ;
        RECT 20.235 -216.405 20.565 -216.075 ;
        RECT 20.235 -217.765 20.565 -217.435 ;
        RECT 20.235 -219.125 20.565 -218.795 ;
        RECT 20.235 -220.485 20.565 -220.155 ;
        RECT 20.235 -221.845 20.565 -221.515 ;
        RECT 20.235 -223.205 20.565 -222.875 ;
        RECT 20.235 -224.565 20.565 -224.235 ;
        RECT 20.235 -225.925 20.565 -225.595 ;
        RECT 20.235 -227.285 20.565 -226.955 ;
        RECT 20.235 -228.645 20.565 -228.315 ;
        RECT 20.235 -230.005 20.565 -229.675 ;
        RECT 20.235 -231.365 20.565 -231.035 ;
        RECT 20.235 -232.725 20.565 -232.395 ;
        RECT 20.235 -234.085 20.565 -233.755 ;
        RECT 20.235 -235.445 20.565 -235.115 ;
        RECT 20.235 -236.805 20.565 -236.475 ;
        RECT 20.235 -238.165 20.565 -237.835 ;
        RECT 20.235 -243.81 20.565 -242.68 ;
        RECT 20.24 -243.925 20.56 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 246.76 21.925 247.89 ;
        RECT 21.595 241.915 21.925 242.245 ;
        RECT 21.595 240.555 21.925 240.885 ;
        RECT 21.595 239.195 21.925 239.525 ;
        RECT 21.595 237.835 21.925 238.165 ;
        RECT 21.6 237.16 21.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 -1.525 21.925 -1.195 ;
        RECT 21.595 -2.885 21.925 -2.555 ;
        RECT 21.6 -3.56 21.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 -122.565 21.925 -122.235 ;
        RECT 21.595 -123.925 21.925 -123.595 ;
        RECT 21.595 -125.285 21.925 -124.955 ;
        RECT 21.595 -126.645 21.925 -126.315 ;
        RECT 21.595 -128.005 21.925 -127.675 ;
        RECT 21.595 -129.365 21.925 -129.035 ;
        RECT 21.595 -130.725 21.925 -130.395 ;
        RECT 21.595 -132.085 21.925 -131.755 ;
        RECT 21.595 -133.445 21.925 -133.115 ;
        RECT 21.595 -134.805 21.925 -134.475 ;
        RECT 21.595 -136.165 21.925 -135.835 ;
        RECT 21.595 -137.525 21.925 -137.195 ;
        RECT 21.595 -138.885 21.925 -138.555 ;
        RECT 21.595 -140.245 21.925 -139.915 ;
        RECT 21.595 -141.605 21.925 -141.275 ;
        RECT 21.595 -142.965 21.925 -142.635 ;
        RECT 21.595 -144.325 21.925 -143.995 ;
        RECT 21.595 -145.685 21.925 -145.355 ;
        RECT 21.595 -147.045 21.925 -146.715 ;
        RECT 21.595 -148.405 21.925 -148.075 ;
        RECT 21.595 -149.765 21.925 -149.435 ;
        RECT 21.595 -151.125 21.925 -150.795 ;
        RECT 21.595 -152.485 21.925 -152.155 ;
        RECT 21.595 -153.845 21.925 -153.515 ;
        RECT 21.595 -155.205 21.925 -154.875 ;
        RECT 21.595 -156.565 21.925 -156.235 ;
        RECT 21.595 -157.925 21.925 -157.595 ;
        RECT 21.595 -159.285 21.925 -158.955 ;
        RECT 21.595 -160.645 21.925 -160.315 ;
        RECT 21.595 -162.005 21.925 -161.675 ;
        RECT 21.595 -163.365 21.925 -163.035 ;
        RECT 21.595 -164.725 21.925 -164.395 ;
        RECT 21.595 -166.085 21.925 -165.755 ;
        RECT 21.595 -167.445 21.925 -167.115 ;
        RECT 21.595 -168.805 21.925 -168.475 ;
        RECT 21.595 -170.165 21.925 -169.835 ;
        RECT 21.595 -171.525 21.925 -171.195 ;
        RECT 21.595 -172.885 21.925 -172.555 ;
        RECT 21.595 -174.245 21.925 -173.915 ;
        RECT 21.595 -175.605 21.925 -175.275 ;
        RECT 21.595 -176.965 21.925 -176.635 ;
        RECT 21.595 -178.325 21.925 -177.995 ;
        RECT 21.595 -179.685 21.925 -179.355 ;
        RECT 21.595 -181.045 21.925 -180.715 ;
        RECT 21.595 -182.405 21.925 -182.075 ;
        RECT 21.595 -183.765 21.925 -183.435 ;
        RECT 21.595 -185.125 21.925 -184.795 ;
        RECT 21.595 -186.485 21.925 -186.155 ;
        RECT 21.595 -187.845 21.925 -187.515 ;
        RECT 21.595 -189.205 21.925 -188.875 ;
        RECT 21.595 -190.565 21.925 -190.235 ;
        RECT 21.595 -191.925 21.925 -191.595 ;
        RECT 21.595 -193.285 21.925 -192.955 ;
        RECT 21.595 -194.645 21.925 -194.315 ;
        RECT 21.595 -196.005 21.925 -195.675 ;
        RECT 21.595 -197.365 21.925 -197.035 ;
        RECT 21.595 -198.725 21.925 -198.395 ;
        RECT 21.595 -200.085 21.925 -199.755 ;
        RECT 21.595 -201.445 21.925 -201.115 ;
        RECT 21.595 -202.805 21.925 -202.475 ;
        RECT 21.595 -204.165 21.925 -203.835 ;
        RECT 21.595 -205.525 21.925 -205.195 ;
        RECT 21.595 -206.885 21.925 -206.555 ;
        RECT 21.595 -208.245 21.925 -207.915 ;
        RECT 21.595 -209.605 21.925 -209.275 ;
        RECT 21.595 -210.965 21.925 -210.635 ;
        RECT 21.595 -212.325 21.925 -211.995 ;
        RECT 21.595 -213.685 21.925 -213.355 ;
        RECT 21.595 -215.045 21.925 -214.715 ;
        RECT 21.595 -216.405 21.925 -216.075 ;
        RECT 21.595 -217.765 21.925 -217.435 ;
        RECT 21.595 -219.125 21.925 -218.795 ;
        RECT 21.595 -220.485 21.925 -220.155 ;
        RECT 21.595 -221.845 21.925 -221.515 ;
        RECT 21.595 -223.205 21.925 -222.875 ;
        RECT 21.595 -224.565 21.925 -224.235 ;
        RECT 21.595 -225.925 21.925 -225.595 ;
        RECT 21.595 -227.285 21.925 -226.955 ;
        RECT 21.595 -228.645 21.925 -228.315 ;
        RECT 21.595 -230.005 21.925 -229.675 ;
        RECT 21.595 -231.365 21.925 -231.035 ;
        RECT 21.595 -232.725 21.925 -232.395 ;
        RECT 21.595 -234.085 21.925 -233.755 ;
        RECT 21.595 -235.445 21.925 -235.115 ;
        RECT 21.595 -236.805 21.925 -236.475 ;
        RECT 21.595 -238.165 21.925 -237.835 ;
        RECT 21.595 -243.81 21.925 -242.68 ;
        RECT 21.6 -243.925 21.92 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 246.76 23.285 247.89 ;
        RECT 22.955 241.915 23.285 242.245 ;
        RECT 22.955 240.555 23.285 240.885 ;
        RECT 22.955 239.195 23.285 239.525 ;
        RECT 22.955 237.835 23.285 238.165 ;
        RECT 22.96 237.16 23.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 -1.525 23.285 -1.195 ;
        RECT 22.955 -2.885 23.285 -2.555 ;
        RECT 22.96 -3.56 23.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 -122.565 23.285 -122.235 ;
        RECT 22.955 -123.925 23.285 -123.595 ;
        RECT 22.955 -125.285 23.285 -124.955 ;
        RECT 22.955 -126.645 23.285 -126.315 ;
        RECT 22.955 -128.005 23.285 -127.675 ;
        RECT 22.955 -129.365 23.285 -129.035 ;
        RECT 22.955 -130.725 23.285 -130.395 ;
        RECT 22.955 -132.085 23.285 -131.755 ;
        RECT 22.955 -133.445 23.285 -133.115 ;
        RECT 22.955 -134.805 23.285 -134.475 ;
        RECT 22.955 -136.165 23.285 -135.835 ;
        RECT 22.955 -137.525 23.285 -137.195 ;
        RECT 22.955 -138.885 23.285 -138.555 ;
        RECT 22.955 -140.245 23.285 -139.915 ;
        RECT 22.955 -141.605 23.285 -141.275 ;
        RECT 22.955 -142.965 23.285 -142.635 ;
        RECT 22.955 -144.325 23.285 -143.995 ;
        RECT 22.955 -145.685 23.285 -145.355 ;
        RECT 22.955 -147.045 23.285 -146.715 ;
        RECT 22.955 -148.405 23.285 -148.075 ;
        RECT 22.955 -149.765 23.285 -149.435 ;
        RECT 22.955 -151.125 23.285 -150.795 ;
        RECT 22.955 -152.485 23.285 -152.155 ;
        RECT 22.955 -153.845 23.285 -153.515 ;
        RECT 22.955 -155.205 23.285 -154.875 ;
        RECT 22.955 -156.565 23.285 -156.235 ;
        RECT 22.955 -157.925 23.285 -157.595 ;
        RECT 22.955 -159.285 23.285 -158.955 ;
        RECT 22.955 -160.645 23.285 -160.315 ;
        RECT 22.955 -162.005 23.285 -161.675 ;
        RECT 22.955 -163.365 23.285 -163.035 ;
        RECT 22.955 -164.725 23.285 -164.395 ;
        RECT 22.955 -166.085 23.285 -165.755 ;
        RECT 22.955 -167.445 23.285 -167.115 ;
        RECT 22.955 -168.805 23.285 -168.475 ;
        RECT 22.955 -170.165 23.285 -169.835 ;
        RECT 22.955 -171.525 23.285 -171.195 ;
        RECT 22.955 -172.885 23.285 -172.555 ;
        RECT 22.955 -174.245 23.285 -173.915 ;
        RECT 22.955 -175.605 23.285 -175.275 ;
        RECT 22.955 -176.965 23.285 -176.635 ;
        RECT 22.955 -178.325 23.285 -177.995 ;
        RECT 22.955 -179.685 23.285 -179.355 ;
        RECT 22.955 -181.045 23.285 -180.715 ;
        RECT 22.955 -182.405 23.285 -182.075 ;
        RECT 22.955 -183.765 23.285 -183.435 ;
        RECT 22.955 -185.125 23.285 -184.795 ;
        RECT 22.955 -186.485 23.285 -186.155 ;
        RECT 22.955 -187.845 23.285 -187.515 ;
        RECT 22.955 -189.205 23.285 -188.875 ;
        RECT 22.955 -190.565 23.285 -190.235 ;
        RECT 22.955 -191.925 23.285 -191.595 ;
        RECT 22.955 -193.285 23.285 -192.955 ;
        RECT 22.955 -194.645 23.285 -194.315 ;
        RECT 22.955 -196.005 23.285 -195.675 ;
        RECT 22.955 -197.365 23.285 -197.035 ;
        RECT 22.955 -198.725 23.285 -198.395 ;
        RECT 22.955 -200.085 23.285 -199.755 ;
        RECT 22.955 -201.445 23.285 -201.115 ;
        RECT 22.955 -202.805 23.285 -202.475 ;
        RECT 22.955 -204.165 23.285 -203.835 ;
        RECT 22.955 -205.525 23.285 -205.195 ;
        RECT 22.955 -206.885 23.285 -206.555 ;
        RECT 22.955 -208.245 23.285 -207.915 ;
        RECT 22.955 -209.605 23.285 -209.275 ;
        RECT 22.955 -210.965 23.285 -210.635 ;
        RECT 22.955 -212.325 23.285 -211.995 ;
        RECT 22.955 -213.685 23.285 -213.355 ;
        RECT 22.955 -215.045 23.285 -214.715 ;
        RECT 22.955 -216.405 23.285 -216.075 ;
        RECT 22.955 -217.765 23.285 -217.435 ;
        RECT 22.955 -219.125 23.285 -218.795 ;
        RECT 22.955 -220.485 23.285 -220.155 ;
        RECT 22.955 -221.845 23.285 -221.515 ;
        RECT 22.955 -223.205 23.285 -222.875 ;
        RECT 22.955 -224.565 23.285 -224.235 ;
        RECT 22.955 -225.925 23.285 -225.595 ;
        RECT 22.955 -227.285 23.285 -226.955 ;
        RECT 22.955 -228.645 23.285 -228.315 ;
        RECT 22.955 -230.005 23.285 -229.675 ;
        RECT 22.955 -231.365 23.285 -231.035 ;
        RECT 22.955 -232.725 23.285 -232.395 ;
        RECT 22.955 -234.085 23.285 -233.755 ;
        RECT 22.955 -235.445 23.285 -235.115 ;
        RECT 22.955 -236.805 23.285 -236.475 ;
        RECT 22.955 -238.165 23.285 -237.835 ;
        RECT 22.955 -243.81 23.285 -242.68 ;
        RECT 22.96 -243.925 23.28 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 246.76 24.645 247.89 ;
        RECT 24.315 241.915 24.645 242.245 ;
        RECT 24.315 240.555 24.645 240.885 ;
        RECT 24.315 239.195 24.645 239.525 ;
        RECT 24.315 237.835 24.645 238.165 ;
        RECT 24.32 237.16 24.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 -126.645 24.645 -126.315 ;
        RECT 24.315 -128.005 24.645 -127.675 ;
        RECT 24.315 -129.365 24.645 -129.035 ;
        RECT 24.315 -130.725 24.645 -130.395 ;
        RECT 24.315 -132.085 24.645 -131.755 ;
        RECT 24.315 -133.445 24.645 -133.115 ;
        RECT 24.315 -134.805 24.645 -134.475 ;
        RECT 24.315 -136.165 24.645 -135.835 ;
        RECT 24.315 -137.525 24.645 -137.195 ;
        RECT 24.315 -138.885 24.645 -138.555 ;
        RECT 24.315 -140.245 24.645 -139.915 ;
        RECT 24.315 -141.605 24.645 -141.275 ;
        RECT 24.315 -142.965 24.645 -142.635 ;
        RECT 24.315 -144.325 24.645 -143.995 ;
        RECT 24.315 -145.685 24.645 -145.355 ;
        RECT 24.315 -147.045 24.645 -146.715 ;
        RECT 24.315 -148.405 24.645 -148.075 ;
        RECT 24.315 -149.765 24.645 -149.435 ;
        RECT 24.315 -151.125 24.645 -150.795 ;
        RECT 24.315 -152.485 24.645 -152.155 ;
        RECT 24.315 -153.845 24.645 -153.515 ;
        RECT 24.315 -155.205 24.645 -154.875 ;
        RECT 24.315 -156.565 24.645 -156.235 ;
        RECT 24.315 -157.925 24.645 -157.595 ;
        RECT 24.315 -159.285 24.645 -158.955 ;
        RECT 24.315 -160.645 24.645 -160.315 ;
        RECT 24.315 -162.005 24.645 -161.675 ;
        RECT 24.315 -163.365 24.645 -163.035 ;
        RECT 24.315 -164.725 24.645 -164.395 ;
        RECT 24.315 -166.085 24.645 -165.755 ;
        RECT 24.315 -167.445 24.645 -167.115 ;
        RECT 24.315 -168.805 24.645 -168.475 ;
        RECT 24.315 -170.165 24.645 -169.835 ;
        RECT 24.315 -171.525 24.645 -171.195 ;
        RECT 24.315 -172.885 24.645 -172.555 ;
        RECT 24.315 -174.245 24.645 -173.915 ;
        RECT 24.315 -175.605 24.645 -175.275 ;
        RECT 24.315 -176.965 24.645 -176.635 ;
        RECT 24.315 -178.325 24.645 -177.995 ;
        RECT 24.315 -179.685 24.645 -179.355 ;
        RECT 24.315 -181.045 24.645 -180.715 ;
        RECT 24.315 -182.405 24.645 -182.075 ;
        RECT 24.315 -183.765 24.645 -183.435 ;
        RECT 24.315 -185.125 24.645 -184.795 ;
        RECT 24.315 -186.485 24.645 -186.155 ;
        RECT 24.315 -187.845 24.645 -187.515 ;
        RECT 24.315 -189.205 24.645 -188.875 ;
        RECT 24.315 -190.565 24.645 -190.235 ;
        RECT 24.315 -191.925 24.645 -191.595 ;
        RECT 24.315 -193.285 24.645 -192.955 ;
        RECT 24.315 -194.645 24.645 -194.315 ;
        RECT 24.315 -196.005 24.645 -195.675 ;
        RECT 24.315 -197.365 24.645 -197.035 ;
        RECT 24.315 -198.725 24.645 -198.395 ;
        RECT 24.315 -200.085 24.645 -199.755 ;
        RECT 24.315 -201.445 24.645 -201.115 ;
        RECT 24.315 -202.805 24.645 -202.475 ;
        RECT 24.315 -204.165 24.645 -203.835 ;
        RECT 24.315 -205.525 24.645 -205.195 ;
        RECT 24.315 -206.885 24.645 -206.555 ;
        RECT 24.315 -208.245 24.645 -207.915 ;
        RECT 24.315 -209.605 24.645 -209.275 ;
        RECT 24.315 -210.965 24.645 -210.635 ;
        RECT 24.315 -212.325 24.645 -211.995 ;
        RECT 24.315 -213.685 24.645 -213.355 ;
        RECT 24.315 -215.045 24.645 -214.715 ;
        RECT 24.315 -216.405 24.645 -216.075 ;
        RECT 24.315 -217.765 24.645 -217.435 ;
        RECT 24.315 -219.125 24.645 -218.795 ;
        RECT 24.315 -220.485 24.645 -220.155 ;
        RECT 24.315 -221.845 24.645 -221.515 ;
        RECT 24.315 -223.205 24.645 -222.875 ;
        RECT 24.315 -224.565 24.645 -224.235 ;
        RECT 24.315 -225.925 24.645 -225.595 ;
        RECT 24.315 -227.285 24.645 -226.955 ;
        RECT 24.315 -228.645 24.645 -228.315 ;
        RECT 24.315 -230.005 24.645 -229.675 ;
        RECT 24.315 -231.365 24.645 -231.035 ;
        RECT 24.315 -232.725 24.645 -232.395 ;
        RECT 24.315 -234.085 24.645 -233.755 ;
        RECT 24.315 -235.445 24.645 -235.115 ;
        RECT 24.315 -236.805 24.645 -236.475 ;
        RECT 24.315 -238.165 24.645 -237.835 ;
        RECT 24.315 -243.81 24.645 -242.68 ;
        RECT 24.32 -243.925 24.64 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.46 -125.535 24.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 246.76 26.005 247.89 ;
        RECT 25.675 241.915 26.005 242.245 ;
        RECT 25.675 240.555 26.005 240.885 ;
        RECT 25.675 239.195 26.005 239.525 ;
        RECT 25.675 237.835 26.005 238.165 ;
        RECT 25.68 237.16 26 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 246.76 27.365 247.89 ;
        RECT 27.035 241.915 27.365 242.245 ;
        RECT 27.035 240.555 27.365 240.885 ;
        RECT 27.035 239.195 27.365 239.525 ;
        RECT 27.035 237.835 27.365 238.165 ;
        RECT 27.04 237.16 27.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 -1.525 27.365 -1.195 ;
        RECT 27.035 -2.885 27.365 -2.555 ;
        RECT 27.04 -3.56 27.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 246.76 28.725 247.89 ;
        RECT 28.395 241.915 28.725 242.245 ;
        RECT 28.395 240.555 28.725 240.885 ;
        RECT 28.395 239.195 28.725 239.525 ;
        RECT 28.395 237.835 28.725 238.165 ;
        RECT 28.4 237.16 28.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -1.525 28.725 -1.195 ;
        RECT 28.395 -2.885 28.725 -2.555 ;
        RECT 28.4 -3.56 28.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -122.565 28.725 -122.235 ;
        RECT 28.395 -123.925 28.725 -123.595 ;
        RECT 28.395 -125.285 28.725 -124.955 ;
        RECT 28.395 -126.645 28.725 -126.315 ;
        RECT 28.395 -128.005 28.725 -127.675 ;
        RECT 28.395 -129.365 28.725 -129.035 ;
        RECT 28.395 -130.725 28.725 -130.395 ;
        RECT 28.395 -132.085 28.725 -131.755 ;
        RECT 28.395 -133.445 28.725 -133.115 ;
        RECT 28.395 -134.805 28.725 -134.475 ;
        RECT 28.395 -136.165 28.725 -135.835 ;
        RECT 28.395 -137.525 28.725 -137.195 ;
        RECT 28.395 -138.885 28.725 -138.555 ;
        RECT 28.395 -140.245 28.725 -139.915 ;
        RECT 28.395 -141.605 28.725 -141.275 ;
        RECT 28.395 -142.965 28.725 -142.635 ;
        RECT 28.395 -144.325 28.725 -143.995 ;
        RECT 28.395 -145.685 28.725 -145.355 ;
        RECT 28.395 -147.045 28.725 -146.715 ;
        RECT 28.395 -148.405 28.725 -148.075 ;
        RECT 28.395 -149.765 28.725 -149.435 ;
        RECT 28.395 -151.125 28.725 -150.795 ;
        RECT 28.395 -152.485 28.725 -152.155 ;
        RECT 28.395 -153.845 28.725 -153.515 ;
        RECT 28.395 -155.205 28.725 -154.875 ;
        RECT 28.395 -156.565 28.725 -156.235 ;
        RECT 28.395 -157.925 28.725 -157.595 ;
        RECT 28.395 -159.285 28.725 -158.955 ;
        RECT 28.395 -160.645 28.725 -160.315 ;
        RECT 28.395 -162.005 28.725 -161.675 ;
        RECT 28.395 -163.365 28.725 -163.035 ;
        RECT 28.395 -164.725 28.725 -164.395 ;
        RECT 28.395 -166.085 28.725 -165.755 ;
        RECT 28.395 -167.445 28.725 -167.115 ;
        RECT 28.395 -168.805 28.725 -168.475 ;
        RECT 28.395 -170.165 28.725 -169.835 ;
        RECT 28.395 -171.525 28.725 -171.195 ;
        RECT 28.395 -172.885 28.725 -172.555 ;
        RECT 28.395 -174.245 28.725 -173.915 ;
        RECT 28.395 -175.605 28.725 -175.275 ;
        RECT 28.395 -176.965 28.725 -176.635 ;
        RECT 28.395 -178.325 28.725 -177.995 ;
        RECT 28.395 -179.685 28.725 -179.355 ;
        RECT 28.395 -181.045 28.725 -180.715 ;
        RECT 28.395 -182.405 28.725 -182.075 ;
        RECT 28.395 -183.765 28.725 -183.435 ;
        RECT 28.395 -185.125 28.725 -184.795 ;
        RECT 28.395 -186.485 28.725 -186.155 ;
        RECT 28.395 -187.845 28.725 -187.515 ;
        RECT 28.395 -189.205 28.725 -188.875 ;
        RECT 28.395 -190.565 28.725 -190.235 ;
        RECT 28.395 -191.925 28.725 -191.595 ;
        RECT 28.395 -193.285 28.725 -192.955 ;
        RECT 28.395 -194.645 28.725 -194.315 ;
        RECT 28.395 -196.005 28.725 -195.675 ;
        RECT 28.395 -197.365 28.725 -197.035 ;
        RECT 28.395 -198.725 28.725 -198.395 ;
        RECT 28.395 -200.085 28.725 -199.755 ;
        RECT 28.395 -201.445 28.725 -201.115 ;
        RECT 28.395 -202.805 28.725 -202.475 ;
        RECT 28.395 -204.165 28.725 -203.835 ;
        RECT 28.395 -205.525 28.725 -205.195 ;
        RECT 28.395 -206.885 28.725 -206.555 ;
        RECT 28.395 -208.245 28.725 -207.915 ;
        RECT 28.395 -209.605 28.725 -209.275 ;
        RECT 28.395 -210.965 28.725 -210.635 ;
        RECT 28.395 -212.325 28.725 -211.995 ;
        RECT 28.395 -213.685 28.725 -213.355 ;
        RECT 28.395 -215.045 28.725 -214.715 ;
        RECT 28.395 -216.405 28.725 -216.075 ;
        RECT 28.395 -217.765 28.725 -217.435 ;
        RECT 28.395 -219.125 28.725 -218.795 ;
        RECT 28.395 -220.485 28.725 -220.155 ;
        RECT 28.395 -221.845 28.725 -221.515 ;
        RECT 28.395 -223.205 28.725 -222.875 ;
        RECT 28.395 -224.565 28.725 -224.235 ;
        RECT 28.395 -225.925 28.725 -225.595 ;
        RECT 28.395 -227.285 28.725 -226.955 ;
        RECT 28.395 -228.645 28.725 -228.315 ;
        RECT 28.395 -230.005 28.725 -229.675 ;
        RECT 28.395 -231.365 28.725 -231.035 ;
        RECT 28.395 -232.725 28.725 -232.395 ;
        RECT 28.395 -234.085 28.725 -233.755 ;
        RECT 28.395 -235.445 28.725 -235.115 ;
        RECT 28.395 -236.805 28.725 -236.475 ;
        RECT 28.395 -238.165 28.725 -237.835 ;
        RECT 28.395 -243.81 28.725 -242.68 ;
        RECT 28.4 -243.925 28.72 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 246.76 30.085 247.89 ;
        RECT 29.755 241.915 30.085 242.245 ;
        RECT 29.755 240.555 30.085 240.885 ;
        RECT 29.755 239.195 30.085 239.525 ;
        RECT 29.755 237.835 30.085 238.165 ;
        RECT 29.76 237.16 30.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -1.525 30.085 -1.195 ;
        RECT 29.755 -2.885 30.085 -2.555 ;
        RECT 29.76 -3.56 30.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -122.565 30.085 -122.235 ;
        RECT 29.755 -123.925 30.085 -123.595 ;
        RECT 29.755 -125.285 30.085 -124.955 ;
        RECT 29.755 -126.645 30.085 -126.315 ;
        RECT 29.755 -128.005 30.085 -127.675 ;
        RECT 29.755 -129.365 30.085 -129.035 ;
        RECT 29.755 -130.725 30.085 -130.395 ;
        RECT 29.755 -132.085 30.085 -131.755 ;
        RECT 29.755 -133.445 30.085 -133.115 ;
        RECT 29.755 -134.805 30.085 -134.475 ;
        RECT 29.755 -136.165 30.085 -135.835 ;
        RECT 29.755 -137.525 30.085 -137.195 ;
        RECT 29.755 -138.885 30.085 -138.555 ;
        RECT 29.755 -140.245 30.085 -139.915 ;
        RECT 29.755 -141.605 30.085 -141.275 ;
        RECT 29.755 -142.965 30.085 -142.635 ;
        RECT 29.755 -144.325 30.085 -143.995 ;
        RECT 29.755 -145.685 30.085 -145.355 ;
        RECT 29.755 -147.045 30.085 -146.715 ;
        RECT 29.755 -148.405 30.085 -148.075 ;
        RECT 29.755 -149.765 30.085 -149.435 ;
        RECT 29.755 -151.125 30.085 -150.795 ;
        RECT 29.755 -152.485 30.085 -152.155 ;
        RECT 29.755 -153.845 30.085 -153.515 ;
        RECT 29.755 -155.205 30.085 -154.875 ;
        RECT 29.755 -156.565 30.085 -156.235 ;
        RECT 29.755 -157.925 30.085 -157.595 ;
        RECT 29.755 -159.285 30.085 -158.955 ;
        RECT 29.755 -160.645 30.085 -160.315 ;
        RECT 29.755 -162.005 30.085 -161.675 ;
        RECT 29.755 -163.365 30.085 -163.035 ;
        RECT 29.755 -164.725 30.085 -164.395 ;
        RECT 29.755 -166.085 30.085 -165.755 ;
        RECT 29.755 -167.445 30.085 -167.115 ;
        RECT 29.755 -168.805 30.085 -168.475 ;
        RECT 29.755 -170.165 30.085 -169.835 ;
        RECT 29.755 -171.525 30.085 -171.195 ;
        RECT 29.755 -172.885 30.085 -172.555 ;
        RECT 29.755 -174.245 30.085 -173.915 ;
        RECT 29.755 -175.605 30.085 -175.275 ;
        RECT 29.755 -176.965 30.085 -176.635 ;
        RECT 29.755 -178.325 30.085 -177.995 ;
        RECT 29.755 -179.685 30.085 -179.355 ;
        RECT 29.755 -181.045 30.085 -180.715 ;
        RECT 29.755 -182.405 30.085 -182.075 ;
        RECT 29.755 -183.765 30.085 -183.435 ;
        RECT 29.755 -185.125 30.085 -184.795 ;
        RECT 29.755 -186.485 30.085 -186.155 ;
        RECT 29.755 -187.845 30.085 -187.515 ;
        RECT 29.755 -189.205 30.085 -188.875 ;
        RECT 29.755 -190.565 30.085 -190.235 ;
        RECT 29.755 -191.925 30.085 -191.595 ;
        RECT 29.755 -193.285 30.085 -192.955 ;
        RECT 29.755 -194.645 30.085 -194.315 ;
        RECT 29.755 -196.005 30.085 -195.675 ;
        RECT 29.755 -197.365 30.085 -197.035 ;
        RECT 29.755 -198.725 30.085 -198.395 ;
        RECT 29.755 -200.085 30.085 -199.755 ;
        RECT 29.755 -201.445 30.085 -201.115 ;
        RECT 29.755 -202.805 30.085 -202.475 ;
        RECT 29.755 -204.165 30.085 -203.835 ;
        RECT 29.755 -205.525 30.085 -205.195 ;
        RECT 29.755 -206.885 30.085 -206.555 ;
        RECT 29.755 -208.245 30.085 -207.915 ;
        RECT 29.755 -209.605 30.085 -209.275 ;
        RECT 29.755 -210.965 30.085 -210.635 ;
        RECT 29.755 -212.325 30.085 -211.995 ;
        RECT 29.755 -213.685 30.085 -213.355 ;
        RECT 29.755 -215.045 30.085 -214.715 ;
        RECT 29.755 -216.405 30.085 -216.075 ;
        RECT 29.755 -217.765 30.085 -217.435 ;
        RECT 29.755 -219.125 30.085 -218.795 ;
        RECT 29.755 -220.485 30.085 -220.155 ;
        RECT 29.755 -221.845 30.085 -221.515 ;
        RECT 29.755 -223.205 30.085 -222.875 ;
        RECT 29.755 -224.565 30.085 -224.235 ;
        RECT 29.755 -225.925 30.085 -225.595 ;
        RECT 29.755 -227.285 30.085 -226.955 ;
        RECT 29.755 -228.645 30.085 -228.315 ;
        RECT 29.755 -230.005 30.085 -229.675 ;
        RECT 29.755 -231.365 30.085 -231.035 ;
        RECT 29.755 -232.725 30.085 -232.395 ;
        RECT 29.755 -234.085 30.085 -233.755 ;
        RECT 29.755 -235.445 30.085 -235.115 ;
        RECT 29.755 -236.805 30.085 -236.475 ;
        RECT 29.755 -238.165 30.085 -237.835 ;
        RECT 29.755 -243.81 30.085 -242.68 ;
        RECT 29.76 -243.925 30.08 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 246.76 31.445 247.89 ;
        RECT 31.115 241.915 31.445 242.245 ;
        RECT 31.115 240.555 31.445 240.885 ;
        RECT 31.115 239.195 31.445 239.525 ;
        RECT 31.115 237.835 31.445 238.165 ;
        RECT 31.12 237.16 31.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -1.525 31.445 -1.195 ;
        RECT 31.115 -2.885 31.445 -2.555 ;
        RECT 31.12 -3.56 31.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -122.565 31.445 -122.235 ;
        RECT 31.115 -123.925 31.445 -123.595 ;
        RECT 31.115 -125.285 31.445 -124.955 ;
        RECT 31.115 -126.645 31.445 -126.315 ;
        RECT 31.115 -128.005 31.445 -127.675 ;
        RECT 31.115 -129.365 31.445 -129.035 ;
        RECT 31.115 -130.725 31.445 -130.395 ;
        RECT 31.115 -132.085 31.445 -131.755 ;
        RECT 31.115 -133.445 31.445 -133.115 ;
        RECT 31.115 -134.805 31.445 -134.475 ;
        RECT 31.115 -136.165 31.445 -135.835 ;
        RECT 31.115 -137.525 31.445 -137.195 ;
        RECT 31.115 -138.885 31.445 -138.555 ;
        RECT 31.115 -140.245 31.445 -139.915 ;
        RECT 31.115 -141.605 31.445 -141.275 ;
        RECT 31.115 -142.965 31.445 -142.635 ;
        RECT 31.115 -144.325 31.445 -143.995 ;
        RECT 31.115 -145.685 31.445 -145.355 ;
        RECT 31.115 -147.045 31.445 -146.715 ;
        RECT 31.115 -148.405 31.445 -148.075 ;
        RECT 31.115 -149.765 31.445 -149.435 ;
        RECT 31.115 -151.125 31.445 -150.795 ;
        RECT 31.115 -152.485 31.445 -152.155 ;
        RECT 31.115 -153.845 31.445 -153.515 ;
        RECT 31.115 -155.205 31.445 -154.875 ;
        RECT 31.115 -156.565 31.445 -156.235 ;
        RECT 31.115 -157.925 31.445 -157.595 ;
        RECT 31.115 -159.285 31.445 -158.955 ;
        RECT 31.115 -160.645 31.445 -160.315 ;
        RECT 31.115 -162.005 31.445 -161.675 ;
        RECT 31.115 -163.365 31.445 -163.035 ;
        RECT 31.115 -164.725 31.445 -164.395 ;
        RECT 31.115 -166.085 31.445 -165.755 ;
        RECT 31.115 -167.445 31.445 -167.115 ;
        RECT 31.115 -168.805 31.445 -168.475 ;
        RECT 31.115 -170.165 31.445 -169.835 ;
        RECT 31.115 -171.525 31.445 -171.195 ;
        RECT 31.115 -172.885 31.445 -172.555 ;
        RECT 31.115 -174.245 31.445 -173.915 ;
        RECT 31.115 -175.605 31.445 -175.275 ;
        RECT 31.115 -176.965 31.445 -176.635 ;
        RECT 31.115 -178.325 31.445 -177.995 ;
        RECT 31.115 -179.685 31.445 -179.355 ;
        RECT 31.115 -181.045 31.445 -180.715 ;
        RECT 31.115 -182.405 31.445 -182.075 ;
        RECT 31.115 -183.765 31.445 -183.435 ;
        RECT 31.115 -185.125 31.445 -184.795 ;
        RECT 31.115 -186.485 31.445 -186.155 ;
        RECT 31.115 -187.845 31.445 -187.515 ;
        RECT 31.115 -189.205 31.445 -188.875 ;
        RECT 31.115 -190.565 31.445 -190.235 ;
        RECT 31.115 -191.925 31.445 -191.595 ;
        RECT 31.115 -193.285 31.445 -192.955 ;
        RECT 31.115 -194.645 31.445 -194.315 ;
        RECT 31.115 -196.005 31.445 -195.675 ;
        RECT 31.115 -197.365 31.445 -197.035 ;
        RECT 31.115 -198.725 31.445 -198.395 ;
        RECT 31.115 -200.085 31.445 -199.755 ;
        RECT 31.115 -201.445 31.445 -201.115 ;
        RECT 31.115 -202.805 31.445 -202.475 ;
        RECT 31.115 -204.165 31.445 -203.835 ;
        RECT 31.115 -205.525 31.445 -205.195 ;
        RECT 31.115 -206.885 31.445 -206.555 ;
        RECT 31.115 -208.245 31.445 -207.915 ;
        RECT 31.115 -209.605 31.445 -209.275 ;
        RECT 31.115 -210.965 31.445 -210.635 ;
        RECT 31.115 -212.325 31.445 -211.995 ;
        RECT 31.115 -213.685 31.445 -213.355 ;
        RECT 31.115 -215.045 31.445 -214.715 ;
        RECT 31.115 -216.405 31.445 -216.075 ;
        RECT 31.115 -217.765 31.445 -217.435 ;
        RECT 31.115 -219.125 31.445 -218.795 ;
        RECT 31.115 -220.485 31.445 -220.155 ;
        RECT 31.115 -221.845 31.445 -221.515 ;
        RECT 31.115 -223.205 31.445 -222.875 ;
        RECT 31.115 -224.565 31.445 -224.235 ;
        RECT 31.115 -225.925 31.445 -225.595 ;
        RECT 31.115 -227.285 31.445 -226.955 ;
        RECT 31.115 -228.645 31.445 -228.315 ;
        RECT 31.115 -230.005 31.445 -229.675 ;
        RECT 31.115 -231.365 31.445 -231.035 ;
        RECT 31.115 -232.725 31.445 -232.395 ;
        RECT 31.115 -234.085 31.445 -233.755 ;
        RECT 31.115 -235.445 31.445 -235.115 ;
        RECT 31.115 -236.805 31.445 -236.475 ;
        RECT 31.115 -238.165 31.445 -237.835 ;
        RECT 31.115 -243.81 31.445 -242.68 ;
        RECT 31.12 -243.925 31.44 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 246.76 32.805 247.89 ;
        RECT 32.475 241.915 32.805 242.245 ;
        RECT 32.475 240.555 32.805 240.885 ;
        RECT 32.475 239.195 32.805 239.525 ;
        RECT 32.475 237.835 32.805 238.165 ;
        RECT 32.48 237.16 32.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -1.525 32.805 -1.195 ;
        RECT 32.475 -2.885 32.805 -2.555 ;
        RECT 32.48 -3.56 32.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -122.565 32.805 -122.235 ;
        RECT 32.475 -123.925 32.805 -123.595 ;
        RECT 32.475 -125.285 32.805 -124.955 ;
        RECT 32.475 -126.645 32.805 -126.315 ;
        RECT 32.475 -128.005 32.805 -127.675 ;
        RECT 32.475 -129.365 32.805 -129.035 ;
        RECT 32.475 -130.725 32.805 -130.395 ;
        RECT 32.475 -132.085 32.805 -131.755 ;
        RECT 32.475 -133.445 32.805 -133.115 ;
        RECT 32.475 -134.805 32.805 -134.475 ;
        RECT 32.475 -136.165 32.805 -135.835 ;
        RECT 32.475 -137.525 32.805 -137.195 ;
        RECT 32.475 -138.885 32.805 -138.555 ;
        RECT 32.475 -140.245 32.805 -139.915 ;
        RECT 32.475 -141.605 32.805 -141.275 ;
        RECT 32.475 -142.965 32.805 -142.635 ;
        RECT 32.475 -144.325 32.805 -143.995 ;
        RECT 32.475 -145.685 32.805 -145.355 ;
        RECT 32.475 -147.045 32.805 -146.715 ;
        RECT 32.475 -148.405 32.805 -148.075 ;
        RECT 32.475 -149.765 32.805 -149.435 ;
        RECT 32.475 -151.125 32.805 -150.795 ;
        RECT 32.475 -152.485 32.805 -152.155 ;
        RECT 32.475 -153.845 32.805 -153.515 ;
        RECT 32.475 -155.205 32.805 -154.875 ;
        RECT 32.475 -156.565 32.805 -156.235 ;
        RECT 32.475 -157.925 32.805 -157.595 ;
        RECT 32.475 -159.285 32.805 -158.955 ;
        RECT 32.475 -160.645 32.805 -160.315 ;
        RECT 32.475 -162.005 32.805 -161.675 ;
        RECT 32.475 -163.365 32.805 -163.035 ;
        RECT 32.475 -164.725 32.805 -164.395 ;
        RECT 32.475 -166.085 32.805 -165.755 ;
        RECT 32.475 -167.445 32.805 -167.115 ;
        RECT 32.475 -168.805 32.805 -168.475 ;
        RECT 32.475 -170.165 32.805 -169.835 ;
        RECT 32.475 -171.525 32.805 -171.195 ;
        RECT 32.475 -172.885 32.805 -172.555 ;
        RECT 32.475 -174.245 32.805 -173.915 ;
        RECT 32.475 -175.605 32.805 -175.275 ;
        RECT 32.475 -176.965 32.805 -176.635 ;
        RECT 32.475 -178.325 32.805 -177.995 ;
        RECT 32.475 -179.685 32.805 -179.355 ;
        RECT 32.475 -181.045 32.805 -180.715 ;
        RECT 32.475 -182.405 32.805 -182.075 ;
        RECT 32.475 -183.765 32.805 -183.435 ;
        RECT 32.475 -185.125 32.805 -184.795 ;
        RECT 32.475 -186.485 32.805 -186.155 ;
        RECT 32.475 -187.845 32.805 -187.515 ;
        RECT 32.475 -189.205 32.805 -188.875 ;
        RECT 32.475 -190.565 32.805 -190.235 ;
        RECT 32.475 -191.925 32.805 -191.595 ;
        RECT 32.475 -193.285 32.805 -192.955 ;
        RECT 32.475 -194.645 32.805 -194.315 ;
        RECT 32.475 -196.005 32.805 -195.675 ;
        RECT 32.475 -197.365 32.805 -197.035 ;
        RECT 32.475 -198.725 32.805 -198.395 ;
        RECT 32.475 -200.085 32.805 -199.755 ;
        RECT 32.475 -201.445 32.805 -201.115 ;
        RECT 32.475 -202.805 32.805 -202.475 ;
        RECT 32.475 -204.165 32.805 -203.835 ;
        RECT 32.475 -205.525 32.805 -205.195 ;
        RECT 32.475 -206.885 32.805 -206.555 ;
        RECT 32.475 -208.245 32.805 -207.915 ;
        RECT 32.475 -209.605 32.805 -209.275 ;
        RECT 32.475 -210.965 32.805 -210.635 ;
        RECT 32.475 -212.325 32.805 -211.995 ;
        RECT 32.475 -213.685 32.805 -213.355 ;
        RECT 32.475 -215.045 32.805 -214.715 ;
        RECT 32.475 -216.405 32.805 -216.075 ;
        RECT 32.475 -217.765 32.805 -217.435 ;
        RECT 32.475 -219.125 32.805 -218.795 ;
        RECT 32.475 -220.485 32.805 -220.155 ;
        RECT 32.475 -221.845 32.805 -221.515 ;
        RECT 32.475 -223.205 32.805 -222.875 ;
        RECT 32.475 -224.565 32.805 -224.235 ;
        RECT 32.475 -225.925 32.805 -225.595 ;
        RECT 32.475 -227.285 32.805 -226.955 ;
        RECT 32.475 -228.645 32.805 -228.315 ;
        RECT 32.475 -230.005 32.805 -229.675 ;
        RECT 32.475 -231.365 32.805 -231.035 ;
        RECT 32.475 -232.725 32.805 -232.395 ;
        RECT 32.475 -234.085 32.805 -233.755 ;
        RECT 32.475 -235.445 32.805 -235.115 ;
        RECT 32.475 -236.805 32.805 -236.475 ;
        RECT 32.475 -238.165 32.805 -237.835 ;
        RECT 32.475 -243.81 32.805 -242.68 ;
        RECT 32.48 -243.925 32.8 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 246.76 34.165 247.89 ;
        RECT 33.835 241.915 34.165 242.245 ;
        RECT 33.835 240.555 34.165 240.885 ;
        RECT 33.835 239.195 34.165 239.525 ;
        RECT 33.835 237.835 34.165 238.165 ;
        RECT 33.84 237.16 34.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 -1.525 34.165 -1.195 ;
        RECT 33.835 -2.885 34.165 -2.555 ;
        RECT 33.84 -3.56 34.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 -122.565 34.165 -122.235 ;
        RECT 33.835 -123.925 34.165 -123.595 ;
        RECT 33.835 -125.285 34.165 -124.955 ;
        RECT 33.835 -126.645 34.165 -126.315 ;
        RECT 33.835 -128.005 34.165 -127.675 ;
        RECT 33.835 -129.365 34.165 -129.035 ;
        RECT 33.835 -130.725 34.165 -130.395 ;
        RECT 33.835 -132.085 34.165 -131.755 ;
        RECT 33.835 -133.445 34.165 -133.115 ;
        RECT 33.835 -134.805 34.165 -134.475 ;
        RECT 33.835 -136.165 34.165 -135.835 ;
        RECT 33.835 -137.525 34.165 -137.195 ;
        RECT 33.835 -138.885 34.165 -138.555 ;
        RECT 33.835 -140.245 34.165 -139.915 ;
        RECT 33.835 -141.605 34.165 -141.275 ;
        RECT 33.835 -142.965 34.165 -142.635 ;
        RECT 33.835 -144.325 34.165 -143.995 ;
        RECT 33.835 -145.685 34.165 -145.355 ;
        RECT 33.835 -147.045 34.165 -146.715 ;
        RECT 33.835 -148.405 34.165 -148.075 ;
        RECT 33.835 -149.765 34.165 -149.435 ;
        RECT 33.835 -151.125 34.165 -150.795 ;
        RECT 33.835 -152.485 34.165 -152.155 ;
        RECT 33.835 -153.845 34.165 -153.515 ;
        RECT 33.835 -155.205 34.165 -154.875 ;
        RECT 33.835 -156.565 34.165 -156.235 ;
        RECT 33.835 -157.925 34.165 -157.595 ;
        RECT 33.835 -159.285 34.165 -158.955 ;
        RECT 33.835 -160.645 34.165 -160.315 ;
        RECT 33.835 -162.005 34.165 -161.675 ;
        RECT 33.835 -163.365 34.165 -163.035 ;
        RECT 33.835 -164.725 34.165 -164.395 ;
        RECT 33.835 -166.085 34.165 -165.755 ;
        RECT 33.835 -167.445 34.165 -167.115 ;
        RECT 33.835 -168.805 34.165 -168.475 ;
        RECT 33.835 -170.165 34.165 -169.835 ;
        RECT 33.835 -171.525 34.165 -171.195 ;
        RECT 33.835 -172.885 34.165 -172.555 ;
        RECT 33.835 -174.245 34.165 -173.915 ;
        RECT 33.835 -175.605 34.165 -175.275 ;
        RECT 33.835 -176.965 34.165 -176.635 ;
        RECT 33.835 -178.325 34.165 -177.995 ;
        RECT 33.835 -179.685 34.165 -179.355 ;
        RECT 33.835 -181.045 34.165 -180.715 ;
        RECT 33.835 -182.405 34.165 -182.075 ;
        RECT 33.835 -183.765 34.165 -183.435 ;
        RECT 33.835 -185.125 34.165 -184.795 ;
        RECT 33.835 -186.485 34.165 -186.155 ;
        RECT 33.835 -187.845 34.165 -187.515 ;
        RECT 33.835 -189.205 34.165 -188.875 ;
        RECT 33.835 -190.565 34.165 -190.235 ;
        RECT 33.835 -191.925 34.165 -191.595 ;
        RECT 33.835 -193.285 34.165 -192.955 ;
        RECT 33.835 -194.645 34.165 -194.315 ;
        RECT 33.835 -196.005 34.165 -195.675 ;
        RECT 33.835 -197.365 34.165 -197.035 ;
        RECT 33.835 -198.725 34.165 -198.395 ;
        RECT 33.835 -200.085 34.165 -199.755 ;
        RECT 33.835 -201.445 34.165 -201.115 ;
        RECT 33.835 -202.805 34.165 -202.475 ;
        RECT 33.835 -204.165 34.165 -203.835 ;
        RECT 33.835 -205.525 34.165 -205.195 ;
        RECT 33.835 -206.885 34.165 -206.555 ;
        RECT 33.835 -208.245 34.165 -207.915 ;
        RECT 33.835 -209.605 34.165 -209.275 ;
        RECT 33.835 -210.965 34.165 -210.635 ;
        RECT 33.835 -212.325 34.165 -211.995 ;
        RECT 33.835 -213.685 34.165 -213.355 ;
        RECT 33.835 -215.045 34.165 -214.715 ;
        RECT 33.835 -216.405 34.165 -216.075 ;
        RECT 33.835 -217.765 34.165 -217.435 ;
        RECT 33.835 -219.125 34.165 -218.795 ;
        RECT 33.835 -220.485 34.165 -220.155 ;
        RECT 33.835 -221.845 34.165 -221.515 ;
        RECT 33.835 -223.205 34.165 -222.875 ;
        RECT 33.835 -224.565 34.165 -224.235 ;
        RECT 33.835 -225.925 34.165 -225.595 ;
        RECT 33.835 -227.285 34.165 -226.955 ;
        RECT 33.835 -228.645 34.165 -228.315 ;
        RECT 33.835 -230.005 34.165 -229.675 ;
        RECT 33.835 -231.365 34.165 -231.035 ;
        RECT 33.835 -232.725 34.165 -232.395 ;
        RECT 33.835 -234.085 34.165 -233.755 ;
        RECT 33.835 -235.445 34.165 -235.115 ;
        RECT 33.835 -236.805 34.165 -236.475 ;
        RECT 33.835 -238.165 34.165 -237.835 ;
        RECT 33.835 -243.81 34.165 -242.68 ;
        RECT 33.84 -243.925 34.16 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 246.76 35.525 247.89 ;
        RECT 35.195 241.915 35.525 242.245 ;
        RECT 35.195 240.555 35.525 240.885 ;
        RECT 35.195 239.195 35.525 239.525 ;
        RECT 35.195 237.835 35.525 238.165 ;
        RECT 35.2 237.16 35.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 -151.125 35.525 -150.795 ;
        RECT 35.195 -152.485 35.525 -152.155 ;
        RECT 35.195 -153.845 35.525 -153.515 ;
        RECT 35.195 -155.205 35.525 -154.875 ;
        RECT 35.195 -156.565 35.525 -156.235 ;
        RECT 35.195 -157.925 35.525 -157.595 ;
        RECT 35.195 -159.285 35.525 -158.955 ;
        RECT 35.195 -160.645 35.525 -160.315 ;
        RECT 35.195 -162.005 35.525 -161.675 ;
        RECT 35.195 -163.365 35.525 -163.035 ;
        RECT 35.195 -164.725 35.525 -164.395 ;
        RECT 35.195 -166.085 35.525 -165.755 ;
        RECT 35.195 -167.445 35.525 -167.115 ;
        RECT 35.195 -168.805 35.525 -168.475 ;
        RECT 35.195 -170.165 35.525 -169.835 ;
        RECT 35.195 -171.525 35.525 -171.195 ;
        RECT 35.195 -172.885 35.525 -172.555 ;
        RECT 35.195 -174.245 35.525 -173.915 ;
        RECT 35.195 -175.605 35.525 -175.275 ;
        RECT 35.195 -176.965 35.525 -176.635 ;
        RECT 35.195 -178.325 35.525 -177.995 ;
        RECT 35.195 -179.685 35.525 -179.355 ;
        RECT 35.195 -181.045 35.525 -180.715 ;
        RECT 35.195 -182.405 35.525 -182.075 ;
        RECT 35.195 -183.765 35.525 -183.435 ;
        RECT 35.195 -185.125 35.525 -184.795 ;
        RECT 35.195 -186.485 35.525 -186.155 ;
        RECT 35.195 -187.845 35.525 -187.515 ;
        RECT 35.195 -189.205 35.525 -188.875 ;
        RECT 35.195 -190.565 35.525 -190.235 ;
        RECT 35.195 -191.925 35.525 -191.595 ;
        RECT 35.195 -193.285 35.525 -192.955 ;
        RECT 35.195 -194.645 35.525 -194.315 ;
        RECT 35.195 -196.005 35.525 -195.675 ;
        RECT 35.195 -197.365 35.525 -197.035 ;
        RECT 35.195 -198.725 35.525 -198.395 ;
        RECT 35.195 -200.085 35.525 -199.755 ;
        RECT 35.195 -201.445 35.525 -201.115 ;
        RECT 35.195 -202.805 35.525 -202.475 ;
        RECT 35.195 -204.165 35.525 -203.835 ;
        RECT 35.195 -205.525 35.525 -205.195 ;
        RECT 35.195 -206.885 35.525 -206.555 ;
        RECT 35.195 -208.245 35.525 -207.915 ;
        RECT 35.195 -209.605 35.525 -209.275 ;
        RECT 35.195 -210.965 35.525 -210.635 ;
        RECT 35.195 -212.325 35.525 -211.995 ;
        RECT 35.195 -213.685 35.525 -213.355 ;
        RECT 35.195 -215.045 35.525 -214.715 ;
        RECT 35.195 -216.405 35.525 -216.075 ;
        RECT 35.195 -217.765 35.525 -217.435 ;
        RECT 35.195 -219.125 35.525 -218.795 ;
        RECT 35.195 -220.485 35.525 -220.155 ;
        RECT 35.195 -221.845 35.525 -221.515 ;
        RECT 35.195 -223.205 35.525 -222.875 ;
        RECT 35.195 -224.565 35.525 -224.235 ;
        RECT 35.195 -225.925 35.525 -225.595 ;
        RECT 35.195 -227.285 35.525 -226.955 ;
        RECT 35.195 -228.645 35.525 -228.315 ;
        RECT 35.195 -230.005 35.525 -229.675 ;
        RECT 35.195 -231.365 35.525 -231.035 ;
        RECT 35.195 -232.725 35.525 -232.395 ;
        RECT 35.195 -234.085 35.525 -233.755 ;
        RECT 35.195 -235.445 35.525 -235.115 ;
        RECT 35.195 -236.805 35.525 -236.475 ;
        RECT 35.195 -238.165 35.525 -237.835 ;
        RECT 35.195 -243.81 35.525 -242.68 ;
        RECT 35.2 -243.925 35.52 -126.315 ;
        RECT 35.195 -126.645 35.525 -126.315 ;
        RECT 35.195 -128.005 35.525 -127.675 ;
        RECT 35.195 -129.365 35.525 -129.035 ;
        RECT 35.195 -130.725 35.525 -130.395 ;
        RECT 35.195 -132.085 35.525 -131.755 ;
        RECT 35.195 -133.445 35.525 -133.115 ;
        RECT 35.195 -134.805 35.525 -134.475 ;
        RECT 35.195 -136.165 35.525 -135.835 ;
        RECT 35.195 -137.525 35.525 -137.195 ;
        RECT 35.195 -138.885 35.525 -138.555 ;
        RECT 35.195 -140.245 35.525 -139.915 ;
        RECT 35.195 -141.605 35.525 -141.275 ;
        RECT 35.195 -142.965 35.525 -142.635 ;
        RECT 35.195 -144.325 35.525 -143.995 ;
        RECT 35.195 -145.685 35.525 -145.355 ;
        RECT 35.195 -147.045 35.525 -146.715 ;
        RECT 35.195 -148.405 35.525 -148.075 ;
        RECT 35.195 -149.765 35.525 -149.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 246.76 0.165 247.89 ;
        RECT -0.165 241.915 0.165 242.245 ;
        RECT -0.165 240.555 0.165 240.885 ;
        RECT -0.165 239.195 0.165 239.525 ;
        RECT -0.165 237.835 0.165 238.165 ;
        RECT -0.16 237.16 0.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -1.525 0.165 -1.195 ;
        RECT -0.165 -2.885 0.165 -2.555 ;
        RECT -0.16 -3.56 0.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -122.565 0.165 -122.235 ;
        RECT -0.165 -123.925 0.165 -123.595 ;
        RECT -0.165 -125.285 0.165 -124.955 ;
        RECT -0.165 -126.645 0.165 -126.315 ;
        RECT -0.165 -128.005 0.165 -127.675 ;
        RECT -0.165 -129.365 0.165 -129.035 ;
        RECT -0.165 -130.725 0.165 -130.395 ;
        RECT -0.165 -132.085 0.165 -131.755 ;
        RECT -0.165 -133.445 0.165 -133.115 ;
        RECT -0.165 -134.805 0.165 -134.475 ;
        RECT -0.165 -136.165 0.165 -135.835 ;
        RECT -0.165 -137.525 0.165 -137.195 ;
        RECT -0.165 -138.885 0.165 -138.555 ;
        RECT -0.165 -140.245 0.165 -139.915 ;
        RECT -0.165 -141.605 0.165 -141.275 ;
        RECT -0.165 -142.965 0.165 -142.635 ;
        RECT -0.165 -144.325 0.165 -143.995 ;
        RECT -0.165 -145.685 0.165 -145.355 ;
        RECT -0.165 -147.045 0.165 -146.715 ;
        RECT -0.165 -148.405 0.165 -148.075 ;
        RECT -0.165 -149.765 0.165 -149.435 ;
        RECT -0.165 -151.125 0.165 -150.795 ;
        RECT -0.165 -152.485 0.165 -152.155 ;
        RECT -0.165 -153.845 0.165 -153.515 ;
        RECT -0.165 -155.205 0.165 -154.875 ;
        RECT -0.165 -156.565 0.165 -156.235 ;
        RECT -0.165 -157.925 0.165 -157.595 ;
        RECT -0.165 -160.645 0.165 -160.315 ;
        RECT -0.165 -162.005 0.165 -161.675 ;
        RECT -0.165 -163.365 0.165 -163.035 ;
        RECT -0.165 -164.725 0.165 -164.395 ;
        RECT -0.165 -166.085 0.165 -165.755 ;
        RECT -0.165 -167.445 0.165 -167.115 ;
        RECT -0.165 -168.805 0.165 -168.475 ;
        RECT -0.165 -170.165 0.165 -169.835 ;
        RECT -0.165 -171.525 0.165 -171.195 ;
        RECT -0.165 -172.885 0.165 -172.555 ;
        RECT -0.165 -174.245 0.165 -173.915 ;
        RECT -0.165 -175.605 0.165 -175.275 ;
        RECT -0.165 -176.965 0.165 -176.635 ;
        RECT -0.165 -178.325 0.165 -177.995 ;
        RECT -0.165 -179.685 0.165 -179.355 ;
        RECT -0.165 -181.045 0.165 -180.715 ;
        RECT -0.165 -182.405 0.165 -182.075 ;
        RECT -0.165 -183.765 0.165 -183.435 ;
        RECT -0.165 -185.125 0.165 -184.795 ;
        RECT -0.165 -186.485 0.165 -186.155 ;
        RECT -0.165 -187.845 0.165 -187.515 ;
        RECT -0.165 -189.205 0.165 -188.875 ;
        RECT -0.165 -190.565 0.165 -190.235 ;
        RECT -0.165 -191.925 0.165 -191.595 ;
        RECT -0.165 -193.285 0.165 -192.955 ;
        RECT -0.165 -194.645 0.165 -194.315 ;
        RECT -0.165 -196.005 0.165 -195.675 ;
        RECT -0.165 -197.365 0.165 -197.035 ;
        RECT -0.165 -198.725 0.165 -198.395 ;
        RECT -0.165 -200.085 0.165 -199.755 ;
        RECT -0.165 -201.445 0.165 -201.115 ;
        RECT -0.165 -202.805 0.165 -202.475 ;
        RECT -0.165 -204.165 0.165 -203.835 ;
        RECT -0.165 -205.525 0.165 -205.195 ;
        RECT -0.165 -206.885 0.165 -206.555 ;
        RECT -0.165 -208.245 0.165 -207.915 ;
        RECT -0.165 -209.605 0.165 -209.275 ;
        RECT -0.165 -210.965 0.165 -210.635 ;
        RECT -0.165 -212.325 0.165 -211.995 ;
        RECT -0.165 -213.685 0.165 -213.355 ;
        RECT -0.165 -215.045 0.165 -214.715 ;
        RECT -0.165 -216.405 0.165 -216.075 ;
        RECT -0.165 -217.765 0.165 -217.435 ;
        RECT -0.165 -219.125 0.165 -218.795 ;
        RECT -0.165 -220.485 0.165 -220.155 ;
        RECT -0.165 -221.845 0.165 -221.515 ;
        RECT -0.165 -223.205 0.165 -222.875 ;
        RECT -0.165 -224.565 0.165 -224.235 ;
        RECT -0.165 -225.925 0.165 -225.595 ;
        RECT -0.165 -227.285 0.165 -226.955 ;
        RECT -0.165 -228.645 0.165 -228.315 ;
        RECT -0.165 -230.005 0.165 -229.675 ;
        RECT -0.165 -231.365 0.165 -231.035 ;
        RECT -0.165 -232.725 0.165 -232.395 ;
        RECT -0.165 -234.085 0.165 -233.755 ;
        RECT -0.165 -235.445 0.165 -235.115 ;
        RECT -0.165 -236.805 0.165 -236.475 ;
        RECT -0.165 -238.165 0.165 -237.835 ;
        RECT -0.165 -243.81 0.165 -242.68 ;
        RECT -0.16 -243.925 0.16 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 246.76 1.525 247.89 ;
        RECT 1.195 241.915 1.525 242.245 ;
        RECT 1.195 240.555 1.525 240.885 ;
        RECT 1.195 239.195 1.525 239.525 ;
        RECT 1.195 237.835 1.525 238.165 ;
        RECT 1.2 237.16 1.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -1.525 1.525 -1.195 ;
        RECT 1.195 -2.885 1.525 -2.555 ;
        RECT 1.2 -3.56 1.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -122.565 1.525 -122.235 ;
        RECT 1.195 -123.925 1.525 -123.595 ;
        RECT 1.195 -125.285 1.525 -124.955 ;
        RECT 1.195 -126.645 1.525 -126.315 ;
        RECT 1.195 -128.005 1.525 -127.675 ;
        RECT 1.195 -129.365 1.525 -129.035 ;
        RECT 1.195 -130.725 1.525 -130.395 ;
        RECT 1.195 -132.085 1.525 -131.755 ;
        RECT 1.195 -133.445 1.525 -133.115 ;
        RECT 1.195 -134.805 1.525 -134.475 ;
        RECT 1.195 -136.165 1.525 -135.835 ;
        RECT 1.195 -137.525 1.525 -137.195 ;
        RECT 1.195 -138.885 1.525 -138.555 ;
        RECT 1.195 -140.245 1.525 -139.915 ;
        RECT 1.195 -141.605 1.525 -141.275 ;
        RECT 1.195 -142.965 1.525 -142.635 ;
        RECT 1.195 -144.325 1.525 -143.995 ;
        RECT 1.195 -145.685 1.525 -145.355 ;
        RECT 1.195 -147.045 1.525 -146.715 ;
        RECT 1.195 -148.405 1.525 -148.075 ;
        RECT 1.195 -149.765 1.525 -149.435 ;
        RECT 1.195 -151.125 1.525 -150.795 ;
        RECT 1.195 -152.485 1.525 -152.155 ;
        RECT 1.195 -153.845 1.525 -153.515 ;
        RECT 1.195 -155.205 1.525 -154.875 ;
        RECT 1.195 -156.565 1.525 -156.235 ;
        RECT 1.195 -157.925 1.525 -157.595 ;
        RECT 1.195 -159.285 1.525 -158.955 ;
        RECT 1.195 -160.645 1.525 -160.315 ;
        RECT 1.195 -162.005 1.525 -161.675 ;
        RECT 1.195 -163.365 1.525 -163.035 ;
        RECT 1.195 -164.725 1.525 -164.395 ;
        RECT 1.195 -166.085 1.525 -165.755 ;
        RECT 1.195 -167.445 1.525 -167.115 ;
        RECT 1.195 -168.805 1.525 -168.475 ;
        RECT 1.195 -170.165 1.525 -169.835 ;
        RECT 1.195 -171.525 1.525 -171.195 ;
        RECT 1.195 -172.885 1.525 -172.555 ;
        RECT 1.195 -174.245 1.525 -173.915 ;
        RECT 1.195 -175.605 1.525 -175.275 ;
        RECT 1.195 -176.965 1.525 -176.635 ;
        RECT 1.195 -178.325 1.525 -177.995 ;
        RECT 1.195 -179.685 1.525 -179.355 ;
        RECT 1.195 -181.045 1.525 -180.715 ;
        RECT 1.195 -182.405 1.525 -182.075 ;
        RECT 1.195 -183.765 1.525 -183.435 ;
        RECT 1.195 -185.125 1.525 -184.795 ;
        RECT 1.195 -186.485 1.525 -186.155 ;
        RECT 1.195 -187.845 1.525 -187.515 ;
        RECT 1.195 -189.205 1.525 -188.875 ;
        RECT 1.195 -190.565 1.525 -190.235 ;
        RECT 1.195 -191.925 1.525 -191.595 ;
        RECT 1.195 -193.285 1.525 -192.955 ;
        RECT 1.195 -194.645 1.525 -194.315 ;
        RECT 1.195 -196.005 1.525 -195.675 ;
        RECT 1.195 -197.365 1.525 -197.035 ;
        RECT 1.195 -198.725 1.525 -198.395 ;
        RECT 1.195 -200.085 1.525 -199.755 ;
        RECT 1.195 -201.445 1.525 -201.115 ;
        RECT 1.195 -202.805 1.525 -202.475 ;
        RECT 1.195 -204.165 1.525 -203.835 ;
        RECT 1.195 -205.525 1.525 -205.195 ;
        RECT 1.195 -206.885 1.525 -206.555 ;
        RECT 1.195 -208.245 1.525 -207.915 ;
        RECT 1.195 -209.605 1.525 -209.275 ;
        RECT 1.195 -210.965 1.525 -210.635 ;
        RECT 1.195 -212.325 1.525 -211.995 ;
        RECT 1.195 -213.685 1.525 -213.355 ;
        RECT 1.195 -215.045 1.525 -214.715 ;
        RECT 1.195 -216.405 1.525 -216.075 ;
        RECT 1.195 -217.765 1.525 -217.435 ;
        RECT 1.195 -219.125 1.525 -218.795 ;
        RECT 1.195 -220.485 1.525 -220.155 ;
        RECT 1.195 -221.845 1.525 -221.515 ;
        RECT 1.195 -223.205 1.525 -222.875 ;
        RECT 1.195 -224.565 1.525 -224.235 ;
        RECT 1.195 -225.925 1.525 -225.595 ;
        RECT 1.195 -227.285 1.525 -226.955 ;
        RECT 1.195 -228.645 1.525 -228.315 ;
        RECT 1.195 -230.005 1.525 -229.675 ;
        RECT 1.195 -231.365 1.525 -231.035 ;
        RECT 1.195 -232.725 1.525 -232.395 ;
        RECT 1.195 -234.085 1.525 -233.755 ;
        RECT 1.195 -235.445 1.525 -235.115 ;
        RECT 1.195 -236.805 1.525 -236.475 ;
        RECT 1.195 -238.165 1.525 -237.835 ;
        RECT 1.195 -243.81 1.525 -242.68 ;
        RECT 1.2 -243.925 1.52 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 246.76 2.885 247.89 ;
        RECT 2.555 241.915 2.885 242.245 ;
        RECT 2.555 240.555 2.885 240.885 ;
        RECT 2.555 239.195 2.885 239.525 ;
        RECT 2.555 237.835 2.885 238.165 ;
        RECT 2.56 237.16 2.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 -126.645 2.885 -126.315 ;
        RECT 2.555 -128.005 2.885 -127.675 ;
        RECT 2.555 -129.365 2.885 -129.035 ;
        RECT 2.555 -130.725 2.885 -130.395 ;
        RECT 2.555 -132.085 2.885 -131.755 ;
        RECT 2.555 -133.445 2.885 -133.115 ;
        RECT 2.555 -134.805 2.885 -134.475 ;
        RECT 2.555 -136.165 2.885 -135.835 ;
        RECT 2.555 -137.525 2.885 -137.195 ;
        RECT 2.555 -138.885 2.885 -138.555 ;
        RECT 2.555 -140.245 2.885 -139.915 ;
        RECT 2.555 -141.605 2.885 -141.275 ;
        RECT 2.555 -142.965 2.885 -142.635 ;
        RECT 2.555 -144.325 2.885 -143.995 ;
        RECT 2.555 -145.685 2.885 -145.355 ;
        RECT 2.555 -147.045 2.885 -146.715 ;
        RECT 2.555 -148.405 2.885 -148.075 ;
        RECT 2.555 -149.765 2.885 -149.435 ;
        RECT 2.555 -151.125 2.885 -150.795 ;
        RECT 2.555 -152.485 2.885 -152.155 ;
        RECT 2.555 -153.845 2.885 -153.515 ;
        RECT 2.555 -155.205 2.885 -154.875 ;
        RECT 2.555 -156.565 2.885 -156.235 ;
        RECT 2.555 -157.925 2.885 -157.595 ;
        RECT 2.555 -159.285 2.885 -158.955 ;
        RECT 2.555 -160.645 2.885 -160.315 ;
        RECT 2.555 -162.005 2.885 -161.675 ;
        RECT 2.555 -163.365 2.885 -163.035 ;
        RECT 2.555 -164.725 2.885 -164.395 ;
        RECT 2.555 -166.085 2.885 -165.755 ;
        RECT 2.555 -167.445 2.885 -167.115 ;
        RECT 2.555 -168.805 2.885 -168.475 ;
        RECT 2.555 -170.165 2.885 -169.835 ;
        RECT 2.555 -171.525 2.885 -171.195 ;
        RECT 2.555 -172.885 2.885 -172.555 ;
        RECT 2.555 -174.245 2.885 -173.915 ;
        RECT 2.555 -175.605 2.885 -175.275 ;
        RECT 2.555 -176.965 2.885 -176.635 ;
        RECT 2.555 -178.325 2.885 -177.995 ;
        RECT 2.555 -179.685 2.885 -179.355 ;
        RECT 2.555 -181.045 2.885 -180.715 ;
        RECT 2.555 -182.405 2.885 -182.075 ;
        RECT 2.555 -183.765 2.885 -183.435 ;
        RECT 2.555 -185.125 2.885 -184.795 ;
        RECT 2.555 -186.485 2.885 -186.155 ;
        RECT 2.555 -187.845 2.885 -187.515 ;
        RECT 2.555 -189.205 2.885 -188.875 ;
        RECT 2.555 -190.565 2.885 -190.235 ;
        RECT 2.555 -191.925 2.885 -191.595 ;
        RECT 2.555 -193.285 2.885 -192.955 ;
        RECT 2.555 -194.645 2.885 -194.315 ;
        RECT 2.555 -196.005 2.885 -195.675 ;
        RECT 2.555 -197.365 2.885 -197.035 ;
        RECT 2.555 -198.725 2.885 -198.395 ;
        RECT 2.555 -200.085 2.885 -199.755 ;
        RECT 2.555 -201.445 2.885 -201.115 ;
        RECT 2.555 -202.805 2.885 -202.475 ;
        RECT 2.555 -204.165 2.885 -203.835 ;
        RECT 2.555 -205.525 2.885 -205.195 ;
        RECT 2.555 -206.885 2.885 -206.555 ;
        RECT 2.555 -208.245 2.885 -207.915 ;
        RECT 2.555 -209.605 2.885 -209.275 ;
        RECT 2.555 -210.965 2.885 -210.635 ;
        RECT 2.555 -212.325 2.885 -211.995 ;
        RECT 2.555 -213.685 2.885 -213.355 ;
        RECT 2.555 -215.045 2.885 -214.715 ;
        RECT 2.555 -216.405 2.885 -216.075 ;
        RECT 2.555 -217.765 2.885 -217.435 ;
        RECT 2.555 -219.125 2.885 -218.795 ;
        RECT 2.555 -220.485 2.885 -220.155 ;
        RECT 2.555 -221.845 2.885 -221.515 ;
        RECT 2.555 -223.205 2.885 -222.875 ;
        RECT 2.555 -224.565 2.885 -224.235 ;
        RECT 2.555 -225.925 2.885 -225.595 ;
        RECT 2.555 -227.285 2.885 -226.955 ;
        RECT 2.555 -228.645 2.885 -228.315 ;
        RECT 2.555 -230.005 2.885 -229.675 ;
        RECT 2.555 -231.365 2.885 -231.035 ;
        RECT 2.555 -232.725 2.885 -232.395 ;
        RECT 2.555 -234.085 2.885 -233.755 ;
        RECT 2.555 -235.445 2.885 -235.115 ;
        RECT 2.555 -236.805 2.885 -236.475 ;
        RECT 2.555 -238.165 2.885 -237.835 ;
        RECT 2.555 -243.81 2.885 -242.68 ;
        RECT 2.56 -243.925 2.88 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.66 -125.535 2.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 246.76 4.245 247.89 ;
        RECT 3.915 241.915 4.245 242.245 ;
        RECT 3.915 240.555 4.245 240.885 ;
        RECT 3.915 239.195 4.245 239.525 ;
        RECT 3.915 237.835 4.245 238.165 ;
        RECT 3.92 237.16 4.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 246.76 5.605 247.89 ;
        RECT 5.275 241.915 5.605 242.245 ;
        RECT 5.275 240.555 5.605 240.885 ;
        RECT 5.275 239.195 5.605 239.525 ;
        RECT 5.275 237.835 5.605 238.165 ;
        RECT 5.28 237.16 5.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 -1.525 5.605 -1.195 ;
        RECT 5.275 -2.885 5.605 -2.555 ;
        RECT 5.28 -3.56 5.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 246.76 6.965 247.89 ;
        RECT 6.635 241.915 6.965 242.245 ;
        RECT 6.635 240.555 6.965 240.885 ;
        RECT 6.635 239.195 6.965 239.525 ;
        RECT 6.635 237.835 6.965 238.165 ;
        RECT 6.64 237.16 6.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 -1.525 6.965 -1.195 ;
        RECT 6.635 -2.885 6.965 -2.555 ;
        RECT 6.64 -3.56 6.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 246.76 8.325 247.89 ;
        RECT 7.995 241.915 8.325 242.245 ;
        RECT 7.995 240.555 8.325 240.885 ;
        RECT 7.995 239.195 8.325 239.525 ;
        RECT 7.995 237.835 8.325 238.165 ;
        RECT 8 237.16 8.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -1.525 8.325 -1.195 ;
        RECT 7.995 -2.885 8.325 -2.555 ;
        RECT 8 -3.56 8.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -122.565 8.325 -122.235 ;
        RECT 7.995 -123.925 8.325 -123.595 ;
        RECT 7.995 -125.285 8.325 -124.955 ;
        RECT 7.995 -126.645 8.325 -126.315 ;
        RECT 7.995 -128.005 8.325 -127.675 ;
        RECT 7.995 -129.365 8.325 -129.035 ;
        RECT 7.995 -130.725 8.325 -130.395 ;
        RECT 7.995 -132.085 8.325 -131.755 ;
        RECT 7.995 -133.445 8.325 -133.115 ;
        RECT 7.995 -134.805 8.325 -134.475 ;
        RECT 7.995 -136.165 8.325 -135.835 ;
        RECT 7.995 -137.525 8.325 -137.195 ;
        RECT 7.995 -138.885 8.325 -138.555 ;
        RECT 7.995 -140.245 8.325 -139.915 ;
        RECT 7.995 -141.605 8.325 -141.275 ;
        RECT 7.995 -142.965 8.325 -142.635 ;
        RECT 7.995 -144.325 8.325 -143.995 ;
        RECT 7.995 -145.685 8.325 -145.355 ;
        RECT 7.995 -147.045 8.325 -146.715 ;
        RECT 7.995 -148.405 8.325 -148.075 ;
        RECT 7.995 -149.765 8.325 -149.435 ;
        RECT 7.995 -151.125 8.325 -150.795 ;
        RECT 7.995 -152.485 8.325 -152.155 ;
        RECT 7.995 -153.845 8.325 -153.515 ;
        RECT 7.995 -155.205 8.325 -154.875 ;
        RECT 7.995 -156.565 8.325 -156.235 ;
        RECT 7.995 -157.925 8.325 -157.595 ;
        RECT 7.995 -159.285 8.325 -158.955 ;
        RECT 7.995 -160.645 8.325 -160.315 ;
        RECT 7.995 -162.005 8.325 -161.675 ;
        RECT 7.995 -163.365 8.325 -163.035 ;
        RECT 7.995 -164.725 8.325 -164.395 ;
        RECT 7.995 -166.085 8.325 -165.755 ;
        RECT 7.995 -167.445 8.325 -167.115 ;
        RECT 7.995 -168.805 8.325 -168.475 ;
        RECT 7.995 -170.165 8.325 -169.835 ;
        RECT 7.995 -171.525 8.325 -171.195 ;
        RECT 7.995 -172.885 8.325 -172.555 ;
        RECT 7.995 -174.245 8.325 -173.915 ;
        RECT 7.995 -175.605 8.325 -175.275 ;
        RECT 7.995 -176.965 8.325 -176.635 ;
        RECT 7.995 -178.325 8.325 -177.995 ;
        RECT 7.995 -179.685 8.325 -179.355 ;
        RECT 7.995 -181.045 8.325 -180.715 ;
        RECT 7.995 -182.405 8.325 -182.075 ;
        RECT 7.995 -183.765 8.325 -183.435 ;
        RECT 7.995 -185.125 8.325 -184.795 ;
        RECT 7.995 -186.485 8.325 -186.155 ;
        RECT 7.995 -187.845 8.325 -187.515 ;
        RECT 7.995 -189.205 8.325 -188.875 ;
        RECT 7.995 -190.565 8.325 -190.235 ;
        RECT 7.995 -191.925 8.325 -191.595 ;
        RECT 7.995 -193.285 8.325 -192.955 ;
        RECT 7.995 -194.645 8.325 -194.315 ;
        RECT 7.995 -196.005 8.325 -195.675 ;
        RECT 7.995 -197.365 8.325 -197.035 ;
        RECT 7.995 -198.725 8.325 -198.395 ;
        RECT 7.995 -200.085 8.325 -199.755 ;
        RECT 7.995 -201.445 8.325 -201.115 ;
        RECT 7.995 -202.805 8.325 -202.475 ;
        RECT 7.995 -204.165 8.325 -203.835 ;
        RECT 7.995 -205.525 8.325 -205.195 ;
        RECT 7.995 -206.885 8.325 -206.555 ;
        RECT 7.995 -208.245 8.325 -207.915 ;
        RECT 7.995 -209.605 8.325 -209.275 ;
        RECT 7.995 -210.965 8.325 -210.635 ;
        RECT 7.995 -212.325 8.325 -211.995 ;
        RECT 7.995 -213.685 8.325 -213.355 ;
        RECT 7.995 -215.045 8.325 -214.715 ;
        RECT 7.995 -216.405 8.325 -216.075 ;
        RECT 7.995 -217.765 8.325 -217.435 ;
        RECT 7.995 -219.125 8.325 -218.795 ;
        RECT 7.995 -220.485 8.325 -220.155 ;
        RECT 7.995 -221.845 8.325 -221.515 ;
        RECT 7.995 -223.205 8.325 -222.875 ;
        RECT 7.995 -224.565 8.325 -224.235 ;
        RECT 7.995 -225.925 8.325 -225.595 ;
        RECT 7.995 -227.285 8.325 -226.955 ;
        RECT 7.995 -228.645 8.325 -228.315 ;
        RECT 7.995 -230.005 8.325 -229.675 ;
        RECT 7.995 -231.365 8.325 -231.035 ;
        RECT 7.995 -232.725 8.325 -232.395 ;
        RECT 7.995 -234.085 8.325 -233.755 ;
        RECT 7.995 -235.445 8.325 -235.115 ;
        RECT 7.995 -236.805 8.325 -236.475 ;
        RECT 7.995 -238.165 8.325 -237.835 ;
        RECT 7.995 -243.81 8.325 -242.68 ;
        RECT 8 -243.925 8.32 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 246.76 9.685 247.89 ;
        RECT 9.355 241.915 9.685 242.245 ;
        RECT 9.355 240.555 9.685 240.885 ;
        RECT 9.355 239.195 9.685 239.525 ;
        RECT 9.355 237.835 9.685 238.165 ;
        RECT 9.36 237.16 9.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 -1.525 9.685 -1.195 ;
        RECT 9.355 -2.885 9.685 -2.555 ;
        RECT 9.36 -3.56 9.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 -122.565 9.685 -122.235 ;
        RECT 9.355 -123.925 9.685 -123.595 ;
        RECT 9.355 -125.285 9.685 -124.955 ;
        RECT 9.355 -126.645 9.685 -126.315 ;
        RECT 9.355 -128.005 9.685 -127.675 ;
        RECT 9.355 -129.365 9.685 -129.035 ;
        RECT 9.355 -130.725 9.685 -130.395 ;
        RECT 9.355 -132.085 9.685 -131.755 ;
        RECT 9.355 -133.445 9.685 -133.115 ;
        RECT 9.355 -134.805 9.685 -134.475 ;
        RECT 9.355 -136.165 9.685 -135.835 ;
        RECT 9.355 -137.525 9.685 -137.195 ;
        RECT 9.355 -138.885 9.685 -138.555 ;
        RECT 9.355 -140.245 9.685 -139.915 ;
        RECT 9.355 -141.605 9.685 -141.275 ;
        RECT 9.355 -142.965 9.685 -142.635 ;
        RECT 9.355 -144.325 9.685 -143.995 ;
        RECT 9.355 -145.685 9.685 -145.355 ;
        RECT 9.355 -147.045 9.685 -146.715 ;
        RECT 9.355 -148.405 9.685 -148.075 ;
        RECT 9.355 -149.765 9.685 -149.435 ;
        RECT 9.355 -151.125 9.685 -150.795 ;
        RECT 9.355 -152.485 9.685 -152.155 ;
        RECT 9.355 -153.845 9.685 -153.515 ;
        RECT 9.355 -155.205 9.685 -154.875 ;
        RECT 9.355 -156.565 9.685 -156.235 ;
        RECT 9.355 -157.925 9.685 -157.595 ;
        RECT 9.355 -159.285 9.685 -158.955 ;
        RECT 9.355 -160.645 9.685 -160.315 ;
        RECT 9.355 -162.005 9.685 -161.675 ;
        RECT 9.355 -163.365 9.685 -163.035 ;
        RECT 9.355 -164.725 9.685 -164.395 ;
        RECT 9.355 -166.085 9.685 -165.755 ;
        RECT 9.355 -167.445 9.685 -167.115 ;
        RECT 9.355 -168.805 9.685 -168.475 ;
        RECT 9.355 -170.165 9.685 -169.835 ;
        RECT 9.355 -171.525 9.685 -171.195 ;
        RECT 9.355 -172.885 9.685 -172.555 ;
        RECT 9.355 -174.245 9.685 -173.915 ;
        RECT 9.355 -175.605 9.685 -175.275 ;
        RECT 9.355 -176.965 9.685 -176.635 ;
        RECT 9.355 -178.325 9.685 -177.995 ;
        RECT 9.355 -179.685 9.685 -179.355 ;
        RECT 9.355 -181.045 9.685 -180.715 ;
        RECT 9.355 -182.405 9.685 -182.075 ;
        RECT 9.355 -183.765 9.685 -183.435 ;
        RECT 9.355 -185.125 9.685 -184.795 ;
        RECT 9.355 -186.485 9.685 -186.155 ;
        RECT 9.355 -187.845 9.685 -187.515 ;
        RECT 9.355 -189.205 9.685 -188.875 ;
        RECT 9.355 -190.565 9.685 -190.235 ;
        RECT 9.355 -191.925 9.685 -191.595 ;
        RECT 9.355 -193.285 9.685 -192.955 ;
        RECT 9.355 -194.645 9.685 -194.315 ;
        RECT 9.355 -196.005 9.685 -195.675 ;
        RECT 9.355 -197.365 9.685 -197.035 ;
        RECT 9.355 -198.725 9.685 -198.395 ;
        RECT 9.355 -200.085 9.685 -199.755 ;
        RECT 9.355 -201.445 9.685 -201.115 ;
        RECT 9.355 -202.805 9.685 -202.475 ;
        RECT 9.355 -204.165 9.685 -203.835 ;
        RECT 9.355 -205.525 9.685 -205.195 ;
        RECT 9.355 -206.885 9.685 -206.555 ;
        RECT 9.355 -208.245 9.685 -207.915 ;
        RECT 9.355 -209.605 9.685 -209.275 ;
        RECT 9.355 -210.965 9.685 -210.635 ;
        RECT 9.355 -212.325 9.685 -211.995 ;
        RECT 9.355 -213.685 9.685 -213.355 ;
        RECT 9.355 -215.045 9.685 -214.715 ;
        RECT 9.355 -216.405 9.685 -216.075 ;
        RECT 9.355 -217.765 9.685 -217.435 ;
        RECT 9.355 -219.125 9.685 -218.795 ;
        RECT 9.355 -220.485 9.685 -220.155 ;
        RECT 9.355 -221.845 9.685 -221.515 ;
        RECT 9.355 -223.205 9.685 -222.875 ;
        RECT 9.355 -224.565 9.685 -224.235 ;
        RECT 9.355 -225.925 9.685 -225.595 ;
        RECT 9.355 -227.285 9.685 -226.955 ;
        RECT 9.355 -228.645 9.685 -228.315 ;
        RECT 9.355 -230.005 9.685 -229.675 ;
        RECT 9.355 -231.365 9.685 -231.035 ;
        RECT 9.355 -232.725 9.685 -232.395 ;
        RECT 9.355 -234.085 9.685 -233.755 ;
        RECT 9.355 -235.445 9.685 -235.115 ;
        RECT 9.355 -236.805 9.685 -236.475 ;
        RECT 9.355 -238.165 9.685 -237.835 ;
        RECT 9.355 -243.81 9.685 -242.68 ;
        RECT 9.36 -243.925 9.68 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 246.76 11.045 247.89 ;
        RECT 10.715 241.915 11.045 242.245 ;
        RECT 10.715 240.555 11.045 240.885 ;
        RECT 10.715 239.195 11.045 239.525 ;
        RECT 10.715 237.835 11.045 238.165 ;
        RECT 10.72 237.16 11.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -1.525 11.045 -1.195 ;
        RECT 10.715 -2.885 11.045 -2.555 ;
        RECT 10.72 -3.56 11.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -122.565 11.045 -122.235 ;
        RECT 10.715 -123.925 11.045 -123.595 ;
        RECT 10.715 -125.285 11.045 -124.955 ;
        RECT 10.715 -126.645 11.045 -126.315 ;
        RECT 10.715 -128.005 11.045 -127.675 ;
        RECT 10.715 -129.365 11.045 -129.035 ;
        RECT 10.715 -130.725 11.045 -130.395 ;
        RECT 10.715 -132.085 11.045 -131.755 ;
        RECT 10.715 -133.445 11.045 -133.115 ;
        RECT 10.715 -134.805 11.045 -134.475 ;
        RECT 10.715 -136.165 11.045 -135.835 ;
        RECT 10.715 -137.525 11.045 -137.195 ;
        RECT 10.715 -138.885 11.045 -138.555 ;
        RECT 10.715 -140.245 11.045 -139.915 ;
        RECT 10.715 -141.605 11.045 -141.275 ;
        RECT 10.715 -142.965 11.045 -142.635 ;
        RECT 10.715 -144.325 11.045 -143.995 ;
        RECT 10.715 -145.685 11.045 -145.355 ;
        RECT 10.715 -147.045 11.045 -146.715 ;
        RECT 10.715 -148.405 11.045 -148.075 ;
        RECT 10.715 -149.765 11.045 -149.435 ;
        RECT 10.715 -151.125 11.045 -150.795 ;
        RECT 10.715 -152.485 11.045 -152.155 ;
        RECT 10.715 -153.845 11.045 -153.515 ;
        RECT 10.715 -155.205 11.045 -154.875 ;
        RECT 10.715 -156.565 11.045 -156.235 ;
        RECT 10.715 -157.925 11.045 -157.595 ;
        RECT 10.715 -159.285 11.045 -158.955 ;
        RECT 10.715 -160.645 11.045 -160.315 ;
        RECT 10.715 -162.005 11.045 -161.675 ;
        RECT 10.715 -163.365 11.045 -163.035 ;
        RECT 10.715 -164.725 11.045 -164.395 ;
        RECT 10.715 -166.085 11.045 -165.755 ;
        RECT 10.715 -167.445 11.045 -167.115 ;
        RECT 10.715 -168.805 11.045 -168.475 ;
        RECT 10.715 -170.165 11.045 -169.835 ;
        RECT 10.715 -171.525 11.045 -171.195 ;
        RECT 10.715 -172.885 11.045 -172.555 ;
        RECT 10.715 -174.245 11.045 -173.915 ;
        RECT 10.715 -175.605 11.045 -175.275 ;
        RECT 10.715 -176.965 11.045 -176.635 ;
        RECT 10.715 -178.325 11.045 -177.995 ;
        RECT 10.715 -179.685 11.045 -179.355 ;
        RECT 10.715 -181.045 11.045 -180.715 ;
        RECT 10.715 -182.405 11.045 -182.075 ;
        RECT 10.715 -183.765 11.045 -183.435 ;
        RECT 10.715 -185.125 11.045 -184.795 ;
        RECT 10.715 -186.485 11.045 -186.155 ;
        RECT 10.715 -187.845 11.045 -187.515 ;
        RECT 10.715 -189.205 11.045 -188.875 ;
        RECT 10.715 -190.565 11.045 -190.235 ;
        RECT 10.715 -191.925 11.045 -191.595 ;
        RECT 10.715 -193.285 11.045 -192.955 ;
        RECT 10.715 -194.645 11.045 -194.315 ;
        RECT 10.715 -196.005 11.045 -195.675 ;
        RECT 10.715 -197.365 11.045 -197.035 ;
        RECT 10.715 -198.725 11.045 -198.395 ;
        RECT 10.715 -200.085 11.045 -199.755 ;
        RECT 10.715 -201.445 11.045 -201.115 ;
        RECT 10.715 -202.805 11.045 -202.475 ;
        RECT 10.715 -204.165 11.045 -203.835 ;
        RECT 10.715 -205.525 11.045 -205.195 ;
        RECT 10.715 -206.885 11.045 -206.555 ;
        RECT 10.715 -208.245 11.045 -207.915 ;
        RECT 10.715 -209.605 11.045 -209.275 ;
        RECT 10.715 -210.965 11.045 -210.635 ;
        RECT 10.715 -212.325 11.045 -211.995 ;
        RECT 10.715 -213.685 11.045 -213.355 ;
        RECT 10.715 -215.045 11.045 -214.715 ;
        RECT 10.715 -216.405 11.045 -216.075 ;
        RECT 10.715 -217.765 11.045 -217.435 ;
        RECT 10.715 -219.125 11.045 -218.795 ;
        RECT 10.715 -220.485 11.045 -220.155 ;
        RECT 10.715 -221.845 11.045 -221.515 ;
        RECT 10.715 -223.205 11.045 -222.875 ;
        RECT 10.715 -224.565 11.045 -224.235 ;
        RECT 10.715 -225.925 11.045 -225.595 ;
        RECT 10.715 -227.285 11.045 -226.955 ;
        RECT 10.715 -228.645 11.045 -228.315 ;
        RECT 10.715 -230.005 11.045 -229.675 ;
        RECT 10.715 -231.365 11.045 -231.035 ;
        RECT 10.715 -232.725 11.045 -232.395 ;
        RECT 10.715 -234.085 11.045 -233.755 ;
        RECT 10.715 -235.445 11.045 -235.115 ;
        RECT 10.715 -236.805 11.045 -236.475 ;
        RECT 10.715 -238.165 11.045 -237.835 ;
        RECT 10.715 -243.81 11.045 -242.68 ;
        RECT 10.72 -243.925 11.04 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 246.76 12.405 247.89 ;
        RECT 12.075 241.915 12.405 242.245 ;
        RECT 12.075 240.555 12.405 240.885 ;
        RECT 12.075 239.195 12.405 239.525 ;
        RECT 12.075 237.835 12.405 238.165 ;
        RECT 12.08 237.16 12.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 -1.525 12.405 -1.195 ;
        RECT 12.075 -2.885 12.405 -2.555 ;
        RECT 12.08 -3.56 12.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 -122.565 12.405 -122.235 ;
        RECT 12.075 -123.925 12.405 -123.595 ;
        RECT 12.075 -125.285 12.405 -124.955 ;
        RECT 12.075 -126.645 12.405 -126.315 ;
        RECT 12.075 -128.005 12.405 -127.675 ;
        RECT 12.075 -129.365 12.405 -129.035 ;
        RECT 12.075 -130.725 12.405 -130.395 ;
        RECT 12.075 -132.085 12.405 -131.755 ;
        RECT 12.075 -133.445 12.405 -133.115 ;
        RECT 12.075 -134.805 12.405 -134.475 ;
        RECT 12.075 -136.165 12.405 -135.835 ;
        RECT 12.075 -137.525 12.405 -137.195 ;
        RECT 12.075 -138.885 12.405 -138.555 ;
        RECT 12.075 -140.245 12.405 -139.915 ;
        RECT 12.075 -141.605 12.405 -141.275 ;
        RECT 12.075 -142.965 12.405 -142.635 ;
        RECT 12.075 -144.325 12.405 -143.995 ;
        RECT 12.075 -145.685 12.405 -145.355 ;
        RECT 12.075 -147.045 12.405 -146.715 ;
        RECT 12.075 -148.405 12.405 -148.075 ;
        RECT 12.075 -149.765 12.405 -149.435 ;
        RECT 12.075 -151.125 12.405 -150.795 ;
        RECT 12.075 -152.485 12.405 -152.155 ;
        RECT 12.075 -153.845 12.405 -153.515 ;
        RECT 12.075 -155.205 12.405 -154.875 ;
        RECT 12.075 -156.565 12.405 -156.235 ;
        RECT 12.075 -157.925 12.405 -157.595 ;
        RECT 12.075 -159.285 12.405 -158.955 ;
        RECT 12.075 -160.645 12.405 -160.315 ;
        RECT 12.075 -162.005 12.405 -161.675 ;
        RECT 12.075 -163.365 12.405 -163.035 ;
        RECT 12.075 -164.725 12.405 -164.395 ;
        RECT 12.075 -166.085 12.405 -165.755 ;
        RECT 12.075 -167.445 12.405 -167.115 ;
        RECT 12.075 -168.805 12.405 -168.475 ;
        RECT 12.075 -170.165 12.405 -169.835 ;
        RECT 12.075 -171.525 12.405 -171.195 ;
        RECT 12.075 -172.885 12.405 -172.555 ;
        RECT 12.075 -174.245 12.405 -173.915 ;
        RECT 12.075 -175.605 12.405 -175.275 ;
        RECT 12.075 -176.965 12.405 -176.635 ;
        RECT 12.075 -178.325 12.405 -177.995 ;
        RECT 12.075 -179.685 12.405 -179.355 ;
        RECT 12.075 -181.045 12.405 -180.715 ;
        RECT 12.075 -182.405 12.405 -182.075 ;
        RECT 12.075 -183.765 12.405 -183.435 ;
        RECT 12.075 -185.125 12.405 -184.795 ;
        RECT 12.075 -186.485 12.405 -186.155 ;
        RECT 12.075 -187.845 12.405 -187.515 ;
        RECT 12.075 -189.205 12.405 -188.875 ;
        RECT 12.075 -190.565 12.405 -190.235 ;
        RECT 12.075 -191.925 12.405 -191.595 ;
        RECT 12.075 -193.285 12.405 -192.955 ;
        RECT 12.075 -194.645 12.405 -194.315 ;
        RECT 12.075 -196.005 12.405 -195.675 ;
        RECT 12.075 -197.365 12.405 -197.035 ;
        RECT 12.075 -198.725 12.405 -198.395 ;
        RECT 12.075 -200.085 12.405 -199.755 ;
        RECT 12.075 -201.445 12.405 -201.115 ;
        RECT 12.075 -202.805 12.405 -202.475 ;
        RECT 12.075 -204.165 12.405 -203.835 ;
        RECT 12.075 -205.525 12.405 -205.195 ;
        RECT 12.075 -206.885 12.405 -206.555 ;
        RECT 12.075 -208.245 12.405 -207.915 ;
        RECT 12.075 -209.605 12.405 -209.275 ;
        RECT 12.075 -210.965 12.405 -210.635 ;
        RECT 12.075 -212.325 12.405 -211.995 ;
        RECT 12.075 -213.685 12.405 -213.355 ;
        RECT 12.075 -215.045 12.405 -214.715 ;
        RECT 12.075 -216.405 12.405 -216.075 ;
        RECT 12.075 -217.765 12.405 -217.435 ;
        RECT 12.075 -219.125 12.405 -218.795 ;
        RECT 12.075 -220.485 12.405 -220.155 ;
        RECT 12.075 -221.845 12.405 -221.515 ;
        RECT 12.075 -223.205 12.405 -222.875 ;
        RECT 12.075 -224.565 12.405 -224.235 ;
        RECT 12.075 -225.925 12.405 -225.595 ;
        RECT 12.075 -227.285 12.405 -226.955 ;
        RECT 12.075 -228.645 12.405 -228.315 ;
        RECT 12.075 -230.005 12.405 -229.675 ;
        RECT 12.075 -231.365 12.405 -231.035 ;
        RECT 12.075 -232.725 12.405 -232.395 ;
        RECT 12.075 -234.085 12.405 -233.755 ;
        RECT 12.075 -235.445 12.405 -235.115 ;
        RECT 12.075 -236.805 12.405 -236.475 ;
        RECT 12.075 -238.165 12.405 -237.835 ;
        RECT 12.075 -243.81 12.405 -242.68 ;
        RECT 12.08 -243.925 12.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 246.76 13.765 247.89 ;
        RECT 13.435 241.915 13.765 242.245 ;
        RECT 13.435 240.555 13.765 240.885 ;
        RECT 13.435 239.195 13.765 239.525 ;
        RECT 13.435 237.835 13.765 238.165 ;
        RECT 13.44 237.16 13.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -126.645 13.765 -126.315 ;
        RECT 13.435 -128.005 13.765 -127.675 ;
        RECT 13.435 -129.365 13.765 -129.035 ;
        RECT 13.435 -130.725 13.765 -130.395 ;
        RECT 13.435 -132.085 13.765 -131.755 ;
        RECT 13.435 -133.445 13.765 -133.115 ;
        RECT 13.435 -134.805 13.765 -134.475 ;
        RECT 13.435 -136.165 13.765 -135.835 ;
        RECT 13.435 -137.525 13.765 -137.195 ;
        RECT 13.435 -138.885 13.765 -138.555 ;
        RECT 13.435 -140.245 13.765 -139.915 ;
        RECT 13.435 -141.605 13.765 -141.275 ;
        RECT 13.435 -142.965 13.765 -142.635 ;
        RECT 13.435 -144.325 13.765 -143.995 ;
        RECT 13.435 -145.685 13.765 -145.355 ;
        RECT 13.435 -147.045 13.765 -146.715 ;
        RECT 13.435 -148.405 13.765 -148.075 ;
        RECT 13.435 -149.765 13.765 -149.435 ;
        RECT 13.435 -151.125 13.765 -150.795 ;
        RECT 13.435 -152.485 13.765 -152.155 ;
        RECT 13.435 -153.845 13.765 -153.515 ;
        RECT 13.435 -155.205 13.765 -154.875 ;
        RECT 13.435 -156.565 13.765 -156.235 ;
        RECT 13.435 -157.925 13.765 -157.595 ;
        RECT 13.435 -159.285 13.765 -158.955 ;
        RECT 13.435 -160.645 13.765 -160.315 ;
        RECT 13.435 -162.005 13.765 -161.675 ;
        RECT 13.435 -163.365 13.765 -163.035 ;
        RECT 13.435 -164.725 13.765 -164.395 ;
        RECT 13.435 -166.085 13.765 -165.755 ;
        RECT 13.435 -167.445 13.765 -167.115 ;
        RECT 13.435 -168.805 13.765 -168.475 ;
        RECT 13.435 -170.165 13.765 -169.835 ;
        RECT 13.435 -171.525 13.765 -171.195 ;
        RECT 13.435 -172.885 13.765 -172.555 ;
        RECT 13.435 -174.245 13.765 -173.915 ;
        RECT 13.435 -175.605 13.765 -175.275 ;
        RECT 13.435 -176.965 13.765 -176.635 ;
        RECT 13.435 -178.325 13.765 -177.995 ;
        RECT 13.435 -179.685 13.765 -179.355 ;
        RECT 13.435 -181.045 13.765 -180.715 ;
        RECT 13.435 -182.405 13.765 -182.075 ;
        RECT 13.435 -183.765 13.765 -183.435 ;
        RECT 13.435 -185.125 13.765 -184.795 ;
        RECT 13.435 -186.485 13.765 -186.155 ;
        RECT 13.435 -187.845 13.765 -187.515 ;
        RECT 13.435 -189.205 13.765 -188.875 ;
        RECT 13.435 -190.565 13.765 -190.235 ;
        RECT 13.435 -191.925 13.765 -191.595 ;
        RECT 13.435 -193.285 13.765 -192.955 ;
        RECT 13.435 -194.645 13.765 -194.315 ;
        RECT 13.435 -196.005 13.765 -195.675 ;
        RECT 13.435 -197.365 13.765 -197.035 ;
        RECT 13.435 -198.725 13.765 -198.395 ;
        RECT 13.435 -200.085 13.765 -199.755 ;
        RECT 13.435 -201.445 13.765 -201.115 ;
        RECT 13.435 -202.805 13.765 -202.475 ;
        RECT 13.435 -204.165 13.765 -203.835 ;
        RECT 13.435 -205.525 13.765 -205.195 ;
        RECT 13.435 -206.885 13.765 -206.555 ;
        RECT 13.435 -208.245 13.765 -207.915 ;
        RECT 13.435 -209.605 13.765 -209.275 ;
        RECT 13.435 -210.965 13.765 -210.635 ;
        RECT 13.435 -212.325 13.765 -211.995 ;
        RECT 13.435 -213.685 13.765 -213.355 ;
        RECT 13.435 -215.045 13.765 -214.715 ;
        RECT 13.435 -216.405 13.765 -216.075 ;
        RECT 13.435 -217.765 13.765 -217.435 ;
        RECT 13.435 -219.125 13.765 -218.795 ;
        RECT 13.435 -220.485 13.765 -220.155 ;
        RECT 13.435 -221.845 13.765 -221.515 ;
        RECT 13.435 -223.205 13.765 -222.875 ;
        RECT 13.435 -224.565 13.765 -224.235 ;
        RECT 13.435 -225.925 13.765 -225.595 ;
        RECT 13.435 -227.285 13.765 -226.955 ;
        RECT 13.435 -228.645 13.765 -228.315 ;
        RECT 13.435 -230.005 13.765 -229.675 ;
        RECT 13.435 -231.365 13.765 -231.035 ;
        RECT 13.435 -232.725 13.765 -232.395 ;
        RECT 13.435 -234.085 13.765 -233.755 ;
        RECT 13.435 -235.445 13.765 -235.115 ;
        RECT 13.435 -236.805 13.765 -236.475 ;
        RECT 13.435 -238.165 13.765 -237.835 ;
        RECT 13.435 -243.81 13.765 -242.68 ;
        RECT 13.44 -243.925 13.76 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.56 -125.535 13.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 246.76 15.125 247.89 ;
        RECT 14.795 241.915 15.125 242.245 ;
        RECT 14.795 240.555 15.125 240.885 ;
        RECT 14.795 239.195 15.125 239.525 ;
        RECT 14.795 237.835 15.125 238.165 ;
        RECT 14.8 237.16 15.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 246.76 16.485 247.89 ;
        RECT 16.155 241.915 16.485 242.245 ;
        RECT 16.155 240.555 16.485 240.885 ;
        RECT 16.155 239.195 16.485 239.525 ;
        RECT 16.155 237.835 16.485 238.165 ;
        RECT 16.16 237.16 16.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 -1.525 16.485 -1.195 ;
        RECT 16.155 -2.885 16.485 -2.555 ;
        RECT 16.16 -3.56 16.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 246.76 17.845 247.89 ;
        RECT 17.515 241.915 17.845 242.245 ;
        RECT 17.515 240.555 17.845 240.885 ;
        RECT 17.515 239.195 17.845 239.525 ;
        RECT 17.515 237.835 17.845 238.165 ;
        RECT 17.52 237.16 17.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -1.525 17.845 -1.195 ;
        RECT 17.515 -2.885 17.845 -2.555 ;
        RECT 17.52 -3.56 17.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -122.565 17.845 -122.235 ;
        RECT 17.515 -123.925 17.845 -123.595 ;
        RECT 17.515 -125.285 17.845 -124.955 ;
        RECT 17.515 -126.645 17.845 -126.315 ;
        RECT 17.515 -128.005 17.845 -127.675 ;
        RECT 17.515 -129.365 17.845 -129.035 ;
        RECT 17.515 -130.725 17.845 -130.395 ;
        RECT 17.515 -132.085 17.845 -131.755 ;
        RECT 17.515 -133.445 17.845 -133.115 ;
        RECT 17.515 -134.805 17.845 -134.475 ;
        RECT 17.515 -136.165 17.845 -135.835 ;
        RECT 17.515 -137.525 17.845 -137.195 ;
        RECT 17.515 -138.885 17.845 -138.555 ;
        RECT 17.515 -140.245 17.845 -139.915 ;
        RECT 17.515 -141.605 17.845 -141.275 ;
        RECT 17.515 -142.965 17.845 -142.635 ;
        RECT 17.515 -144.325 17.845 -143.995 ;
        RECT 17.515 -145.685 17.845 -145.355 ;
        RECT 17.515 -147.045 17.845 -146.715 ;
        RECT 17.515 -148.405 17.845 -148.075 ;
        RECT 17.515 -149.765 17.845 -149.435 ;
        RECT 17.515 -151.125 17.845 -150.795 ;
        RECT 17.515 -152.485 17.845 -152.155 ;
        RECT 17.515 -153.845 17.845 -153.515 ;
        RECT 17.515 -155.205 17.845 -154.875 ;
        RECT 17.515 -156.565 17.845 -156.235 ;
        RECT 17.515 -157.925 17.845 -157.595 ;
        RECT 17.515 -159.285 17.845 -158.955 ;
        RECT 17.515 -160.645 17.845 -160.315 ;
        RECT 17.515 -162.005 17.845 -161.675 ;
        RECT 17.515 -163.365 17.845 -163.035 ;
        RECT 17.515 -164.725 17.845 -164.395 ;
        RECT 17.515 -166.085 17.845 -165.755 ;
        RECT 17.515 -167.445 17.845 -167.115 ;
        RECT 17.515 -168.805 17.845 -168.475 ;
        RECT 17.515 -170.165 17.845 -169.835 ;
        RECT 17.515 -171.525 17.845 -171.195 ;
        RECT 17.515 -172.885 17.845 -172.555 ;
        RECT 17.515 -174.245 17.845 -173.915 ;
        RECT 17.515 -175.605 17.845 -175.275 ;
        RECT 17.515 -176.965 17.845 -176.635 ;
        RECT 17.515 -178.325 17.845 -177.995 ;
        RECT 17.515 -179.685 17.845 -179.355 ;
        RECT 17.515 -181.045 17.845 -180.715 ;
        RECT 17.515 -182.405 17.845 -182.075 ;
        RECT 17.515 -183.765 17.845 -183.435 ;
        RECT 17.515 -185.125 17.845 -184.795 ;
        RECT 17.515 -186.485 17.845 -186.155 ;
        RECT 17.515 -187.845 17.845 -187.515 ;
        RECT 17.515 -189.205 17.845 -188.875 ;
        RECT 17.515 -190.565 17.845 -190.235 ;
        RECT 17.515 -191.925 17.845 -191.595 ;
        RECT 17.515 -193.285 17.845 -192.955 ;
        RECT 17.515 -194.645 17.845 -194.315 ;
        RECT 17.515 -196.005 17.845 -195.675 ;
        RECT 17.515 -197.365 17.845 -197.035 ;
        RECT 17.515 -198.725 17.845 -198.395 ;
        RECT 17.515 -200.085 17.845 -199.755 ;
        RECT 17.515 -201.445 17.845 -201.115 ;
        RECT 17.515 -202.805 17.845 -202.475 ;
        RECT 17.515 -204.165 17.845 -203.835 ;
        RECT 17.515 -205.525 17.845 -205.195 ;
        RECT 17.515 -206.885 17.845 -206.555 ;
        RECT 17.515 -208.245 17.845 -207.915 ;
        RECT 17.515 -209.605 17.845 -209.275 ;
        RECT 17.515 -210.965 17.845 -210.635 ;
        RECT 17.515 -212.325 17.845 -211.995 ;
        RECT 17.515 -213.685 17.845 -213.355 ;
        RECT 17.515 -215.045 17.845 -214.715 ;
        RECT 17.515 -216.405 17.845 -216.075 ;
        RECT 17.515 -217.765 17.845 -217.435 ;
        RECT 17.515 -219.125 17.845 -218.795 ;
        RECT 17.515 -220.485 17.845 -220.155 ;
        RECT 17.515 -221.845 17.845 -221.515 ;
        RECT 17.515 -223.205 17.845 -222.875 ;
        RECT 17.515 -224.565 17.845 -224.235 ;
        RECT 17.515 -225.925 17.845 -225.595 ;
        RECT 17.515 -227.285 17.845 -226.955 ;
        RECT 17.515 -228.645 17.845 -228.315 ;
        RECT 17.515 -230.005 17.845 -229.675 ;
        RECT 17.515 -231.365 17.845 -231.035 ;
        RECT 17.515 -232.725 17.845 -232.395 ;
        RECT 17.515 -234.085 17.845 -233.755 ;
        RECT 17.515 -235.445 17.845 -235.115 ;
        RECT 17.515 -236.805 17.845 -236.475 ;
        RECT 17.515 -238.165 17.845 -237.835 ;
        RECT 17.515 -243.81 17.845 -242.68 ;
        RECT 17.52 -243.925 17.84 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 246.76 19.205 247.89 ;
        RECT 18.875 241.915 19.205 242.245 ;
        RECT 18.875 240.555 19.205 240.885 ;
        RECT 18.875 239.195 19.205 239.525 ;
        RECT 18.875 237.835 19.205 238.165 ;
        RECT 18.88 237.16 19.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -1.525 19.205 -1.195 ;
        RECT 18.875 -2.885 19.205 -2.555 ;
        RECT 18.88 -3.56 19.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -182.405 19.205 -182.075 ;
        RECT 18.875 -183.765 19.205 -183.435 ;
        RECT 18.875 -185.125 19.205 -184.795 ;
        RECT 18.875 -186.485 19.205 -186.155 ;
        RECT 18.875 -187.845 19.205 -187.515 ;
        RECT 18.875 -189.205 19.205 -188.875 ;
        RECT 18.875 -190.565 19.205 -190.235 ;
        RECT 18.875 -191.925 19.205 -191.595 ;
        RECT 18.875 -193.285 19.205 -192.955 ;
        RECT 18.875 -194.645 19.205 -194.315 ;
        RECT 18.875 -196.005 19.205 -195.675 ;
        RECT 18.875 -197.365 19.205 -197.035 ;
        RECT 18.875 -198.725 19.205 -198.395 ;
        RECT 18.875 -200.085 19.205 -199.755 ;
        RECT 18.875 -201.445 19.205 -201.115 ;
        RECT 18.875 -202.805 19.205 -202.475 ;
        RECT 18.875 -204.165 19.205 -203.835 ;
        RECT 18.875 -205.525 19.205 -205.195 ;
        RECT 18.875 -206.885 19.205 -206.555 ;
        RECT 18.875 -208.245 19.205 -207.915 ;
        RECT 18.875 -209.605 19.205 -209.275 ;
        RECT 18.875 -210.965 19.205 -210.635 ;
        RECT 18.875 -212.325 19.205 -211.995 ;
        RECT 18.875 -213.685 19.205 -213.355 ;
        RECT 18.875 -215.045 19.205 -214.715 ;
        RECT 18.875 -216.405 19.205 -216.075 ;
        RECT 18.875 -217.765 19.205 -217.435 ;
        RECT 18.875 -219.125 19.205 -218.795 ;
        RECT 18.875 -220.485 19.205 -220.155 ;
        RECT 18.875 -221.845 19.205 -221.515 ;
        RECT 18.875 -223.205 19.205 -222.875 ;
        RECT 18.875 -224.565 19.205 -224.235 ;
        RECT 18.875 -225.925 19.205 -225.595 ;
        RECT 18.875 -227.285 19.205 -226.955 ;
        RECT 18.875 -228.645 19.205 -228.315 ;
        RECT 18.875 -230.005 19.205 -229.675 ;
        RECT 18.875 -231.365 19.205 -231.035 ;
        RECT 18.875 -232.725 19.205 -232.395 ;
        RECT 18.875 -234.085 19.205 -233.755 ;
        RECT 18.875 -235.445 19.205 -235.115 ;
        RECT 18.875 -236.805 19.205 -236.475 ;
        RECT 18.875 -238.165 19.205 -237.835 ;
        RECT 18.875 -243.81 19.205 -242.68 ;
        RECT 18.88 -243.925 19.2 -122.235 ;
        RECT 18.875 -122.565 19.205 -122.235 ;
        RECT 18.875 -123.925 19.205 -123.595 ;
        RECT 18.875 -125.285 19.205 -124.955 ;
        RECT 18.875 -126.645 19.205 -126.315 ;
        RECT 18.875 -128.005 19.205 -127.675 ;
        RECT 18.875 -129.365 19.205 -129.035 ;
        RECT 18.875 -130.725 19.205 -130.395 ;
        RECT 18.875 -132.085 19.205 -131.755 ;
        RECT 18.875 -133.445 19.205 -133.115 ;
        RECT 18.875 -134.805 19.205 -134.475 ;
        RECT 18.875 -136.165 19.205 -135.835 ;
        RECT 18.875 -137.525 19.205 -137.195 ;
        RECT 18.875 -138.885 19.205 -138.555 ;
        RECT 18.875 -140.245 19.205 -139.915 ;
        RECT 18.875 -141.605 19.205 -141.275 ;
        RECT 18.875 -142.965 19.205 -142.635 ;
        RECT 18.875 -144.325 19.205 -143.995 ;
        RECT 18.875 -145.685 19.205 -145.355 ;
        RECT 18.875 -147.045 19.205 -146.715 ;
        RECT 18.875 -148.405 19.205 -148.075 ;
        RECT 18.875 -149.765 19.205 -149.435 ;
        RECT 18.875 -151.125 19.205 -150.795 ;
        RECT 18.875 -152.485 19.205 -152.155 ;
        RECT 18.875 -153.845 19.205 -153.515 ;
        RECT 18.875 -155.205 19.205 -154.875 ;
        RECT 18.875 -156.565 19.205 -156.235 ;
        RECT 18.875 -157.925 19.205 -157.595 ;
        RECT 18.875 -159.285 19.205 -158.955 ;
        RECT 18.875 -160.645 19.205 -160.315 ;
        RECT 18.875 -162.005 19.205 -161.675 ;
        RECT 18.875 -163.365 19.205 -163.035 ;
        RECT 18.875 -164.725 19.205 -164.395 ;
        RECT 18.875 -166.085 19.205 -165.755 ;
        RECT 18.875 -167.445 19.205 -167.115 ;
        RECT 18.875 -168.805 19.205 -168.475 ;
        RECT 18.875 -170.165 19.205 -169.835 ;
        RECT 18.875 -171.525 19.205 -171.195 ;
        RECT 18.875 -172.885 19.205 -172.555 ;
        RECT 18.875 -174.245 19.205 -173.915 ;
        RECT 18.875 -175.605 19.205 -175.275 ;
        RECT 18.875 -176.965 19.205 -176.635 ;
        RECT 18.875 -178.325 19.205 -177.995 ;
        RECT 18.875 -179.685 19.205 -179.355 ;
        RECT 18.875 -181.045 19.205 -180.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.245 246.76 -3.915 247.89 ;
        RECT -4.245 241.915 -3.915 242.245 ;
        RECT -4.245 240.555 -3.915 240.885 ;
        RECT -4.245 239.195 -3.915 239.525 ;
        RECT -4.245 237.835 -3.915 238.165 ;
        RECT -4.245 235.17 -3.915 235.5 ;
        RECT -4.245 232.995 -3.915 233.325 ;
        RECT -4.245 231.415 -3.915 231.745 ;
        RECT -4.245 230.565 -3.915 230.895 ;
        RECT -4.245 228.255 -3.915 228.585 ;
        RECT -4.245 227.405 -3.915 227.735 ;
        RECT -4.245 225.095 -3.915 225.425 ;
        RECT -4.245 224.245 -3.915 224.575 ;
        RECT -4.245 221.935 -3.915 222.265 ;
        RECT -4.245 221.085 -3.915 221.415 ;
        RECT -4.245 218.775 -3.915 219.105 ;
        RECT -4.245 217.195 -3.915 217.525 ;
        RECT -4.245 216.345 -3.915 216.675 ;
        RECT -4.245 214.035 -3.915 214.365 ;
        RECT -4.245 213.185 -3.915 213.515 ;
        RECT -4.245 210.875 -3.915 211.205 ;
        RECT -4.245 210.025 -3.915 210.355 ;
        RECT -4.245 207.715 -3.915 208.045 ;
        RECT -4.245 206.865 -3.915 207.195 ;
        RECT -4.245 204.555 -3.915 204.885 ;
        RECT -4.245 202.975 -3.915 203.305 ;
        RECT -4.245 202.125 -3.915 202.455 ;
        RECT -4.245 199.815 -3.915 200.145 ;
        RECT -4.245 198.965 -3.915 199.295 ;
        RECT -4.245 196.655 -3.915 196.985 ;
        RECT -4.245 195.805 -3.915 196.135 ;
        RECT -4.245 193.495 -3.915 193.825 ;
        RECT -4.245 192.645 -3.915 192.975 ;
        RECT -4.245 190.335 -3.915 190.665 ;
        RECT -4.245 188.755 -3.915 189.085 ;
        RECT -4.245 187.905 -3.915 188.235 ;
        RECT -4.245 185.595 -3.915 185.925 ;
        RECT -4.245 184.745 -3.915 185.075 ;
        RECT -4.245 182.435 -3.915 182.765 ;
        RECT -4.245 181.585 -3.915 181.915 ;
        RECT -4.245 179.275 -3.915 179.605 ;
        RECT -4.245 178.425 -3.915 178.755 ;
        RECT -4.245 176.115 -3.915 176.445 ;
        RECT -4.245 174.535 -3.915 174.865 ;
        RECT -4.245 173.685 -3.915 174.015 ;
        RECT -4.245 171.375 -3.915 171.705 ;
        RECT -4.245 170.525 -3.915 170.855 ;
        RECT -4.245 168.215 -3.915 168.545 ;
        RECT -4.245 167.365 -3.915 167.695 ;
        RECT -4.245 165.055 -3.915 165.385 ;
        RECT -4.245 164.205 -3.915 164.535 ;
        RECT -4.245 161.895 -3.915 162.225 ;
        RECT -4.245 160.315 -3.915 160.645 ;
        RECT -4.245 159.465 -3.915 159.795 ;
        RECT -4.245 157.155 -3.915 157.485 ;
        RECT -4.245 156.305 -3.915 156.635 ;
        RECT -4.245 153.995 -3.915 154.325 ;
        RECT -4.245 153.145 -3.915 153.475 ;
        RECT -4.245 150.835 -3.915 151.165 ;
        RECT -4.245 149.985 -3.915 150.315 ;
        RECT -4.245 147.675 -3.915 148.005 ;
        RECT -4.245 146.095 -3.915 146.425 ;
        RECT -4.245 145.245 -3.915 145.575 ;
        RECT -4.245 142.935 -3.915 143.265 ;
        RECT -4.245 142.085 -3.915 142.415 ;
        RECT -4.245 139.775 -3.915 140.105 ;
        RECT -4.245 138.925 -3.915 139.255 ;
        RECT -4.245 136.615 -3.915 136.945 ;
        RECT -4.245 135.765 -3.915 136.095 ;
        RECT -4.245 133.455 -3.915 133.785 ;
        RECT -4.245 131.875 -3.915 132.205 ;
        RECT -4.245 131.025 -3.915 131.355 ;
        RECT -4.245 128.715 -3.915 129.045 ;
        RECT -4.245 127.865 -3.915 128.195 ;
        RECT -4.245 125.555 -3.915 125.885 ;
        RECT -4.245 124.705 -3.915 125.035 ;
        RECT -4.245 122.395 -3.915 122.725 ;
        RECT -4.245 121.545 -3.915 121.875 ;
        RECT -4.245 119.235 -3.915 119.565 ;
        RECT -4.245 117.655 -3.915 117.985 ;
        RECT -4.245 116.805 -3.915 117.135 ;
        RECT -4.245 114.495 -3.915 114.825 ;
        RECT -4.245 113.645 -3.915 113.975 ;
        RECT -4.245 111.335 -3.915 111.665 ;
        RECT -4.245 110.485 -3.915 110.815 ;
        RECT -4.245 108.175 -3.915 108.505 ;
        RECT -4.245 107.325 -3.915 107.655 ;
        RECT -4.245 105.015 -3.915 105.345 ;
        RECT -4.245 103.435 -3.915 103.765 ;
        RECT -4.245 102.585 -3.915 102.915 ;
        RECT -4.245 100.275 -3.915 100.605 ;
        RECT -4.245 99.425 -3.915 99.755 ;
        RECT -4.245 97.115 -3.915 97.445 ;
        RECT -4.245 96.265 -3.915 96.595 ;
        RECT -4.245 93.955 -3.915 94.285 ;
        RECT -4.245 93.105 -3.915 93.435 ;
        RECT -4.245 90.795 -3.915 91.125 ;
        RECT -4.245 89.215 -3.915 89.545 ;
        RECT -4.245 88.365 -3.915 88.695 ;
        RECT -4.245 86.055 -3.915 86.385 ;
        RECT -4.245 85.205 -3.915 85.535 ;
        RECT -4.245 82.895 -3.915 83.225 ;
        RECT -4.245 82.045 -3.915 82.375 ;
        RECT -4.245 79.735 -3.915 80.065 ;
        RECT -4.245 78.885 -3.915 79.215 ;
        RECT -4.245 76.575 -3.915 76.905 ;
        RECT -4.245 74.995 -3.915 75.325 ;
        RECT -4.245 74.145 -3.915 74.475 ;
        RECT -4.245 71.835 -3.915 72.165 ;
        RECT -4.245 70.985 -3.915 71.315 ;
        RECT -4.245 68.675 -3.915 69.005 ;
        RECT -4.245 67.825 -3.915 68.155 ;
        RECT -4.245 65.515 -3.915 65.845 ;
        RECT -4.245 64.665 -3.915 64.995 ;
        RECT -4.245 62.355 -3.915 62.685 ;
        RECT -4.245 60.775 -3.915 61.105 ;
        RECT -4.245 59.925 -3.915 60.255 ;
        RECT -4.245 57.615 -3.915 57.945 ;
        RECT -4.245 56.765 -3.915 57.095 ;
        RECT -4.245 54.455 -3.915 54.785 ;
        RECT -4.245 53.605 -3.915 53.935 ;
        RECT -4.245 51.295 -3.915 51.625 ;
        RECT -4.245 50.445 -3.915 50.775 ;
        RECT -4.245 48.135 -3.915 48.465 ;
        RECT -4.245 46.555 -3.915 46.885 ;
        RECT -4.245 45.705 -3.915 46.035 ;
        RECT -4.245 43.395 -3.915 43.725 ;
        RECT -4.245 42.545 -3.915 42.875 ;
        RECT -4.245 40.235 -3.915 40.565 ;
        RECT -4.245 39.385 -3.915 39.715 ;
        RECT -4.245 37.075 -3.915 37.405 ;
        RECT -4.245 36.225 -3.915 36.555 ;
        RECT -4.245 33.915 -3.915 34.245 ;
        RECT -4.245 32.335 -3.915 32.665 ;
        RECT -4.245 31.485 -3.915 31.815 ;
        RECT -4.245 29.175 -3.915 29.505 ;
        RECT -4.245 28.325 -3.915 28.655 ;
        RECT -4.245 26.015 -3.915 26.345 ;
        RECT -4.245 25.165 -3.915 25.495 ;
        RECT -4.245 22.855 -3.915 23.185 ;
        RECT -4.245 22.005 -3.915 22.335 ;
        RECT -4.245 19.695 -3.915 20.025 ;
        RECT -4.245 18.115 -3.915 18.445 ;
        RECT -4.245 17.265 -3.915 17.595 ;
        RECT -4.245 14.955 -3.915 15.285 ;
        RECT -4.245 14.105 -3.915 14.435 ;
        RECT -4.245 11.795 -3.915 12.125 ;
        RECT -4.245 10.945 -3.915 11.275 ;
        RECT -4.245 8.635 -3.915 8.965 ;
        RECT -4.245 7.785 -3.915 8.115 ;
        RECT -4.245 5.475 -3.915 5.805 ;
        RECT -4.245 3.895 -3.915 4.225 ;
        RECT -4.245 3.045 -3.915 3.375 ;
        RECT -4.245 0.87 -3.915 1.2 ;
        RECT -4.245 -1.525 -3.915 -1.195 ;
        RECT -4.245 -2.885 -3.915 -2.555 ;
        RECT -4.245 -4.245 -3.915 -3.915 ;
        RECT -4.245 -5.605 -3.915 -5.275 ;
        RECT -4.245 -6.965 -3.915 -6.635 ;
        RECT -4.245 -8.325 -3.915 -7.995 ;
        RECT -4.245 -9.685 -3.915 -9.355 ;
        RECT -4.245 -12.405 -3.915 -12.075 ;
        RECT -4.245 -13.765 -3.915 -13.435 ;
        RECT -4.245 -15.125 -3.915 -14.795 ;
        RECT -4.245 -16.485 -3.915 -16.155 ;
        RECT -4.245 -17.845 -3.915 -17.515 ;
        RECT -4.245 -19.205 -3.915 -18.875 ;
        RECT -4.245 -20.565 -3.915 -20.235 ;
        RECT -4.245 -21.925 -3.915 -21.595 ;
        RECT -4.245 -23.285 -3.915 -22.955 ;
        RECT -4.245 -24.645 -3.915 -24.315 ;
        RECT -4.245 -26.005 -3.915 -25.675 ;
        RECT -4.245 -27.365 -3.915 -27.035 ;
        RECT -4.245 -28.725 -3.915 -28.395 ;
        RECT -4.245 -30.085 -3.915 -29.755 ;
        RECT -4.245 -31.445 -3.915 -31.115 ;
        RECT -4.245 -32.805 -3.915 -32.475 ;
        RECT -4.245 -34.165 -3.915 -33.835 ;
        RECT -4.245 -35.525 -3.915 -35.195 ;
        RECT -4.245 -36.885 -3.915 -36.555 ;
        RECT -4.245 -38.245 -3.915 -37.915 ;
        RECT -4.245 -39.605 -3.915 -39.275 ;
        RECT -4.245 -40.965 -3.915 -40.635 ;
        RECT -4.245 -42.325 -3.915 -41.995 ;
        RECT -4.245 -43.685 -3.915 -43.355 ;
        RECT -4.245 -45.045 -3.915 -44.715 ;
        RECT -4.245 -46.405 -3.915 -46.075 ;
        RECT -4.245 -47.765 -3.915 -47.435 ;
        RECT -4.245 -49.125 -3.915 -48.795 ;
        RECT -4.245 -50.485 -3.915 -50.155 ;
        RECT -4.245 -51.845 -3.915 -51.515 ;
        RECT -4.245 -53.205 -3.915 -52.875 ;
        RECT -4.245 -54.565 -3.915 -54.235 ;
        RECT -4.245 -55.925 -3.915 -55.595 ;
        RECT -4.245 -57.285 -3.915 -56.955 ;
        RECT -4.245 -58.645 -3.915 -58.315 ;
        RECT -4.245 -60.005 -3.915 -59.675 ;
        RECT -4.245 -61.365 -3.915 -61.035 ;
        RECT -4.245 -68.165 -3.915 -67.835 ;
        RECT -4.245 -69.525 -3.915 -69.195 ;
        RECT -4.245 -70.885 -3.915 -70.555 ;
        RECT -4.245 -72.245 -3.915 -71.915 ;
        RECT -4.245 -73.605 -3.915 -73.275 ;
        RECT -4.245 -74.965 -3.915 -74.635 ;
        RECT -4.245 -76.325 -3.915 -75.995 ;
        RECT -4.245 -77.685 -3.915 -77.355 ;
        RECT -4.245 -79.045 -3.915 -78.715 ;
        RECT -4.245 -80.405 -3.915 -80.075 ;
        RECT -4.245 -81.765 -3.915 -81.435 ;
        RECT -4.245 -83.125 -3.915 -82.795 ;
        RECT -4.245 -84.485 -3.915 -84.155 ;
        RECT -4.245 -85.845 -3.915 -85.515 ;
        RECT -4.245 -87.205 -3.915 -86.875 ;
        RECT -4.245 -88.565 -3.915 -88.235 ;
        RECT -4.245 -89.925 -3.915 -89.595 ;
        RECT -4.245 -91.285 -3.915 -90.955 ;
        RECT -4.245 -92.645 -3.915 -92.315 ;
        RECT -4.245 -94.005 -3.915 -93.675 ;
        RECT -4.245 -95.365 -3.915 -95.035 ;
        RECT -4.245 -96.725 -3.915 -96.395 ;
        RECT -4.245 -98.085 -3.915 -97.755 ;
        RECT -4.245 -99.445 -3.915 -99.115 ;
        RECT -4.245 -100.805 -3.915 -100.475 ;
        RECT -4.245 -102.165 -3.915 -101.835 ;
        RECT -4.245 -103.525 -3.915 -103.195 ;
        RECT -4.245 -104.885 -3.915 -104.555 ;
        RECT -4.245 -106.245 -3.915 -105.915 ;
        RECT -4.245 -107.605 -3.915 -107.275 ;
        RECT -4.245 -108.965 -3.915 -108.635 ;
        RECT -4.245 -110.325 -3.915 -109.995 ;
        RECT -4.245 -111.685 -3.915 -111.355 ;
        RECT -4.245 -113.045 -3.915 -112.715 ;
        RECT -4.245 -114.405 -3.915 -114.075 ;
        RECT -4.245 -115.765 -3.915 -115.435 ;
        RECT -4.245 -117.125 -3.915 -116.795 ;
        RECT -4.245 -118.485 -3.915 -118.155 ;
        RECT -4.245 -119.845 -3.915 -119.515 ;
        RECT -4.245 -121.205 -3.915 -120.875 ;
        RECT -4.245 -122.565 -3.915 -122.235 ;
        RECT -4.245 -123.925 -3.915 -123.595 ;
        RECT -4.245 -125.285 -3.915 -124.955 ;
        RECT -4.245 -126.645 -3.915 -126.315 ;
        RECT -4.245 -128.005 -3.915 -127.675 ;
        RECT -4.245 -129.365 -3.915 -129.035 ;
        RECT -4.245 -130.725 -3.915 -130.395 ;
        RECT -4.245 -132.085 -3.915 -131.755 ;
        RECT -4.245 -133.445 -3.915 -133.115 ;
        RECT -4.245 -140.245 -3.915 -139.915 ;
        RECT -4.245 -141.605 -3.915 -141.275 ;
        RECT -4.245 -142.965 -3.915 -142.635 ;
        RECT -4.245 -144.325 -3.915 -143.995 ;
        RECT -4.245 -145.685 -3.915 -145.355 ;
        RECT -4.245 -147.045 -3.915 -146.715 ;
        RECT -4.245 -148.405 -3.915 -148.075 ;
        RECT -4.245 -149.765 -3.915 -149.435 ;
        RECT -4.245 -151.125 -3.915 -150.795 ;
        RECT -4.245 -152.485 -3.915 -152.155 ;
        RECT -4.245 -153.845 -3.915 -153.515 ;
        RECT -4.245 -155.205 -3.915 -154.875 ;
        RECT -4.245 -156.565 -3.915 -156.235 ;
        RECT -4.245 -157.925 -3.915 -157.595 ;
        RECT -4.245 -160.645 -3.915 -160.315 ;
        RECT -4.245 -162.005 -3.915 -161.675 ;
        RECT -4.245 -163.365 -3.915 -163.035 ;
        RECT -4.245 -164.725 -3.915 -164.395 ;
        RECT -4.245 -166.085 -3.915 -165.755 ;
        RECT -4.245 -167.445 -3.915 -167.115 ;
        RECT -4.245 -168.805 -3.915 -168.475 ;
        RECT -4.245 -170.165 -3.915 -169.835 ;
        RECT -4.245 -171.525 -3.915 -171.195 ;
        RECT -4.245 -172.885 -3.915 -172.555 ;
        RECT -4.245 -174.245 -3.915 -173.915 ;
        RECT -4.245 -175.605 -3.915 -175.275 ;
        RECT -4.245 -176.965 -3.915 -176.635 ;
        RECT -4.245 -178.325 -3.915 -177.995 ;
        RECT -4.245 -179.685 -3.915 -179.355 ;
        RECT -4.245 -181.045 -3.915 -180.715 ;
        RECT -4.245 -182.405 -3.915 -182.075 ;
        RECT -4.245 -183.765 -3.915 -183.435 ;
        RECT -4.245 -185.125 -3.915 -184.795 ;
        RECT -4.245 -186.485 -3.915 -186.155 ;
        RECT -4.245 -187.845 -3.915 -187.515 ;
        RECT -4.245 -189.205 -3.915 -188.875 ;
        RECT -4.245 -190.565 -3.915 -190.235 ;
        RECT -4.245 -191.925 -3.915 -191.595 ;
        RECT -4.245 -193.285 -3.915 -192.955 ;
        RECT -4.245 -194.645 -3.915 -194.315 ;
        RECT -4.245 -196.005 -3.915 -195.675 ;
        RECT -4.245 -197.365 -3.915 -197.035 ;
        RECT -4.245 -198.725 -3.915 -198.395 ;
        RECT -4.245 -200.085 -3.915 -199.755 ;
        RECT -4.245 -201.445 -3.915 -201.115 ;
        RECT -4.245 -202.805 -3.915 -202.475 ;
        RECT -4.245 -204.165 -3.915 -203.835 ;
        RECT -4.245 -205.525 -3.915 -205.195 ;
        RECT -4.245 -206.885 -3.915 -206.555 ;
        RECT -4.245 -208.245 -3.915 -207.915 ;
        RECT -4.245 -209.605 -3.915 -209.275 ;
        RECT -4.245 -210.965 -3.915 -210.635 ;
        RECT -4.245 -212.325 -3.915 -211.995 ;
        RECT -4.245 -213.685 -3.915 -213.355 ;
        RECT -4.245 -215.045 -3.915 -214.715 ;
        RECT -4.245 -216.405 -3.915 -216.075 ;
        RECT -4.245 -217.765 -3.915 -217.435 ;
        RECT -4.245 -219.125 -3.915 -218.795 ;
        RECT -4.245 -220.485 -3.915 -220.155 ;
        RECT -4.245 -221.845 -3.915 -221.515 ;
        RECT -4.245 -223.205 -3.915 -222.875 ;
        RECT -4.245 -224.565 -3.915 -224.235 ;
        RECT -4.245 -225.925 -3.915 -225.595 ;
        RECT -4.245 -227.285 -3.915 -226.955 ;
        RECT -4.245 -228.645 -3.915 -228.315 ;
        RECT -4.245 -230.005 -3.915 -229.675 ;
        RECT -4.245 -231.365 -3.915 -231.035 ;
        RECT -4.245 -232.725 -3.915 -232.395 ;
        RECT -4.245 -234.085 -3.915 -233.755 ;
        RECT -4.245 -235.445 -3.915 -235.115 ;
        RECT -4.245 -236.805 -3.915 -236.475 ;
        RECT -4.245 -238.165 -3.915 -237.835 ;
        RECT -4.245 -243.81 -3.915 -242.68 ;
        RECT -4.24 -243.925 -3.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.885 246.76 -2.555 247.89 ;
        RECT -2.885 241.915 -2.555 242.245 ;
        RECT -2.885 240.555 -2.555 240.885 ;
        RECT -2.885 239.195 -2.555 239.525 ;
        RECT -2.885 237.835 -2.555 238.165 ;
        RECT -2.885 235.17 -2.555 235.5 ;
        RECT -2.885 232.995 -2.555 233.325 ;
        RECT -2.885 231.415 -2.555 231.745 ;
        RECT -2.885 230.565 -2.555 230.895 ;
        RECT -2.885 228.255 -2.555 228.585 ;
        RECT -2.885 227.405 -2.555 227.735 ;
        RECT -2.885 225.095 -2.555 225.425 ;
        RECT -2.885 224.245 -2.555 224.575 ;
        RECT -2.885 221.935 -2.555 222.265 ;
        RECT -2.885 221.085 -2.555 221.415 ;
        RECT -2.885 218.775 -2.555 219.105 ;
        RECT -2.885 217.195 -2.555 217.525 ;
        RECT -2.885 216.345 -2.555 216.675 ;
        RECT -2.885 214.035 -2.555 214.365 ;
        RECT -2.885 213.185 -2.555 213.515 ;
        RECT -2.885 210.875 -2.555 211.205 ;
        RECT -2.885 210.025 -2.555 210.355 ;
        RECT -2.885 207.715 -2.555 208.045 ;
        RECT -2.885 206.865 -2.555 207.195 ;
        RECT -2.885 204.555 -2.555 204.885 ;
        RECT -2.885 202.975 -2.555 203.305 ;
        RECT -2.885 202.125 -2.555 202.455 ;
        RECT -2.885 199.815 -2.555 200.145 ;
        RECT -2.885 198.965 -2.555 199.295 ;
        RECT -2.885 196.655 -2.555 196.985 ;
        RECT -2.885 195.805 -2.555 196.135 ;
        RECT -2.885 193.495 -2.555 193.825 ;
        RECT -2.885 192.645 -2.555 192.975 ;
        RECT -2.885 190.335 -2.555 190.665 ;
        RECT -2.885 188.755 -2.555 189.085 ;
        RECT -2.885 187.905 -2.555 188.235 ;
        RECT -2.885 185.595 -2.555 185.925 ;
        RECT -2.885 184.745 -2.555 185.075 ;
        RECT -2.885 182.435 -2.555 182.765 ;
        RECT -2.885 181.585 -2.555 181.915 ;
        RECT -2.885 179.275 -2.555 179.605 ;
        RECT -2.885 178.425 -2.555 178.755 ;
        RECT -2.885 176.115 -2.555 176.445 ;
        RECT -2.885 174.535 -2.555 174.865 ;
        RECT -2.885 173.685 -2.555 174.015 ;
        RECT -2.885 171.375 -2.555 171.705 ;
        RECT -2.885 170.525 -2.555 170.855 ;
        RECT -2.885 168.215 -2.555 168.545 ;
        RECT -2.885 167.365 -2.555 167.695 ;
        RECT -2.885 165.055 -2.555 165.385 ;
        RECT -2.885 164.205 -2.555 164.535 ;
        RECT -2.885 161.895 -2.555 162.225 ;
        RECT -2.885 160.315 -2.555 160.645 ;
        RECT -2.885 159.465 -2.555 159.795 ;
        RECT -2.885 157.155 -2.555 157.485 ;
        RECT -2.885 156.305 -2.555 156.635 ;
        RECT -2.885 153.995 -2.555 154.325 ;
        RECT -2.885 153.145 -2.555 153.475 ;
        RECT -2.885 150.835 -2.555 151.165 ;
        RECT -2.885 149.985 -2.555 150.315 ;
        RECT -2.885 147.675 -2.555 148.005 ;
        RECT -2.885 146.095 -2.555 146.425 ;
        RECT -2.885 145.245 -2.555 145.575 ;
        RECT -2.885 142.935 -2.555 143.265 ;
        RECT -2.885 142.085 -2.555 142.415 ;
        RECT -2.885 139.775 -2.555 140.105 ;
        RECT -2.885 138.925 -2.555 139.255 ;
        RECT -2.885 136.615 -2.555 136.945 ;
        RECT -2.885 135.765 -2.555 136.095 ;
        RECT -2.885 133.455 -2.555 133.785 ;
        RECT -2.885 131.875 -2.555 132.205 ;
        RECT -2.885 131.025 -2.555 131.355 ;
        RECT -2.885 128.715 -2.555 129.045 ;
        RECT -2.885 127.865 -2.555 128.195 ;
        RECT -2.885 125.555 -2.555 125.885 ;
        RECT -2.885 124.705 -2.555 125.035 ;
        RECT -2.885 122.395 -2.555 122.725 ;
        RECT -2.885 121.545 -2.555 121.875 ;
        RECT -2.885 119.235 -2.555 119.565 ;
        RECT -2.885 117.655 -2.555 117.985 ;
        RECT -2.885 116.805 -2.555 117.135 ;
        RECT -2.885 114.495 -2.555 114.825 ;
        RECT -2.885 113.645 -2.555 113.975 ;
        RECT -2.885 111.335 -2.555 111.665 ;
        RECT -2.885 110.485 -2.555 110.815 ;
        RECT -2.885 108.175 -2.555 108.505 ;
        RECT -2.885 107.325 -2.555 107.655 ;
        RECT -2.885 105.015 -2.555 105.345 ;
        RECT -2.885 103.435 -2.555 103.765 ;
        RECT -2.885 102.585 -2.555 102.915 ;
        RECT -2.885 100.275 -2.555 100.605 ;
        RECT -2.885 99.425 -2.555 99.755 ;
        RECT -2.885 97.115 -2.555 97.445 ;
        RECT -2.885 96.265 -2.555 96.595 ;
        RECT -2.885 93.955 -2.555 94.285 ;
        RECT -2.885 93.105 -2.555 93.435 ;
        RECT -2.885 90.795 -2.555 91.125 ;
        RECT -2.885 89.215 -2.555 89.545 ;
        RECT -2.885 88.365 -2.555 88.695 ;
        RECT -2.885 86.055 -2.555 86.385 ;
        RECT -2.885 85.205 -2.555 85.535 ;
        RECT -2.885 82.895 -2.555 83.225 ;
        RECT -2.885 82.045 -2.555 82.375 ;
        RECT -2.885 79.735 -2.555 80.065 ;
        RECT -2.885 78.885 -2.555 79.215 ;
        RECT -2.885 76.575 -2.555 76.905 ;
        RECT -2.885 74.995 -2.555 75.325 ;
        RECT -2.885 74.145 -2.555 74.475 ;
        RECT -2.885 71.835 -2.555 72.165 ;
        RECT -2.885 70.985 -2.555 71.315 ;
        RECT -2.885 68.675 -2.555 69.005 ;
        RECT -2.885 67.825 -2.555 68.155 ;
        RECT -2.885 65.515 -2.555 65.845 ;
        RECT -2.885 64.665 -2.555 64.995 ;
        RECT -2.885 62.355 -2.555 62.685 ;
        RECT -2.885 60.775 -2.555 61.105 ;
        RECT -2.885 59.925 -2.555 60.255 ;
        RECT -2.885 57.615 -2.555 57.945 ;
        RECT -2.885 56.765 -2.555 57.095 ;
        RECT -2.885 54.455 -2.555 54.785 ;
        RECT -2.885 53.605 -2.555 53.935 ;
        RECT -2.885 51.295 -2.555 51.625 ;
        RECT -2.885 50.445 -2.555 50.775 ;
        RECT -2.885 48.135 -2.555 48.465 ;
        RECT -2.885 46.555 -2.555 46.885 ;
        RECT -2.885 45.705 -2.555 46.035 ;
        RECT -2.885 43.395 -2.555 43.725 ;
        RECT -2.885 42.545 -2.555 42.875 ;
        RECT -2.885 40.235 -2.555 40.565 ;
        RECT -2.885 39.385 -2.555 39.715 ;
        RECT -2.885 37.075 -2.555 37.405 ;
        RECT -2.885 36.225 -2.555 36.555 ;
        RECT -2.885 33.915 -2.555 34.245 ;
        RECT -2.885 32.335 -2.555 32.665 ;
        RECT -2.885 31.485 -2.555 31.815 ;
        RECT -2.885 29.175 -2.555 29.505 ;
        RECT -2.885 28.325 -2.555 28.655 ;
        RECT -2.885 26.015 -2.555 26.345 ;
        RECT -2.885 25.165 -2.555 25.495 ;
        RECT -2.885 22.855 -2.555 23.185 ;
        RECT -2.885 22.005 -2.555 22.335 ;
        RECT -2.885 19.695 -2.555 20.025 ;
        RECT -2.885 18.115 -2.555 18.445 ;
        RECT -2.885 17.265 -2.555 17.595 ;
        RECT -2.885 14.955 -2.555 15.285 ;
        RECT -2.885 14.105 -2.555 14.435 ;
        RECT -2.885 11.795 -2.555 12.125 ;
        RECT -2.885 10.945 -2.555 11.275 ;
        RECT -2.885 8.635 -2.555 8.965 ;
        RECT -2.885 7.785 -2.555 8.115 ;
        RECT -2.885 5.475 -2.555 5.805 ;
        RECT -2.885 3.895 -2.555 4.225 ;
        RECT -2.885 3.045 -2.555 3.375 ;
        RECT -2.885 0.87 -2.555 1.2 ;
        RECT -2.885 -1.525 -2.555 -1.195 ;
        RECT -2.885 -2.885 -2.555 -2.555 ;
        RECT -2.885 -4.245 -2.555 -3.915 ;
        RECT -2.885 -5.605 -2.555 -5.275 ;
        RECT -2.885 -6.965 -2.555 -6.635 ;
        RECT -2.885 -8.325 -2.555 -7.995 ;
        RECT -2.885 -9.685 -2.555 -9.355 ;
        RECT -2.885 -12.405 -2.555 -12.075 ;
        RECT -2.885 -13.765 -2.555 -13.435 ;
        RECT -2.885 -15.125 -2.555 -14.795 ;
        RECT -2.885 -16.485 -2.555 -16.155 ;
        RECT -2.885 -17.845 -2.555 -17.515 ;
        RECT -2.885 -19.205 -2.555 -18.875 ;
        RECT -2.88 -21.92 -2.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.885 -138.885 -2.555 -138.555 ;
        RECT -2.885 -140.245 -2.555 -139.915 ;
        RECT -2.885 -141.605 -2.555 -141.275 ;
        RECT -2.885 -142.965 -2.555 -142.635 ;
        RECT -2.885 -144.325 -2.555 -143.995 ;
        RECT -2.885 -145.685 -2.555 -145.355 ;
        RECT -2.885 -147.045 -2.555 -146.715 ;
        RECT -2.885 -148.405 -2.555 -148.075 ;
        RECT -2.885 -149.765 -2.555 -149.435 ;
        RECT -2.885 -151.125 -2.555 -150.795 ;
        RECT -2.885 -152.485 -2.555 -152.155 ;
        RECT -2.885 -153.845 -2.555 -153.515 ;
        RECT -2.885 -155.205 -2.555 -154.875 ;
        RECT -2.885 -156.565 -2.555 -156.235 ;
        RECT -2.885 -157.925 -2.555 -157.595 ;
        RECT -2.885 -160.645 -2.555 -160.315 ;
        RECT -2.885 -162.005 -2.555 -161.675 ;
        RECT -2.885 -163.365 -2.555 -163.035 ;
        RECT -2.885 -164.725 -2.555 -164.395 ;
        RECT -2.885 -166.085 -2.555 -165.755 ;
        RECT -2.885 -167.445 -2.555 -167.115 ;
        RECT -2.885 -168.805 -2.555 -168.475 ;
        RECT -2.885 -170.165 -2.555 -169.835 ;
        RECT -2.885 -171.525 -2.555 -171.195 ;
        RECT -2.885 -172.885 -2.555 -172.555 ;
        RECT -2.885 -174.245 -2.555 -173.915 ;
        RECT -2.885 -175.605 -2.555 -175.275 ;
        RECT -2.885 -176.965 -2.555 -176.635 ;
        RECT -2.885 -178.325 -2.555 -177.995 ;
        RECT -2.885 -179.685 -2.555 -179.355 ;
        RECT -2.885 -181.045 -2.555 -180.715 ;
        RECT -2.885 -182.405 -2.555 -182.075 ;
        RECT -2.885 -183.765 -2.555 -183.435 ;
        RECT -2.885 -185.125 -2.555 -184.795 ;
        RECT -2.885 -186.485 -2.555 -186.155 ;
        RECT -2.885 -187.845 -2.555 -187.515 ;
        RECT -2.885 -189.205 -2.555 -188.875 ;
        RECT -2.885 -190.565 -2.555 -190.235 ;
        RECT -2.885 -191.925 -2.555 -191.595 ;
        RECT -2.885 -193.285 -2.555 -192.955 ;
        RECT -2.885 -194.645 -2.555 -194.315 ;
        RECT -2.885 -196.005 -2.555 -195.675 ;
        RECT -2.885 -197.365 -2.555 -197.035 ;
        RECT -2.885 -198.725 -2.555 -198.395 ;
        RECT -2.885 -200.085 -2.555 -199.755 ;
        RECT -2.885 -201.445 -2.555 -201.115 ;
        RECT -2.885 -202.805 -2.555 -202.475 ;
        RECT -2.885 -204.165 -2.555 -203.835 ;
        RECT -2.885 -205.525 -2.555 -205.195 ;
        RECT -2.885 -206.885 -2.555 -206.555 ;
        RECT -2.885 -208.245 -2.555 -207.915 ;
        RECT -2.885 -209.605 -2.555 -209.275 ;
        RECT -2.885 -210.965 -2.555 -210.635 ;
        RECT -2.885 -212.325 -2.555 -211.995 ;
        RECT -2.885 -213.685 -2.555 -213.355 ;
        RECT -2.885 -215.045 -2.555 -214.715 ;
        RECT -2.885 -216.405 -2.555 -216.075 ;
        RECT -2.885 -217.765 -2.555 -217.435 ;
        RECT -2.885 -219.125 -2.555 -218.795 ;
        RECT -2.885 -220.485 -2.555 -220.155 ;
        RECT -2.885 -221.845 -2.555 -221.515 ;
        RECT -2.885 -223.205 -2.555 -222.875 ;
        RECT -2.885 -224.565 -2.555 -224.235 ;
        RECT -2.885 -225.925 -2.555 -225.595 ;
        RECT -2.885 -227.285 -2.555 -226.955 ;
        RECT -2.885 -228.645 -2.555 -228.315 ;
        RECT -2.885 -230.005 -2.555 -229.675 ;
        RECT -2.885 -231.365 -2.555 -231.035 ;
        RECT -2.885 -232.725 -2.555 -232.395 ;
        RECT -2.885 -234.085 -2.555 -233.755 ;
        RECT -2.885 -235.445 -2.555 -235.115 ;
        RECT -2.885 -236.805 -2.555 -236.475 ;
        RECT -2.885 -238.165 -2.555 -237.835 ;
        RECT -2.885 -243.81 -2.555 -242.68 ;
        RECT -2.88 -243.925 -2.56 -137.88 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 246.76 -1.195 247.89 ;
        RECT -1.525 241.915 -1.195 242.245 ;
        RECT -1.525 240.555 -1.195 240.885 ;
        RECT -1.525 239.195 -1.195 239.525 ;
        RECT -1.525 237.835 -1.195 238.165 ;
        RECT -1.525 235.17 -1.195 235.5 ;
        RECT -1.525 232.995 -1.195 233.325 ;
        RECT -1.525 231.415 -1.195 231.745 ;
        RECT -1.525 230.565 -1.195 230.895 ;
        RECT -1.525 228.255 -1.195 228.585 ;
        RECT -1.525 227.405 -1.195 227.735 ;
        RECT -1.525 225.095 -1.195 225.425 ;
        RECT -1.525 224.245 -1.195 224.575 ;
        RECT -1.525 221.935 -1.195 222.265 ;
        RECT -1.525 221.085 -1.195 221.415 ;
        RECT -1.525 218.775 -1.195 219.105 ;
        RECT -1.525 217.195 -1.195 217.525 ;
        RECT -1.525 216.345 -1.195 216.675 ;
        RECT -1.525 214.035 -1.195 214.365 ;
        RECT -1.525 213.185 -1.195 213.515 ;
        RECT -1.525 210.875 -1.195 211.205 ;
        RECT -1.525 210.025 -1.195 210.355 ;
        RECT -1.525 207.715 -1.195 208.045 ;
        RECT -1.525 206.865 -1.195 207.195 ;
        RECT -1.525 204.555 -1.195 204.885 ;
        RECT -1.525 202.975 -1.195 203.305 ;
        RECT -1.525 202.125 -1.195 202.455 ;
        RECT -1.525 199.815 -1.195 200.145 ;
        RECT -1.525 198.965 -1.195 199.295 ;
        RECT -1.525 196.655 -1.195 196.985 ;
        RECT -1.525 195.805 -1.195 196.135 ;
        RECT -1.525 193.495 -1.195 193.825 ;
        RECT -1.525 192.645 -1.195 192.975 ;
        RECT -1.525 190.335 -1.195 190.665 ;
        RECT -1.525 188.755 -1.195 189.085 ;
        RECT -1.525 187.905 -1.195 188.235 ;
        RECT -1.525 185.595 -1.195 185.925 ;
        RECT -1.525 184.745 -1.195 185.075 ;
        RECT -1.525 182.435 -1.195 182.765 ;
        RECT -1.525 181.585 -1.195 181.915 ;
        RECT -1.525 179.275 -1.195 179.605 ;
        RECT -1.525 178.425 -1.195 178.755 ;
        RECT -1.525 176.115 -1.195 176.445 ;
        RECT -1.525 174.535 -1.195 174.865 ;
        RECT -1.525 173.685 -1.195 174.015 ;
        RECT -1.525 171.375 -1.195 171.705 ;
        RECT -1.525 170.525 -1.195 170.855 ;
        RECT -1.525 168.215 -1.195 168.545 ;
        RECT -1.525 167.365 -1.195 167.695 ;
        RECT -1.525 165.055 -1.195 165.385 ;
        RECT -1.525 164.205 -1.195 164.535 ;
        RECT -1.525 161.895 -1.195 162.225 ;
        RECT -1.525 160.315 -1.195 160.645 ;
        RECT -1.525 159.465 -1.195 159.795 ;
        RECT -1.525 157.155 -1.195 157.485 ;
        RECT -1.525 156.305 -1.195 156.635 ;
        RECT -1.525 153.995 -1.195 154.325 ;
        RECT -1.525 153.145 -1.195 153.475 ;
        RECT -1.525 150.835 -1.195 151.165 ;
        RECT -1.525 149.985 -1.195 150.315 ;
        RECT -1.525 147.675 -1.195 148.005 ;
        RECT -1.525 146.095 -1.195 146.425 ;
        RECT -1.525 145.245 -1.195 145.575 ;
        RECT -1.525 142.935 -1.195 143.265 ;
        RECT -1.525 142.085 -1.195 142.415 ;
        RECT -1.525 139.775 -1.195 140.105 ;
        RECT -1.525 138.925 -1.195 139.255 ;
        RECT -1.525 136.615 -1.195 136.945 ;
        RECT -1.525 135.765 -1.195 136.095 ;
        RECT -1.525 133.455 -1.195 133.785 ;
        RECT -1.525 131.875 -1.195 132.205 ;
        RECT -1.525 131.025 -1.195 131.355 ;
        RECT -1.525 128.715 -1.195 129.045 ;
        RECT -1.525 127.865 -1.195 128.195 ;
        RECT -1.525 125.555 -1.195 125.885 ;
        RECT -1.525 124.705 -1.195 125.035 ;
        RECT -1.525 122.395 -1.195 122.725 ;
        RECT -1.525 121.545 -1.195 121.875 ;
        RECT -1.525 119.235 -1.195 119.565 ;
        RECT -1.525 117.655 -1.195 117.985 ;
        RECT -1.525 116.805 -1.195 117.135 ;
        RECT -1.525 114.495 -1.195 114.825 ;
        RECT -1.525 113.645 -1.195 113.975 ;
        RECT -1.525 111.335 -1.195 111.665 ;
        RECT -1.525 110.485 -1.195 110.815 ;
        RECT -1.525 108.175 -1.195 108.505 ;
        RECT -1.525 107.325 -1.195 107.655 ;
        RECT -1.525 105.015 -1.195 105.345 ;
        RECT -1.525 103.435 -1.195 103.765 ;
        RECT -1.525 102.585 -1.195 102.915 ;
        RECT -1.525 100.275 -1.195 100.605 ;
        RECT -1.525 99.425 -1.195 99.755 ;
        RECT -1.525 97.115 -1.195 97.445 ;
        RECT -1.525 96.265 -1.195 96.595 ;
        RECT -1.525 93.955 -1.195 94.285 ;
        RECT -1.525 93.105 -1.195 93.435 ;
        RECT -1.525 90.795 -1.195 91.125 ;
        RECT -1.525 89.215 -1.195 89.545 ;
        RECT -1.525 88.365 -1.195 88.695 ;
        RECT -1.525 86.055 -1.195 86.385 ;
        RECT -1.525 85.205 -1.195 85.535 ;
        RECT -1.525 82.895 -1.195 83.225 ;
        RECT -1.525 82.045 -1.195 82.375 ;
        RECT -1.525 79.735 -1.195 80.065 ;
        RECT -1.525 78.885 -1.195 79.215 ;
        RECT -1.525 76.575 -1.195 76.905 ;
        RECT -1.525 74.995 -1.195 75.325 ;
        RECT -1.525 74.145 -1.195 74.475 ;
        RECT -1.525 71.835 -1.195 72.165 ;
        RECT -1.525 70.985 -1.195 71.315 ;
        RECT -1.525 68.675 -1.195 69.005 ;
        RECT -1.525 67.825 -1.195 68.155 ;
        RECT -1.525 65.515 -1.195 65.845 ;
        RECT -1.525 64.665 -1.195 64.995 ;
        RECT -1.525 62.355 -1.195 62.685 ;
        RECT -1.525 60.775 -1.195 61.105 ;
        RECT -1.525 59.925 -1.195 60.255 ;
        RECT -1.525 57.615 -1.195 57.945 ;
        RECT -1.525 56.765 -1.195 57.095 ;
        RECT -1.525 54.455 -1.195 54.785 ;
        RECT -1.525 53.605 -1.195 53.935 ;
        RECT -1.525 51.295 -1.195 51.625 ;
        RECT -1.525 50.445 -1.195 50.775 ;
        RECT -1.525 48.135 -1.195 48.465 ;
        RECT -1.525 46.555 -1.195 46.885 ;
        RECT -1.525 45.705 -1.195 46.035 ;
        RECT -1.525 43.395 -1.195 43.725 ;
        RECT -1.525 42.545 -1.195 42.875 ;
        RECT -1.525 40.235 -1.195 40.565 ;
        RECT -1.525 39.385 -1.195 39.715 ;
        RECT -1.525 37.075 -1.195 37.405 ;
        RECT -1.525 36.225 -1.195 36.555 ;
        RECT -1.525 33.915 -1.195 34.245 ;
        RECT -1.525 32.335 -1.195 32.665 ;
        RECT -1.525 31.485 -1.195 31.815 ;
        RECT -1.525 29.175 -1.195 29.505 ;
        RECT -1.525 28.325 -1.195 28.655 ;
        RECT -1.525 26.015 -1.195 26.345 ;
        RECT -1.525 25.165 -1.195 25.495 ;
        RECT -1.525 22.855 -1.195 23.185 ;
        RECT -1.525 22.005 -1.195 22.335 ;
        RECT -1.525 19.695 -1.195 20.025 ;
        RECT -1.525 18.115 -1.195 18.445 ;
        RECT -1.525 17.265 -1.195 17.595 ;
        RECT -1.525 14.955 -1.195 15.285 ;
        RECT -1.525 14.105 -1.195 14.435 ;
        RECT -1.525 11.795 -1.195 12.125 ;
        RECT -1.525 10.945 -1.195 11.275 ;
        RECT -1.525 8.635 -1.195 8.965 ;
        RECT -1.525 7.785 -1.195 8.115 ;
        RECT -1.525 5.475 -1.195 5.805 ;
        RECT -1.525 3.895 -1.195 4.225 ;
        RECT -1.525 3.045 -1.195 3.375 ;
        RECT -1.525 0.87 -1.195 1.2 ;
        RECT -1.525 -1.525 -1.195 -1.195 ;
        RECT -1.525 -2.885 -1.195 -2.555 ;
        RECT -1.525 -4.245 -1.195 -3.915 ;
        RECT -1.525 -5.605 -1.195 -5.275 ;
        RECT -1.525 -6.965 -1.195 -6.635 ;
        RECT -1.525 -8.325 -1.195 -7.995 ;
        RECT -1.525 -9.685 -1.195 -9.355 ;
        RECT -1.525 -12.405 -1.195 -12.075 ;
        RECT -1.525 -13.765 -1.195 -13.435 ;
        RECT -1.525 -15.125 -1.195 -14.795 ;
        RECT -1.525 -16.485 -1.195 -16.155 ;
        RECT -1.525 -17.845 -1.195 -17.515 ;
        RECT -1.525 -19.205 -1.195 -18.875 ;
        RECT -1.52 -24.64 -1.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -200.085 -1.195 -199.755 ;
        RECT -1.525 -201.445 -1.195 -201.115 ;
        RECT -1.525 -202.805 -1.195 -202.475 ;
        RECT -1.525 -204.165 -1.195 -203.835 ;
        RECT -1.525 -205.525 -1.195 -205.195 ;
        RECT -1.525 -206.885 -1.195 -206.555 ;
        RECT -1.525 -208.245 -1.195 -207.915 ;
        RECT -1.525 -209.605 -1.195 -209.275 ;
        RECT -1.525 -210.965 -1.195 -210.635 ;
        RECT -1.525 -212.325 -1.195 -211.995 ;
        RECT -1.525 -213.685 -1.195 -213.355 ;
        RECT -1.525 -215.045 -1.195 -214.715 ;
        RECT -1.525 -216.405 -1.195 -216.075 ;
        RECT -1.525 -217.765 -1.195 -217.435 ;
        RECT -1.525 -219.125 -1.195 -218.795 ;
        RECT -1.525 -220.485 -1.195 -220.155 ;
        RECT -1.525 -221.845 -1.195 -221.515 ;
        RECT -1.525 -223.205 -1.195 -222.875 ;
        RECT -1.525 -224.565 -1.195 -224.235 ;
        RECT -1.525 -225.925 -1.195 -225.595 ;
        RECT -1.525 -227.285 -1.195 -226.955 ;
        RECT -1.525 -228.645 -1.195 -228.315 ;
        RECT -1.525 -230.005 -1.195 -229.675 ;
        RECT -1.525 -231.365 -1.195 -231.035 ;
        RECT -1.525 -232.725 -1.195 -232.395 ;
        RECT -1.525 -234.085 -1.195 -233.755 ;
        RECT -1.525 -235.445 -1.195 -235.115 ;
        RECT -1.525 -236.805 -1.195 -236.475 ;
        RECT -1.525 -238.165 -1.195 -237.835 ;
        RECT -1.525 -243.81 -1.195 -242.68 ;
        RECT -1.52 -243.925 -1.2 -135.16 ;
        RECT -1.525 -136.165 -1.195 -135.835 ;
        RECT -1.525 -137.525 -1.195 -137.195 ;
        RECT -1.525 -138.885 -1.195 -138.555 ;
        RECT -1.525 -140.245 -1.195 -139.915 ;
        RECT -1.525 -141.605 -1.195 -141.275 ;
        RECT -1.525 -142.965 -1.195 -142.635 ;
        RECT -1.525 -144.325 -1.195 -143.995 ;
        RECT -1.525 -145.685 -1.195 -145.355 ;
        RECT -1.525 -147.045 -1.195 -146.715 ;
        RECT -1.525 -148.405 -1.195 -148.075 ;
        RECT -1.525 -149.765 -1.195 -149.435 ;
        RECT -1.525 -151.125 -1.195 -150.795 ;
        RECT -1.525 -152.485 -1.195 -152.155 ;
        RECT -1.525 -153.845 -1.195 -153.515 ;
        RECT -1.525 -155.205 -1.195 -154.875 ;
        RECT -1.525 -156.565 -1.195 -156.235 ;
        RECT -1.525 -157.925 -1.195 -157.595 ;
        RECT -1.525 -160.645 -1.195 -160.315 ;
        RECT -1.525 -162.005 -1.195 -161.675 ;
        RECT -1.525 -163.365 -1.195 -163.035 ;
        RECT -1.525 -164.725 -1.195 -164.395 ;
        RECT -1.525 -166.085 -1.195 -165.755 ;
        RECT -1.525 -167.445 -1.195 -167.115 ;
        RECT -1.525 -168.805 -1.195 -168.475 ;
        RECT -1.525 -170.165 -1.195 -169.835 ;
        RECT -1.525 -171.525 -1.195 -171.195 ;
        RECT -1.525 -172.885 -1.195 -172.555 ;
        RECT -1.525 -174.245 -1.195 -173.915 ;
        RECT -1.525 -175.605 -1.195 -175.275 ;
        RECT -1.525 -176.965 -1.195 -176.635 ;
        RECT -1.525 -178.325 -1.195 -177.995 ;
        RECT -1.525 -179.685 -1.195 -179.355 ;
        RECT -1.525 -181.045 -1.195 -180.715 ;
        RECT -1.525 -182.405 -1.195 -182.075 ;
        RECT -1.525 -183.765 -1.195 -183.435 ;
        RECT -1.525 -185.125 -1.195 -184.795 ;
        RECT -1.525 -186.485 -1.195 -186.155 ;
        RECT -1.525 -187.845 -1.195 -187.515 ;
        RECT -1.525 -189.205 -1.195 -188.875 ;
        RECT -1.525 -190.565 -1.195 -190.235 ;
        RECT -1.525 -191.925 -1.195 -191.595 ;
        RECT -1.525 -193.285 -1.195 -192.955 ;
        RECT -1.525 -194.645 -1.195 -194.315 ;
        RECT -1.525 -196.005 -1.195 -195.675 ;
        RECT -1.525 -197.365 -1.195 -197.035 ;
        RECT -1.525 -198.725 -1.195 -198.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 246.76 -10.715 247.89 ;
        RECT -11.045 241.915 -10.715 242.245 ;
        RECT -11.045 240.555 -10.715 240.885 ;
        RECT -11.045 239.195 -10.715 239.525 ;
        RECT -11.045 237.835 -10.715 238.165 ;
        RECT -11.045 236.475 -10.715 236.805 ;
        RECT -11.045 235.115 -10.715 235.445 ;
        RECT -11.045 233.755 -10.715 234.085 ;
        RECT -11.045 232.395 -10.715 232.725 ;
        RECT -11.045 231.035 -10.715 231.365 ;
        RECT -11.045 221.515 -10.715 221.845 ;
        RECT -11.045 217.435 -10.715 217.765 ;
        RECT -11.045 213.355 -10.715 213.685 ;
        RECT -11.045 210.635 -10.715 210.965 ;
        RECT -11.045 203.835 -10.715 204.165 ;
        RECT -11.045 202.475 -10.715 202.805 ;
        RECT -11.045 199.755 -10.715 200.085 ;
        RECT -11.045 192.955 -10.715 193.285 ;
        RECT -11.045 190.235 -10.715 190.565 ;
        RECT -11.045 188.875 -10.715 189.205 ;
        RECT -11.045 184.795 -10.715 185.125 ;
        RECT -11.045 182.075 -10.715 182.405 ;
        RECT -11.045 175.275 -10.715 175.605 ;
        RECT -11.045 173.915 -10.715 174.245 ;
        RECT -11.045 171.195 -10.715 171.525 ;
        RECT -11.045 164.395 -10.715 164.725 ;
        RECT -11.045 161.675 -10.715 162.005 ;
        RECT -11.045 160.315 -10.715 160.645 ;
        RECT -11.045 153.515 -10.715 153.845 ;
        RECT -11.045 150.795 -10.715 151.125 ;
        RECT -11.045 146.715 -10.715 147.045 ;
        RECT -11.045 145.355 -10.715 145.685 ;
        RECT -11.045 142.635 -10.715 142.965 ;
        RECT -11.045 135.835 -10.715 136.165 ;
        RECT -11.045 133.115 -10.715 133.445 ;
        RECT -11.045 131.755 -10.715 132.085 ;
        RECT -11.045 124.955 -10.715 125.285 ;
        RECT -11.045 122.235 -10.715 122.565 ;
        RECT -11.045 118.155 -10.715 118.485 ;
        RECT -11.045 114.075 -10.715 114.405 ;
        RECT -11.045 104.555 -10.715 104.885 ;
        RECT -11.045 103.195 -10.715 103.525 ;
        RECT -11.045 96.395 -10.715 96.725 ;
        RECT -11.045 93.675 -10.715 94.005 ;
        RECT -11.045 89.595 -10.715 89.925 ;
        RECT -11.045 85.515 -10.715 85.845 ;
        RECT -11.045 82.795 -10.715 83.125 ;
        RECT -11.045 75.995 -10.715 76.325 ;
        RECT -11.045 74.635 -10.715 74.965 ;
        RECT -11.045 65.115 -10.715 65.445 ;
        RECT -11.045 61.035 -10.715 61.365 ;
        RECT -11.045 56.955 -10.715 57.285 ;
        RECT -11.045 54.235 -10.715 54.565 ;
        RECT -11.045 47.435 -10.715 47.765 ;
        RECT -11.045 46.075 -10.715 46.405 ;
        RECT -11.045 43.355 -10.715 43.685 ;
        RECT -11.045 36.555 -10.715 36.885 ;
        RECT -11.045 33.835 -10.715 34.165 ;
        RECT -11.045 32.475 -10.715 32.805 ;
        RECT -11.045 28.395 -10.715 28.725 ;
        RECT -11.045 25.675 -10.715 26.005 ;
        RECT -11.045 18.875 -10.715 19.205 ;
        RECT -11.045 17.515 -10.715 17.845 ;
        RECT -11.045 14.795 -10.715 15.125 ;
        RECT -11.045 7.995 -10.715 8.325 ;
        RECT -11.045 5.275 -10.715 5.605 ;
        RECT -11.045 3.915 -10.715 4.245 ;
        RECT -11.045 2.555 -10.715 2.885 ;
        RECT -11.045 1.195 -10.715 1.525 ;
        RECT -11.045 -0.165 -10.715 0.165 ;
        RECT -11.045 -1.525 -10.715 -1.195 ;
        RECT -11.045 -2.885 -10.715 -2.555 ;
        RECT -11.045 -4.245 -10.715 -3.915 ;
        RECT -11.045 -5.605 -10.715 -5.275 ;
        RECT -11.045 -6.965 -10.715 -6.635 ;
        RECT -11.045 -8.325 -10.715 -7.995 ;
        RECT -11.045 -9.48 -10.715 -9.15 ;
        RECT -11.045 -12.405 -10.715 -12.075 ;
        RECT -11.045 -15.125 -10.715 -14.795 ;
        RECT -11.045 -16.67 -10.715 -16.34 ;
        RECT -11.045 -17.845 -10.715 -17.515 ;
        RECT -11.045 -24.645 -10.715 -24.315 ;
        RECT -11.045 -26.005 -10.715 -25.675 ;
        RECT -11.045 -27.365 -10.715 -27.035 ;
        RECT -11.045 -28.725 -10.715 -28.395 ;
        RECT -11.045 -30.66 -10.715 -30.33 ;
        RECT -11.045 -31.445 -10.715 -31.115 ;
        RECT -11.045 -32.805 -10.715 -32.475 ;
        RECT -11.045 -34.165 -10.715 -33.835 ;
        RECT -11.045 -36.885 -10.715 -36.555 ;
        RECT -11.045 -37.85 -10.715 -37.52 ;
        RECT -11.045 -40.965 -10.715 -40.635 ;
        RECT -11.045 -46.405 -10.715 -46.075 ;
        RECT -11.045 -47.765 -10.715 -47.435 ;
        RECT -11.045 -49.125 -10.715 -48.795 ;
        RECT -11.045 -50.485 -10.715 -50.155 ;
        RECT -11.045 -51.845 -10.715 -51.515 ;
        RECT -11.045 -53.205 -10.715 -52.875 ;
        RECT -11.045 -54.565 -10.715 -54.235 ;
        RECT -11.045 -55.925 -10.715 -55.595 ;
        RECT -11.045 -57.285 -10.715 -56.955 ;
        RECT -11.045 -58.645 -10.715 -58.315 ;
        RECT -11.045 -60.005 -10.715 -59.675 ;
        RECT -11.045 -61.365 -10.715 -61.035 ;
        RECT -11.045 -68.165 -10.715 -67.835 ;
        RECT -11.045 -69.525 -10.715 -69.195 ;
        RECT -11.045 -70.79 -10.715 -70.46 ;
        RECT -11.045 -72.245 -10.715 -71.915 ;
        RECT -11.045 -73.605 -10.715 -73.275 ;
        RECT -11.045 -74.965 -10.715 -74.635 ;
        RECT -11.045 -76.325 -10.715 -75.995 ;
        RECT -11.045 -77.685 -10.715 -77.355 ;
        RECT -11.045 -79.045 -10.715 -78.715 ;
        RECT -11.045 -81.765 -10.715 -81.435 ;
        RECT -11.045 -83.125 -10.715 -82.795 ;
        RECT -11.045 -84.485 -10.715 -84.155 ;
        RECT -11.045 -85.845 -10.715 -85.515 ;
        RECT -11.045 -87.205 -10.715 -86.875 ;
        RECT -11.045 -88.565 -10.715 -88.235 ;
        RECT -11.045 -89.33 -10.715 -89 ;
        RECT -11.045 -91.285 -10.715 -90.955 ;
        RECT -11.045 -92.645 -10.715 -92.315 ;
        RECT -11.045 -94.005 -10.715 -93.675 ;
        RECT -11.045 -95.365 -10.715 -95.035 ;
        RECT -11.045 -96.725 -10.715 -96.395 ;
        RECT -11.045 -98.085 -10.715 -97.755 ;
        RECT -11.045 -100.805 -10.715 -100.475 ;
        RECT -11.045 -102.165 -10.715 -101.835 ;
        RECT -11.045 -103.525 -10.715 -103.195 ;
        RECT -11.045 -106.245 -10.715 -105.915 ;
        RECT -11.045 -107.605 -10.715 -107.275 ;
        RECT -11.045 -108.965 -10.715 -108.635 ;
        RECT -11.045 -110.325 -10.715 -109.995 ;
        RECT -11.045 -111.685 -10.715 -111.355 ;
        RECT -11.045 -113.045 -10.715 -112.715 ;
        RECT -11.045 -114.97 -10.715 -114.64 ;
        RECT -11.045 -115.765 -10.715 -115.435 ;
        RECT -11.045 -117.125 -10.715 -116.795 ;
        RECT -11.045 -118.485 -10.715 -118.155 ;
        RECT -11.045 -119.845 -10.715 -119.515 ;
        RECT -11.045 -121.205 -10.715 -120.875 ;
        RECT -11.045 -122.565 -10.715 -122.235 ;
        RECT -11.045 -125.285 -10.715 -124.955 ;
        RECT -11.045 -126.645 -10.715 -126.315 ;
        RECT -11.045 -128.005 -10.715 -127.675 ;
        RECT -11.045 -129.365 -10.715 -129.035 ;
        RECT -11.045 -130.725 -10.715 -130.395 ;
        RECT -11.045 -132.085 -10.715 -131.755 ;
        RECT -11.045 -133.51 -10.715 -133.18 ;
        RECT -11.045 -140.245 -10.715 -139.915 ;
        RECT -11.045 -141.605 -10.715 -141.275 ;
        RECT -11.045 -144.325 -10.715 -143.995 ;
        RECT -11.045 -145.685 -10.715 -145.355 ;
        RECT -11.045 -147.045 -10.715 -146.715 ;
        RECT -11.045 -152.485 -10.715 -152.155 ;
        RECT -11.045 -153.845 -10.715 -153.515 ;
        RECT -11.045 -155.205 -10.715 -154.875 ;
        RECT -11.045 -156.565 -10.715 -156.235 ;
        RECT -11.045 -157.925 -10.715 -157.595 ;
        RECT -11.045 -160.645 -10.715 -160.315 ;
        RECT -11.045 -162.005 -10.715 -161.675 ;
        RECT -11.045 -164.725 -10.715 -164.395 ;
        RECT -11.045 -167.445 -10.715 -167.115 ;
        RECT -11.045 -168.805 -10.715 -168.475 ;
        RECT -11.045 -171.525 -10.715 -171.195 ;
        RECT -11.045 -172.885 -10.715 -172.555 ;
        RECT -11.045 -174.245 -10.715 -173.915 ;
        RECT -11.045 -175.605 -10.715 -175.275 ;
        RECT -11.045 -176.965 -10.715 -176.635 ;
        RECT -11.045 -178.325 -10.715 -177.995 ;
        RECT -11.045 -179.685 -10.715 -179.355 ;
        RECT -11.045 -181.045 -10.715 -180.715 ;
        RECT -11.045 -182.405 -10.715 -182.075 ;
        RECT -11.045 -183.765 -10.715 -183.435 ;
        RECT -11.045 -185.125 -10.715 -184.795 ;
        RECT -11.045 -186.485 -10.715 -186.155 ;
        RECT -11.045 -187.845 -10.715 -187.515 ;
        RECT -11.045 -189.205 -10.715 -188.875 ;
        RECT -11.045 -190.565 -10.715 -190.235 ;
        RECT -11.045 -191.925 -10.715 -191.595 ;
        RECT -11.045 -193.285 -10.715 -192.955 ;
        RECT -11.045 -194.645 -10.715 -194.315 ;
        RECT -11.045 -196.005 -10.715 -195.675 ;
        RECT -11.045 -197.365 -10.715 -197.035 ;
        RECT -11.045 -198.725 -10.715 -198.395 ;
        RECT -11.045 -201.445 -10.715 -201.115 ;
        RECT -11.045 -204.165 -10.715 -203.835 ;
        RECT -11.045 -205.525 -10.715 -205.195 ;
        RECT -11.045 -206.885 -10.715 -206.555 ;
        RECT -11.045 -208.245 -10.715 -207.915 ;
        RECT -11.045 -209.605 -10.715 -209.275 ;
        RECT -11.045 -210.965 -10.715 -210.635 ;
        RECT -11.045 -212.325 -10.715 -211.995 ;
        RECT -11.045 -213.685 -10.715 -213.355 ;
        RECT -11.045 -215.045 -10.715 -214.715 ;
        RECT -11.045 -216.405 -10.715 -216.075 ;
        RECT -11.045 -217.765 -10.715 -217.435 ;
        RECT -11.045 -219.125 -10.715 -218.795 ;
        RECT -11.045 -220.485 -10.715 -220.155 ;
        RECT -11.045 -221.845 -10.715 -221.515 ;
        RECT -11.045 -223.205 -10.715 -222.875 ;
        RECT -11.04 -224.56 -10.72 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 -234.085 -10.715 -233.755 ;
        RECT -11.045 -235.445 -10.715 -235.115 ;
        RECT -11.045 -236.805 -10.715 -236.475 ;
        RECT -11.045 -238.165 -10.715 -237.835 ;
        RECT -11.045 -243.81 -10.715 -242.68 ;
        RECT -11.04 -243.925 -10.72 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.685 246.76 -9.355 247.89 ;
        RECT -9.685 241.915 -9.355 242.245 ;
        RECT -9.685 240.555 -9.355 240.885 ;
        RECT -9.685 239.195 -9.355 239.525 ;
        RECT -9.685 237.835 -9.355 238.165 ;
        RECT -9.685 236.475 -9.355 236.805 ;
        RECT -9.685 235.115 -9.355 235.445 ;
        RECT -9.685 233.755 -9.355 234.085 ;
        RECT -9.685 232.395 -9.355 232.725 ;
        RECT -9.685 231.035 -9.355 231.365 ;
        RECT -9.685 221.515 -9.355 221.845 ;
        RECT -9.685 217.435 -9.355 217.765 ;
        RECT -9.685 213.355 -9.355 213.685 ;
        RECT -9.685 210.635 -9.355 210.965 ;
        RECT -9.685 203.835 -9.355 204.165 ;
        RECT -9.685 202.475 -9.355 202.805 ;
        RECT -9.685 199.755 -9.355 200.085 ;
        RECT -9.685 192.955 -9.355 193.285 ;
        RECT -9.685 190.235 -9.355 190.565 ;
        RECT -9.685 188.875 -9.355 189.205 ;
        RECT -9.685 184.795 -9.355 185.125 ;
        RECT -9.685 182.075 -9.355 182.405 ;
        RECT -9.685 175.275 -9.355 175.605 ;
        RECT -9.685 173.915 -9.355 174.245 ;
        RECT -9.685 171.195 -9.355 171.525 ;
        RECT -9.685 164.395 -9.355 164.725 ;
        RECT -9.685 161.675 -9.355 162.005 ;
        RECT -9.685 160.315 -9.355 160.645 ;
        RECT -9.685 153.515 -9.355 153.845 ;
        RECT -9.685 150.795 -9.355 151.125 ;
        RECT -9.685 146.715 -9.355 147.045 ;
        RECT -9.685 145.355 -9.355 145.685 ;
        RECT -9.685 142.635 -9.355 142.965 ;
        RECT -9.685 135.835 -9.355 136.165 ;
        RECT -9.685 133.115 -9.355 133.445 ;
        RECT -9.685 131.755 -9.355 132.085 ;
        RECT -9.685 124.955 -9.355 125.285 ;
        RECT -9.685 122.235 -9.355 122.565 ;
        RECT -9.685 118.155 -9.355 118.485 ;
        RECT -9.685 114.075 -9.355 114.405 ;
        RECT -9.685 104.555 -9.355 104.885 ;
        RECT -9.685 103.195 -9.355 103.525 ;
        RECT -9.685 96.395 -9.355 96.725 ;
        RECT -9.685 93.675 -9.355 94.005 ;
        RECT -9.685 89.595 -9.355 89.925 ;
        RECT -9.685 85.515 -9.355 85.845 ;
        RECT -9.685 82.795 -9.355 83.125 ;
        RECT -9.685 75.995 -9.355 76.325 ;
        RECT -9.685 74.635 -9.355 74.965 ;
        RECT -9.685 65.115 -9.355 65.445 ;
        RECT -9.685 61.035 -9.355 61.365 ;
        RECT -9.685 56.955 -9.355 57.285 ;
        RECT -9.685 54.235 -9.355 54.565 ;
        RECT -9.685 47.435 -9.355 47.765 ;
        RECT -9.685 46.075 -9.355 46.405 ;
        RECT -9.685 43.355 -9.355 43.685 ;
        RECT -9.685 36.555 -9.355 36.885 ;
        RECT -9.685 33.835 -9.355 34.165 ;
        RECT -9.685 32.475 -9.355 32.805 ;
        RECT -9.685 28.395 -9.355 28.725 ;
        RECT -9.685 25.675 -9.355 26.005 ;
        RECT -9.685 18.875 -9.355 19.205 ;
        RECT -9.685 17.515 -9.355 17.845 ;
        RECT -9.685 14.795 -9.355 15.125 ;
        RECT -9.685 7.995 -9.355 8.325 ;
        RECT -9.685 5.275 -9.355 5.605 ;
        RECT -9.685 3.915 -9.355 4.245 ;
        RECT -9.685 2.555 -9.355 2.885 ;
        RECT -9.685 1.195 -9.355 1.525 ;
        RECT -9.685 -0.165 -9.355 0.165 ;
        RECT -9.685 -1.525 -9.355 -1.195 ;
        RECT -9.685 -2.885 -9.355 -2.555 ;
        RECT -9.685 -4.245 -9.355 -3.915 ;
        RECT -9.685 -5.605 -9.355 -5.275 ;
        RECT -9.685 -6.965 -9.355 -6.635 ;
        RECT -9.685 -8.325 -9.355 -7.995 ;
        RECT -9.685 -9.685 -9.355 -9.355 ;
        RECT -9.685 -12.405 -9.355 -12.075 ;
        RECT -9.685 -13.765 -9.355 -13.435 ;
        RECT -9.685 -15.125 -9.355 -14.795 ;
        RECT -9.685 -16.485 -9.355 -16.155 ;
        RECT -9.685 -17.845 -9.355 -17.515 ;
        RECT -9.685 -19.205 -9.355 -18.875 ;
        RECT -9.685 -20.565 -9.355 -20.235 ;
        RECT -9.685 -21.925 -9.355 -21.595 ;
        RECT -9.685 -23.285 -9.355 -22.955 ;
        RECT -9.685 -24.645 -9.355 -24.315 ;
        RECT -9.685 -26.005 -9.355 -25.675 ;
        RECT -9.685 -27.365 -9.355 -27.035 ;
        RECT -9.685 -28.725 -9.355 -28.395 ;
        RECT -9.685 -30.085 -9.355 -29.755 ;
        RECT -9.685 -31.445 -9.355 -31.115 ;
        RECT -9.685 -32.805 -9.355 -32.475 ;
        RECT -9.685 -34.165 -9.355 -33.835 ;
        RECT -9.685 -35.525 -9.355 -35.195 ;
        RECT -9.685 -36.885 -9.355 -36.555 ;
        RECT -9.685 -38.245 -9.355 -37.915 ;
        RECT -9.685 -39.605 -9.355 -39.275 ;
        RECT -9.685 -40.965 -9.355 -40.635 ;
        RECT -9.685 -42.325 -9.355 -41.995 ;
        RECT -9.685 -43.685 -9.355 -43.355 ;
        RECT -9.685 -45.045 -9.355 -44.715 ;
        RECT -9.685 -46.405 -9.355 -46.075 ;
        RECT -9.685 -47.765 -9.355 -47.435 ;
        RECT -9.685 -49.125 -9.355 -48.795 ;
        RECT -9.685 -50.485 -9.355 -50.155 ;
        RECT -9.685 -51.845 -9.355 -51.515 ;
        RECT -9.685 -53.205 -9.355 -52.875 ;
        RECT -9.685 -54.565 -9.355 -54.235 ;
        RECT -9.685 -55.925 -9.355 -55.595 ;
        RECT -9.685 -57.285 -9.355 -56.955 ;
        RECT -9.685 -58.645 -9.355 -58.315 ;
        RECT -9.685 -60.005 -9.355 -59.675 ;
        RECT -9.685 -61.365 -9.355 -61.035 ;
        RECT -9.685 -68.165 -9.355 -67.835 ;
        RECT -9.685 -69.525 -9.355 -69.195 ;
        RECT -9.685 -70.885 -9.355 -70.555 ;
        RECT -9.685 -72.245 -9.355 -71.915 ;
        RECT -9.685 -73.605 -9.355 -73.275 ;
        RECT -9.685 -74.965 -9.355 -74.635 ;
        RECT -9.685 -76.325 -9.355 -75.995 ;
        RECT -9.685 -77.685 -9.355 -77.355 ;
        RECT -9.685 -79.045 -9.355 -78.715 ;
        RECT -9.685 -80.405 -9.355 -80.075 ;
        RECT -9.685 -81.765 -9.355 -81.435 ;
        RECT -9.685 -83.125 -9.355 -82.795 ;
        RECT -9.685 -84.485 -9.355 -84.155 ;
        RECT -9.685 -85.845 -9.355 -85.515 ;
        RECT -9.685 -87.205 -9.355 -86.875 ;
        RECT -9.685 -88.565 -9.355 -88.235 ;
        RECT -9.685 -89.925 -9.355 -89.595 ;
        RECT -9.685 -91.285 -9.355 -90.955 ;
        RECT -9.685 -92.645 -9.355 -92.315 ;
        RECT -9.685 -94.005 -9.355 -93.675 ;
        RECT -9.685 -95.365 -9.355 -95.035 ;
        RECT -9.685 -96.725 -9.355 -96.395 ;
        RECT -9.685 -98.085 -9.355 -97.755 ;
        RECT -9.685 -99.445 -9.355 -99.115 ;
        RECT -9.685 -100.805 -9.355 -100.475 ;
        RECT -9.685 -102.165 -9.355 -101.835 ;
        RECT -9.685 -103.525 -9.355 -103.195 ;
        RECT -9.685 -104.885 -9.355 -104.555 ;
        RECT -9.685 -106.245 -9.355 -105.915 ;
        RECT -9.685 -107.605 -9.355 -107.275 ;
        RECT -9.685 -108.965 -9.355 -108.635 ;
        RECT -9.685 -110.325 -9.355 -109.995 ;
        RECT -9.685 -111.685 -9.355 -111.355 ;
        RECT -9.685 -113.045 -9.355 -112.715 ;
        RECT -9.685 -114.405 -9.355 -114.075 ;
        RECT -9.685 -115.765 -9.355 -115.435 ;
        RECT -9.685 -117.125 -9.355 -116.795 ;
        RECT -9.685 -118.485 -9.355 -118.155 ;
        RECT -9.685 -119.845 -9.355 -119.515 ;
        RECT -9.685 -121.205 -9.355 -120.875 ;
        RECT -9.685 -122.565 -9.355 -122.235 ;
        RECT -9.685 -123.925 -9.355 -123.595 ;
        RECT -9.685 -125.285 -9.355 -124.955 ;
        RECT -9.685 -126.645 -9.355 -126.315 ;
        RECT -9.685 -128.005 -9.355 -127.675 ;
        RECT -9.685 -129.365 -9.355 -129.035 ;
        RECT -9.685 -130.725 -9.355 -130.395 ;
        RECT -9.685 -132.085 -9.355 -131.755 ;
        RECT -9.685 -133.445 -9.355 -133.115 ;
        RECT -9.685 -140.245 -9.355 -139.915 ;
        RECT -9.685 -141.605 -9.355 -141.275 ;
        RECT -9.685 -142.965 -9.355 -142.635 ;
        RECT -9.685 -144.325 -9.355 -143.995 ;
        RECT -9.685 -145.685 -9.355 -145.355 ;
        RECT -9.685 -147.045 -9.355 -146.715 ;
        RECT -9.685 -148.405 -9.355 -148.075 ;
        RECT -9.685 -149.765 -9.355 -149.435 ;
        RECT -9.685 -151.125 -9.355 -150.795 ;
        RECT -9.685 -152.485 -9.355 -152.155 ;
        RECT -9.685 -153.845 -9.355 -153.515 ;
        RECT -9.685 -155.205 -9.355 -154.875 ;
        RECT -9.685 -156.565 -9.355 -156.235 ;
        RECT -9.685 -157.925 -9.355 -157.595 ;
        RECT -9.685 -160.645 -9.355 -160.315 ;
        RECT -9.685 -162.005 -9.355 -161.675 ;
        RECT -9.685 -163.365 -9.355 -163.035 ;
        RECT -9.685 -164.725 -9.355 -164.395 ;
        RECT -9.685 -166.085 -9.355 -165.755 ;
        RECT -9.685 -167.445 -9.355 -167.115 ;
        RECT -9.685 -168.805 -9.355 -168.475 ;
        RECT -9.685 -170.165 -9.355 -169.835 ;
        RECT -9.685 -171.525 -9.355 -171.195 ;
        RECT -9.685 -172.885 -9.355 -172.555 ;
        RECT -9.685 -174.245 -9.355 -173.915 ;
        RECT -9.685 -175.605 -9.355 -175.275 ;
        RECT -9.685 -176.965 -9.355 -176.635 ;
        RECT -9.685 -178.325 -9.355 -177.995 ;
        RECT -9.685 -179.685 -9.355 -179.355 ;
        RECT -9.685 -181.045 -9.355 -180.715 ;
        RECT -9.685 -182.405 -9.355 -182.075 ;
        RECT -9.685 -183.765 -9.355 -183.435 ;
        RECT -9.685 -185.125 -9.355 -184.795 ;
        RECT -9.685 -186.485 -9.355 -186.155 ;
        RECT -9.685 -187.845 -9.355 -187.515 ;
        RECT -9.685 -189.205 -9.355 -188.875 ;
        RECT -9.685 -190.565 -9.355 -190.235 ;
        RECT -9.685 -191.925 -9.355 -191.595 ;
        RECT -9.685 -193.285 -9.355 -192.955 ;
        RECT -9.685 -194.645 -9.355 -194.315 ;
        RECT -9.685 -196.005 -9.355 -195.675 ;
        RECT -9.685 -197.365 -9.355 -197.035 ;
        RECT -9.685 -198.725 -9.355 -198.395 ;
        RECT -9.685 -200.085 -9.355 -199.755 ;
        RECT -9.685 -201.445 -9.355 -201.115 ;
        RECT -9.685 -202.805 -9.355 -202.475 ;
        RECT -9.685 -204.165 -9.355 -203.835 ;
        RECT -9.685 -205.525 -9.355 -205.195 ;
        RECT -9.685 -206.885 -9.355 -206.555 ;
        RECT -9.685 -208.245 -9.355 -207.915 ;
        RECT -9.685 -209.605 -9.355 -209.275 ;
        RECT -9.685 -210.965 -9.355 -210.635 ;
        RECT -9.685 -212.325 -9.355 -211.995 ;
        RECT -9.685 -213.685 -9.355 -213.355 ;
        RECT -9.685 -215.045 -9.355 -214.715 ;
        RECT -9.685 -216.405 -9.355 -216.075 ;
        RECT -9.685 -217.765 -9.355 -217.435 ;
        RECT -9.685 -219.125 -9.355 -218.795 ;
        RECT -9.685 -220.485 -9.355 -220.155 ;
        RECT -9.685 -221.845 -9.355 -221.515 ;
        RECT -9.685 -223.205 -9.355 -222.875 ;
        RECT -9.68 -223.88 -9.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 246.76 -7.995 247.89 ;
        RECT -8.325 241.915 -7.995 242.245 ;
        RECT -8.325 240.555 -7.995 240.885 ;
        RECT -8.325 239.195 -7.995 239.525 ;
        RECT -8.325 237.835 -7.995 238.165 ;
        RECT -8.325 236.475 -7.995 236.805 ;
        RECT -8.325 235.115 -7.995 235.445 ;
        RECT -8.325 233.755 -7.995 234.085 ;
        RECT -8.325 232.395 -7.995 232.725 ;
        RECT -8.325 231.035 -7.995 231.365 ;
        RECT -8.325 221.515 -7.995 221.845 ;
        RECT -8.325 217.435 -7.995 217.765 ;
        RECT -8.325 213.355 -7.995 213.685 ;
        RECT -8.325 210.635 -7.995 210.965 ;
        RECT -8.325 203.835 -7.995 204.165 ;
        RECT -8.325 202.475 -7.995 202.805 ;
        RECT -8.325 199.755 -7.995 200.085 ;
        RECT -8.325 192.955 -7.995 193.285 ;
        RECT -8.325 190.235 -7.995 190.565 ;
        RECT -8.325 188.875 -7.995 189.205 ;
        RECT -8.325 184.795 -7.995 185.125 ;
        RECT -8.325 182.075 -7.995 182.405 ;
        RECT -8.325 175.275 -7.995 175.605 ;
        RECT -8.325 173.915 -7.995 174.245 ;
        RECT -8.325 171.195 -7.995 171.525 ;
        RECT -8.325 164.395 -7.995 164.725 ;
        RECT -8.325 161.675 -7.995 162.005 ;
        RECT -8.325 160.315 -7.995 160.645 ;
        RECT -8.325 153.515 -7.995 153.845 ;
        RECT -8.325 150.795 -7.995 151.125 ;
        RECT -8.325 146.715 -7.995 147.045 ;
        RECT -8.325 145.355 -7.995 145.685 ;
        RECT -8.325 142.635 -7.995 142.965 ;
        RECT -8.325 135.835 -7.995 136.165 ;
        RECT -8.325 133.115 -7.995 133.445 ;
        RECT -8.325 131.755 -7.995 132.085 ;
        RECT -8.325 124.955 -7.995 125.285 ;
        RECT -8.325 122.235 -7.995 122.565 ;
        RECT -8.325 118.155 -7.995 118.485 ;
        RECT -8.325 114.075 -7.995 114.405 ;
        RECT -8.325 104.555 -7.995 104.885 ;
        RECT -8.325 103.195 -7.995 103.525 ;
        RECT -8.325 96.395 -7.995 96.725 ;
        RECT -8.325 93.675 -7.995 94.005 ;
        RECT -8.325 89.595 -7.995 89.925 ;
        RECT -8.325 85.515 -7.995 85.845 ;
        RECT -8.325 82.795 -7.995 83.125 ;
        RECT -8.325 75.995 -7.995 76.325 ;
        RECT -8.325 74.635 -7.995 74.965 ;
        RECT -8.325 65.115 -7.995 65.445 ;
        RECT -8.325 61.035 -7.995 61.365 ;
        RECT -8.325 56.955 -7.995 57.285 ;
        RECT -8.325 54.235 -7.995 54.565 ;
        RECT -8.325 47.435 -7.995 47.765 ;
        RECT -8.325 46.075 -7.995 46.405 ;
        RECT -8.325 43.355 -7.995 43.685 ;
        RECT -8.325 36.555 -7.995 36.885 ;
        RECT -8.325 33.835 -7.995 34.165 ;
        RECT -8.325 32.475 -7.995 32.805 ;
        RECT -8.325 28.395 -7.995 28.725 ;
        RECT -8.325 25.675 -7.995 26.005 ;
        RECT -8.325 18.875 -7.995 19.205 ;
        RECT -8.325 17.515 -7.995 17.845 ;
        RECT -8.325 14.795 -7.995 15.125 ;
        RECT -8.325 7.995 -7.995 8.325 ;
        RECT -8.325 5.275 -7.995 5.605 ;
        RECT -8.325 3.915 -7.995 4.245 ;
        RECT -8.325 2.555 -7.995 2.885 ;
        RECT -8.325 1.195 -7.995 1.525 ;
        RECT -8.325 -0.165 -7.995 0.165 ;
        RECT -8.325 -1.525 -7.995 -1.195 ;
        RECT -8.325 -2.885 -7.995 -2.555 ;
        RECT -8.325 -4.245 -7.995 -3.915 ;
        RECT -8.325 -5.605 -7.995 -5.275 ;
        RECT -8.325 -6.965 -7.995 -6.635 ;
        RECT -8.325 -8.325 -7.995 -7.995 ;
        RECT -8.325 -9.685 -7.995 -9.355 ;
        RECT -8.325 -12.405 -7.995 -12.075 ;
        RECT -8.325 -13.765 -7.995 -13.435 ;
        RECT -8.325 -15.125 -7.995 -14.795 ;
        RECT -8.325 -16.485 -7.995 -16.155 ;
        RECT -8.325 -17.845 -7.995 -17.515 ;
        RECT -8.325 -19.205 -7.995 -18.875 ;
        RECT -8.325 -20.565 -7.995 -20.235 ;
        RECT -8.325 -21.925 -7.995 -21.595 ;
        RECT -8.325 -23.285 -7.995 -22.955 ;
        RECT -8.325 -24.645 -7.995 -24.315 ;
        RECT -8.325 -26.005 -7.995 -25.675 ;
        RECT -8.325 -27.365 -7.995 -27.035 ;
        RECT -8.325 -28.725 -7.995 -28.395 ;
        RECT -8.325 -30.085 -7.995 -29.755 ;
        RECT -8.325 -31.445 -7.995 -31.115 ;
        RECT -8.325 -32.805 -7.995 -32.475 ;
        RECT -8.325 -34.165 -7.995 -33.835 ;
        RECT -8.325 -35.525 -7.995 -35.195 ;
        RECT -8.325 -36.885 -7.995 -36.555 ;
        RECT -8.325 -38.245 -7.995 -37.915 ;
        RECT -8.325 -39.605 -7.995 -39.275 ;
        RECT -8.325 -40.965 -7.995 -40.635 ;
        RECT -8.325 -42.325 -7.995 -41.995 ;
        RECT -8.325 -43.685 -7.995 -43.355 ;
        RECT -8.325 -45.045 -7.995 -44.715 ;
        RECT -8.325 -46.405 -7.995 -46.075 ;
        RECT -8.325 -47.765 -7.995 -47.435 ;
        RECT -8.325 -49.125 -7.995 -48.795 ;
        RECT -8.325 -50.485 -7.995 -50.155 ;
        RECT -8.325 -51.845 -7.995 -51.515 ;
        RECT -8.325 -53.205 -7.995 -52.875 ;
        RECT -8.325 -54.565 -7.995 -54.235 ;
        RECT -8.325 -55.925 -7.995 -55.595 ;
        RECT -8.325 -57.285 -7.995 -56.955 ;
        RECT -8.325 -58.645 -7.995 -58.315 ;
        RECT -8.325 -60.005 -7.995 -59.675 ;
        RECT -8.325 -61.365 -7.995 -61.035 ;
        RECT -8.325 -68.165 -7.995 -67.835 ;
        RECT -8.325 -69.525 -7.995 -69.195 ;
        RECT -8.325 -70.885 -7.995 -70.555 ;
        RECT -8.325 -72.245 -7.995 -71.915 ;
        RECT -8.325 -73.605 -7.995 -73.275 ;
        RECT -8.325 -74.965 -7.995 -74.635 ;
        RECT -8.325 -76.325 -7.995 -75.995 ;
        RECT -8.325 -77.685 -7.995 -77.355 ;
        RECT -8.325 -79.045 -7.995 -78.715 ;
        RECT -8.325 -80.405 -7.995 -80.075 ;
        RECT -8.325 -81.765 -7.995 -81.435 ;
        RECT -8.325 -83.125 -7.995 -82.795 ;
        RECT -8.325 -84.485 -7.995 -84.155 ;
        RECT -8.325 -85.845 -7.995 -85.515 ;
        RECT -8.325 -87.205 -7.995 -86.875 ;
        RECT -8.325 -88.565 -7.995 -88.235 ;
        RECT -8.325 -89.925 -7.995 -89.595 ;
        RECT -8.325 -91.285 -7.995 -90.955 ;
        RECT -8.325 -92.645 -7.995 -92.315 ;
        RECT -8.325 -94.005 -7.995 -93.675 ;
        RECT -8.325 -95.365 -7.995 -95.035 ;
        RECT -8.325 -96.725 -7.995 -96.395 ;
        RECT -8.325 -98.085 -7.995 -97.755 ;
        RECT -8.325 -99.445 -7.995 -99.115 ;
        RECT -8.325 -100.805 -7.995 -100.475 ;
        RECT -8.325 -102.165 -7.995 -101.835 ;
        RECT -8.325 -103.525 -7.995 -103.195 ;
        RECT -8.325 -104.885 -7.995 -104.555 ;
        RECT -8.325 -106.245 -7.995 -105.915 ;
        RECT -8.325 -107.605 -7.995 -107.275 ;
        RECT -8.325 -108.965 -7.995 -108.635 ;
        RECT -8.325 -110.325 -7.995 -109.995 ;
        RECT -8.325 -111.685 -7.995 -111.355 ;
        RECT -8.325 -113.045 -7.995 -112.715 ;
        RECT -8.325 -114.405 -7.995 -114.075 ;
        RECT -8.325 -115.765 -7.995 -115.435 ;
        RECT -8.325 -117.125 -7.995 -116.795 ;
        RECT -8.325 -118.485 -7.995 -118.155 ;
        RECT -8.325 -119.845 -7.995 -119.515 ;
        RECT -8.325 -121.205 -7.995 -120.875 ;
        RECT -8.325 -122.565 -7.995 -122.235 ;
        RECT -8.325 -123.925 -7.995 -123.595 ;
        RECT -8.325 -125.285 -7.995 -124.955 ;
        RECT -8.325 -126.645 -7.995 -126.315 ;
        RECT -8.325 -128.005 -7.995 -127.675 ;
        RECT -8.325 -129.365 -7.995 -129.035 ;
        RECT -8.325 -130.725 -7.995 -130.395 ;
        RECT -8.325 -132.085 -7.995 -131.755 ;
        RECT -8.325 -133.445 -7.995 -133.115 ;
        RECT -8.325 -140.245 -7.995 -139.915 ;
        RECT -8.325 -141.605 -7.995 -141.275 ;
        RECT -8.325 -142.965 -7.995 -142.635 ;
        RECT -8.325 -144.325 -7.995 -143.995 ;
        RECT -8.325 -145.685 -7.995 -145.355 ;
        RECT -8.325 -147.045 -7.995 -146.715 ;
        RECT -8.325 -148.405 -7.995 -148.075 ;
        RECT -8.325 -149.765 -7.995 -149.435 ;
        RECT -8.325 -151.125 -7.995 -150.795 ;
        RECT -8.325 -152.485 -7.995 -152.155 ;
        RECT -8.325 -153.845 -7.995 -153.515 ;
        RECT -8.325 -155.205 -7.995 -154.875 ;
        RECT -8.325 -156.565 -7.995 -156.235 ;
        RECT -8.325 -157.925 -7.995 -157.595 ;
        RECT -8.325 -160.645 -7.995 -160.315 ;
        RECT -8.325 -162.005 -7.995 -161.675 ;
        RECT -8.325 -163.365 -7.995 -163.035 ;
        RECT -8.325 -164.725 -7.995 -164.395 ;
        RECT -8.325 -166.085 -7.995 -165.755 ;
        RECT -8.325 -167.445 -7.995 -167.115 ;
        RECT -8.325 -168.805 -7.995 -168.475 ;
        RECT -8.325 -170.165 -7.995 -169.835 ;
        RECT -8.325 -171.525 -7.995 -171.195 ;
        RECT -8.325 -172.885 -7.995 -172.555 ;
        RECT -8.325 -174.245 -7.995 -173.915 ;
        RECT -8.325 -175.605 -7.995 -175.275 ;
        RECT -8.325 -176.965 -7.995 -176.635 ;
        RECT -8.325 -178.325 -7.995 -177.995 ;
        RECT -8.325 -179.685 -7.995 -179.355 ;
        RECT -8.325 -181.045 -7.995 -180.715 ;
        RECT -8.325 -182.405 -7.995 -182.075 ;
        RECT -8.325 -183.765 -7.995 -183.435 ;
        RECT -8.325 -185.125 -7.995 -184.795 ;
        RECT -8.325 -186.485 -7.995 -186.155 ;
        RECT -8.325 -187.845 -7.995 -187.515 ;
        RECT -8.325 -189.205 -7.995 -188.875 ;
        RECT -8.325 -190.565 -7.995 -190.235 ;
        RECT -8.325 -191.925 -7.995 -191.595 ;
        RECT -8.325 -193.285 -7.995 -192.955 ;
        RECT -8.325 -194.645 -7.995 -194.315 ;
        RECT -8.325 -196.005 -7.995 -195.675 ;
        RECT -8.325 -197.365 -7.995 -197.035 ;
        RECT -8.325 -198.725 -7.995 -198.395 ;
        RECT -8.325 -200.085 -7.995 -199.755 ;
        RECT -8.325 -201.445 -7.995 -201.115 ;
        RECT -8.325 -202.805 -7.995 -202.475 ;
        RECT -8.325 -204.165 -7.995 -203.835 ;
        RECT -8.325 -205.525 -7.995 -205.195 ;
        RECT -8.325 -206.885 -7.995 -206.555 ;
        RECT -8.325 -208.245 -7.995 -207.915 ;
        RECT -8.325 -209.605 -7.995 -209.275 ;
        RECT -8.325 -210.965 -7.995 -210.635 ;
        RECT -8.325 -212.325 -7.995 -211.995 ;
        RECT -8.325 -213.685 -7.995 -213.355 ;
        RECT -8.325 -215.045 -7.995 -214.715 ;
        RECT -8.325 -216.405 -7.995 -216.075 ;
        RECT -8.325 -217.765 -7.995 -217.435 ;
        RECT -8.325 -219.125 -7.995 -218.795 ;
        RECT -8.325 -220.485 -7.995 -220.155 ;
        RECT -8.325 -221.845 -7.995 -221.515 ;
        RECT -8.325 -223.205 -7.995 -222.875 ;
        RECT -8.325 -224.565 -7.995 -224.235 ;
        RECT -8.325 -225.925 -7.995 -225.595 ;
        RECT -8.325 -227.285 -7.995 -226.955 ;
        RECT -8.325 -228.645 -7.995 -228.315 ;
        RECT -8.325 -230.005 -7.995 -229.675 ;
        RECT -8.325 -231.365 -7.995 -231.035 ;
        RECT -8.325 -232.725 -7.995 -232.395 ;
        RECT -8.325 -234.085 -7.995 -233.755 ;
        RECT -8.325 -235.445 -7.995 -235.115 ;
        RECT -8.325 -236.805 -7.995 -236.475 ;
        RECT -8.325 -238.165 -7.995 -237.835 ;
        RECT -8.325 -243.81 -7.995 -242.68 ;
        RECT -8.32 -243.925 -8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.965 246.76 -6.635 247.89 ;
        RECT -6.965 241.915 -6.635 242.245 ;
        RECT -6.965 240.555 -6.635 240.885 ;
        RECT -6.965 239.195 -6.635 239.525 ;
        RECT -6.965 237.835 -6.635 238.165 ;
        RECT -6.965 236.475 -6.635 236.805 ;
        RECT -6.965 235.115 -6.635 235.445 ;
        RECT -6.965 233.755 -6.635 234.085 ;
        RECT -6.965 232.395 -6.635 232.725 ;
        RECT -6.965 231.035 -6.635 231.365 ;
        RECT -6.965 221.515 -6.635 221.845 ;
        RECT -6.965 217.435 -6.635 217.765 ;
        RECT -6.965 213.355 -6.635 213.685 ;
        RECT -6.965 210.635 -6.635 210.965 ;
        RECT -6.965 203.835 -6.635 204.165 ;
        RECT -6.965 202.475 -6.635 202.805 ;
        RECT -6.965 199.755 -6.635 200.085 ;
        RECT -6.965 192.955 -6.635 193.285 ;
        RECT -6.965 190.235 -6.635 190.565 ;
        RECT -6.965 188.875 -6.635 189.205 ;
        RECT -6.965 184.795 -6.635 185.125 ;
        RECT -6.965 182.075 -6.635 182.405 ;
        RECT -6.965 175.275 -6.635 175.605 ;
        RECT -6.965 173.915 -6.635 174.245 ;
        RECT -6.965 171.195 -6.635 171.525 ;
        RECT -6.965 164.395 -6.635 164.725 ;
        RECT -6.965 161.675 -6.635 162.005 ;
        RECT -6.965 160.315 -6.635 160.645 ;
        RECT -6.965 153.515 -6.635 153.845 ;
        RECT -6.965 150.795 -6.635 151.125 ;
        RECT -6.965 146.715 -6.635 147.045 ;
        RECT -6.965 145.355 -6.635 145.685 ;
        RECT -6.965 142.635 -6.635 142.965 ;
        RECT -6.965 135.835 -6.635 136.165 ;
        RECT -6.965 133.115 -6.635 133.445 ;
        RECT -6.965 131.755 -6.635 132.085 ;
        RECT -6.965 124.955 -6.635 125.285 ;
        RECT -6.965 122.235 -6.635 122.565 ;
        RECT -6.965 118.155 -6.635 118.485 ;
        RECT -6.965 114.075 -6.635 114.405 ;
        RECT -6.965 104.555 -6.635 104.885 ;
        RECT -6.965 103.195 -6.635 103.525 ;
        RECT -6.965 96.395 -6.635 96.725 ;
        RECT -6.965 93.675 -6.635 94.005 ;
        RECT -6.965 89.595 -6.635 89.925 ;
        RECT -6.965 85.515 -6.635 85.845 ;
        RECT -6.965 82.795 -6.635 83.125 ;
        RECT -6.965 75.995 -6.635 76.325 ;
        RECT -6.965 74.635 -6.635 74.965 ;
        RECT -6.965 65.115 -6.635 65.445 ;
        RECT -6.965 61.035 -6.635 61.365 ;
        RECT -6.965 56.955 -6.635 57.285 ;
        RECT -6.965 54.235 -6.635 54.565 ;
        RECT -6.965 47.435 -6.635 47.765 ;
        RECT -6.965 46.075 -6.635 46.405 ;
        RECT -6.965 43.355 -6.635 43.685 ;
        RECT -6.965 36.555 -6.635 36.885 ;
        RECT -6.965 33.835 -6.635 34.165 ;
        RECT -6.965 32.475 -6.635 32.805 ;
        RECT -6.965 28.395 -6.635 28.725 ;
        RECT -6.965 25.675 -6.635 26.005 ;
        RECT -6.965 18.875 -6.635 19.205 ;
        RECT -6.965 17.515 -6.635 17.845 ;
        RECT -6.965 14.795 -6.635 15.125 ;
        RECT -6.965 7.995 -6.635 8.325 ;
        RECT -6.965 5.275 -6.635 5.605 ;
        RECT -6.965 3.915 -6.635 4.245 ;
        RECT -6.965 2.555 -6.635 2.885 ;
        RECT -6.965 1.195 -6.635 1.525 ;
        RECT -6.965 -0.165 -6.635 0.165 ;
        RECT -6.965 -1.525 -6.635 -1.195 ;
        RECT -6.965 -2.885 -6.635 -2.555 ;
        RECT -6.965 -4.245 -6.635 -3.915 ;
        RECT -6.965 -5.605 -6.635 -5.275 ;
        RECT -6.965 -6.965 -6.635 -6.635 ;
        RECT -6.965 -8.325 -6.635 -7.995 ;
        RECT -6.965 -9.685 -6.635 -9.355 ;
        RECT -6.965 -12.405 -6.635 -12.075 ;
        RECT -6.965 -13.765 -6.635 -13.435 ;
        RECT -6.965 -15.125 -6.635 -14.795 ;
        RECT -6.965 -16.485 -6.635 -16.155 ;
        RECT -6.965 -17.845 -6.635 -17.515 ;
        RECT -6.965 -19.205 -6.635 -18.875 ;
        RECT -6.965 -20.565 -6.635 -20.235 ;
        RECT -6.965 -21.925 -6.635 -21.595 ;
        RECT -6.965 -23.285 -6.635 -22.955 ;
        RECT -6.965 -24.645 -6.635 -24.315 ;
        RECT -6.965 -26.005 -6.635 -25.675 ;
        RECT -6.965 -27.365 -6.635 -27.035 ;
        RECT -6.965 -28.725 -6.635 -28.395 ;
        RECT -6.965 -30.085 -6.635 -29.755 ;
        RECT -6.965 -31.445 -6.635 -31.115 ;
        RECT -6.965 -32.805 -6.635 -32.475 ;
        RECT -6.965 -34.165 -6.635 -33.835 ;
        RECT -6.965 -35.525 -6.635 -35.195 ;
        RECT -6.965 -36.885 -6.635 -36.555 ;
        RECT -6.965 -38.245 -6.635 -37.915 ;
        RECT -6.965 -39.605 -6.635 -39.275 ;
        RECT -6.965 -40.965 -6.635 -40.635 ;
        RECT -6.965 -42.325 -6.635 -41.995 ;
        RECT -6.965 -43.685 -6.635 -43.355 ;
        RECT -6.965 -45.045 -6.635 -44.715 ;
        RECT -6.965 -46.405 -6.635 -46.075 ;
        RECT -6.965 -47.765 -6.635 -47.435 ;
        RECT -6.965 -49.125 -6.635 -48.795 ;
        RECT -6.965 -50.485 -6.635 -50.155 ;
        RECT -6.965 -51.845 -6.635 -51.515 ;
        RECT -6.965 -53.205 -6.635 -52.875 ;
        RECT -6.965 -54.565 -6.635 -54.235 ;
        RECT -6.965 -55.925 -6.635 -55.595 ;
        RECT -6.965 -57.285 -6.635 -56.955 ;
        RECT -6.965 -58.645 -6.635 -58.315 ;
        RECT -6.965 -60.005 -6.635 -59.675 ;
        RECT -6.965 -61.365 -6.635 -61.035 ;
        RECT -6.965 -68.165 -6.635 -67.835 ;
        RECT -6.965 -69.525 -6.635 -69.195 ;
        RECT -6.965 -70.885 -6.635 -70.555 ;
        RECT -6.965 -72.245 -6.635 -71.915 ;
        RECT -6.965 -73.605 -6.635 -73.275 ;
        RECT -6.965 -74.965 -6.635 -74.635 ;
        RECT -6.965 -76.325 -6.635 -75.995 ;
        RECT -6.965 -77.685 -6.635 -77.355 ;
        RECT -6.965 -79.045 -6.635 -78.715 ;
        RECT -6.965 -80.405 -6.635 -80.075 ;
        RECT -6.965 -81.765 -6.635 -81.435 ;
        RECT -6.965 -83.125 -6.635 -82.795 ;
        RECT -6.965 -84.485 -6.635 -84.155 ;
        RECT -6.965 -85.845 -6.635 -85.515 ;
        RECT -6.965 -87.205 -6.635 -86.875 ;
        RECT -6.965 -88.565 -6.635 -88.235 ;
        RECT -6.965 -89.925 -6.635 -89.595 ;
        RECT -6.965 -91.285 -6.635 -90.955 ;
        RECT -6.965 -92.645 -6.635 -92.315 ;
        RECT -6.965 -94.005 -6.635 -93.675 ;
        RECT -6.965 -95.365 -6.635 -95.035 ;
        RECT -6.965 -96.725 -6.635 -96.395 ;
        RECT -6.965 -98.085 -6.635 -97.755 ;
        RECT -6.965 -99.445 -6.635 -99.115 ;
        RECT -6.965 -100.805 -6.635 -100.475 ;
        RECT -6.965 -102.165 -6.635 -101.835 ;
        RECT -6.965 -103.525 -6.635 -103.195 ;
        RECT -6.965 -104.885 -6.635 -104.555 ;
        RECT -6.965 -106.245 -6.635 -105.915 ;
        RECT -6.965 -107.605 -6.635 -107.275 ;
        RECT -6.965 -108.965 -6.635 -108.635 ;
        RECT -6.965 -110.325 -6.635 -109.995 ;
        RECT -6.965 -111.685 -6.635 -111.355 ;
        RECT -6.965 -113.045 -6.635 -112.715 ;
        RECT -6.965 -114.405 -6.635 -114.075 ;
        RECT -6.965 -115.765 -6.635 -115.435 ;
        RECT -6.965 -117.125 -6.635 -116.795 ;
        RECT -6.965 -118.485 -6.635 -118.155 ;
        RECT -6.965 -119.845 -6.635 -119.515 ;
        RECT -6.965 -121.205 -6.635 -120.875 ;
        RECT -6.965 -122.565 -6.635 -122.235 ;
        RECT -6.965 -123.925 -6.635 -123.595 ;
        RECT -6.965 -125.285 -6.635 -124.955 ;
        RECT -6.965 -126.645 -6.635 -126.315 ;
        RECT -6.965 -128.005 -6.635 -127.675 ;
        RECT -6.965 -129.365 -6.635 -129.035 ;
        RECT -6.965 -130.725 -6.635 -130.395 ;
        RECT -6.965 -132.085 -6.635 -131.755 ;
        RECT -6.965 -133.445 -6.635 -133.115 ;
        RECT -6.965 -140.245 -6.635 -139.915 ;
        RECT -6.965 -141.605 -6.635 -141.275 ;
        RECT -6.965 -142.965 -6.635 -142.635 ;
        RECT -6.965 -144.325 -6.635 -143.995 ;
        RECT -6.965 -145.685 -6.635 -145.355 ;
        RECT -6.965 -147.045 -6.635 -146.715 ;
        RECT -6.965 -148.405 -6.635 -148.075 ;
        RECT -6.965 -149.765 -6.635 -149.435 ;
        RECT -6.965 -151.125 -6.635 -150.795 ;
        RECT -6.965 -152.485 -6.635 -152.155 ;
        RECT -6.965 -153.845 -6.635 -153.515 ;
        RECT -6.965 -155.205 -6.635 -154.875 ;
        RECT -6.965 -156.565 -6.635 -156.235 ;
        RECT -6.965 -157.925 -6.635 -157.595 ;
        RECT -6.965 -160.645 -6.635 -160.315 ;
        RECT -6.965 -162.005 -6.635 -161.675 ;
        RECT -6.965 -163.365 -6.635 -163.035 ;
        RECT -6.965 -164.725 -6.635 -164.395 ;
        RECT -6.965 -166.085 -6.635 -165.755 ;
        RECT -6.965 -167.445 -6.635 -167.115 ;
        RECT -6.965 -168.805 -6.635 -168.475 ;
        RECT -6.965 -170.165 -6.635 -169.835 ;
        RECT -6.965 -171.525 -6.635 -171.195 ;
        RECT -6.965 -172.885 -6.635 -172.555 ;
        RECT -6.965 -174.245 -6.635 -173.915 ;
        RECT -6.965 -175.605 -6.635 -175.275 ;
        RECT -6.965 -176.965 -6.635 -176.635 ;
        RECT -6.965 -178.325 -6.635 -177.995 ;
        RECT -6.965 -179.685 -6.635 -179.355 ;
        RECT -6.965 -181.045 -6.635 -180.715 ;
        RECT -6.965 -182.405 -6.635 -182.075 ;
        RECT -6.965 -183.765 -6.635 -183.435 ;
        RECT -6.965 -185.125 -6.635 -184.795 ;
        RECT -6.965 -186.485 -6.635 -186.155 ;
        RECT -6.965 -187.845 -6.635 -187.515 ;
        RECT -6.965 -189.205 -6.635 -188.875 ;
        RECT -6.965 -190.565 -6.635 -190.235 ;
        RECT -6.965 -191.925 -6.635 -191.595 ;
        RECT -6.965 -193.285 -6.635 -192.955 ;
        RECT -6.965 -194.645 -6.635 -194.315 ;
        RECT -6.965 -196.005 -6.635 -195.675 ;
        RECT -6.965 -197.365 -6.635 -197.035 ;
        RECT -6.965 -198.725 -6.635 -198.395 ;
        RECT -6.965 -200.085 -6.635 -199.755 ;
        RECT -6.965 -201.445 -6.635 -201.115 ;
        RECT -6.965 -202.805 -6.635 -202.475 ;
        RECT -6.965 -204.165 -6.635 -203.835 ;
        RECT -6.965 -205.525 -6.635 -205.195 ;
        RECT -6.965 -206.885 -6.635 -206.555 ;
        RECT -6.965 -208.245 -6.635 -207.915 ;
        RECT -6.965 -209.605 -6.635 -209.275 ;
        RECT -6.965 -210.965 -6.635 -210.635 ;
        RECT -6.965 -212.325 -6.635 -211.995 ;
        RECT -6.965 -213.685 -6.635 -213.355 ;
        RECT -6.965 -215.045 -6.635 -214.715 ;
        RECT -6.965 -216.405 -6.635 -216.075 ;
        RECT -6.965 -217.765 -6.635 -217.435 ;
        RECT -6.965 -219.125 -6.635 -218.795 ;
        RECT -6.965 -220.485 -6.635 -220.155 ;
        RECT -6.965 -221.845 -6.635 -221.515 ;
        RECT -6.965 -223.205 -6.635 -222.875 ;
        RECT -6.965 -224.565 -6.635 -224.235 ;
        RECT -6.965 -225.925 -6.635 -225.595 ;
        RECT -6.965 -227.285 -6.635 -226.955 ;
        RECT -6.965 -228.645 -6.635 -228.315 ;
        RECT -6.965 -230.005 -6.635 -229.675 ;
        RECT -6.965 -231.365 -6.635 -231.035 ;
        RECT -6.965 -232.725 -6.635 -232.395 ;
        RECT -6.965 -234.085 -6.635 -233.755 ;
        RECT -6.965 -235.445 -6.635 -235.115 ;
        RECT -6.965 -236.805 -6.635 -236.475 ;
        RECT -6.965 -238.165 -6.635 -237.835 ;
        RECT -6.965 -243.81 -6.635 -242.68 ;
        RECT -6.96 -243.925 -6.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.605 -121.205 -5.275 -120.875 ;
        RECT -5.605 -122.565 -5.275 -122.235 ;
        RECT -5.605 -123.925 -5.275 -123.595 ;
        RECT -5.605 -125.285 -5.275 -124.955 ;
        RECT -5.605 -126.645 -5.275 -126.315 ;
        RECT -5.605 -128.005 -5.275 -127.675 ;
        RECT -5.605 -129.365 -5.275 -129.035 ;
        RECT -5.605 -130.725 -5.275 -130.395 ;
        RECT -5.605 -132.085 -5.275 -131.755 ;
        RECT -5.605 -133.445 -5.275 -133.115 ;
        RECT -5.605 -140.245 -5.275 -139.915 ;
        RECT -5.605 -141.605 -5.275 -141.275 ;
        RECT -5.605 -142.965 -5.275 -142.635 ;
        RECT -5.605 -144.325 -5.275 -143.995 ;
        RECT -5.605 -145.685 -5.275 -145.355 ;
        RECT -5.605 -147.045 -5.275 -146.715 ;
        RECT -5.605 -148.405 -5.275 -148.075 ;
        RECT -5.605 -149.765 -5.275 -149.435 ;
        RECT -5.605 -151.125 -5.275 -150.795 ;
        RECT -5.605 -152.485 -5.275 -152.155 ;
        RECT -5.605 -153.845 -5.275 -153.515 ;
        RECT -5.605 -155.205 -5.275 -154.875 ;
        RECT -5.605 -156.565 -5.275 -156.235 ;
        RECT -5.605 -157.925 -5.275 -157.595 ;
        RECT -5.605 -160.645 -5.275 -160.315 ;
        RECT -5.605 -162.005 -5.275 -161.675 ;
        RECT -5.605 -163.365 -5.275 -163.035 ;
        RECT -5.605 -164.725 -5.275 -164.395 ;
        RECT -5.605 -166.085 -5.275 -165.755 ;
        RECT -5.605 -167.445 -5.275 -167.115 ;
        RECT -5.605 -168.805 -5.275 -168.475 ;
        RECT -5.605 -170.165 -5.275 -169.835 ;
        RECT -5.605 -171.525 -5.275 -171.195 ;
        RECT -5.605 -172.885 -5.275 -172.555 ;
        RECT -5.605 -174.245 -5.275 -173.915 ;
        RECT -5.605 -175.605 -5.275 -175.275 ;
        RECT -5.605 -176.965 -5.275 -176.635 ;
        RECT -5.605 -178.325 -5.275 -177.995 ;
        RECT -5.605 -179.685 -5.275 -179.355 ;
        RECT -5.605 -181.045 -5.275 -180.715 ;
        RECT -5.605 -182.405 -5.275 -182.075 ;
        RECT -5.605 -183.765 -5.275 -183.435 ;
        RECT -5.605 -185.125 -5.275 -184.795 ;
        RECT -5.605 -186.485 -5.275 -186.155 ;
        RECT -5.605 -187.845 -5.275 -187.515 ;
        RECT -5.605 -189.205 -5.275 -188.875 ;
        RECT -5.605 -190.565 -5.275 -190.235 ;
        RECT -5.605 -191.925 -5.275 -191.595 ;
        RECT -5.605 -193.285 -5.275 -192.955 ;
        RECT -5.605 -194.645 -5.275 -194.315 ;
        RECT -5.605 -196.005 -5.275 -195.675 ;
        RECT -5.605 -197.365 -5.275 -197.035 ;
        RECT -5.605 -198.725 -5.275 -198.395 ;
        RECT -5.605 -200.085 -5.275 -199.755 ;
        RECT -5.605 -201.445 -5.275 -201.115 ;
        RECT -5.605 -202.805 -5.275 -202.475 ;
        RECT -5.605 -204.165 -5.275 -203.835 ;
        RECT -5.605 -205.525 -5.275 -205.195 ;
        RECT -5.605 -206.885 -5.275 -206.555 ;
        RECT -5.605 -208.245 -5.275 -207.915 ;
        RECT -5.605 -209.605 -5.275 -209.275 ;
        RECT -5.605 -210.965 -5.275 -210.635 ;
        RECT -5.605 -212.325 -5.275 -211.995 ;
        RECT -5.605 -213.685 -5.275 -213.355 ;
        RECT -5.605 -215.045 -5.275 -214.715 ;
        RECT -5.605 -216.405 -5.275 -216.075 ;
        RECT -5.605 -217.765 -5.275 -217.435 ;
        RECT -5.605 -219.125 -5.275 -218.795 ;
        RECT -5.605 -220.485 -5.275 -220.155 ;
        RECT -5.605 -221.845 -5.275 -221.515 ;
        RECT -5.605 -223.205 -5.275 -222.875 ;
        RECT -5.605 -224.565 -5.275 -224.235 ;
        RECT -5.605 -225.925 -5.275 -225.595 ;
        RECT -5.605 -227.285 -5.275 -226.955 ;
        RECT -5.605 -228.645 -5.275 -228.315 ;
        RECT -5.605 -230.005 -5.275 -229.675 ;
        RECT -5.605 -231.365 -5.275 -231.035 ;
        RECT -5.605 -232.725 -5.275 -232.395 ;
        RECT -5.605 -234.085 -5.275 -233.755 ;
        RECT -5.605 -235.445 -5.275 -235.115 ;
        RECT -5.605 -236.805 -5.275 -236.475 ;
        RECT -5.605 -238.165 -5.275 -237.835 ;
        RECT -5.605 -243.81 -5.275 -242.68 ;
        RECT -5.6 -243.925 -5.28 248.005 ;
        RECT -5.605 246.76 -5.275 247.89 ;
        RECT -5.605 241.915 -5.275 242.245 ;
        RECT -5.605 240.555 -5.275 240.885 ;
        RECT -5.605 239.195 -5.275 239.525 ;
        RECT -5.605 237.835 -5.275 238.165 ;
        RECT -5.605 235.17 -5.275 235.5 ;
        RECT -5.605 232.995 -5.275 233.325 ;
        RECT -5.605 231.415 -5.275 231.745 ;
        RECT -5.605 230.565 -5.275 230.895 ;
        RECT -5.605 228.255 -5.275 228.585 ;
        RECT -5.605 227.405 -5.275 227.735 ;
        RECT -5.605 225.095 -5.275 225.425 ;
        RECT -5.605 224.245 -5.275 224.575 ;
        RECT -5.605 221.935 -5.275 222.265 ;
        RECT -5.605 221.085 -5.275 221.415 ;
        RECT -5.605 218.775 -5.275 219.105 ;
        RECT -5.605 217.195 -5.275 217.525 ;
        RECT -5.605 216.345 -5.275 216.675 ;
        RECT -5.605 214.035 -5.275 214.365 ;
        RECT -5.605 213.185 -5.275 213.515 ;
        RECT -5.605 210.875 -5.275 211.205 ;
        RECT -5.605 210.025 -5.275 210.355 ;
        RECT -5.605 207.715 -5.275 208.045 ;
        RECT -5.605 206.865 -5.275 207.195 ;
        RECT -5.605 204.555 -5.275 204.885 ;
        RECT -5.605 202.975 -5.275 203.305 ;
        RECT -5.605 202.125 -5.275 202.455 ;
        RECT -5.605 199.815 -5.275 200.145 ;
        RECT -5.605 198.965 -5.275 199.295 ;
        RECT -5.605 196.655 -5.275 196.985 ;
        RECT -5.605 195.805 -5.275 196.135 ;
        RECT -5.605 193.495 -5.275 193.825 ;
        RECT -5.605 192.645 -5.275 192.975 ;
        RECT -5.605 190.335 -5.275 190.665 ;
        RECT -5.605 188.755 -5.275 189.085 ;
        RECT -5.605 187.905 -5.275 188.235 ;
        RECT -5.605 185.595 -5.275 185.925 ;
        RECT -5.605 184.745 -5.275 185.075 ;
        RECT -5.605 182.435 -5.275 182.765 ;
        RECT -5.605 181.585 -5.275 181.915 ;
        RECT -5.605 179.275 -5.275 179.605 ;
        RECT -5.605 178.425 -5.275 178.755 ;
        RECT -5.605 176.115 -5.275 176.445 ;
        RECT -5.605 174.535 -5.275 174.865 ;
        RECT -5.605 173.685 -5.275 174.015 ;
        RECT -5.605 171.375 -5.275 171.705 ;
        RECT -5.605 170.525 -5.275 170.855 ;
        RECT -5.605 168.215 -5.275 168.545 ;
        RECT -5.605 167.365 -5.275 167.695 ;
        RECT -5.605 165.055 -5.275 165.385 ;
        RECT -5.605 164.205 -5.275 164.535 ;
        RECT -5.605 161.895 -5.275 162.225 ;
        RECT -5.605 160.315 -5.275 160.645 ;
        RECT -5.605 159.465 -5.275 159.795 ;
        RECT -5.605 157.155 -5.275 157.485 ;
        RECT -5.605 156.305 -5.275 156.635 ;
        RECT -5.605 153.995 -5.275 154.325 ;
        RECT -5.605 153.145 -5.275 153.475 ;
        RECT -5.605 150.835 -5.275 151.165 ;
        RECT -5.605 149.985 -5.275 150.315 ;
        RECT -5.605 147.675 -5.275 148.005 ;
        RECT -5.605 146.095 -5.275 146.425 ;
        RECT -5.605 145.245 -5.275 145.575 ;
        RECT -5.605 142.935 -5.275 143.265 ;
        RECT -5.605 142.085 -5.275 142.415 ;
        RECT -5.605 139.775 -5.275 140.105 ;
        RECT -5.605 138.925 -5.275 139.255 ;
        RECT -5.605 136.615 -5.275 136.945 ;
        RECT -5.605 135.765 -5.275 136.095 ;
        RECT -5.605 133.455 -5.275 133.785 ;
        RECT -5.605 131.875 -5.275 132.205 ;
        RECT -5.605 131.025 -5.275 131.355 ;
        RECT -5.605 128.715 -5.275 129.045 ;
        RECT -5.605 127.865 -5.275 128.195 ;
        RECT -5.605 125.555 -5.275 125.885 ;
        RECT -5.605 124.705 -5.275 125.035 ;
        RECT -5.605 122.395 -5.275 122.725 ;
        RECT -5.605 121.545 -5.275 121.875 ;
        RECT -5.605 119.235 -5.275 119.565 ;
        RECT -5.605 117.655 -5.275 117.985 ;
        RECT -5.605 116.805 -5.275 117.135 ;
        RECT -5.605 114.495 -5.275 114.825 ;
        RECT -5.605 113.645 -5.275 113.975 ;
        RECT -5.605 111.335 -5.275 111.665 ;
        RECT -5.605 110.485 -5.275 110.815 ;
        RECT -5.605 108.175 -5.275 108.505 ;
        RECT -5.605 107.325 -5.275 107.655 ;
        RECT -5.605 105.015 -5.275 105.345 ;
        RECT -5.605 103.435 -5.275 103.765 ;
        RECT -5.605 102.585 -5.275 102.915 ;
        RECT -5.605 100.275 -5.275 100.605 ;
        RECT -5.605 99.425 -5.275 99.755 ;
        RECT -5.605 97.115 -5.275 97.445 ;
        RECT -5.605 96.265 -5.275 96.595 ;
        RECT -5.605 93.955 -5.275 94.285 ;
        RECT -5.605 93.105 -5.275 93.435 ;
        RECT -5.605 90.795 -5.275 91.125 ;
        RECT -5.605 89.215 -5.275 89.545 ;
        RECT -5.605 88.365 -5.275 88.695 ;
        RECT -5.605 86.055 -5.275 86.385 ;
        RECT -5.605 85.205 -5.275 85.535 ;
        RECT -5.605 82.895 -5.275 83.225 ;
        RECT -5.605 82.045 -5.275 82.375 ;
        RECT -5.605 79.735 -5.275 80.065 ;
        RECT -5.605 78.885 -5.275 79.215 ;
        RECT -5.605 76.575 -5.275 76.905 ;
        RECT -5.605 74.995 -5.275 75.325 ;
        RECT -5.605 74.145 -5.275 74.475 ;
        RECT -5.605 71.835 -5.275 72.165 ;
        RECT -5.605 70.985 -5.275 71.315 ;
        RECT -5.605 68.675 -5.275 69.005 ;
        RECT -5.605 67.825 -5.275 68.155 ;
        RECT -5.605 65.515 -5.275 65.845 ;
        RECT -5.605 64.665 -5.275 64.995 ;
        RECT -5.605 62.355 -5.275 62.685 ;
        RECT -5.605 60.775 -5.275 61.105 ;
        RECT -5.605 59.925 -5.275 60.255 ;
        RECT -5.605 57.615 -5.275 57.945 ;
        RECT -5.605 56.765 -5.275 57.095 ;
        RECT -5.605 54.455 -5.275 54.785 ;
        RECT -5.605 53.605 -5.275 53.935 ;
        RECT -5.605 51.295 -5.275 51.625 ;
        RECT -5.605 50.445 -5.275 50.775 ;
        RECT -5.605 48.135 -5.275 48.465 ;
        RECT -5.605 46.555 -5.275 46.885 ;
        RECT -5.605 45.705 -5.275 46.035 ;
        RECT -5.605 43.395 -5.275 43.725 ;
        RECT -5.605 42.545 -5.275 42.875 ;
        RECT -5.605 40.235 -5.275 40.565 ;
        RECT -5.605 39.385 -5.275 39.715 ;
        RECT -5.605 37.075 -5.275 37.405 ;
        RECT -5.605 36.225 -5.275 36.555 ;
        RECT -5.605 33.915 -5.275 34.245 ;
        RECT -5.605 32.335 -5.275 32.665 ;
        RECT -5.605 31.485 -5.275 31.815 ;
        RECT -5.605 29.175 -5.275 29.505 ;
        RECT -5.605 28.325 -5.275 28.655 ;
        RECT -5.605 26.015 -5.275 26.345 ;
        RECT -5.605 25.165 -5.275 25.495 ;
        RECT -5.605 22.855 -5.275 23.185 ;
        RECT -5.605 22.005 -5.275 22.335 ;
        RECT -5.605 19.695 -5.275 20.025 ;
        RECT -5.605 18.115 -5.275 18.445 ;
        RECT -5.605 17.265 -5.275 17.595 ;
        RECT -5.605 14.955 -5.275 15.285 ;
        RECT -5.605 14.105 -5.275 14.435 ;
        RECT -5.605 11.795 -5.275 12.125 ;
        RECT -5.605 10.945 -5.275 11.275 ;
        RECT -5.605 8.635 -5.275 8.965 ;
        RECT -5.605 7.785 -5.275 8.115 ;
        RECT -5.605 5.475 -5.275 5.805 ;
        RECT -5.605 3.895 -5.275 4.225 ;
        RECT -5.605 3.045 -5.275 3.375 ;
        RECT -5.605 0.87 -5.275 1.2 ;
        RECT -5.605 -1.525 -5.275 -1.195 ;
        RECT -5.605 -2.885 -5.275 -2.555 ;
        RECT -5.605 -4.245 -5.275 -3.915 ;
        RECT -5.605 -5.605 -5.275 -5.275 ;
        RECT -5.605 -6.965 -5.275 -6.635 ;
        RECT -5.605 -8.325 -5.275 -7.995 ;
        RECT -5.605 -9.685 -5.275 -9.355 ;
        RECT -5.605 -12.405 -5.275 -12.075 ;
        RECT -5.605 -13.765 -5.275 -13.435 ;
        RECT -5.605 -15.125 -5.275 -14.795 ;
        RECT -5.605 -16.485 -5.275 -16.155 ;
        RECT -5.605 -17.845 -5.275 -17.515 ;
        RECT -5.605 -19.205 -5.275 -18.875 ;
        RECT -5.605 -20.565 -5.275 -20.235 ;
        RECT -5.605 -21.925 -5.275 -21.595 ;
        RECT -5.605 -23.285 -5.275 -22.955 ;
        RECT -5.605 -24.645 -5.275 -24.315 ;
        RECT -5.605 -26.005 -5.275 -25.675 ;
        RECT -5.605 -27.365 -5.275 -27.035 ;
        RECT -5.605 -28.725 -5.275 -28.395 ;
        RECT -5.605 -30.085 -5.275 -29.755 ;
        RECT -5.605 -31.445 -5.275 -31.115 ;
        RECT -5.605 -32.805 -5.275 -32.475 ;
        RECT -5.605 -34.165 -5.275 -33.835 ;
        RECT -5.605 -35.525 -5.275 -35.195 ;
        RECT -5.605 -36.885 -5.275 -36.555 ;
        RECT -5.605 -38.245 -5.275 -37.915 ;
        RECT -5.605 -39.605 -5.275 -39.275 ;
        RECT -5.605 -40.965 -5.275 -40.635 ;
        RECT -5.605 -42.325 -5.275 -41.995 ;
        RECT -5.605 -43.685 -5.275 -43.355 ;
        RECT -5.605 -45.045 -5.275 -44.715 ;
        RECT -5.605 -46.405 -5.275 -46.075 ;
        RECT -5.605 -47.765 -5.275 -47.435 ;
        RECT -5.605 -49.125 -5.275 -48.795 ;
        RECT -5.605 -50.485 -5.275 -50.155 ;
        RECT -5.605 -51.845 -5.275 -51.515 ;
        RECT -5.605 -53.205 -5.275 -52.875 ;
        RECT -5.605 -54.565 -5.275 -54.235 ;
        RECT -5.605 -55.925 -5.275 -55.595 ;
        RECT -5.605 -57.285 -5.275 -56.955 ;
        RECT -5.605 -58.645 -5.275 -58.315 ;
        RECT -5.605 -60.005 -5.275 -59.675 ;
        RECT -5.605 -61.365 -5.275 -61.035 ;
        RECT -5.605 -68.165 -5.275 -67.835 ;
        RECT -5.605 -69.525 -5.275 -69.195 ;
        RECT -5.605 -70.885 -5.275 -70.555 ;
        RECT -5.605 -72.245 -5.275 -71.915 ;
        RECT -5.605 -73.605 -5.275 -73.275 ;
        RECT -5.605 -74.965 -5.275 -74.635 ;
        RECT -5.605 -76.325 -5.275 -75.995 ;
        RECT -5.605 -77.685 -5.275 -77.355 ;
        RECT -5.605 -79.045 -5.275 -78.715 ;
        RECT -5.605 -80.405 -5.275 -80.075 ;
        RECT -5.605 -81.765 -5.275 -81.435 ;
        RECT -5.605 -83.125 -5.275 -82.795 ;
        RECT -5.605 -84.485 -5.275 -84.155 ;
        RECT -5.605 -85.845 -5.275 -85.515 ;
        RECT -5.605 -87.205 -5.275 -86.875 ;
        RECT -5.605 -88.565 -5.275 -88.235 ;
        RECT -5.605 -89.925 -5.275 -89.595 ;
        RECT -5.605 -91.285 -5.275 -90.955 ;
        RECT -5.605 -92.645 -5.275 -92.315 ;
        RECT -5.605 -94.005 -5.275 -93.675 ;
        RECT -5.605 -95.365 -5.275 -95.035 ;
        RECT -5.605 -96.725 -5.275 -96.395 ;
        RECT -5.605 -98.085 -5.275 -97.755 ;
        RECT -5.605 -99.445 -5.275 -99.115 ;
        RECT -5.605 -100.805 -5.275 -100.475 ;
        RECT -5.605 -102.165 -5.275 -101.835 ;
        RECT -5.605 -103.525 -5.275 -103.195 ;
        RECT -5.605 -104.885 -5.275 -104.555 ;
        RECT -5.605 -106.245 -5.275 -105.915 ;
        RECT -5.605 -107.605 -5.275 -107.275 ;
        RECT -5.605 -108.965 -5.275 -108.635 ;
        RECT -5.605 -110.325 -5.275 -109.995 ;
        RECT -5.605 -111.685 -5.275 -111.355 ;
        RECT -5.605 -113.045 -5.275 -112.715 ;
        RECT -5.605 -114.405 -5.275 -114.075 ;
        RECT -5.605 -115.765 -5.275 -115.435 ;
        RECT -5.605 -117.125 -5.275 -116.795 ;
        RECT -5.605 -118.485 -5.275 -118.155 ;
        RECT -5.605 -119.845 -5.275 -119.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -164.725 -16.155 -164.395 ;
        RECT -16.485 -167.445 -16.155 -167.115 ;
        RECT -16.485 -168.805 -16.155 -168.475 ;
        RECT -16.485 -170.165 -16.155 -169.835 ;
        RECT -16.485 -171.525 -16.155 -171.195 ;
        RECT -16.485 -175.605 -16.155 -175.275 ;
        RECT -16.485 -176.965 -16.155 -176.635 ;
        RECT -16.485 -178.325 -16.155 -177.995 ;
        RECT -16.485 -179.685 -16.155 -179.355 ;
        RECT -16.485 -181.045 -16.155 -180.715 ;
        RECT -16.485 -182.405 -16.155 -182.075 ;
        RECT -16.485 -185.125 -16.155 -184.795 ;
        RECT -16.485 -194.645 -16.155 -194.315 ;
        RECT -16.485 -196.005 -16.155 -195.675 ;
        RECT -16.485 -198.725 -16.155 -198.395 ;
        RECT -16.485 -201.445 -16.155 -201.115 ;
        RECT -16.485 -202.805 -16.155 -202.475 ;
        RECT -16.485 -209.605 -16.155 -209.275 ;
        RECT -16.485 -213.685 -16.155 -213.355 ;
        RECT -16.485 -215.045 -16.155 -214.715 ;
        RECT -16.485 -216.405 -16.155 -216.075 ;
        RECT -16.485 -217.765 -16.155 -217.435 ;
        RECT -16.485 -219.125 -16.155 -218.795 ;
        RECT -16.485 -220.485 -16.155 -220.155 ;
        RECT -16.485 -221.845 -16.155 -221.515 ;
        RECT -16.485 -223.205 -16.155 -222.875 ;
        RECT -16.48 -223.88 -16.16 -161.68 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -234.085 -16.155 -233.755 ;
        RECT -16.485 -235.445 -16.155 -235.115 ;
        RECT -16.485 -236.805 -16.155 -236.475 ;
        RECT -16.485 -238.165 -16.155 -237.835 ;
        RECT -16.485 -243.81 -16.155 -242.68 ;
        RECT -16.48 -243.925 -16.16 -231.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 246.76 -14.795 247.89 ;
        RECT -15.125 241.915 -14.795 242.245 ;
        RECT -15.125 240.555 -14.795 240.885 ;
        RECT -15.125 239.195 -14.795 239.525 ;
        RECT -15.125 237.835 -14.795 238.165 ;
        RECT -15.125 236.475 -14.795 236.805 ;
        RECT -15.125 235.115 -14.795 235.445 ;
        RECT -15.125 233.755 -14.795 234.085 ;
        RECT -15.125 232.395 -14.795 232.725 ;
        RECT -15.125 231.035 -14.795 231.365 ;
        RECT -15.125 229.675 -14.795 230.005 ;
        RECT -15.125 228.315 -14.795 228.645 ;
        RECT -15.125 226.955 -14.795 227.285 ;
        RECT -15.125 225.595 -14.795 225.925 ;
        RECT -15.125 224.235 -14.795 224.565 ;
        RECT -15.125 222.875 -14.795 223.205 ;
        RECT -15.125 221.515 -14.795 221.845 ;
        RECT -15.125 220.155 -14.795 220.485 ;
        RECT -15.125 218.795 -14.795 219.125 ;
        RECT -15.125 217.435 -14.795 217.765 ;
        RECT -15.125 216.075 -14.795 216.405 ;
        RECT -15.125 214.715 -14.795 215.045 ;
        RECT -15.125 213.355 -14.795 213.685 ;
        RECT -15.125 211.995 -14.795 212.325 ;
        RECT -15.125 210.635 -14.795 210.965 ;
        RECT -15.125 209.275 -14.795 209.605 ;
        RECT -15.125 207.915 -14.795 208.245 ;
        RECT -15.125 206.555 -14.795 206.885 ;
        RECT -15.125 205.195 -14.795 205.525 ;
        RECT -15.125 203.835 -14.795 204.165 ;
        RECT -15.125 202.475 -14.795 202.805 ;
        RECT -15.125 201.115 -14.795 201.445 ;
        RECT -15.125 199.755 -14.795 200.085 ;
        RECT -15.125 198.395 -14.795 198.725 ;
        RECT -15.125 197.035 -14.795 197.365 ;
        RECT -15.125 195.675 -14.795 196.005 ;
        RECT -15.125 194.315 -14.795 194.645 ;
        RECT -15.125 192.955 -14.795 193.285 ;
        RECT -15.125 191.595 -14.795 191.925 ;
        RECT -15.125 190.235 -14.795 190.565 ;
        RECT -15.125 188.875 -14.795 189.205 ;
        RECT -15.125 187.515 -14.795 187.845 ;
        RECT -15.125 186.155 -14.795 186.485 ;
        RECT -15.125 184.795 -14.795 185.125 ;
        RECT -15.125 183.435 -14.795 183.765 ;
        RECT -15.125 182.075 -14.795 182.405 ;
        RECT -15.125 180.715 -14.795 181.045 ;
        RECT -15.125 179.355 -14.795 179.685 ;
        RECT -15.125 177.995 -14.795 178.325 ;
        RECT -15.125 176.635 -14.795 176.965 ;
        RECT -15.125 175.275 -14.795 175.605 ;
        RECT -15.125 173.915 -14.795 174.245 ;
        RECT -15.125 172.555 -14.795 172.885 ;
        RECT -15.125 171.195 -14.795 171.525 ;
        RECT -15.125 169.835 -14.795 170.165 ;
        RECT -15.125 168.475 -14.795 168.805 ;
        RECT -15.125 167.115 -14.795 167.445 ;
        RECT -15.125 165.755 -14.795 166.085 ;
        RECT -15.125 164.395 -14.795 164.725 ;
        RECT -15.125 163.035 -14.795 163.365 ;
        RECT -15.125 161.675 -14.795 162.005 ;
        RECT -15.125 160.315 -14.795 160.645 ;
        RECT -15.125 158.955 -14.795 159.285 ;
        RECT -15.125 157.595 -14.795 157.925 ;
        RECT -15.125 156.235 -14.795 156.565 ;
        RECT -15.125 154.875 -14.795 155.205 ;
        RECT -15.125 153.515 -14.795 153.845 ;
        RECT -15.125 152.155 -14.795 152.485 ;
        RECT -15.125 150.795 -14.795 151.125 ;
        RECT -15.125 149.435 -14.795 149.765 ;
        RECT -15.125 148.075 -14.795 148.405 ;
        RECT -15.125 146.715 -14.795 147.045 ;
        RECT -15.125 145.355 -14.795 145.685 ;
        RECT -15.125 143.995 -14.795 144.325 ;
        RECT -15.125 142.635 -14.795 142.965 ;
        RECT -15.125 141.275 -14.795 141.605 ;
        RECT -15.125 139.915 -14.795 140.245 ;
        RECT -15.125 138.555 -14.795 138.885 ;
        RECT -15.125 137.195 -14.795 137.525 ;
        RECT -15.125 135.835 -14.795 136.165 ;
        RECT -15.125 134.475 -14.795 134.805 ;
        RECT -15.125 133.115 -14.795 133.445 ;
        RECT -15.125 131.755 -14.795 132.085 ;
        RECT -15.125 130.395 -14.795 130.725 ;
        RECT -15.125 129.035 -14.795 129.365 ;
        RECT -15.125 127.675 -14.795 128.005 ;
        RECT -15.125 126.315 -14.795 126.645 ;
        RECT -15.125 124.955 -14.795 125.285 ;
        RECT -15.125 123.595 -14.795 123.925 ;
        RECT -15.125 122.235 -14.795 122.565 ;
        RECT -15.125 120.875 -14.795 121.205 ;
        RECT -15.125 119.515 -14.795 119.845 ;
        RECT -15.125 118.155 -14.795 118.485 ;
        RECT -15.125 116.795 -14.795 117.125 ;
        RECT -15.125 115.435 -14.795 115.765 ;
        RECT -15.125 114.075 -14.795 114.405 ;
        RECT -15.125 112.715 -14.795 113.045 ;
        RECT -15.125 111.355 -14.795 111.685 ;
        RECT -15.125 109.995 -14.795 110.325 ;
        RECT -15.125 108.635 -14.795 108.965 ;
        RECT -15.125 107.275 -14.795 107.605 ;
        RECT -15.125 105.915 -14.795 106.245 ;
        RECT -15.125 104.555 -14.795 104.885 ;
        RECT -15.125 103.195 -14.795 103.525 ;
        RECT -15.125 101.835 -14.795 102.165 ;
        RECT -15.125 100.475 -14.795 100.805 ;
        RECT -15.125 99.115 -14.795 99.445 ;
        RECT -15.125 97.755 -14.795 98.085 ;
        RECT -15.125 96.395 -14.795 96.725 ;
        RECT -15.125 95.035 -14.795 95.365 ;
        RECT -15.125 93.675 -14.795 94.005 ;
        RECT -15.125 92.315 -14.795 92.645 ;
        RECT -15.125 90.955 -14.795 91.285 ;
        RECT -15.125 89.595 -14.795 89.925 ;
        RECT -15.125 88.235 -14.795 88.565 ;
        RECT -15.125 86.875 -14.795 87.205 ;
        RECT -15.125 85.515 -14.795 85.845 ;
        RECT -15.125 84.155 -14.795 84.485 ;
        RECT -15.125 82.795 -14.795 83.125 ;
        RECT -15.125 81.435 -14.795 81.765 ;
        RECT -15.125 80.075 -14.795 80.405 ;
        RECT -15.125 78.715 -14.795 79.045 ;
        RECT -15.125 77.355 -14.795 77.685 ;
        RECT -15.125 75.995 -14.795 76.325 ;
        RECT -15.125 74.635 -14.795 74.965 ;
        RECT -15.125 73.275 -14.795 73.605 ;
        RECT -15.125 71.915 -14.795 72.245 ;
        RECT -15.125 70.555 -14.795 70.885 ;
        RECT -15.125 69.195 -14.795 69.525 ;
        RECT -15.125 67.835 -14.795 68.165 ;
        RECT -15.125 66.475 -14.795 66.805 ;
        RECT -15.125 65.115 -14.795 65.445 ;
        RECT -15.125 63.755 -14.795 64.085 ;
        RECT -15.125 62.395 -14.795 62.725 ;
        RECT -15.125 61.035 -14.795 61.365 ;
        RECT -15.125 59.675 -14.795 60.005 ;
        RECT -15.125 58.315 -14.795 58.645 ;
        RECT -15.125 56.955 -14.795 57.285 ;
        RECT -15.125 55.595 -14.795 55.925 ;
        RECT -15.125 54.235 -14.795 54.565 ;
        RECT -15.125 52.875 -14.795 53.205 ;
        RECT -15.125 51.515 -14.795 51.845 ;
        RECT -15.125 50.155 -14.795 50.485 ;
        RECT -15.125 48.795 -14.795 49.125 ;
        RECT -15.125 47.435 -14.795 47.765 ;
        RECT -15.125 46.075 -14.795 46.405 ;
        RECT -15.125 44.715 -14.795 45.045 ;
        RECT -15.125 43.355 -14.795 43.685 ;
        RECT -15.125 41.995 -14.795 42.325 ;
        RECT -15.125 40.635 -14.795 40.965 ;
        RECT -15.125 39.275 -14.795 39.605 ;
        RECT -15.125 37.915 -14.795 38.245 ;
        RECT -15.125 36.555 -14.795 36.885 ;
        RECT -15.125 35.195 -14.795 35.525 ;
        RECT -15.125 33.835 -14.795 34.165 ;
        RECT -15.125 32.475 -14.795 32.805 ;
        RECT -15.125 31.115 -14.795 31.445 ;
        RECT -15.125 29.755 -14.795 30.085 ;
        RECT -15.125 28.395 -14.795 28.725 ;
        RECT -15.125 27.035 -14.795 27.365 ;
        RECT -15.125 25.675 -14.795 26.005 ;
        RECT -15.125 24.315 -14.795 24.645 ;
        RECT -15.125 22.955 -14.795 23.285 ;
        RECT -15.125 21.595 -14.795 21.925 ;
        RECT -15.125 20.235 -14.795 20.565 ;
        RECT -15.125 18.875 -14.795 19.205 ;
        RECT -15.125 17.515 -14.795 17.845 ;
        RECT -15.125 16.155 -14.795 16.485 ;
        RECT -15.125 14.795 -14.795 15.125 ;
        RECT -15.125 13.435 -14.795 13.765 ;
        RECT -15.125 12.075 -14.795 12.405 ;
        RECT -15.125 10.715 -14.795 11.045 ;
        RECT -15.125 9.355 -14.795 9.685 ;
        RECT -15.125 7.995 -14.795 8.325 ;
        RECT -15.125 6.635 -14.795 6.965 ;
        RECT -15.125 5.275 -14.795 5.605 ;
        RECT -15.125 3.915 -14.795 4.245 ;
        RECT -15.125 2.555 -14.795 2.885 ;
        RECT -15.125 1.195 -14.795 1.525 ;
        RECT -15.125 -0.165 -14.795 0.165 ;
        RECT -15.125 -1.525 -14.795 -1.195 ;
        RECT -15.125 -2.885 -14.795 -2.555 ;
        RECT -15.125 -4.245 -14.795 -3.915 ;
        RECT -15.125 -5.605 -14.795 -5.275 ;
        RECT -15.125 -6.965 -14.795 -6.635 ;
        RECT -15.125 -8.325 -14.795 -7.995 ;
        RECT -15.125 -9.48 -14.795 -9.15 ;
        RECT -15.125 -12.405 -14.795 -12.075 ;
        RECT -15.125 -15.125 -14.795 -14.795 ;
        RECT -15.125 -16.67 -14.795 -16.34 ;
        RECT -15.125 -17.845 -14.795 -17.515 ;
        RECT -15.125 -24.645 -14.795 -24.315 ;
        RECT -15.125 -26.005 -14.795 -25.675 ;
        RECT -15.125 -27.365 -14.795 -27.035 ;
        RECT -15.125 -30.66 -14.795 -30.33 ;
        RECT -15.125 -31.445 -14.795 -31.115 ;
        RECT -15.125 -32.805 -14.795 -32.475 ;
        RECT -15.125 -34.165 -14.795 -33.835 ;
        RECT -15.125 -36.885 -14.795 -36.555 ;
        RECT -15.125 -37.85 -14.795 -37.52 ;
        RECT -15.125 -40.965 -14.795 -40.635 ;
        RECT -15.125 -46.405 -14.795 -46.075 ;
        RECT -15.125 -47.765 -14.795 -47.435 ;
        RECT -15.125 -49.125 -14.795 -48.795 ;
        RECT -15.125 -50.485 -14.795 -50.155 ;
        RECT -15.125 -51.845 -14.795 -51.515 ;
        RECT -15.125 -53.205 -14.795 -52.875 ;
        RECT -15.125 -54.565 -14.795 -54.235 ;
        RECT -15.125 -55.925 -14.795 -55.595 ;
        RECT -15.125 -57.285 -14.795 -56.955 ;
        RECT -15.125 -58.645 -14.795 -58.315 ;
        RECT -15.125 -60.005 -14.795 -59.675 ;
        RECT -15.125 -61.365 -14.795 -61.035 ;
        RECT -15.125 -62.725 -14.795 -62.395 ;
        RECT -15.125 -68.165 -14.795 -67.835 ;
        RECT -15.125 -69.525 -14.795 -69.195 ;
        RECT -15.125 -70.79 -14.795 -70.46 ;
        RECT -15.125 -72.245 -14.795 -71.915 ;
        RECT -15.125 -73.605 -14.795 -73.275 ;
        RECT -15.125 -74.965 -14.795 -74.635 ;
        RECT -15.125 -76.325 -14.795 -75.995 ;
        RECT -15.125 -77.685 -14.795 -77.355 ;
        RECT -15.125 -79.045 -14.795 -78.715 ;
        RECT -15.125 -81.765 -14.795 -81.435 ;
        RECT -15.125 -83.125 -14.795 -82.795 ;
        RECT -15.125 -84.485 -14.795 -84.155 ;
        RECT -15.125 -85.845 -14.795 -85.515 ;
        RECT -15.125 -87.205 -14.795 -86.875 ;
        RECT -15.125 -88.565 -14.795 -88.235 ;
        RECT -15.125 -89.33 -14.795 -89 ;
        RECT -15.125 -91.285 -14.795 -90.955 ;
        RECT -15.125 -92.645 -14.795 -92.315 ;
        RECT -15.125 -94.005 -14.795 -93.675 ;
        RECT -15.125 -95.365 -14.795 -95.035 ;
        RECT -15.125 -96.725 -14.795 -96.395 ;
        RECT -15.125 -98.085 -14.795 -97.755 ;
        RECT -15.125 -100.805 -14.795 -100.475 ;
        RECT -15.125 -102.165 -14.795 -101.835 ;
        RECT -15.125 -103.525 -14.795 -103.195 ;
        RECT -15.125 -106.245 -14.795 -105.915 ;
        RECT -15.125 -107.605 -14.795 -107.275 ;
        RECT -15.125 -108.965 -14.795 -108.635 ;
        RECT -15.125 -110.325 -14.795 -109.995 ;
        RECT -15.125 -111.685 -14.795 -111.355 ;
        RECT -15.125 -113.045 -14.795 -112.715 ;
        RECT -15.125 -114.97 -14.795 -114.64 ;
        RECT -15.125 -115.765 -14.795 -115.435 ;
        RECT -15.125 -117.125 -14.795 -116.795 ;
        RECT -15.125 -118.485 -14.795 -118.155 ;
        RECT -15.125 -119.845 -14.795 -119.515 ;
        RECT -15.125 -121.205 -14.795 -120.875 ;
        RECT -15.125 -122.565 -14.795 -122.235 ;
        RECT -15.125 -125.285 -14.795 -124.955 ;
        RECT -15.125 -126.645 -14.795 -126.315 ;
        RECT -15.125 -128.005 -14.795 -127.675 ;
        RECT -15.125 -129.365 -14.795 -129.035 ;
        RECT -15.125 -130.725 -14.795 -130.395 ;
        RECT -15.125 -132.085 -14.795 -131.755 ;
        RECT -15.125 -133.51 -14.795 -133.18 ;
        RECT -15.125 -138.885 -14.795 -138.555 ;
        RECT -15.125 -140.245 -14.795 -139.915 ;
        RECT -15.125 -141.605 -14.795 -141.275 ;
        RECT -15.125 -144.325 -14.795 -143.995 ;
        RECT -15.125 -145.685 -14.795 -145.355 ;
        RECT -15.125 -147.045 -14.795 -146.715 ;
        RECT -15.125 -152.485 -14.795 -152.155 ;
        RECT -15.125 -153.845 -14.795 -153.515 ;
        RECT -15.125 -155.205 -14.795 -154.875 ;
        RECT -15.125 -156.565 -14.795 -156.235 ;
        RECT -15.125 -157.925 -14.795 -157.595 ;
        RECT -15.125 -164.725 -14.795 -164.395 ;
        RECT -15.125 -167.445 -14.795 -167.115 ;
        RECT -15.125 -168.805 -14.795 -168.475 ;
        RECT -15.125 -170.165 -14.795 -169.835 ;
        RECT -15.125 -171.525 -14.795 -171.195 ;
        RECT -15.125 -175.605 -14.795 -175.275 ;
        RECT -15.125 -176.965 -14.795 -176.635 ;
        RECT -15.125 -178.325 -14.795 -177.995 ;
        RECT -15.125 -179.685 -14.795 -179.355 ;
        RECT -15.125 -181.045 -14.795 -180.715 ;
        RECT -15.125 -182.405 -14.795 -182.075 ;
        RECT -15.125 -185.125 -14.795 -184.795 ;
        RECT -15.125 -189.205 -14.795 -188.875 ;
        RECT -15.125 -190.565 -14.795 -190.235 ;
        RECT -15.125 -194.645 -14.795 -194.315 ;
        RECT -15.125 -196.005 -14.795 -195.675 ;
        RECT -15.125 -198.725 -14.795 -198.395 ;
        RECT -15.125 -202.805 -14.795 -202.475 ;
        RECT -15.125 -204.165 -14.795 -203.835 ;
        RECT -15.125 -209.605 -14.795 -209.275 ;
        RECT -15.125 -213.685 -14.795 -213.355 ;
        RECT -15.125 -215.045 -14.795 -214.715 ;
        RECT -15.125 -216.405 -14.795 -216.075 ;
        RECT -15.125 -217.765 -14.795 -217.435 ;
        RECT -15.125 -219.125 -14.795 -218.795 ;
        RECT -15.125 -220.485 -14.795 -220.155 ;
        RECT -15.125 -221.845 -14.795 -221.515 ;
        RECT -15.125 -223.205 -14.795 -222.875 ;
        RECT -15.125 -224.565 -14.795 -224.235 ;
        RECT -15.125 -226.155 -14.795 -225.825 ;
        RECT -15.125 -227.285 -14.795 -226.955 ;
        RECT -15.125 -228.645 -14.795 -228.315 ;
        RECT -15.125 -231.365 -14.795 -231.035 ;
        RECT -15.125 -234.085 -14.795 -233.755 ;
        RECT -15.125 -235.445 -14.795 -235.115 ;
        RECT -15.125 -236.805 -14.795 -236.475 ;
        RECT -15.125 -238.165 -14.795 -237.835 ;
        RECT -15.125 -243.81 -14.795 -242.68 ;
        RECT -15.12 -243.925 -14.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 246.76 -13.435 247.89 ;
        RECT -13.765 241.915 -13.435 242.245 ;
        RECT -13.765 240.555 -13.435 240.885 ;
        RECT -13.765 239.195 -13.435 239.525 ;
        RECT -13.765 237.835 -13.435 238.165 ;
        RECT -13.765 236.475 -13.435 236.805 ;
        RECT -13.765 235.115 -13.435 235.445 ;
        RECT -13.765 233.755 -13.435 234.085 ;
        RECT -13.765 232.395 -13.435 232.725 ;
        RECT -13.765 231.035 -13.435 231.365 ;
        RECT -13.765 229.675 -13.435 230.005 ;
        RECT -13.765 228.315 -13.435 228.645 ;
        RECT -13.765 226.955 -13.435 227.285 ;
        RECT -13.765 225.595 -13.435 225.925 ;
        RECT -13.765 224.235 -13.435 224.565 ;
        RECT -13.765 222.875 -13.435 223.205 ;
        RECT -13.765 221.515 -13.435 221.845 ;
        RECT -13.765 220.155 -13.435 220.485 ;
        RECT -13.765 218.795 -13.435 219.125 ;
        RECT -13.765 217.435 -13.435 217.765 ;
        RECT -13.765 216.075 -13.435 216.405 ;
        RECT -13.765 214.715 -13.435 215.045 ;
        RECT -13.765 213.355 -13.435 213.685 ;
        RECT -13.765 211.995 -13.435 212.325 ;
        RECT -13.765 210.635 -13.435 210.965 ;
        RECT -13.765 209.275 -13.435 209.605 ;
        RECT -13.765 207.915 -13.435 208.245 ;
        RECT -13.765 206.555 -13.435 206.885 ;
        RECT -13.765 205.195 -13.435 205.525 ;
        RECT -13.765 203.835 -13.435 204.165 ;
        RECT -13.765 202.475 -13.435 202.805 ;
        RECT -13.765 201.115 -13.435 201.445 ;
        RECT -13.765 199.755 -13.435 200.085 ;
        RECT -13.765 198.395 -13.435 198.725 ;
        RECT -13.765 197.035 -13.435 197.365 ;
        RECT -13.765 195.675 -13.435 196.005 ;
        RECT -13.765 194.315 -13.435 194.645 ;
        RECT -13.765 192.955 -13.435 193.285 ;
        RECT -13.765 191.595 -13.435 191.925 ;
        RECT -13.765 190.235 -13.435 190.565 ;
        RECT -13.765 188.875 -13.435 189.205 ;
        RECT -13.765 187.515 -13.435 187.845 ;
        RECT -13.765 186.155 -13.435 186.485 ;
        RECT -13.765 184.795 -13.435 185.125 ;
        RECT -13.765 183.435 -13.435 183.765 ;
        RECT -13.765 182.075 -13.435 182.405 ;
        RECT -13.765 180.715 -13.435 181.045 ;
        RECT -13.765 179.355 -13.435 179.685 ;
        RECT -13.765 177.995 -13.435 178.325 ;
        RECT -13.765 176.635 -13.435 176.965 ;
        RECT -13.765 175.275 -13.435 175.605 ;
        RECT -13.765 173.915 -13.435 174.245 ;
        RECT -13.765 172.555 -13.435 172.885 ;
        RECT -13.765 171.195 -13.435 171.525 ;
        RECT -13.765 169.835 -13.435 170.165 ;
        RECT -13.765 168.475 -13.435 168.805 ;
        RECT -13.765 167.115 -13.435 167.445 ;
        RECT -13.765 165.755 -13.435 166.085 ;
        RECT -13.765 164.395 -13.435 164.725 ;
        RECT -13.765 163.035 -13.435 163.365 ;
        RECT -13.765 161.675 -13.435 162.005 ;
        RECT -13.765 160.315 -13.435 160.645 ;
        RECT -13.765 158.955 -13.435 159.285 ;
        RECT -13.765 157.595 -13.435 157.925 ;
        RECT -13.765 156.235 -13.435 156.565 ;
        RECT -13.765 154.875 -13.435 155.205 ;
        RECT -13.765 153.515 -13.435 153.845 ;
        RECT -13.765 152.155 -13.435 152.485 ;
        RECT -13.765 150.795 -13.435 151.125 ;
        RECT -13.765 149.435 -13.435 149.765 ;
        RECT -13.765 148.075 -13.435 148.405 ;
        RECT -13.765 146.715 -13.435 147.045 ;
        RECT -13.765 145.355 -13.435 145.685 ;
        RECT -13.765 143.995 -13.435 144.325 ;
        RECT -13.765 142.635 -13.435 142.965 ;
        RECT -13.765 141.275 -13.435 141.605 ;
        RECT -13.765 139.915 -13.435 140.245 ;
        RECT -13.765 138.555 -13.435 138.885 ;
        RECT -13.765 137.195 -13.435 137.525 ;
        RECT -13.765 135.835 -13.435 136.165 ;
        RECT -13.765 134.475 -13.435 134.805 ;
        RECT -13.765 133.115 -13.435 133.445 ;
        RECT -13.765 131.755 -13.435 132.085 ;
        RECT -13.765 130.395 -13.435 130.725 ;
        RECT -13.765 129.035 -13.435 129.365 ;
        RECT -13.765 127.675 -13.435 128.005 ;
        RECT -13.765 126.315 -13.435 126.645 ;
        RECT -13.765 124.955 -13.435 125.285 ;
        RECT -13.765 123.595 -13.435 123.925 ;
        RECT -13.765 122.235 -13.435 122.565 ;
        RECT -13.765 120.875 -13.435 121.205 ;
        RECT -13.765 119.515 -13.435 119.845 ;
        RECT -13.765 118.155 -13.435 118.485 ;
        RECT -13.765 116.795 -13.435 117.125 ;
        RECT -13.765 115.435 -13.435 115.765 ;
        RECT -13.765 114.075 -13.435 114.405 ;
        RECT -13.765 112.715 -13.435 113.045 ;
        RECT -13.765 111.355 -13.435 111.685 ;
        RECT -13.765 109.995 -13.435 110.325 ;
        RECT -13.765 108.635 -13.435 108.965 ;
        RECT -13.765 107.275 -13.435 107.605 ;
        RECT -13.765 105.915 -13.435 106.245 ;
        RECT -13.765 104.555 -13.435 104.885 ;
        RECT -13.765 103.195 -13.435 103.525 ;
        RECT -13.765 101.835 -13.435 102.165 ;
        RECT -13.765 100.475 -13.435 100.805 ;
        RECT -13.765 99.115 -13.435 99.445 ;
        RECT -13.765 97.755 -13.435 98.085 ;
        RECT -13.765 96.395 -13.435 96.725 ;
        RECT -13.765 95.035 -13.435 95.365 ;
        RECT -13.765 93.675 -13.435 94.005 ;
        RECT -13.765 92.315 -13.435 92.645 ;
        RECT -13.765 90.955 -13.435 91.285 ;
        RECT -13.765 89.595 -13.435 89.925 ;
        RECT -13.765 88.235 -13.435 88.565 ;
        RECT -13.765 86.875 -13.435 87.205 ;
        RECT -13.765 85.515 -13.435 85.845 ;
        RECT -13.765 84.155 -13.435 84.485 ;
        RECT -13.765 82.795 -13.435 83.125 ;
        RECT -13.765 81.435 -13.435 81.765 ;
        RECT -13.765 80.075 -13.435 80.405 ;
        RECT -13.765 78.715 -13.435 79.045 ;
        RECT -13.765 77.355 -13.435 77.685 ;
        RECT -13.765 75.995 -13.435 76.325 ;
        RECT -13.765 74.635 -13.435 74.965 ;
        RECT -13.765 73.275 -13.435 73.605 ;
        RECT -13.765 71.915 -13.435 72.245 ;
        RECT -13.765 70.555 -13.435 70.885 ;
        RECT -13.765 69.195 -13.435 69.525 ;
        RECT -13.765 67.835 -13.435 68.165 ;
        RECT -13.765 66.475 -13.435 66.805 ;
        RECT -13.765 65.115 -13.435 65.445 ;
        RECT -13.765 63.755 -13.435 64.085 ;
        RECT -13.765 62.395 -13.435 62.725 ;
        RECT -13.765 61.035 -13.435 61.365 ;
        RECT -13.765 59.675 -13.435 60.005 ;
        RECT -13.765 58.315 -13.435 58.645 ;
        RECT -13.765 56.955 -13.435 57.285 ;
        RECT -13.765 55.595 -13.435 55.925 ;
        RECT -13.765 54.235 -13.435 54.565 ;
        RECT -13.765 52.875 -13.435 53.205 ;
        RECT -13.765 51.515 -13.435 51.845 ;
        RECT -13.765 50.155 -13.435 50.485 ;
        RECT -13.765 48.795 -13.435 49.125 ;
        RECT -13.765 47.435 -13.435 47.765 ;
        RECT -13.765 46.075 -13.435 46.405 ;
        RECT -13.765 44.715 -13.435 45.045 ;
        RECT -13.765 43.355 -13.435 43.685 ;
        RECT -13.765 41.995 -13.435 42.325 ;
        RECT -13.765 40.635 -13.435 40.965 ;
        RECT -13.765 39.275 -13.435 39.605 ;
        RECT -13.765 37.915 -13.435 38.245 ;
        RECT -13.765 36.555 -13.435 36.885 ;
        RECT -13.765 35.195 -13.435 35.525 ;
        RECT -13.765 33.835 -13.435 34.165 ;
        RECT -13.765 32.475 -13.435 32.805 ;
        RECT -13.765 31.115 -13.435 31.445 ;
        RECT -13.765 29.755 -13.435 30.085 ;
        RECT -13.765 28.395 -13.435 28.725 ;
        RECT -13.765 27.035 -13.435 27.365 ;
        RECT -13.765 25.675 -13.435 26.005 ;
        RECT -13.765 24.315 -13.435 24.645 ;
        RECT -13.765 22.955 -13.435 23.285 ;
        RECT -13.765 21.595 -13.435 21.925 ;
        RECT -13.765 20.235 -13.435 20.565 ;
        RECT -13.765 18.875 -13.435 19.205 ;
        RECT -13.765 17.515 -13.435 17.845 ;
        RECT -13.765 16.155 -13.435 16.485 ;
        RECT -13.765 14.795 -13.435 15.125 ;
        RECT -13.765 13.435 -13.435 13.765 ;
        RECT -13.765 12.075 -13.435 12.405 ;
        RECT -13.765 10.715 -13.435 11.045 ;
        RECT -13.765 9.355 -13.435 9.685 ;
        RECT -13.765 7.995 -13.435 8.325 ;
        RECT -13.765 6.635 -13.435 6.965 ;
        RECT -13.765 5.275 -13.435 5.605 ;
        RECT -13.765 3.915 -13.435 4.245 ;
        RECT -13.765 2.555 -13.435 2.885 ;
        RECT -13.765 1.195 -13.435 1.525 ;
        RECT -13.765 -0.165 -13.435 0.165 ;
        RECT -13.765 -1.525 -13.435 -1.195 ;
        RECT -13.765 -2.885 -13.435 -2.555 ;
        RECT -13.765 -4.245 -13.435 -3.915 ;
        RECT -13.765 -5.605 -13.435 -5.275 ;
        RECT -13.765 -6.965 -13.435 -6.635 ;
        RECT -13.765 -8.325 -13.435 -7.995 ;
        RECT -13.765 -9.48 -13.435 -9.15 ;
        RECT -13.765 -12.405 -13.435 -12.075 ;
        RECT -13.765 -15.125 -13.435 -14.795 ;
        RECT -13.765 -16.67 -13.435 -16.34 ;
        RECT -13.765 -17.845 -13.435 -17.515 ;
        RECT -13.765 -24.645 -13.435 -24.315 ;
        RECT -13.765 -26.005 -13.435 -25.675 ;
        RECT -13.765 -27.365 -13.435 -27.035 ;
        RECT -13.765 -30.66 -13.435 -30.33 ;
        RECT -13.765 -31.445 -13.435 -31.115 ;
        RECT -13.765 -32.805 -13.435 -32.475 ;
        RECT -13.765 -34.165 -13.435 -33.835 ;
        RECT -13.765 -36.885 -13.435 -36.555 ;
        RECT -13.765 -37.85 -13.435 -37.52 ;
        RECT -13.765 -40.965 -13.435 -40.635 ;
        RECT -13.765 -46.405 -13.435 -46.075 ;
        RECT -13.765 -47.765 -13.435 -47.435 ;
        RECT -13.765 -49.125 -13.435 -48.795 ;
        RECT -13.765 -50.485 -13.435 -50.155 ;
        RECT -13.765 -51.845 -13.435 -51.515 ;
        RECT -13.765 -53.205 -13.435 -52.875 ;
        RECT -13.765 -54.565 -13.435 -54.235 ;
        RECT -13.765 -55.925 -13.435 -55.595 ;
        RECT -13.765 -57.285 -13.435 -56.955 ;
        RECT -13.765 -58.645 -13.435 -58.315 ;
        RECT -13.765 -60.005 -13.435 -59.675 ;
        RECT -13.765 -61.365 -13.435 -61.035 ;
        RECT -13.765 -62.725 -13.435 -62.395 ;
        RECT -13.765 -68.165 -13.435 -67.835 ;
        RECT -13.765 -69.525 -13.435 -69.195 ;
        RECT -13.765 -70.79 -13.435 -70.46 ;
        RECT -13.765 -72.245 -13.435 -71.915 ;
        RECT -13.765 -73.605 -13.435 -73.275 ;
        RECT -13.765 -74.965 -13.435 -74.635 ;
        RECT -13.765 -76.325 -13.435 -75.995 ;
        RECT -13.765 -77.685 -13.435 -77.355 ;
        RECT -13.765 -79.045 -13.435 -78.715 ;
        RECT -13.765 -81.765 -13.435 -81.435 ;
        RECT -13.765 -83.125 -13.435 -82.795 ;
        RECT -13.765 -84.485 -13.435 -84.155 ;
        RECT -13.765 -85.845 -13.435 -85.515 ;
        RECT -13.765 -87.205 -13.435 -86.875 ;
        RECT -13.765 -88.565 -13.435 -88.235 ;
        RECT -13.765 -89.33 -13.435 -89 ;
        RECT -13.765 -91.285 -13.435 -90.955 ;
        RECT -13.765 -92.645 -13.435 -92.315 ;
        RECT -13.765 -94.005 -13.435 -93.675 ;
        RECT -13.765 -95.365 -13.435 -95.035 ;
        RECT -13.765 -96.725 -13.435 -96.395 ;
        RECT -13.765 -98.085 -13.435 -97.755 ;
        RECT -13.765 -100.805 -13.435 -100.475 ;
        RECT -13.765 -102.165 -13.435 -101.835 ;
        RECT -13.765 -103.525 -13.435 -103.195 ;
        RECT -13.765 -106.245 -13.435 -105.915 ;
        RECT -13.765 -107.605 -13.435 -107.275 ;
        RECT -13.765 -108.965 -13.435 -108.635 ;
        RECT -13.765 -110.325 -13.435 -109.995 ;
        RECT -13.765 -111.685 -13.435 -111.355 ;
        RECT -13.765 -113.045 -13.435 -112.715 ;
        RECT -13.765 -114.97 -13.435 -114.64 ;
        RECT -13.765 -115.765 -13.435 -115.435 ;
        RECT -13.765 -117.125 -13.435 -116.795 ;
        RECT -13.765 -118.485 -13.435 -118.155 ;
        RECT -13.765 -119.845 -13.435 -119.515 ;
        RECT -13.765 -121.205 -13.435 -120.875 ;
        RECT -13.765 -122.565 -13.435 -122.235 ;
        RECT -13.765 -125.285 -13.435 -124.955 ;
        RECT -13.765 -126.645 -13.435 -126.315 ;
        RECT -13.765 -128.005 -13.435 -127.675 ;
        RECT -13.765 -129.365 -13.435 -129.035 ;
        RECT -13.765 -130.725 -13.435 -130.395 ;
        RECT -13.765 -132.085 -13.435 -131.755 ;
        RECT -13.765 -133.51 -13.435 -133.18 ;
        RECT -13.765 -140.245 -13.435 -139.915 ;
        RECT -13.765 -141.605 -13.435 -141.275 ;
        RECT -13.765 -144.325 -13.435 -143.995 ;
        RECT -13.765 -145.685 -13.435 -145.355 ;
        RECT -13.765 -147.045 -13.435 -146.715 ;
        RECT -13.765 -152.485 -13.435 -152.155 ;
        RECT -13.765 -153.845 -13.435 -153.515 ;
        RECT -13.765 -155.205 -13.435 -154.875 ;
        RECT -13.765 -156.565 -13.435 -156.235 ;
        RECT -13.765 -157.925 -13.435 -157.595 ;
        RECT -13.765 -160.645 -13.435 -160.315 ;
        RECT -13.765 -164.725 -13.435 -164.395 ;
        RECT -13.765 -167.445 -13.435 -167.115 ;
        RECT -13.765 -168.805 -13.435 -168.475 ;
        RECT -13.765 -175.605 -13.435 -175.275 ;
        RECT -13.765 -176.965 -13.435 -176.635 ;
        RECT -13.765 -178.325 -13.435 -177.995 ;
        RECT -13.765 -179.685 -13.435 -179.355 ;
        RECT -13.765 -181.045 -13.435 -180.715 ;
        RECT -13.765 -182.405 -13.435 -182.075 ;
        RECT -13.765 -189.205 -13.435 -188.875 ;
        RECT -13.765 -190.565 -13.435 -190.235 ;
        RECT -13.765 -191.925 -13.435 -191.595 ;
        RECT -13.765 -194.645 -13.435 -194.315 ;
        RECT -13.765 -196.005 -13.435 -195.675 ;
        RECT -13.765 -197.365 -13.435 -197.035 ;
        RECT -13.765 -198.725 -13.435 -198.395 ;
        RECT -13.765 -204.165 -13.435 -203.835 ;
        RECT -13.765 -206.885 -13.435 -206.555 ;
        RECT -13.765 -209.605 -13.435 -209.275 ;
        RECT -13.765 -213.685 -13.435 -213.355 ;
        RECT -13.765 -215.045 -13.435 -214.715 ;
        RECT -13.765 -216.405 -13.435 -216.075 ;
        RECT -13.765 -217.765 -13.435 -217.435 ;
        RECT -13.765 -219.125 -13.435 -218.795 ;
        RECT -13.765 -220.485 -13.435 -220.155 ;
        RECT -13.765 -221.845 -13.435 -221.515 ;
        RECT -13.765 -223.205 -13.435 -222.875 ;
        RECT -13.765 -224.565 -13.435 -224.235 ;
        RECT -13.765 -226.155 -13.435 -225.825 ;
        RECT -13.765 -227.285 -13.435 -226.955 ;
        RECT -13.765 -228.645 -13.435 -228.315 ;
        RECT -13.765 -230.005 -13.435 -229.675 ;
        RECT -13.765 -231.365 -13.435 -231.035 ;
        RECT -13.765 -234.085 -13.435 -233.755 ;
        RECT -13.765 -235.445 -13.435 -235.115 ;
        RECT -13.765 -236.805 -13.435 -236.475 ;
        RECT -13.765 -238.165 -13.435 -237.835 ;
        RECT -13.765 -243.81 -13.435 -242.68 ;
        RECT -13.76 -243.925 -13.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 246.76 -12.075 247.89 ;
        RECT -12.405 241.915 -12.075 242.245 ;
        RECT -12.405 240.555 -12.075 240.885 ;
        RECT -12.405 239.195 -12.075 239.525 ;
        RECT -12.405 237.835 -12.075 238.165 ;
        RECT -12.405 236.475 -12.075 236.805 ;
        RECT -12.405 235.115 -12.075 235.445 ;
        RECT -12.405 233.755 -12.075 234.085 ;
        RECT -12.405 232.395 -12.075 232.725 ;
        RECT -12.405 231.035 -12.075 231.365 ;
        RECT -12.405 229.675 -12.075 230.005 ;
        RECT -12.405 228.315 -12.075 228.645 ;
        RECT -12.405 226.955 -12.075 227.285 ;
        RECT -12.405 225.595 -12.075 225.925 ;
        RECT -12.405 224.235 -12.075 224.565 ;
        RECT -12.405 222.875 -12.075 223.205 ;
        RECT -12.405 221.515 -12.075 221.845 ;
        RECT -12.405 220.155 -12.075 220.485 ;
        RECT -12.405 218.795 -12.075 219.125 ;
        RECT -12.405 217.435 -12.075 217.765 ;
        RECT -12.405 216.075 -12.075 216.405 ;
        RECT -12.405 214.715 -12.075 215.045 ;
        RECT -12.405 213.355 -12.075 213.685 ;
        RECT -12.405 211.995 -12.075 212.325 ;
        RECT -12.405 210.635 -12.075 210.965 ;
        RECT -12.405 209.275 -12.075 209.605 ;
        RECT -12.405 207.915 -12.075 208.245 ;
        RECT -12.405 206.555 -12.075 206.885 ;
        RECT -12.405 205.195 -12.075 205.525 ;
        RECT -12.405 203.835 -12.075 204.165 ;
        RECT -12.405 202.475 -12.075 202.805 ;
        RECT -12.405 201.115 -12.075 201.445 ;
        RECT -12.405 199.755 -12.075 200.085 ;
        RECT -12.405 198.395 -12.075 198.725 ;
        RECT -12.405 197.035 -12.075 197.365 ;
        RECT -12.405 195.675 -12.075 196.005 ;
        RECT -12.405 194.315 -12.075 194.645 ;
        RECT -12.405 192.955 -12.075 193.285 ;
        RECT -12.405 191.595 -12.075 191.925 ;
        RECT -12.405 190.235 -12.075 190.565 ;
        RECT -12.405 188.875 -12.075 189.205 ;
        RECT -12.405 187.515 -12.075 187.845 ;
        RECT -12.405 186.155 -12.075 186.485 ;
        RECT -12.405 184.795 -12.075 185.125 ;
        RECT -12.405 183.435 -12.075 183.765 ;
        RECT -12.405 182.075 -12.075 182.405 ;
        RECT -12.405 180.715 -12.075 181.045 ;
        RECT -12.405 179.355 -12.075 179.685 ;
        RECT -12.405 177.995 -12.075 178.325 ;
        RECT -12.405 176.635 -12.075 176.965 ;
        RECT -12.405 175.275 -12.075 175.605 ;
        RECT -12.405 173.915 -12.075 174.245 ;
        RECT -12.405 172.555 -12.075 172.885 ;
        RECT -12.405 171.195 -12.075 171.525 ;
        RECT -12.405 169.835 -12.075 170.165 ;
        RECT -12.405 168.475 -12.075 168.805 ;
        RECT -12.405 167.115 -12.075 167.445 ;
        RECT -12.405 165.755 -12.075 166.085 ;
        RECT -12.405 164.395 -12.075 164.725 ;
        RECT -12.405 163.035 -12.075 163.365 ;
        RECT -12.405 161.675 -12.075 162.005 ;
        RECT -12.405 160.315 -12.075 160.645 ;
        RECT -12.405 158.955 -12.075 159.285 ;
        RECT -12.405 157.595 -12.075 157.925 ;
        RECT -12.405 156.235 -12.075 156.565 ;
        RECT -12.405 154.875 -12.075 155.205 ;
        RECT -12.405 153.515 -12.075 153.845 ;
        RECT -12.405 152.155 -12.075 152.485 ;
        RECT -12.405 150.795 -12.075 151.125 ;
        RECT -12.405 149.435 -12.075 149.765 ;
        RECT -12.405 148.075 -12.075 148.405 ;
        RECT -12.405 146.715 -12.075 147.045 ;
        RECT -12.405 145.355 -12.075 145.685 ;
        RECT -12.405 143.995 -12.075 144.325 ;
        RECT -12.405 142.635 -12.075 142.965 ;
        RECT -12.405 141.275 -12.075 141.605 ;
        RECT -12.405 139.915 -12.075 140.245 ;
        RECT -12.405 138.555 -12.075 138.885 ;
        RECT -12.405 137.195 -12.075 137.525 ;
        RECT -12.405 135.835 -12.075 136.165 ;
        RECT -12.405 134.475 -12.075 134.805 ;
        RECT -12.405 133.115 -12.075 133.445 ;
        RECT -12.405 131.755 -12.075 132.085 ;
        RECT -12.405 130.395 -12.075 130.725 ;
        RECT -12.405 129.035 -12.075 129.365 ;
        RECT -12.405 127.675 -12.075 128.005 ;
        RECT -12.405 126.315 -12.075 126.645 ;
        RECT -12.405 124.955 -12.075 125.285 ;
        RECT -12.405 123.595 -12.075 123.925 ;
        RECT -12.405 122.235 -12.075 122.565 ;
        RECT -12.405 120.875 -12.075 121.205 ;
        RECT -12.405 119.515 -12.075 119.845 ;
        RECT -12.405 118.155 -12.075 118.485 ;
        RECT -12.405 116.795 -12.075 117.125 ;
        RECT -12.405 115.435 -12.075 115.765 ;
        RECT -12.405 114.075 -12.075 114.405 ;
        RECT -12.405 112.715 -12.075 113.045 ;
        RECT -12.405 111.355 -12.075 111.685 ;
        RECT -12.405 109.995 -12.075 110.325 ;
        RECT -12.405 108.635 -12.075 108.965 ;
        RECT -12.405 107.275 -12.075 107.605 ;
        RECT -12.405 105.915 -12.075 106.245 ;
        RECT -12.405 104.555 -12.075 104.885 ;
        RECT -12.405 103.195 -12.075 103.525 ;
        RECT -12.405 101.835 -12.075 102.165 ;
        RECT -12.405 100.475 -12.075 100.805 ;
        RECT -12.405 99.115 -12.075 99.445 ;
        RECT -12.405 97.755 -12.075 98.085 ;
        RECT -12.405 96.395 -12.075 96.725 ;
        RECT -12.405 95.035 -12.075 95.365 ;
        RECT -12.405 93.675 -12.075 94.005 ;
        RECT -12.405 92.315 -12.075 92.645 ;
        RECT -12.405 90.955 -12.075 91.285 ;
        RECT -12.405 89.595 -12.075 89.925 ;
        RECT -12.405 88.235 -12.075 88.565 ;
        RECT -12.405 86.875 -12.075 87.205 ;
        RECT -12.405 85.515 -12.075 85.845 ;
        RECT -12.405 84.155 -12.075 84.485 ;
        RECT -12.405 82.795 -12.075 83.125 ;
        RECT -12.405 81.435 -12.075 81.765 ;
        RECT -12.405 80.075 -12.075 80.405 ;
        RECT -12.405 78.715 -12.075 79.045 ;
        RECT -12.405 77.355 -12.075 77.685 ;
        RECT -12.405 75.995 -12.075 76.325 ;
        RECT -12.405 74.635 -12.075 74.965 ;
        RECT -12.405 73.275 -12.075 73.605 ;
        RECT -12.405 71.915 -12.075 72.245 ;
        RECT -12.405 70.555 -12.075 70.885 ;
        RECT -12.405 69.195 -12.075 69.525 ;
        RECT -12.405 67.835 -12.075 68.165 ;
        RECT -12.405 66.475 -12.075 66.805 ;
        RECT -12.405 65.115 -12.075 65.445 ;
        RECT -12.405 63.755 -12.075 64.085 ;
        RECT -12.405 62.395 -12.075 62.725 ;
        RECT -12.405 61.035 -12.075 61.365 ;
        RECT -12.405 59.675 -12.075 60.005 ;
        RECT -12.405 58.315 -12.075 58.645 ;
        RECT -12.405 56.955 -12.075 57.285 ;
        RECT -12.405 55.595 -12.075 55.925 ;
        RECT -12.405 54.235 -12.075 54.565 ;
        RECT -12.405 52.875 -12.075 53.205 ;
        RECT -12.405 51.515 -12.075 51.845 ;
        RECT -12.405 50.155 -12.075 50.485 ;
        RECT -12.405 48.795 -12.075 49.125 ;
        RECT -12.405 47.435 -12.075 47.765 ;
        RECT -12.405 46.075 -12.075 46.405 ;
        RECT -12.405 44.715 -12.075 45.045 ;
        RECT -12.405 43.355 -12.075 43.685 ;
        RECT -12.405 41.995 -12.075 42.325 ;
        RECT -12.405 40.635 -12.075 40.965 ;
        RECT -12.405 39.275 -12.075 39.605 ;
        RECT -12.405 37.915 -12.075 38.245 ;
        RECT -12.405 36.555 -12.075 36.885 ;
        RECT -12.405 35.195 -12.075 35.525 ;
        RECT -12.405 33.835 -12.075 34.165 ;
        RECT -12.405 32.475 -12.075 32.805 ;
        RECT -12.405 31.115 -12.075 31.445 ;
        RECT -12.405 29.755 -12.075 30.085 ;
        RECT -12.405 28.395 -12.075 28.725 ;
        RECT -12.405 27.035 -12.075 27.365 ;
        RECT -12.405 25.675 -12.075 26.005 ;
        RECT -12.405 24.315 -12.075 24.645 ;
        RECT -12.405 22.955 -12.075 23.285 ;
        RECT -12.405 21.595 -12.075 21.925 ;
        RECT -12.405 20.235 -12.075 20.565 ;
        RECT -12.405 18.875 -12.075 19.205 ;
        RECT -12.405 17.515 -12.075 17.845 ;
        RECT -12.405 16.155 -12.075 16.485 ;
        RECT -12.405 14.795 -12.075 15.125 ;
        RECT -12.405 13.435 -12.075 13.765 ;
        RECT -12.405 12.075 -12.075 12.405 ;
        RECT -12.405 10.715 -12.075 11.045 ;
        RECT -12.405 9.355 -12.075 9.685 ;
        RECT -12.405 7.995 -12.075 8.325 ;
        RECT -12.405 6.635 -12.075 6.965 ;
        RECT -12.405 5.275 -12.075 5.605 ;
        RECT -12.405 3.915 -12.075 4.245 ;
        RECT -12.405 2.555 -12.075 2.885 ;
        RECT -12.405 1.195 -12.075 1.525 ;
        RECT -12.405 -0.165 -12.075 0.165 ;
        RECT -12.405 -1.525 -12.075 -1.195 ;
        RECT -12.405 -2.885 -12.075 -2.555 ;
        RECT -12.405 -4.245 -12.075 -3.915 ;
        RECT -12.405 -5.605 -12.075 -5.275 ;
        RECT -12.405 -6.965 -12.075 -6.635 ;
        RECT -12.405 -8.325 -12.075 -7.995 ;
        RECT -12.405 -9.48 -12.075 -9.15 ;
        RECT -12.4 -10.36 -12.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 -183.765 -12.075 -183.435 ;
        RECT -12.405 -186.485 -12.075 -186.155 ;
        RECT -12.405 -189.205 -12.075 -188.875 ;
        RECT -12.405 -190.565 -12.075 -190.235 ;
        RECT -12.405 -191.925 -12.075 -191.595 ;
        RECT -12.405 -193.285 -12.075 -192.955 ;
        RECT -12.405 -194.645 -12.075 -194.315 ;
        RECT -12.405 -196.005 -12.075 -195.675 ;
        RECT -12.405 -197.365 -12.075 -197.035 ;
        RECT -12.405 -198.725 -12.075 -198.395 ;
        RECT -12.405 -201.445 -12.075 -201.115 ;
        RECT -12.405 -204.165 -12.075 -203.835 ;
        RECT -12.405 -205.525 -12.075 -205.195 ;
        RECT -12.405 -206.885 -12.075 -206.555 ;
        RECT -12.405 -208.245 -12.075 -207.915 ;
        RECT -12.405 -209.605 -12.075 -209.275 ;
        RECT -12.405 -210.965 -12.075 -210.635 ;
        RECT -12.405 -212.325 -12.075 -211.995 ;
        RECT -12.405 -213.685 -12.075 -213.355 ;
        RECT -12.405 -215.045 -12.075 -214.715 ;
        RECT -12.405 -216.405 -12.075 -216.075 ;
        RECT -12.405 -217.765 -12.075 -217.435 ;
        RECT -12.405 -219.125 -12.075 -218.795 ;
        RECT -12.405 -220.485 -12.075 -220.155 ;
        RECT -12.405 -221.845 -12.075 -221.515 ;
        RECT -12.405 -223.205 -12.075 -222.875 ;
        RECT -12.405 -226.155 -12.075 -225.825 ;
        RECT -12.405 -227.285 -12.075 -226.955 ;
        RECT -12.405 -228.645 -12.075 -228.315 ;
        RECT -12.405 -230.005 -12.075 -229.675 ;
        RECT -12.405 -231.365 -12.075 -231.035 ;
        RECT -12.405 -234.085 -12.075 -233.755 ;
        RECT -12.405 -235.445 -12.075 -235.115 ;
        RECT -12.405 -236.805 -12.075 -236.475 ;
        RECT -12.405 -238.165 -12.075 -237.835 ;
        RECT -12.405 -243.81 -12.075 -242.68 ;
        RECT -12.4 -243.925 -12.08 -161.68 ;
        RECT -12.405 -164.725 -12.075 -164.395 ;
        RECT -12.405 -167.445 -12.075 -167.115 ;
        RECT -12.405 -174.245 -12.075 -173.915 ;
        RECT -12.405 -175.605 -12.075 -175.275 ;
        RECT -12.405 -176.965 -12.075 -176.635 ;
        RECT -12.405 -178.325 -12.075 -177.995 ;
        RECT -12.405 -179.685 -12.075 -179.355 ;
        RECT -12.405 -181.045 -12.075 -180.715 ;
        RECT -12.405 -182.405 -12.075 -182.075 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 -129.365 -21.595 -129.035 ;
        RECT -21.925 -130.725 -21.595 -130.395 ;
        RECT -21.925 -132.085 -21.595 -131.755 ;
        RECT -21.925 -133.51 -21.595 -133.18 ;
        RECT -21.925 -137.525 -21.595 -137.195 ;
        RECT -21.925 -138.885 -21.595 -138.555 ;
        RECT -21.925 -140.245 -21.595 -139.915 ;
        RECT -21.925 -141.605 -21.595 -141.275 ;
        RECT -21.925 -144.325 -21.595 -143.995 ;
        RECT -21.925 -145.685 -21.595 -145.355 ;
        RECT -21.925 -147.045 -21.595 -146.715 ;
        RECT -21.92 -150.44 -21.6 -123.6 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 -226.155 -21.595 -225.825 ;
        RECT -21.92 -229.32 -21.6 -224.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 246.76 -20.235 247.89 ;
        RECT -20.565 241.915 -20.235 242.245 ;
        RECT -20.565 240.555 -20.235 240.885 ;
        RECT -20.565 239.195 -20.235 239.525 ;
        RECT -20.565 237.835 -20.235 238.165 ;
        RECT -20.565 236.475 -20.235 236.805 ;
        RECT -20.565 235.115 -20.235 235.445 ;
        RECT -20.565 233.755 -20.235 234.085 ;
        RECT -20.565 232.395 -20.235 232.725 ;
        RECT -20.565 231.035 -20.235 231.365 ;
        RECT -20.565 229.675 -20.235 230.005 ;
        RECT -20.565 228.315 -20.235 228.645 ;
        RECT -20.565 226.955 -20.235 227.285 ;
        RECT -20.565 225.595 -20.235 225.925 ;
        RECT -20.565 224.235 -20.235 224.565 ;
        RECT -20.565 222.875 -20.235 223.205 ;
        RECT -20.565 221.515 -20.235 221.845 ;
        RECT -20.565 220.155 -20.235 220.485 ;
        RECT -20.565 218.795 -20.235 219.125 ;
        RECT -20.565 217.435 -20.235 217.765 ;
        RECT -20.565 216.075 -20.235 216.405 ;
        RECT -20.565 214.715 -20.235 215.045 ;
        RECT -20.565 213.355 -20.235 213.685 ;
        RECT -20.565 211.995 -20.235 212.325 ;
        RECT -20.565 210.635 -20.235 210.965 ;
        RECT -20.565 209.275 -20.235 209.605 ;
        RECT -20.565 207.915 -20.235 208.245 ;
        RECT -20.565 206.555 -20.235 206.885 ;
        RECT -20.565 205.195 -20.235 205.525 ;
        RECT -20.565 203.835 -20.235 204.165 ;
        RECT -20.565 202.475 -20.235 202.805 ;
        RECT -20.565 201.115 -20.235 201.445 ;
        RECT -20.565 199.755 -20.235 200.085 ;
        RECT -20.565 198.395 -20.235 198.725 ;
        RECT -20.565 197.035 -20.235 197.365 ;
        RECT -20.565 195.675 -20.235 196.005 ;
        RECT -20.565 194.315 -20.235 194.645 ;
        RECT -20.565 192.955 -20.235 193.285 ;
        RECT -20.565 191.595 -20.235 191.925 ;
        RECT -20.565 190.235 -20.235 190.565 ;
        RECT -20.565 188.875 -20.235 189.205 ;
        RECT -20.565 187.515 -20.235 187.845 ;
        RECT -20.565 186.155 -20.235 186.485 ;
        RECT -20.565 184.795 -20.235 185.125 ;
        RECT -20.565 183.435 -20.235 183.765 ;
        RECT -20.565 182.075 -20.235 182.405 ;
        RECT -20.565 180.715 -20.235 181.045 ;
        RECT -20.565 179.355 -20.235 179.685 ;
        RECT -20.565 177.995 -20.235 178.325 ;
        RECT -20.565 176.635 -20.235 176.965 ;
        RECT -20.565 175.275 -20.235 175.605 ;
        RECT -20.565 173.915 -20.235 174.245 ;
        RECT -20.565 172.555 -20.235 172.885 ;
        RECT -20.565 171.195 -20.235 171.525 ;
        RECT -20.565 169.835 -20.235 170.165 ;
        RECT -20.565 168.475 -20.235 168.805 ;
        RECT -20.565 167.115 -20.235 167.445 ;
        RECT -20.565 165.755 -20.235 166.085 ;
        RECT -20.565 164.395 -20.235 164.725 ;
        RECT -20.565 163.035 -20.235 163.365 ;
        RECT -20.565 161.675 -20.235 162.005 ;
        RECT -20.565 160.315 -20.235 160.645 ;
        RECT -20.565 158.955 -20.235 159.285 ;
        RECT -20.565 157.595 -20.235 157.925 ;
        RECT -20.565 156.235 -20.235 156.565 ;
        RECT -20.565 154.875 -20.235 155.205 ;
        RECT -20.565 153.515 -20.235 153.845 ;
        RECT -20.565 152.155 -20.235 152.485 ;
        RECT -20.565 150.795 -20.235 151.125 ;
        RECT -20.565 149.435 -20.235 149.765 ;
        RECT -20.565 148.075 -20.235 148.405 ;
        RECT -20.565 146.715 -20.235 147.045 ;
        RECT -20.565 145.355 -20.235 145.685 ;
        RECT -20.565 143.995 -20.235 144.325 ;
        RECT -20.565 142.635 -20.235 142.965 ;
        RECT -20.565 141.275 -20.235 141.605 ;
        RECT -20.565 139.915 -20.235 140.245 ;
        RECT -20.565 138.555 -20.235 138.885 ;
        RECT -20.565 137.195 -20.235 137.525 ;
        RECT -20.565 135.835 -20.235 136.165 ;
        RECT -20.565 134.475 -20.235 134.805 ;
        RECT -20.565 133.115 -20.235 133.445 ;
        RECT -20.565 131.755 -20.235 132.085 ;
        RECT -20.565 130.395 -20.235 130.725 ;
        RECT -20.565 129.035 -20.235 129.365 ;
        RECT -20.565 127.675 -20.235 128.005 ;
        RECT -20.565 126.315 -20.235 126.645 ;
        RECT -20.565 124.955 -20.235 125.285 ;
        RECT -20.565 123.595 -20.235 123.925 ;
        RECT -20.565 122.235 -20.235 122.565 ;
        RECT -20.565 120.875 -20.235 121.205 ;
        RECT -20.565 119.515 -20.235 119.845 ;
        RECT -20.565 118.155 -20.235 118.485 ;
        RECT -20.565 116.795 -20.235 117.125 ;
        RECT -20.565 115.435 -20.235 115.765 ;
        RECT -20.565 114.075 -20.235 114.405 ;
        RECT -20.565 112.715 -20.235 113.045 ;
        RECT -20.565 111.355 -20.235 111.685 ;
        RECT -20.565 109.995 -20.235 110.325 ;
        RECT -20.565 108.635 -20.235 108.965 ;
        RECT -20.565 107.275 -20.235 107.605 ;
        RECT -20.565 105.915 -20.235 106.245 ;
        RECT -20.565 104.555 -20.235 104.885 ;
        RECT -20.565 103.195 -20.235 103.525 ;
        RECT -20.565 101.835 -20.235 102.165 ;
        RECT -20.565 100.475 -20.235 100.805 ;
        RECT -20.565 99.115 -20.235 99.445 ;
        RECT -20.565 97.755 -20.235 98.085 ;
        RECT -20.565 96.395 -20.235 96.725 ;
        RECT -20.565 95.035 -20.235 95.365 ;
        RECT -20.565 93.675 -20.235 94.005 ;
        RECT -20.565 92.315 -20.235 92.645 ;
        RECT -20.565 90.955 -20.235 91.285 ;
        RECT -20.565 89.595 -20.235 89.925 ;
        RECT -20.565 88.235 -20.235 88.565 ;
        RECT -20.565 86.875 -20.235 87.205 ;
        RECT -20.565 85.515 -20.235 85.845 ;
        RECT -20.565 84.155 -20.235 84.485 ;
        RECT -20.565 82.795 -20.235 83.125 ;
        RECT -20.565 81.435 -20.235 81.765 ;
        RECT -20.565 80.075 -20.235 80.405 ;
        RECT -20.565 78.715 -20.235 79.045 ;
        RECT -20.565 77.355 -20.235 77.685 ;
        RECT -20.565 75.995 -20.235 76.325 ;
        RECT -20.565 74.635 -20.235 74.965 ;
        RECT -20.565 73.275 -20.235 73.605 ;
        RECT -20.565 71.915 -20.235 72.245 ;
        RECT -20.565 70.555 -20.235 70.885 ;
        RECT -20.565 69.195 -20.235 69.525 ;
        RECT -20.565 67.835 -20.235 68.165 ;
        RECT -20.565 66.475 -20.235 66.805 ;
        RECT -20.565 65.115 -20.235 65.445 ;
        RECT -20.565 63.755 -20.235 64.085 ;
        RECT -20.565 62.395 -20.235 62.725 ;
        RECT -20.565 61.035 -20.235 61.365 ;
        RECT -20.565 59.675 -20.235 60.005 ;
        RECT -20.565 58.315 -20.235 58.645 ;
        RECT -20.565 56.955 -20.235 57.285 ;
        RECT -20.565 55.595 -20.235 55.925 ;
        RECT -20.565 54.235 -20.235 54.565 ;
        RECT -20.565 52.875 -20.235 53.205 ;
        RECT -20.565 51.515 -20.235 51.845 ;
        RECT -20.565 50.155 -20.235 50.485 ;
        RECT -20.565 48.795 -20.235 49.125 ;
        RECT -20.565 47.435 -20.235 47.765 ;
        RECT -20.565 46.075 -20.235 46.405 ;
        RECT -20.565 44.715 -20.235 45.045 ;
        RECT -20.565 43.355 -20.235 43.685 ;
        RECT -20.565 41.995 -20.235 42.325 ;
        RECT -20.565 40.635 -20.235 40.965 ;
        RECT -20.565 39.275 -20.235 39.605 ;
        RECT -20.565 37.915 -20.235 38.245 ;
        RECT -20.565 36.555 -20.235 36.885 ;
        RECT -20.565 35.195 -20.235 35.525 ;
        RECT -20.565 33.835 -20.235 34.165 ;
        RECT -20.565 32.475 -20.235 32.805 ;
        RECT -20.565 31.115 -20.235 31.445 ;
        RECT -20.565 29.755 -20.235 30.085 ;
        RECT -20.565 28.395 -20.235 28.725 ;
        RECT -20.565 27.035 -20.235 27.365 ;
        RECT -20.565 25.675 -20.235 26.005 ;
        RECT -20.565 24.315 -20.235 24.645 ;
        RECT -20.565 22.955 -20.235 23.285 ;
        RECT -20.565 21.595 -20.235 21.925 ;
        RECT -20.565 20.235 -20.235 20.565 ;
        RECT -20.565 18.875 -20.235 19.205 ;
        RECT -20.565 17.515 -20.235 17.845 ;
        RECT -20.565 16.155 -20.235 16.485 ;
        RECT -20.565 14.795 -20.235 15.125 ;
        RECT -20.565 13.435 -20.235 13.765 ;
        RECT -20.565 12.075 -20.235 12.405 ;
        RECT -20.565 10.715 -20.235 11.045 ;
        RECT -20.565 9.355 -20.235 9.685 ;
        RECT -20.565 7.995 -20.235 8.325 ;
        RECT -20.565 6.635 -20.235 6.965 ;
        RECT -20.565 5.275 -20.235 5.605 ;
        RECT -20.565 3.915 -20.235 4.245 ;
        RECT -20.565 2.555 -20.235 2.885 ;
        RECT -20.565 1.195 -20.235 1.525 ;
        RECT -20.565 -0.165 -20.235 0.165 ;
        RECT -20.565 -1.525 -20.235 -1.195 ;
        RECT -20.565 -2.885 -20.235 -2.555 ;
        RECT -20.565 -4.245 -20.235 -3.915 ;
        RECT -20.565 -6.965 -20.235 -6.635 ;
        RECT -20.565 -8.325 -20.235 -7.995 ;
        RECT -20.565 -9.48 -20.235 -9.15 ;
        RECT -20.565 -12.405 -20.235 -12.075 ;
        RECT -20.565 -15.125 -20.235 -14.795 ;
        RECT -20.565 -16.67 -20.235 -16.34 ;
        RECT -20.565 -17.845 -20.235 -17.515 ;
        RECT -20.56 -21.24 -20.24 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -129.365 -20.235 -129.035 ;
        RECT -20.565 -130.725 -20.235 -130.395 ;
        RECT -20.565 -132.085 -20.235 -131.755 ;
        RECT -20.565 -133.51 -20.235 -133.18 ;
        RECT -20.565 -137.525 -20.235 -137.195 ;
        RECT -20.565 -138.885 -20.235 -138.555 ;
        RECT -20.565 -140.245 -20.235 -139.915 ;
        RECT -20.565 -141.605 -20.235 -141.275 ;
        RECT -20.565 -144.325 -20.235 -143.995 ;
        RECT -20.565 -145.685 -20.235 -145.355 ;
        RECT -20.565 -147.045 -20.235 -146.715 ;
        RECT -20.56 -149.08 -20.24 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -234.085 -20.235 -233.755 ;
        RECT -20.565 -235.445 -20.235 -235.115 ;
        RECT -20.565 -236.805 -20.235 -236.475 ;
        RECT -20.565 -238.165 -20.235 -237.835 ;
        RECT -20.565 -243.81 -20.235 -242.68 ;
        RECT -20.56 -243.925 -20.24 -231.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 246.76 -18.875 247.89 ;
        RECT -19.205 241.915 -18.875 242.245 ;
        RECT -19.205 240.555 -18.875 240.885 ;
        RECT -19.205 239.195 -18.875 239.525 ;
        RECT -19.205 237.835 -18.875 238.165 ;
        RECT -19.205 236.475 -18.875 236.805 ;
        RECT -19.205 235.115 -18.875 235.445 ;
        RECT -19.205 233.755 -18.875 234.085 ;
        RECT -19.205 232.395 -18.875 232.725 ;
        RECT -19.205 231.035 -18.875 231.365 ;
        RECT -19.205 229.675 -18.875 230.005 ;
        RECT -19.205 228.315 -18.875 228.645 ;
        RECT -19.205 226.955 -18.875 227.285 ;
        RECT -19.205 225.595 -18.875 225.925 ;
        RECT -19.205 224.235 -18.875 224.565 ;
        RECT -19.205 222.875 -18.875 223.205 ;
        RECT -19.205 221.515 -18.875 221.845 ;
        RECT -19.205 220.155 -18.875 220.485 ;
        RECT -19.205 218.795 -18.875 219.125 ;
        RECT -19.205 217.435 -18.875 217.765 ;
        RECT -19.205 216.075 -18.875 216.405 ;
        RECT -19.205 214.715 -18.875 215.045 ;
        RECT -19.205 213.355 -18.875 213.685 ;
        RECT -19.205 211.995 -18.875 212.325 ;
        RECT -19.205 210.635 -18.875 210.965 ;
        RECT -19.205 209.275 -18.875 209.605 ;
        RECT -19.205 207.915 -18.875 208.245 ;
        RECT -19.205 206.555 -18.875 206.885 ;
        RECT -19.205 205.195 -18.875 205.525 ;
        RECT -19.205 203.835 -18.875 204.165 ;
        RECT -19.205 202.475 -18.875 202.805 ;
        RECT -19.205 201.115 -18.875 201.445 ;
        RECT -19.205 199.755 -18.875 200.085 ;
        RECT -19.205 198.395 -18.875 198.725 ;
        RECT -19.205 197.035 -18.875 197.365 ;
        RECT -19.205 195.675 -18.875 196.005 ;
        RECT -19.205 194.315 -18.875 194.645 ;
        RECT -19.205 192.955 -18.875 193.285 ;
        RECT -19.205 191.595 -18.875 191.925 ;
        RECT -19.205 190.235 -18.875 190.565 ;
        RECT -19.205 188.875 -18.875 189.205 ;
        RECT -19.205 187.515 -18.875 187.845 ;
        RECT -19.205 186.155 -18.875 186.485 ;
        RECT -19.205 184.795 -18.875 185.125 ;
        RECT -19.205 183.435 -18.875 183.765 ;
        RECT -19.205 182.075 -18.875 182.405 ;
        RECT -19.205 180.715 -18.875 181.045 ;
        RECT -19.205 179.355 -18.875 179.685 ;
        RECT -19.205 177.995 -18.875 178.325 ;
        RECT -19.205 176.635 -18.875 176.965 ;
        RECT -19.205 175.275 -18.875 175.605 ;
        RECT -19.205 173.915 -18.875 174.245 ;
        RECT -19.205 172.555 -18.875 172.885 ;
        RECT -19.205 171.195 -18.875 171.525 ;
        RECT -19.205 169.835 -18.875 170.165 ;
        RECT -19.205 168.475 -18.875 168.805 ;
        RECT -19.205 167.115 -18.875 167.445 ;
        RECT -19.205 165.755 -18.875 166.085 ;
        RECT -19.205 164.395 -18.875 164.725 ;
        RECT -19.205 163.035 -18.875 163.365 ;
        RECT -19.205 161.675 -18.875 162.005 ;
        RECT -19.205 160.315 -18.875 160.645 ;
        RECT -19.205 158.955 -18.875 159.285 ;
        RECT -19.205 157.595 -18.875 157.925 ;
        RECT -19.205 156.235 -18.875 156.565 ;
        RECT -19.205 154.875 -18.875 155.205 ;
        RECT -19.205 153.515 -18.875 153.845 ;
        RECT -19.205 152.155 -18.875 152.485 ;
        RECT -19.205 150.795 -18.875 151.125 ;
        RECT -19.205 149.435 -18.875 149.765 ;
        RECT -19.205 148.075 -18.875 148.405 ;
        RECT -19.205 146.715 -18.875 147.045 ;
        RECT -19.205 145.355 -18.875 145.685 ;
        RECT -19.205 143.995 -18.875 144.325 ;
        RECT -19.205 142.635 -18.875 142.965 ;
        RECT -19.205 141.275 -18.875 141.605 ;
        RECT -19.205 139.915 -18.875 140.245 ;
        RECT -19.205 138.555 -18.875 138.885 ;
        RECT -19.205 137.195 -18.875 137.525 ;
        RECT -19.205 135.835 -18.875 136.165 ;
        RECT -19.205 134.475 -18.875 134.805 ;
        RECT -19.205 133.115 -18.875 133.445 ;
        RECT -19.205 131.755 -18.875 132.085 ;
        RECT -19.205 130.395 -18.875 130.725 ;
        RECT -19.205 129.035 -18.875 129.365 ;
        RECT -19.205 127.675 -18.875 128.005 ;
        RECT -19.205 126.315 -18.875 126.645 ;
        RECT -19.205 124.955 -18.875 125.285 ;
        RECT -19.205 123.595 -18.875 123.925 ;
        RECT -19.205 122.235 -18.875 122.565 ;
        RECT -19.205 120.875 -18.875 121.205 ;
        RECT -19.205 119.515 -18.875 119.845 ;
        RECT -19.205 118.155 -18.875 118.485 ;
        RECT -19.205 116.795 -18.875 117.125 ;
        RECT -19.205 115.435 -18.875 115.765 ;
        RECT -19.205 114.075 -18.875 114.405 ;
        RECT -19.205 112.715 -18.875 113.045 ;
        RECT -19.205 111.355 -18.875 111.685 ;
        RECT -19.205 109.995 -18.875 110.325 ;
        RECT -19.205 108.635 -18.875 108.965 ;
        RECT -19.205 107.275 -18.875 107.605 ;
        RECT -19.205 105.915 -18.875 106.245 ;
        RECT -19.205 104.555 -18.875 104.885 ;
        RECT -19.205 103.195 -18.875 103.525 ;
        RECT -19.205 101.835 -18.875 102.165 ;
        RECT -19.205 100.475 -18.875 100.805 ;
        RECT -19.205 99.115 -18.875 99.445 ;
        RECT -19.205 97.755 -18.875 98.085 ;
        RECT -19.205 96.395 -18.875 96.725 ;
        RECT -19.205 95.035 -18.875 95.365 ;
        RECT -19.205 93.675 -18.875 94.005 ;
        RECT -19.205 92.315 -18.875 92.645 ;
        RECT -19.205 90.955 -18.875 91.285 ;
        RECT -19.205 89.595 -18.875 89.925 ;
        RECT -19.205 88.235 -18.875 88.565 ;
        RECT -19.205 86.875 -18.875 87.205 ;
        RECT -19.205 85.515 -18.875 85.845 ;
        RECT -19.205 84.155 -18.875 84.485 ;
        RECT -19.205 82.795 -18.875 83.125 ;
        RECT -19.205 81.435 -18.875 81.765 ;
        RECT -19.205 80.075 -18.875 80.405 ;
        RECT -19.205 78.715 -18.875 79.045 ;
        RECT -19.205 77.355 -18.875 77.685 ;
        RECT -19.205 75.995 -18.875 76.325 ;
        RECT -19.205 74.635 -18.875 74.965 ;
        RECT -19.205 73.275 -18.875 73.605 ;
        RECT -19.205 71.915 -18.875 72.245 ;
        RECT -19.205 70.555 -18.875 70.885 ;
        RECT -19.205 69.195 -18.875 69.525 ;
        RECT -19.205 67.835 -18.875 68.165 ;
        RECT -19.205 66.475 -18.875 66.805 ;
        RECT -19.205 65.115 -18.875 65.445 ;
        RECT -19.205 63.755 -18.875 64.085 ;
        RECT -19.205 62.395 -18.875 62.725 ;
        RECT -19.205 61.035 -18.875 61.365 ;
        RECT -19.205 59.675 -18.875 60.005 ;
        RECT -19.205 58.315 -18.875 58.645 ;
        RECT -19.205 56.955 -18.875 57.285 ;
        RECT -19.205 55.595 -18.875 55.925 ;
        RECT -19.205 54.235 -18.875 54.565 ;
        RECT -19.205 52.875 -18.875 53.205 ;
        RECT -19.205 51.515 -18.875 51.845 ;
        RECT -19.205 50.155 -18.875 50.485 ;
        RECT -19.205 48.795 -18.875 49.125 ;
        RECT -19.205 47.435 -18.875 47.765 ;
        RECT -19.205 46.075 -18.875 46.405 ;
        RECT -19.205 44.715 -18.875 45.045 ;
        RECT -19.205 43.355 -18.875 43.685 ;
        RECT -19.205 41.995 -18.875 42.325 ;
        RECT -19.205 40.635 -18.875 40.965 ;
        RECT -19.205 39.275 -18.875 39.605 ;
        RECT -19.205 37.915 -18.875 38.245 ;
        RECT -19.205 36.555 -18.875 36.885 ;
        RECT -19.205 35.195 -18.875 35.525 ;
        RECT -19.205 33.835 -18.875 34.165 ;
        RECT -19.205 32.475 -18.875 32.805 ;
        RECT -19.205 31.115 -18.875 31.445 ;
        RECT -19.205 29.755 -18.875 30.085 ;
        RECT -19.205 28.395 -18.875 28.725 ;
        RECT -19.205 27.035 -18.875 27.365 ;
        RECT -19.205 25.675 -18.875 26.005 ;
        RECT -19.205 24.315 -18.875 24.645 ;
        RECT -19.205 22.955 -18.875 23.285 ;
        RECT -19.205 21.595 -18.875 21.925 ;
        RECT -19.205 20.235 -18.875 20.565 ;
        RECT -19.205 18.875 -18.875 19.205 ;
        RECT -19.205 17.515 -18.875 17.845 ;
        RECT -19.205 16.155 -18.875 16.485 ;
        RECT -19.205 14.795 -18.875 15.125 ;
        RECT -19.205 13.435 -18.875 13.765 ;
        RECT -19.205 12.075 -18.875 12.405 ;
        RECT -19.205 10.715 -18.875 11.045 ;
        RECT -19.205 9.355 -18.875 9.685 ;
        RECT -19.205 7.995 -18.875 8.325 ;
        RECT -19.205 6.635 -18.875 6.965 ;
        RECT -19.205 5.275 -18.875 5.605 ;
        RECT -19.205 3.915 -18.875 4.245 ;
        RECT -19.205 2.555 -18.875 2.885 ;
        RECT -19.205 1.195 -18.875 1.525 ;
        RECT -19.205 -0.165 -18.875 0.165 ;
        RECT -19.205 -1.525 -18.875 -1.195 ;
        RECT -19.205 -2.885 -18.875 -2.555 ;
        RECT -19.205 -4.245 -18.875 -3.915 ;
        RECT -19.205 -6.965 -18.875 -6.635 ;
        RECT -19.205 -8.325 -18.875 -7.995 ;
        RECT -19.205 -9.48 -18.875 -9.15 ;
        RECT -19.205 -12.405 -18.875 -12.075 ;
        RECT -19.205 -15.125 -18.875 -14.795 ;
        RECT -19.205 -16.67 -18.875 -16.34 ;
        RECT -19.205 -17.845 -18.875 -17.515 ;
        RECT -19.2 -19.88 -18.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -129.365 -18.875 -129.035 ;
        RECT -19.205 -130.725 -18.875 -130.395 ;
        RECT -19.205 -132.085 -18.875 -131.755 ;
        RECT -19.205 -133.51 -18.875 -133.18 ;
        RECT -19.205 -137.525 -18.875 -137.195 ;
        RECT -19.205 -138.885 -18.875 -138.555 ;
        RECT -19.205 -140.245 -18.875 -139.915 ;
        RECT -19.205 -141.605 -18.875 -141.275 ;
        RECT -19.205 -144.325 -18.875 -143.995 ;
        RECT -19.205 -145.685 -18.875 -145.355 ;
        RECT -19.205 -147.045 -18.875 -146.715 ;
        RECT -19.2 -148.4 -18.88 -127.68 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -230.005 -18.875 -229.675 ;
        RECT -19.205 -231.365 -18.875 -231.035 ;
        RECT -19.205 -234.085 -18.875 -233.755 ;
        RECT -19.205 -235.445 -18.875 -235.115 ;
        RECT -19.205 -236.805 -18.875 -236.475 ;
        RECT -19.205 -238.165 -18.875 -237.835 ;
        RECT -19.205 -243.81 -18.875 -242.68 ;
        RECT -19.2 -243.925 -18.88 -228.32 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 246.76 -17.515 247.89 ;
        RECT -17.845 241.915 -17.515 242.245 ;
        RECT -17.845 240.555 -17.515 240.885 ;
        RECT -17.845 239.195 -17.515 239.525 ;
        RECT -17.845 237.835 -17.515 238.165 ;
        RECT -17.845 236.475 -17.515 236.805 ;
        RECT -17.845 235.115 -17.515 235.445 ;
        RECT -17.845 233.755 -17.515 234.085 ;
        RECT -17.845 232.395 -17.515 232.725 ;
        RECT -17.845 231.035 -17.515 231.365 ;
        RECT -17.845 229.675 -17.515 230.005 ;
        RECT -17.845 228.315 -17.515 228.645 ;
        RECT -17.845 226.955 -17.515 227.285 ;
        RECT -17.845 225.595 -17.515 225.925 ;
        RECT -17.845 224.235 -17.515 224.565 ;
        RECT -17.845 222.875 -17.515 223.205 ;
        RECT -17.845 221.515 -17.515 221.845 ;
        RECT -17.845 220.155 -17.515 220.485 ;
        RECT -17.845 218.795 -17.515 219.125 ;
        RECT -17.845 217.435 -17.515 217.765 ;
        RECT -17.845 216.075 -17.515 216.405 ;
        RECT -17.845 214.715 -17.515 215.045 ;
        RECT -17.845 213.355 -17.515 213.685 ;
        RECT -17.845 211.995 -17.515 212.325 ;
        RECT -17.845 210.635 -17.515 210.965 ;
        RECT -17.845 209.275 -17.515 209.605 ;
        RECT -17.845 207.915 -17.515 208.245 ;
        RECT -17.845 206.555 -17.515 206.885 ;
        RECT -17.845 205.195 -17.515 205.525 ;
        RECT -17.845 203.835 -17.515 204.165 ;
        RECT -17.845 202.475 -17.515 202.805 ;
        RECT -17.845 201.115 -17.515 201.445 ;
        RECT -17.845 199.755 -17.515 200.085 ;
        RECT -17.845 198.395 -17.515 198.725 ;
        RECT -17.845 197.035 -17.515 197.365 ;
        RECT -17.845 195.675 -17.515 196.005 ;
        RECT -17.845 194.315 -17.515 194.645 ;
        RECT -17.845 192.955 -17.515 193.285 ;
        RECT -17.845 191.595 -17.515 191.925 ;
        RECT -17.845 190.235 -17.515 190.565 ;
        RECT -17.845 188.875 -17.515 189.205 ;
        RECT -17.845 187.515 -17.515 187.845 ;
        RECT -17.845 186.155 -17.515 186.485 ;
        RECT -17.845 184.795 -17.515 185.125 ;
        RECT -17.845 183.435 -17.515 183.765 ;
        RECT -17.845 182.075 -17.515 182.405 ;
        RECT -17.845 180.715 -17.515 181.045 ;
        RECT -17.845 179.355 -17.515 179.685 ;
        RECT -17.845 177.995 -17.515 178.325 ;
        RECT -17.845 176.635 -17.515 176.965 ;
        RECT -17.845 175.275 -17.515 175.605 ;
        RECT -17.845 173.915 -17.515 174.245 ;
        RECT -17.845 172.555 -17.515 172.885 ;
        RECT -17.845 171.195 -17.515 171.525 ;
        RECT -17.845 169.835 -17.515 170.165 ;
        RECT -17.845 168.475 -17.515 168.805 ;
        RECT -17.845 167.115 -17.515 167.445 ;
        RECT -17.845 165.755 -17.515 166.085 ;
        RECT -17.845 164.395 -17.515 164.725 ;
        RECT -17.845 163.035 -17.515 163.365 ;
        RECT -17.845 161.675 -17.515 162.005 ;
        RECT -17.845 160.315 -17.515 160.645 ;
        RECT -17.845 158.955 -17.515 159.285 ;
        RECT -17.845 157.595 -17.515 157.925 ;
        RECT -17.845 156.235 -17.515 156.565 ;
        RECT -17.845 154.875 -17.515 155.205 ;
        RECT -17.845 153.515 -17.515 153.845 ;
        RECT -17.845 152.155 -17.515 152.485 ;
        RECT -17.845 150.795 -17.515 151.125 ;
        RECT -17.845 149.435 -17.515 149.765 ;
        RECT -17.845 148.075 -17.515 148.405 ;
        RECT -17.845 146.715 -17.515 147.045 ;
        RECT -17.845 145.355 -17.515 145.685 ;
        RECT -17.845 143.995 -17.515 144.325 ;
        RECT -17.845 142.635 -17.515 142.965 ;
        RECT -17.845 141.275 -17.515 141.605 ;
        RECT -17.845 139.915 -17.515 140.245 ;
        RECT -17.845 138.555 -17.515 138.885 ;
        RECT -17.845 137.195 -17.515 137.525 ;
        RECT -17.845 135.835 -17.515 136.165 ;
        RECT -17.845 134.475 -17.515 134.805 ;
        RECT -17.845 133.115 -17.515 133.445 ;
        RECT -17.845 131.755 -17.515 132.085 ;
        RECT -17.845 130.395 -17.515 130.725 ;
        RECT -17.845 129.035 -17.515 129.365 ;
        RECT -17.845 127.675 -17.515 128.005 ;
        RECT -17.845 126.315 -17.515 126.645 ;
        RECT -17.845 124.955 -17.515 125.285 ;
        RECT -17.845 123.595 -17.515 123.925 ;
        RECT -17.845 122.235 -17.515 122.565 ;
        RECT -17.845 120.875 -17.515 121.205 ;
        RECT -17.845 119.515 -17.515 119.845 ;
        RECT -17.845 118.155 -17.515 118.485 ;
        RECT -17.845 116.795 -17.515 117.125 ;
        RECT -17.845 115.435 -17.515 115.765 ;
        RECT -17.845 114.075 -17.515 114.405 ;
        RECT -17.845 112.715 -17.515 113.045 ;
        RECT -17.845 111.355 -17.515 111.685 ;
        RECT -17.845 109.995 -17.515 110.325 ;
        RECT -17.845 108.635 -17.515 108.965 ;
        RECT -17.845 107.275 -17.515 107.605 ;
        RECT -17.845 105.915 -17.515 106.245 ;
        RECT -17.845 104.555 -17.515 104.885 ;
        RECT -17.845 103.195 -17.515 103.525 ;
        RECT -17.845 101.835 -17.515 102.165 ;
        RECT -17.845 100.475 -17.515 100.805 ;
        RECT -17.845 99.115 -17.515 99.445 ;
        RECT -17.845 97.755 -17.515 98.085 ;
        RECT -17.845 96.395 -17.515 96.725 ;
        RECT -17.845 95.035 -17.515 95.365 ;
        RECT -17.845 93.675 -17.515 94.005 ;
        RECT -17.845 92.315 -17.515 92.645 ;
        RECT -17.845 90.955 -17.515 91.285 ;
        RECT -17.845 89.595 -17.515 89.925 ;
        RECT -17.845 88.235 -17.515 88.565 ;
        RECT -17.845 86.875 -17.515 87.205 ;
        RECT -17.845 85.515 -17.515 85.845 ;
        RECT -17.845 84.155 -17.515 84.485 ;
        RECT -17.845 82.795 -17.515 83.125 ;
        RECT -17.845 81.435 -17.515 81.765 ;
        RECT -17.845 80.075 -17.515 80.405 ;
        RECT -17.845 78.715 -17.515 79.045 ;
        RECT -17.845 77.355 -17.515 77.685 ;
        RECT -17.845 75.995 -17.515 76.325 ;
        RECT -17.845 74.635 -17.515 74.965 ;
        RECT -17.845 73.275 -17.515 73.605 ;
        RECT -17.845 71.915 -17.515 72.245 ;
        RECT -17.845 70.555 -17.515 70.885 ;
        RECT -17.845 69.195 -17.515 69.525 ;
        RECT -17.845 67.835 -17.515 68.165 ;
        RECT -17.845 66.475 -17.515 66.805 ;
        RECT -17.845 65.115 -17.515 65.445 ;
        RECT -17.845 63.755 -17.515 64.085 ;
        RECT -17.845 62.395 -17.515 62.725 ;
        RECT -17.845 61.035 -17.515 61.365 ;
        RECT -17.845 59.675 -17.515 60.005 ;
        RECT -17.845 58.315 -17.515 58.645 ;
        RECT -17.845 56.955 -17.515 57.285 ;
        RECT -17.845 55.595 -17.515 55.925 ;
        RECT -17.845 54.235 -17.515 54.565 ;
        RECT -17.845 52.875 -17.515 53.205 ;
        RECT -17.845 51.515 -17.515 51.845 ;
        RECT -17.845 50.155 -17.515 50.485 ;
        RECT -17.845 48.795 -17.515 49.125 ;
        RECT -17.845 47.435 -17.515 47.765 ;
        RECT -17.845 46.075 -17.515 46.405 ;
        RECT -17.845 44.715 -17.515 45.045 ;
        RECT -17.845 43.355 -17.515 43.685 ;
        RECT -17.845 41.995 -17.515 42.325 ;
        RECT -17.845 40.635 -17.515 40.965 ;
        RECT -17.845 39.275 -17.515 39.605 ;
        RECT -17.845 37.915 -17.515 38.245 ;
        RECT -17.845 36.555 -17.515 36.885 ;
        RECT -17.845 35.195 -17.515 35.525 ;
        RECT -17.845 33.835 -17.515 34.165 ;
        RECT -17.845 32.475 -17.515 32.805 ;
        RECT -17.845 31.115 -17.515 31.445 ;
        RECT -17.845 29.755 -17.515 30.085 ;
        RECT -17.845 28.395 -17.515 28.725 ;
        RECT -17.845 27.035 -17.515 27.365 ;
        RECT -17.845 25.675 -17.515 26.005 ;
        RECT -17.845 24.315 -17.515 24.645 ;
        RECT -17.845 22.955 -17.515 23.285 ;
        RECT -17.845 21.595 -17.515 21.925 ;
        RECT -17.845 20.235 -17.515 20.565 ;
        RECT -17.845 18.875 -17.515 19.205 ;
        RECT -17.845 17.515 -17.515 17.845 ;
        RECT -17.845 16.155 -17.515 16.485 ;
        RECT -17.845 14.795 -17.515 15.125 ;
        RECT -17.845 13.435 -17.515 13.765 ;
        RECT -17.845 12.075 -17.515 12.405 ;
        RECT -17.845 10.715 -17.515 11.045 ;
        RECT -17.845 9.355 -17.515 9.685 ;
        RECT -17.845 7.995 -17.515 8.325 ;
        RECT -17.845 6.635 -17.515 6.965 ;
        RECT -17.845 5.275 -17.515 5.605 ;
        RECT -17.845 3.915 -17.515 4.245 ;
        RECT -17.845 2.555 -17.515 2.885 ;
        RECT -17.845 1.195 -17.515 1.525 ;
        RECT -17.845 -0.165 -17.515 0.165 ;
        RECT -17.845 -1.525 -17.515 -1.195 ;
        RECT -17.845 -2.885 -17.515 -2.555 ;
        RECT -17.845 -4.245 -17.515 -3.915 ;
        RECT -17.845 -6.965 -17.515 -6.635 ;
        RECT -17.845 -8.325 -17.515 -7.995 ;
        RECT -17.845 -9.48 -17.515 -9.15 ;
        RECT -17.845 -12.405 -17.515 -12.075 ;
        RECT -17.845 -15.125 -17.515 -14.795 ;
        RECT -17.845 -16.67 -17.515 -16.34 ;
        RECT -17.845 -17.845 -17.515 -17.515 ;
        RECT -17.845 -24.645 -17.515 -24.315 ;
        RECT -17.845 -26.005 -17.515 -25.675 ;
        RECT -17.845 -30.66 -17.515 -30.33 ;
        RECT -17.845 -31.445 -17.515 -31.115 ;
        RECT -17.845 -32.805 -17.515 -32.475 ;
        RECT -17.845 -34.165 -17.515 -33.835 ;
        RECT -17.845 -36.885 -17.515 -36.555 ;
        RECT -17.845 -37.85 -17.515 -37.52 ;
        RECT -17.845 -40.965 -17.515 -40.635 ;
        RECT -17.845 -46.405 -17.515 -46.075 ;
        RECT -17.845 -47.765 -17.515 -47.435 ;
        RECT -17.845 -49.125 -17.515 -48.795 ;
        RECT -17.845 -50.485 -17.515 -50.155 ;
        RECT -17.845 -51.845 -17.515 -51.515 ;
        RECT -17.845 -53.205 -17.515 -52.875 ;
        RECT -17.845 -54.565 -17.515 -54.235 ;
        RECT -17.845 -55.925 -17.515 -55.595 ;
        RECT -17.845 -57.285 -17.515 -56.955 ;
        RECT -17.845 -58.645 -17.515 -58.315 ;
        RECT -17.845 -60.005 -17.515 -59.675 ;
        RECT -17.845 -61.365 -17.515 -61.035 ;
        RECT -17.845 -62.725 -17.515 -62.395 ;
        RECT -17.845 -68.165 -17.515 -67.835 ;
        RECT -17.845 -69.525 -17.515 -69.195 ;
        RECT -17.845 -70.79 -17.515 -70.46 ;
        RECT -17.845 -72.245 -17.515 -71.915 ;
        RECT -17.845 -73.605 -17.515 -73.275 ;
        RECT -17.845 -74.965 -17.515 -74.635 ;
        RECT -17.845 -76.325 -17.515 -75.995 ;
        RECT -17.845 -77.685 -17.515 -77.355 ;
        RECT -17.845 -79.045 -17.515 -78.715 ;
        RECT -17.845 -81.765 -17.515 -81.435 ;
        RECT -17.845 -83.125 -17.515 -82.795 ;
        RECT -17.845 -84.485 -17.515 -84.155 ;
        RECT -17.845 -85.845 -17.515 -85.515 ;
        RECT -17.845 -87.205 -17.515 -86.875 ;
        RECT -17.845 -88.565 -17.515 -88.235 ;
        RECT -17.845 -89.33 -17.515 -89 ;
        RECT -17.845 -91.285 -17.515 -90.955 ;
        RECT -17.845 -92.645 -17.515 -92.315 ;
        RECT -17.845 -94.005 -17.515 -93.675 ;
        RECT -17.845 -95.365 -17.515 -95.035 ;
        RECT -17.845 -96.725 -17.515 -96.395 ;
        RECT -17.845 -98.085 -17.515 -97.755 ;
        RECT -17.845 -100.805 -17.515 -100.475 ;
        RECT -17.845 -102.165 -17.515 -101.835 ;
        RECT -17.845 -103.525 -17.515 -103.195 ;
        RECT -17.845 -106.245 -17.515 -105.915 ;
        RECT -17.845 -107.605 -17.515 -107.275 ;
        RECT -17.845 -108.965 -17.515 -108.635 ;
        RECT -17.845 -110.325 -17.515 -109.995 ;
        RECT -17.845 -111.685 -17.515 -111.355 ;
        RECT -17.845 -113.045 -17.515 -112.715 ;
        RECT -17.845 -114.97 -17.515 -114.64 ;
        RECT -17.845 -115.765 -17.515 -115.435 ;
        RECT -17.845 -117.125 -17.515 -116.795 ;
        RECT -17.845 -118.485 -17.515 -118.155 ;
        RECT -17.845 -119.845 -17.515 -119.515 ;
        RECT -17.845 -121.205 -17.515 -120.875 ;
        RECT -17.845 -122.565 -17.515 -122.235 ;
        RECT -17.845 -125.285 -17.515 -124.955 ;
        RECT -17.845 -126.645 -17.515 -126.315 ;
        RECT -17.845 -128.005 -17.515 -127.675 ;
        RECT -17.845 -129.365 -17.515 -129.035 ;
        RECT -17.845 -130.725 -17.515 -130.395 ;
        RECT -17.845 -132.085 -17.515 -131.755 ;
        RECT -17.845 -133.51 -17.515 -133.18 ;
        RECT -17.845 -138.885 -17.515 -138.555 ;
        RECT -17.845 -140.245 -17.515 -139.915 ;
        RECT -17.845 -141.605 -17.515 -141.275 ;
        RECT -17.845 -144.325 -17.515 -143.995 ;
        RECT -17.845 -145.685 -17.515 -145.355 ;
        RECT -17.845 -147.045 -17.515 -146.715 ;
        RECT -17.845 -152.485 -17.515 -152.155 ;
        RECT -17.845 -153.845 -17.515 -153.515 ;
        RECT -17.845 -155.205 -17.515 -154.875 ;
        RECT -17.845 -156.565 -17.515 -156.235 ;
        RECT -17.845 -157.925 -17.515 -157.595 ;
        RECT -17.845 -164.725 -17.515 -164.395 ;
        RECT -17.845 -167.445 -17.515 -167.115 ;
        RECT -17.845 -168.805 -17.515 -168.475 ;
        RECT -17.845 -170.165 -17.515 -169.835 ;
        RECT -17.845 -171.525 -17.515 -171.195 ;
        RECT -17.845 -175.605 -17.515 -175.275 ;
        RECT -17.845 -176.965 -17.515 -176.635 ;
        RECT -17.845 -178.325 -17.515 -177.995 ;
        RECT -17.845 -179.685 -17.515 -179.355 ;
        RECT -17.845 -181.045 -17.515 -180.715 ;
        RECT -17.845 -182.405 -17.515 -182.075 ;
        RECT -17.845 -185.125 -17.515 -184.795 ;
        RECT -17.845 -194.645 -17.515 -194.315 ;
        RECT -17.845 -196.005 -17.515 -195.675 ;
        RECT -17.845 -201.445 -17.515 -201.115 ;
        RECT -17.845 -202.805 -17.515 -202.475 ;
        RECT -17.845 -209.605 -17.515 -209.275 ;
        RECT -17.845 -213.685 -17.515 -213.355 ;
        RECT -17.845 -215.045 -17.515 -214.715 ;
        RECT -17.845 -216.405 -17.515 -216.075 ;
        RECT -17.845 -217.765 -17.515 -217.435 ;
        RECT -17.845 -219.125 -17.515 -218.795 ;
        RECT -17.845 -220.485 -17.515 -220.155 ;
        RECT -17.845 -221.845 -17.515 -221.515 ;
        RECT -17.845 -223.205 -17.515 -222.875 ;
        RECT -17.845 -226.155 -17.515 -225.825 ;
        RECT -17.845 -227.285 -17.515 -226.955 ;
        RECT -17.845 -228.645 -17.515 -228.315 ;
        RECT -17.845 -230.005 -17.515 -229.675 ;
        RECT -17.845 -234.085 -17.515 -233.755 ;
        RECT -17.845 -235.445 -17.515 -235.115 ;
        RECT -17.845 -236.805 -17.515 -236.475 ;
        RECT -17.845 -238.165 -17.515 -237.835 ;
        RECT -17.845 -243.81 -17.515 -242.68 ;
        RECT -17.84 -243.925 -17.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 74.635 -16.155 74.965 ;
        RECT -16.485 73.275 -16.155 73.605 ;
        RECT -16.485 71.915 -16.155 72.245 ;
        RECT -16.485 70.555 -16.155 70.885 ;
        RECT -16.485 69.195 -16.155 69.525 ;
        RECT -16.485 67.835 -16.155 68.165 ;
        RECT -16.485 66.475 -16.155 66.805 ;
        RECT -16.485 65.115 -16.155 65.445 ;
        RECT -16.485 63.755 -16.155 64.085 ;
        RECT -16.485 62.395 -16.155 62.725 ;
        RECT -16.485 61.035 -16.155 61.365 ;
        RECT -16.485 59.675 -16.155 60.005 ;
        RECT -16.485 58.315 -16.155 58.645 ;
        RECT -16.485 56.955 -16.155 57.285 ;
        RECT -16.485 55.595 -16.155 55.925 ;
        RECT -16.485 54.235 -16.155 54.565 ;
        RECT -16.485 52.875 -16.155 53.205 ;
        RECT -16.485 51.515 -16.155 51.845 ;
        RECT -16.485 50.155 -16.155 50.485 ;
        RECT -16.485 48.795 -16.155 49.125 ;
        RECT -16.485 47.435 -16.155 47.765 ;
        RECT -16.485 46.075 -16.155 46.405 ;
        RECT -16.485 44.715 -16.155 45.045 ;
        RECT -16.485 43.355 -16.155 43.685 ;
        RECT -16.485 41.995 -16.155 42.325 ;
        RECT -16.485 40.635 -16.155 40.965 ;
        RECT -16.485 39.275 -16.155 39.605 ;
        RECT -16.485 37.915 -16.155 38.245 ;
        RECT -16.485 36.555 -16.155 36.885 ;
        RECT -16.485 35.195 -16.155 35.525 ;
        RECT -16.485 33.835 -16.155 34.165 ;
        RECT -16.485 32.475 -16.155 32.805 ;
        RECT -16.485 31.115 -16.155 31.445 ;
        RECT -16.485 29.755 -16.155 30.085 ;
        RECT -16.485 28.395 -16.155 28.725 ;
        RECT -16.485 27.035 -16.155 27.365 ;
        RECT -16.485 25.675 -16.155 26.005 ;
        RECT -16.485 24.315 -16.155 24.645 ;
        RECT -16.485 22.955 -16.155 23.285 ;
        RECT -16.485 21.595 -16.155 21.925 ;
        RECT -16.485 20.235 -16.155 20.565 ;
        RECT -16.485 18.875 -16.155 19.205 ;
        RECT -16.485 17.515 -16.155 17.845 ;
        RECT -16.485 16.155 -16.155 16.485 ;
        RECT -16.485 14.795 -16.155 15.125 ;
        RECT -16.485 13.435 -16.155 13.765 ;
        RECT -16.485 12.075 -16.155 12.405 ;
        RECT -16.485 10.715 -16.155 11.045 ;
        RECT -16.485 9.355 -16.155 9.685 ;
        RECT -16.485 7.995 -16.155 8.325 ;
        RECT -16.485 6.635 -16.155 6.965 ;
        RECT -16.485 5.275 -16.155 5.605 ;
        RECT -16.485 3.915 -16.155 4.245 ;
        RECT -16.485 2.555 -16.155 2.885 ;
        RECT -16.485 1.195 -16.155 1.525 ;
        RECT -16.485 -0.165 -16.155 0.165 ;
        RECT -16.485 -1.525 -16.155 -1.195 ;
        RECT -16.485 -2.885 -16.155 -2.555 ;
        RECT -16.485 -4.245 -16.155 -3.915 ;
        RECT -16.485 -5.605 -16.155 -5.275 ;
        RECT -16.485 -6.965 -16.155 -6.635 ;
        RECT -16.485 -8.325 -16.155 -7.995 ;
        RECT -16.485 -9.48 -16.155 -9.15 ;
        RECT -16.485 -12.405 -16.155 -12.075 ;
        RECT -16.485 -15.125 -16.155 -14.795 ;
        RECT -16.485 -16.67 -16.155 -16.34 ;
        RECT -16.485 -17.845 -16.155 -17.515 ;
        RECT -16.485 -24.645 -16.155 -24.315 ;
        RECT -16.485 -26.005 -16.155 -25.675 ;
        RECT -16.485 -27.365 -16.155 -27.035 ;
        RECT -16.485 -30.66 -16.155 -30.33 ;
        RECT -16.485 -31.445 -16.155 -31.115 ;
        RECT -16.485 -32.805 -16.155 -32.475 ;
        RECT -16.485 -34.165 -16.155 -33.835 ;
        RECT -16.485 -36.885 -16.155 -36.555 ;
        RECT -16.485 -37.85 -16.155 -37.52 ;
        RECT -16.485 -40.965 -16.155 -40.635 ;
        RECT -16.485 -46.405 -16.155 -46.075 ;
        RECT -16.485 -47.765 -16.155 -47.435 ;
        RECT -16.485 -49.125 -16.155 -48.795 ;
        RECT -16.485 -50.485 -16.155 -50.155 ;
        RECT -16.485 -51.845 -16.155 -51.515 ;
        RECT -16.485 -53.205 -16.155 -52.875 ;
        RECT -16.485 -54.565 -16.155 -54.235 ;
        RECT -16.485 -55.925 -16.155 -55.595 ;
        RECT -16.485 -57.285 -16.155 -56.955 ;
        RECT -16.485 -58.645 -16.155 -58.315 ;
        RECT -16.485 -60.005 -16.155 -59.675 ;
        RECT -16.485 -61.365 -16.155 -61.035 ;
        RECT -16.485 -62.725 -16.155 -62.395 ;
        RECT -16.485 -68.165 -16.155 -67.835 ;
        RECT -16.485 -69.525 -16.155 -69.195 ;
        RECT -16.485 -70.79 -16.155 -70.46 ;
        RECT -16.48 -70.88 -16.16 248.005 ;
        RECT -16.485 246.76 -16.155 247.89 ;
        RECT -16.485 241.915 -16.155 242.245 ;
        RECT -16.485 240.555 -16.155 240.885 ;
        RECT -16.485 239.195 -16.155 239.525 ;
        RECT -16.485 237.835 -16.155 238.165 ;
        RECT -16.485 236.475 -16.155 236.805 ;
        RECT -16.485 235.115 -16.155 235.445 ;
        RECT -16.485 233.755 -16.155 234.085 ;
        RECT -16.485 232.395 -16.155 232.725 ;
        RECT -16.485 231.035 -16.155 231.365 ;
        RECT -16.485 229.675 -16.155 230.005 ;
        RECT -16.485 228.315 -16.155 228.645 ;
        RECT -16.485 226.955 -16.155 227.285 ;
        RECT -16.485 225.595 -16.155 225.925 ;
        RECT -16.485 224.235 -16.155 224.565 ;
        RECT -16.485 222.875 -16.155 223.205 ;
        RECT -16.485 221.515 -16.155 221.845 ;
        RECT -16.485 220.155 -16.155 220.485 ;
        RECT -16.485 218.795 -16.155 219.125 ;
        RECT -16.485 217.435 -16.155 217.765 ;
        RECT -16.485 216.075 -16.155 216.405 ;
        RECT -16.485 214.715 -16.155 215.045 ;
        RECT -16.485 213.355 -16.155 213.685 ;
        RECT -16.485 211.995 -16.155 212.325 ;
        RECT -16.485 210.635 -16.155 210.965 ;
        RECT -16.485 209.275 -16.155 209.605 ;
        RECT -16.485 207.915 -16.155 208.245 ;
        RECT -16.485 206.555 -16.155 206.885 ;
        RECT -16.485 205.195 -16.155 205.525 ;
        RECT -16.485 203.835 -16.155 204.165 ;
        RECT -16.485 202.475 -16.155 202.805 ;
        RECT -16.485 201.115 -16.155 201.445 ;
        RECT -16.485 199.755 -16.155 200.085 ;
        RECT -16.485 198.395 -16.155 198.725 ;
        RECT -16.485 197.035 -16.155 197.365 ;
        RECT -16.485 195.675 -16.155 196.005 ;
        RECT -16.485 194.315 -16.155 194.645 ;
        RECT -16.485 192.955 -16.155 193.285 ;
        RECT -16.485 191.595 -16.155 191.925 ;
        RECT -16.485 190.235 -16.155 190.565 ;
        RECT -16.485 188.875 -16.155 189.205 ;
        RECT -16.485 187.515 -16.155 187.845 ;
        RECT -16.485 186.155 -16.155 186.485 ;
        RECT -16.485 184.795 -16.155 185.125 ;
        RECT -16.485 183.435 -16.155 183.765 ;
        RECT -16.485 182.075 -16.155 182.405 ;
        RECT -16.485 180.715 -16.155 181.045 ;
        RECT -16.485 179.355 -16.155 179.685 ;
        RECT -16.485 177.995 -16.155 178.325 ;
        RECT -16.485 176.635 -16.155 176.965 ;
        RECT -16.485 175.275 -16.155 175.605 ;
        RECT -16.485 173.915 -16.155 174.245 ;
        RECT -16.485 172.555 -16.155 172.885 ;
        RECT -16.485 171.195 -16.155 171.525 ;
        RECT -16.485 169.835 -16.155 170.165 ;
        RECT -16.485 168.475 -16.155 168.805 ;
        RECT -16.485 167.115 -16.155 167.445 ;
        RECT -16.485 165.755 -16.155 166.085 ;
        RECT -16.485 164.395 -16.155 164.725 ;
        RECT -16.485 163.035 -16.155 163.365 ;
        RECT -16.485 161.675 -16.155 162.005 ;
        RECT -16.485 160.315 -16.155 160.645 ;
        RECT -16.485 158.955 -16.155 159.285 ;
        RECT -16.485 157.595 -16.155 157.925 ;
        RECT -16.485 156.235 -16.155 156.565 ;
        RECT -16.485 154.875 -16.155 155.205 ;
        RECT -16.485 153.515 -16.155 153.845 ;
        RECT -16.485 152.155 -16.155 152.485 ;
        RECT -16.485 150.795 -16.155 151.125 ;
        RECT -16.485 149.435 -16.155 149.765 ;
        RECT -16.485 148.075 -16.155 148.405 ;
        RECT -16.485 146.715 -16.155 147.045 ;
        RECT -16.485 145.355 -16.155 145.685 ;
        RECT -16.485 143.995 -16.155 144.325 ;
        RECT -16.485 142.635 -16.155 142.965 ;
        RECT -16.485 141.275 -16.155 141.605 ;
        RECT -16.485 139.915 -16.155 140.245 ;
        RECT -16.485 138.555 -16.155 138.885 ;
        RECT -16.485 137.195 -16.155 137.525 ;
        RECT -16.485 135.835 -16.155 136.165 ;
        RECT -16.485 134.475 -16.155 134.805 ;
        RECT -16.485 133.115 -16.155 133.445 ;
        RECT -16.485 131.755 -16.155 132.085 ;
        RECT -16.485 130.395 -16.155 130.725 ;
        RECT -16.485 129.035 -16.155 129.365 ;
        RECT -16.485 127.675 -16.155 128.005 ;
        RECT -16.485 126.315 -16.155 126.645 ;
        RECT -16.485 124.955 -16.155 125.285 ;
        RECT -16.485 123.595 -16.155 123.925 ;
        RECT -16.485 122.235 -16.155 122.565 ;
        RECT -16.485 120.875 -16.155 121.205 ;
        RECT -16.485 119.515 -16.155 119.845 ;
        RECT -16.485 118.155 -16.155 118.485 ;
        RECT -16.485 116.795 -16.155 117.125 ;
        RECT -16.485 115.435 -16.155 115.765 ;
        RECT -16.485 114.075 -16.155 114.405 ;
        RECT -16.485 112.715 -16.155 113.045 ;
        RECT -16.485 111.355 -16.155 111.685 ;
        RECT -16.485 109.995 -16.155 110.325 ;
        RECT -16.485 108.635 -16.155 108.965 ;
        RECT -16.485 107.275 -16.155 107.605 ;
        RECT -16.485 105.915 -16.155 106.245 ;
        RECT -16.485 104.555 -16.155 104.885 ;
        RECT -16.485 103.195 -16.155 103.525 ;
        RECT -16.485 101.835 -16.155 102.165 ;
        RECT -16.485 100.475 -16.155 100.805 ;
        RECT -16.485 99.115 -16.155 99.445 ;
        RECT -16.485 97.755 -16.155 98.085 ;
        RECT -16.485 96.395 -16.155 96.725 ;
        RECT -16.485 95.035 -16.155 95.365 ;
        RECT -16.485 93.675 -16.155 94.005 ;
        RECT -16.485 92.315 -16.155 92.645 ;
        RECT -16.485 90.955 -16.155 91.285 ;
        RECT -16.485 89.595 -16.155 89.925 ;
        RECT -16.485 88.235 -16.155 88.565 ;
        RECT -16.485 86.875 -16.155 87.205 ;
        RECT -16.485 85.515 -16.155 85.845 ;
        RECT -16.485 84.155 -16.155 84.485 ;
        RECT -16.485 82.795 -16.155 83.125 ;
        RECT -16.485 81.435 -16.155 81.765 ;
        RECT -16.485 80.075 -16.155 80.405 ;
        RECT -16.485 78.715 -16.155 79.045 ;
        RECT -16.485 77.355 -16.155 77.685 ;
        RECT -16.485 75.995 -16.155 76.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.005 246.76 -25.675 247.89 ;
        RECT -26.005 241.915 -25.675 242.245 ;
        RECT -26.005 240.555 -25.675 240.885 ;
        RECT -26.005 239.195 -25.675 239.525 ;
        RECT -26.005 237.835 -25.675 238.165 ;
        RECT -26.005 236.475 -25.675 236.805 ;
        RECT -26.005 235.115 -25.675 235.445 ;
        RECT -26.005 233.755 -25.675 234.085 ;
        RECT -26.005 232.395 -25.675 232.725 ;
        RECT -26.005 231.035 -25.675 231.365 ;
        RECT -26.005 229.675 -25.675 230.005 ;
        RECT -26.005 228.315 -25.675 228.645 ;
        RECT -26.005 226.955 -25.675 227.285 ;
        RECT -26.005 225.595 -25.675 225.925 ;
        RECT -26.005 224.235 -25.675 224.565 ;
        RECT -26.005 222.875 -25.675 223.205 ;
        RECT -26.005 221.515 -25.675 221.845 ;
        RECT -26.005 220.155 -25.675 220.485 ;
        RECT -26.005 218.795 -25.675 219.125 ;
        RECT -26.005 217.435 -25.675 217.765 ;
        RECT -26.005 216.075 -25.675 216.405 ;
        RECT -26.005 214.715 -25.675 215.045 ;
        RECT -26.005 213.355 -25.675 213.685 ;
        RECT -26.005 211.995 -25.675 212.325 ;
        RECT -26.005 210.635 -25.675 210.965 ;
        RECT -26.005 209.275 -25.675 209.605 ;
        RECT -26.005 207.915 -25.675 208.245 ;
        RECT -26.005 206.555 -25.675 206.885 ;
        RECT -26.005 205.195 -25.675 205.525 ;
        RECT -26.005 203.835 -25.675 204.165 ;
        RECT -26.005 202.475 -25.675 202.805 ;
        RECT -26.005 201.115 -25.675 201.445 ;
        RECT -26.005 199.755 -25.675 200.085 ;
        RECT -26.005 198.395 -25.675 198.725 ;
        RECT -26.005 197.035 -25.675 197.365 ;
        RECT -26.005 195.675 -25.675 196.005 ;
        RECT -26.005 194.315 -25.675 194.645 ;
        RECT -26.005 192.955 -25.675 193.285 ;
        RECT -26.005 191.595 -25.675 191.925 ;
        RECT -26.005 190.235 -25.675 190.565 ;
        RECT -26.005 188.875 -25.675 189.205 ;
        RECT -26.005 187.515 -25.675 187.845 ;
        RECT -26.005 186.155 -25.675 186.485 ;
        RECT -26.005 184.795 -25.675 185.125 ;
        RECT -26.005 183.435 -25.675 183.765 ;
        RECT -26.005 182.075 -25.675 182.405 ;
        RECT -26.005 180.715 -25.675 181.045 ;
        RECT -26.005 179.355 -25.675 179.685 ;
        RECT -26.005 177.995 -25.675 178.325 ;
        RECT -26.005 176.635 -25.675 176.965 ;
        RECT -26.005 175.275 -25.675 175.605 ;
        RECT -26.005 173.915 -25.675 174.245 ;
        RECT -26.005 172.555 -25.675 172.885 ;
        RECT -26.005 171.195 -25.675 171.525 ;
        RECT -26.005 169.835 -25.675 170.165 ;
        RECT -26.005 168.475 -25.675 168.805 ;
        RECT -26.005 167.115 -25.675 167.445 ;
        RECT -26.005 165.755 -25.675 166.085 ;
        RECT -26.005 164.395 -25.675 164.725 ;
        RECT -26.005 163.035 -25.675 163.365 ;
        RECT -26.005 161.675 -25.675 162.005 ;
        RECT -26.005 160.315 -25.675 160.645 ;
        RECT -26.005 158.955 -25.675 159.285 ;
        RECT -26.005 157.595 -25.675 157.925 ;
        RECT -26.005 156.235 -25.675 156.565 ;
        RECT -26.005 154.875 -25.675 155.205 ;
        RECT -26.005 153.515 -25.675 153.845 ;
        RECT -26.005 152.155 -25.675 152.485 ;
        RECT -26.005 150.795 -25.675 151.125 ;
        RECT -26.005 149.435 -25.675 149.765 ;
        RECT -26.005 148.075 -25.675 148.405 ;
        RECT -26.005 146.715 -25.675 147.045 ;
        RECT -26.005 145.355 -25.675 145.685 ;
        RECT -26.005 143.995 -25.675 144.325 ;
        RECT -26.005 142.635 -25.675 142.965 ;
        RECT -26.005 141.275 -25.675 141.605 ;
        RECT -26.005 139.915 -25.675 140.245 ;
        RECT -26.005 138.555 -25.675 138.885 ;
        RECT -26.005 137.195 -25.675 137.525 ;
        RECT -26.005 135.835 -25.675 136.165 ;
        RECT -26.005 134.475 -25.675 134.805 ;
        RECT -26.005 133.115 -25.675 133.445 ;
        RECT -26.005 131.755 -25.675 132.085 ;
        RECT -26.005 130.395 -25.675 130.725 ;
        RECT -26.005 129.035 -25.675 129.365 ;
        RECT -26.005 127.675 -25.675 128.005 ;
        RECT -26.005 126.315 -25.675 126.645 ;
        RECT -26.005 124.955 -25.675 125.285 ;
        RECT -26.005 123.595 -25.675 123.925 ;
        RECT -26.005 122.235 -25.675 122.565 ;
        RECT -26.005 120.875 -25.675 121.205 ;
        RECT -26.005 119.515 -25.675 119.845 ;
        RECT -26.005 118.155 -25.675 118.485 ;
        RECT -26.005 116.795 -25.675 117.125 ;
        RECT -26.005 115.435 -25.675 115.765 ;
        RECT -26.005 114.075 -25.675 114.405 ;
        RECT -26.005 112.715 -25.675 113.045 ;
        RECT -26.005 111.355 -25.675 111.685 ;
        RECT -26.005 109.995 -25.675 110.325 ;
        RECT -26.005 108.635 -25.675 108.965 ;
        RECT -26.005 107.275 -25.675 107.605 ;
        RECT -26.005 105.915 -25.675 106.245 ;
        RECT -26.005 104.555 -25.675 104.885 ;
        RECT -26.005 103.195 -25.675 103.525 ;
        RECT -26.005 101.835 -25.675 102.165 ;
        RECT -26.005 100.475 -25.675 100.805 ;
        RECT -26.005 99.115 -25.675 99.445 ;
        RECT -26.005 97.755 -25.675 98.085 ;
        RECT -26.005 96.395 -25.675 96.725 ;
        RECT -26.005 95.035 -25.675 95.365 ;
        RECT -26.005 93.675 -25.675 94.005 ;
        RECT -26.005 92.315 -25.675 92.645 ;
        RECT -26.005 90.955 -25.675 91.285 ;
        RECT -26.005 89.595 -25.675 89.925 ;
        RECT -26.005 88.235 -25.675 88.565 ;
        RECT -26.005 86.875 -25.675 87.205 ;
        RECT -26.005 85.515 -25.675 85.845 ;
        RECT -26.005 84.155 -25.675 84.485 ;
        RECT -26.005 82.795 -25.675 83.125 ;
        RECT -26.005 81.435 -25.675 81.765 ;
        RECT -26.005 80.075 -25.675 80.405 ;
        RECT -26.005 78.715 -25.675 79.045 ;
        RECT -26.005 77.355 -25.675 77.685 ;
        RECT -26.005 75.995 -25.675 76.325 ;
        RECT -26.005 74.635 -25.675 74.965 ;
        RECT -26.005 73.275 -25.675 73.605 ;
        RECT -26.005 71.915 -25.675 72.245 ;
        RECT -26.005 70.555 -25.675 70.885 ;
        RECT -26.005 69.195 -25.675 69.525 ;
        RECT -26.005 67.835 -25.675 68.165 ;
        RECT -26.005 66.475 -25.675 66.805 ;
        RECT -26.005 65.115 -25.675 65.445 ;
        RECT -26.005 63.755 -25.675 64.085 ;
        RECT -26.005 62.395 -25.675 62.725 ;
        RECT -26.005 61.035 -25.675 61.365 ;
        RECT -26.005 59.675 -25.675 60.005 ;
        RECT -26.005 58.315 -25.675 58.645 ;
        RECT -26.005 56.955 -25.675 57.285 ;
        RECT -26.005 55.595 -25.675 55.925 ;
        RECT -26.005 54.235 -25.675 54.565 ;
        RECT -26.005 52.875 -25.675 53.205 ;
        RECT -26.005 51.515 -25.675 51.845 ;
        RECT -26.005 50.155 -25.675 50.485 ;
        RECT -26.005 48.795 -25.675 49.125 ;
        RECT -26.005 47.435 -25.675 47.765 ;
        RECT -26.005 46.075 -25.675 46.405 ;
        RECT -26.005 44.715 -25.675 45.045 ;
        RECT -26.005 43.355 -25.675 43.685 ;
        RECT -26.005 41.995 -25.675 42.325 ;
        RECT -26.005 40.635 -25.675 40.965 ;
        RECT -26.005 39.275 -25.675 39.605 ;
        RECT -26.005 37.915 -25.675 38.245 ;
        RECT -26.005 36.555 -25.675 36.885 ;
        RECT -26.005 35.195 -25.675 35.525 ;
        RECT -26.005 33.835 -25.675 34.165 ;
        RECT -26.005 32.475 -25.675 32.805 ;
        RECT -26.005 31.115 -25.675 31.445 ;
        RECT -26.005 29.755 -25.675 30.085 ;
        RECT -26.005 28.395 -25.675 28.725 ;
        RECT -26.005 27.035 -25.675 27.365 ;
        RECT -26.005 25.675 -25.675 26.005 ;
        RECT -26.005 24.315 -25.675 24.645 ;
        RECT -26.005 22.955 -25.675 23.285 ;
        RECT -26.005 21.595 -25.675 21.925 ;
        RECT -26.005 20.235 -25.675 20.565 ;
        RECT -26.005 18.875 -25.675 19.205 ;
        RECT -26.005 17.515 -25.675 17.845 ;
        RECT -26.005 16.155 -25.675 16.485 ;
        RECT -26.005 14.795 -25.675 15.125 ;
        RECT -26.005 13.435 -25.675 13.765 ;
        RECT -26.005 12.075 -25.675 12.405 ;
        RECT -26.005 10.715 -25.675 11.045 ;
        RECT -26.005 9.355 -25.675 9.685 ;
        RECT -26.005 7.995 -25.675 8.325 ;
        RECT -26.005 6.635 -25.675 6.965 ;
        RECT -26.005 5.275 -25.675 5.605 ;
        RECT -26.005 3.915 -25.675 4.245 ;
        RECT -26.005 2.555 -25.675 2.885 ;
        RECT -26.005 1.195 -25.675 1.525 ;
        RECT -26.005 -0.165 -25.675 0.165 ;
        RECT -26.005 -1.525 -25.675 -1.195 ;
        RECT -26.005 -2.885 -25.675 -2.555 ;
        RECT -26.005 -6.965 -25.675 -6.635 ;
        RECT -26.005 -8.325 -25.675 -7.995 ;
        RECT -26.005 -9.48 -25.675 -9.15 ;
        RECT -26.005 -12.405 -25.675 -12.075 ;
        RECT -26.005 -15.125 -25.675 -14.795 ;
        RECT -26.005 -16.67 -25.675 -16.34 ;
        RECT -26.005 -17.845 -25.675 -17.515 ;
        RECT -26.005 -24.645 -25.675 -24.315 ;
        RECT -26.005 -30.66 -25.675 -30.33 ;
        RECT -26.005 -31.445 -25.675 -31.115 ;
        RECT -26.005 -32.805 -25.675 -32.475 ;
        RECT -26.005 -34.165 -25.675 -33.835 ;
        RECT -26.005 -36.885 -25.675 -36.555 ;
        RECT -26.005 -37.85 -25.675 -37.52 ;
        RECT -26.005 -40.965 -25.675 -40.635 ;
        RECT -26.005 -46.405 -25.675 -46.075 ;
        RECT -26.005 -49.125 -25.675 -48.795 ;
        RECT -26.005 -50.485 -25.675 -50.155 ;
        RECT -26.005 -53.205 -25.675 -52.875 ;
        RECT -26.005 -55.925 -25.675 -55.595 ;
        RECT -26.005 -61.365 -25.675 -61.035 ;
        RECT -26.005 -62.725 -25.675 -62.395 ;
        RECT -26.005 -64.085 -25.675 -63.755 ;
        RECT -26.005 -65.445 -25.675 -65.115 ;
        RECT -26.005 -68.165 -25.675 -67.835 ;
        RECT -26.005 -69.525 -25.675 -69.195 ;
        RECT -26.005 -70.79 -25.675 -70.46 ;
        RECT -26.005 -72.245 -25.675 -71.915 ;
        RECT -26.005 -73.605 -25.675 -73.275 ;
        RECT -26.005 -74.965 -25.675 -74.635 ;
        RECT -26.005 -76.325 -25.675 -75.995 ;
        RECT -26.005 -77.685 -25.675 -77.355 ;
        RECT -26.005 -79.045 -25.675 -78.715 ;
        RECT -26.005 -81.765 -25.675 -81.435 ;
        RECT -26.005 -83.125 -25.675 -82.795 ;
        RECT -26.005 -84.485 -25.675 -84.155 ;
        RECT -26.005 -85.845 -25.675 -85.515 ;
        RECT -26.005 -87.205 -25.675 -86.875 ;
        RECT -26.005 -88.565 -25.675 -88.235 ;
        RECT -26.005 -89.33 -25.675 -89 ;
        RECT -26.005 -91.285 -25.675 -90.955 ;
        RECT -26.005 -92.645 -25.675 -92.315 ;
        RECT -26.005 -94.005 -25.675 -93.675 ;
        RECT -26.005 -95.365 -25.675 -95.035 ;
        RECT -26.005 -96.725 -25.675 -96.395 ;
        RECT -26.005 -98.085 -25.675 -97.755 ;
        RECT -26.005 -100.805 -25.675 -100.475 ;
        RECT -26.005 -102.165 -25.675 -101.835 ;
        RECT -26.005 -103.525 -25.675 -103.195 ;
        RECT -26.005 -106.245 -25.675 -105.915 ;
        RECT -26.005 -107.605 -25.675 -107.275 ;
        RECT -26.005 -108.965 -25.675 -108.635 ;
        RECT -26.005 -110.325 -25.675 -109.995 ;
        RECT -26.005 -111.685 -25.675 -111.355 ;
        RECT -26.005 -113.045 -25.675 -112.715 ;
        RECT -26.005 -114.97 -25.675 -114.64 ;
        RECT -26.005 -115.765 -25.675 -115.435 ;
        RECT -26.005 -117.125 -25.675 -116.795 ;
        RECT -26.005 -118.485 -25.675 -118.155 ;
        RECT -26.005 -119.845 -25.675 -119.515 ;
        RECT -26.005 -121.205 -25.675 -120.875 ;
        RECT -26.005 -122.565 -25.675 -122.235 ;
        RECT -26.005 -129.365 -25.675 -129.035 ;
        RECT -26.005 -130.725 -25.675 -130.395 ;
        RECT -26.005 -132.085 -25.675 -131.755 ;
        RECT -26.005 -133.51 -25.675 -133.18 ;
        RECT -26.005 -136.165 -25.675 -135.835 ;
        RECT -26.005 -137.525 -25.675 -137.195 ;
        RECT -26.005 -138.885 -25.675 -138.555 ;
        RECT -26.005 -140.245 -25.675 -139.915 ;
        RECT -26.005 -141.605 -25.675 -141.275 ;
        RECT -26.005 -144.325 -25.675 -143.995 ;
        RECT -26.005 -145.685 -25.675 -145.355 ;
        RECT -26.005 -147.045 -25.675 -146.715 ;
        RECT -26.005 -152.485 -25.675 -152.155 ;
        RECT -26.005 -153.845 -25.675 -153.515 ;
        RECT -26.005 -155.205 -25.675 -154.875 ;
        RECT -26.005 -156.565 -25.675 -156.235 ;
        RECT -26.005 -157.925 -25.675 -157.595 ;
        RECT -26.005 -159.285 -25.675 -158.955 ;
        RECT -26.005 -162.005 -25.675 -161.675 ;
        RECT -26.005 -163.365 -25.675 -163.035 ;
        RECT -26.005 -164.725 -25.675 -164.395 ;
        RECT -26.005 -166.085 -25.675 -165.755 ;
        RECT -26.005 -167.445 -25.675 -167.115 ;
        RECT -26.005 -168.805 -25.675 -168.475 ;
        RECT -26.005 -170.165 -25.675 -169.835 ;
        RECT -26.005 -171.525 -25.675 -171.195 ;
        RECT -26.005 -172.885 -25.675 -172.555 ;
        RECT -26.005 -174.245 -25.675 -173.915 ;
        RECT -26.005 -175.605 -25.675 -175.275 ;
        RECT -26.005 -176.965 -25.675 -176.635 ;
        RECT -26.005 -178.325 -25.675 -177.995 ;
        RECT -26.005 -179.685 -25.675 -179.355 ;
        RECT -26.005 -181.045 -25.675 -180.715 ;
        RECT -26.005 -182.405 -25.675 -182.075 ;
        RECT -26.005 -185.125 -25.675 -184.795 ;
        RECT -26.005 -186.485 -25.675 -186.155 ;
        RECT -26.005 -191.925 -25.675 -191.595 ;
        RECT -26.005 -193.285 -25.675 -192.955 ;
        RECT -26.005 -194.645 -25.675 -194.315 ;
        RECT -26.005 -196.005 -25.675 -195.675 ;
        RECT -26.005 -198.725 -25.675 -198.395 ;
        RECT -26.005 -200.085 -25.675 -199.755 ;
        RECT -26.005 -201.445 -25.675 -201.115 ;
        RECT -26.005 -204.165 -25.675 -203.835 ;
        RECT -26.005 -205.525 -25.675 -205.195 ;
        RECT -26.005 -209.605 -25.675 -209.275 ;
        RECT -26.005 -215.045 -25.675 -214.715 ;
        RECT -26.005 -216.405 -25.675 -216.075 ;
        RECT -26.005 -217.765 -25.675 -217.435 ;
        RECT -26.005 -219.125 -25.675 -218.795 ;
        RECT -26.005 -220.485 -25.675 -220.155 ;
        RECT -26.005 -221.845 -25.675 -221.515 ;
        RECT -26.005 -223.205 -25.675 -222.875 ;
        RECT -26.005 -224.565 -25.675 -224.235 ;
        RECT -26.005 -226.155 -25.675 -225.825 ;
        RECT -26.005 -227.285 -25.675 -226.955 ;
        RECT -26.005 -230.005 -25.675 -229.675 ;
        RECT -26.005 -231.365 -25.675 -231.035 ;
        RECT -26.005 -234.085 -25.675 -233.755 ;
        RECT -26.005 -235.445 -25.675 -235.115 ;
        RECT -26.005 -236.805 -25.675 -236.475 ;
        RECT -26.005 -238.165 -25.675 -237.835 ;
        RECT -26.005 -243.81 -25.675 -242.68 ;
        RECT -26 -243.925 -25.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.645 246.76 -24.315 247.89 ;
        RECT -24.645 241.915 -24.315 242.245 ;
        RECT -24.645 240.555 -24.315 240.885 ;
        RECT -24.645 239.195 -24.315 239.525 ;
        RECT -24.645 237.835 -24.315 238.165 ;
        RECT -24.645 236.475 -24.315 236.805 ;
        RECT -24.645 235.115 -24.315 235.445 ;
        RECT -24.645 233.755 -24.315 234.085 ;
        RECT -24.645 232.395 -24.315 232.725 ;
        RECT -24.645 231.035 -24.315 231.365 ;
        RECT -24.645 229.675 -24.315 230.005 ;
        RECT -24.645 228.315 -24.315 228.645 ;
        RECT -24.645 226.955 -24.315 227.285 ;
        RECT -24.645 225.595 -24.315 225.925 ;
        RECT -24.645 224.235 -24.315 224.565 ;
        RECT -24.645 222.875 -24.315 223.205 ;
        RECT -24.645 221.515 -24.315 221.845 ;
        RECT -24.645 220.155 -24.315 220.485 ;
        RECT -24.645 218.795 -24.315 219.125 ;
        RECT -24.645 217.435 -24.315 217.765 ;
        RECT -24.645 216.075 -24.315 216.405 ;
        RECT -24.645 214.715 -24.315 215.045 ;
        RECT -24.645 213.355 -24.315 213.685 ;
        RECT -24.645 211.995 -24.315 212.325 ;
        RECT -24.645 210.635 -24.315 210.965 ;
        RECT -24.645 209.275 -24.315 209.605 ;
        RECT -24.645 207.915 -24.315 208.245 ;
        RECT -24.645 206.555 -24.315 206.885 ;
        RECT -24.645 205.195 -24.315 205.525 ;
        RECT -24.645 203.835 -24.315 204.165 ;
        RECT -24.645 202.475 -24.315 202.805 ;
        RECT -24.645 201.115 -24.315 201.445 ;
        RECT -24.645 199.755 -24.315 200.085 ;
        RECT -24.645 198.395 -24.315 198.725 ;
        RECT -24.645 197.035 -24.315 197.365 ;
        RECT -24.645 195.675 -24.315 196.005 ;
        RECT -24.645 194.315 -24.315 194.645 ;
        RECT -24.645 192.955 -24.315 193.285 ;
        RECT -24.645 191.595 -24.315 191.925 ;
        RECT -24.645 190.235 -24.315 190.565 ;
        RECT -24.645 188.875 -24.315 189.205 ;
        RECT -24.645 187.515 -24.315 187.845 ;
        RECT -24.645 186.155 -24.315 186.485 ;
        RECT -24.645 184.795 -24.315 185.125 ;
        RECT -24.645 183.435 -24.315 183.765 ;
        RECT -24.645 182.075 -24.315 182.405 ;
        RECT -24.645 180.715 -24.315 181.045 ;
        RECT -24.645 179.355 -24.315 179.685 ;
        RECT -24.645 177.995 -24.315 178.325 ;
        RECT -24.645 176.635 -24.315 176.965 ;
        RECT -24.645 175.275 -24.315 175.605 ;
        RECT -24.645 173.915 -24.315 174.245 ;
        RECT -24.645 172.555 -24.315 172.885 ;
        RECT -24.645 171.195 -24.315 171.525 ;
        RECT -24.645 169.835 -24.315 170.165 ;
        RECT -24.645 168.475 -24.315 168.805 ;
        RECT -24.645 167.115 -24.315 167.445 ;
        RECT -24.645 165.755 -24.315 166.085 ;
        RECT -24.645 164.395 -24.315 164.725 ;
        RECT -24.645 163.035 -24.315 163.365 ;
        RECT -24.645 161.675 -24.315 162.005 ;
        RECT -24.645 160.315 -24.315 160.645 ;
        RECT -24.645 158.955 -24.315 159.285 ;
        RECT -24.645 157.595 -24.315 157.925 ;
        RECT -24.645 156.235 -24.315 156.565 ;
        RECT -24.645 154.875 -24.315 155.205 ;
        RECT -24.645 153.515 -24.315 153.845 ;
        RECT -24.645 152.155 -24.315 152.485 ;
        RECT -24.645 150.795 -24.315 151.125 ;
        RECT -24.645 149.435 -24.315 149.765 ;
        RECT -24.645 148.075 -24.315 148.405 ;
        RECT -24.645 146.715 -24.315 147.045 ;
        RECT -24.645 145.355 -24.315 145.685 ;
        RECT -24.645 143.995 -24.315 144.325 ;
        RECT -24.645 142.635 -24.315 142.965 ;
        RECT -24.645 141.275 -24.315 141.605 ;
        RECT -24.645 139.915 -24.315 140.245 ;
        RECT -24.645 138.555 -24.315 138.885 ;
        RECT -24.645 137.195 -24.315 137.525 ;
        RECT -24.645 135.835 -24.315 136.165 ;
        RECT -24.645 134.475 -24.315 134.805 ;
        RECT -24.645 133.115 -24.315 133.445 ;
        RECT -24.645 131.755 -24.315 132.085 ;
        RECT -24.645 130.395 -24.315 130.725 ;
        RECT -24.645 129.035 -24.315 129.365 ;
        RECT -24.645 127.675 -24.315 128.005 ;
        RECT -24.645 126.315 -24.315 126.645 ;
        RECT -24.645 124.955 -24.315 125.285 ;
        RECT -24.645 123.595 -24.315 123.925 ;
        RECT -24.645 122.235 -24.315 122.565 ;
        RECT -24.645 120.875 -24.315 121.205 ;
        RECT -24.645 119.515 -24.315 119.845 ;
        RECT -24.645 118.155 -24.315 118.485 ;
        RECT -24.645 116.795 -24.315 117.125 ;
        RECT -24.645 115.435 -24.315 115.765 ;
        RECT -24.645 114.075 -24.315 114.405 ;
        RECT -24.645 112.715 -24.315 113.045 ;
        RECT -24.645 111.355 -24.315 111.685 ;
        RECT -24.645 109.995 -24.315 110.325 ;
        RECT -24.645 108.635 -24.315 108.965 ;
        RECT -24.645 107.275 -24.315 107.605 ;
        RECT -24.645 105.915 -24.315 106.245 ;
        RECT -24.645 104.555 -24.315 104.885 ;
        RECT -24.645 103.195 -24.315 103.525 ;
        RECT -24.645 101.835 -24.315 102.165 ;
        RECT -24.645 100.475 -24.315 100.805 ;
        RECT -24.645 99.115 -24.315 99.445 ;
        RECT -24.645 97.755 -24.315 98.085 ;
        RECT -24.645 96.395 -24.315 96.725 ;
        RECT -24.645 95.035 -24.315 95.365 ;
        RECT -24.645 93.675 -24.315 94.005 ;
        RECT -24.645 92.315 -24.315 92.645 ;
        RECT -24.645 90.955 -24.315 91.285 ;
        RECT -24.645 89.595 -24.315 89.925 ;
        RECT -24.645 88.235 -24.315 88.565 ;
        RECT -24.645 86.875 -24.315 87.205 ;
        RECT -24.645 85.515 -24.315 85.845 ;
        RECT -24.645 84.155 -24.315 84.485 ;
        RECT -24.645 82.795 -24.315 83.125 ;
        RECT -24.645 81.435 -24.315 81.765 ;
        RECT -24.645 80.075 -24.315 80.405 ;
        RECT -24.645 78.715 -24.315 79.045 ;
        RECT -24.645 77.355 -24.315 77.685 ;
        RECT -24.645 75.995 -24.315 76.325 ;
        RECT -24.645 74.635 -24.315 74.965 ;
        RECT -24.645 73.275 -24.315 73.605 ;
        RECT -24.645 71.915 -24.315 72.245 ;
        RECT -24.645 70.555 -24.315 70.885 ;
        RECT -24.645 69.195 -24.315 69.525 ;
        RECT -24.645 67.835 -24.315 68.165 ;
        RECT -24.645 66.475 -24.315 66.805 ;
        RECT -24.645 65.115 -24.315 65.445 ;
        RECT -24.645 63.755 -24.315 64.085 ;
        RECT -24.645 62.395 -24.315 62.725 ;
        RECT -24.645 61.035 -24.315 61.365 ;
        RECT -24.645 59.675 -24.315 60.005 ;
        RECT -24.645 58.315 -24.315 58.645 ;
        RECT -24.645 56.955 -24.315 57.285 ;
        RECT -24.645 55.595 -24.315 55.925 ;
        RECT -24.645 54.235 -24.315 54.565 ;
        RECT -24.645 52.875 -24.315 53.205 ;
        RECT -24.645 51.515 -24.315 51.845 ;
        RECT -24.645 50.155 -24.315 50.485 ;
        RECT -24.645 48.795 -24.315 49.125 ;
        RECT -24.645 47.435 -24.315 47.765 ;
        RECT -24.645 46.075 -24.315 46.405 ;
        RECT -24.645 44.715 -24.315 45.045 ;
        RECT -24.645 43.355 -24.315 43.685 ;
        RECT -24.645 41.995 -24.315 42.325 ;
        RECT -24.645 40.635 -24.315 40.965 ;
        RECT -24.645 39.275 -24.315 39.605 ;
        RECT -24.645 37.915 -24.315 38.245 ;
        RECT -24.645 36.555 -24.315 36.885 ;
        RECT -24.645 35.195 -24.315 35.525 ;
        RECT -24.645 33.835 -24.315 34.165 ;
        RECT -24.645 32.475 -24.315 32.805 ;
        RECT -24.645 31.115 -24.315 31.445 ;
        RECT -24.645 29.755 -24.315 30.085 ;
        RECT -24.645 28.395 -24.315 28.725 ;
        RECT -24.645 27.035 -24.315 27.365 ;
        RECT -24.645 25.675 -24.315 26.005 ;
        RECT -24.645 24.315 -24.315 24.645 ;
        RECT -24.645 22.955 -24.315 23.285 ;
        RECT -24.645 21.595 -24.315 21.925 ;
        RECT -24.645 20.235 -24.315 20.565 ;
        RECT -24.645 18.875 -24.315 19.205 ;
        RECT -24.645 17.515 -24.315 17.845 ;
        RECT -24.645 16.155 -24.315 16.485 ;
        RECT -24.645 14.795 -24.315 15.125 ;
        RECT -24.645 13.435 -24.315 13.765 ;
        RECT -24.645 12.075 -24.315 12.405 ;
        RECT -24.645 10.715 -24.315 11.045 ;
        RECT -24.645 9.355 -24.315 9.685 ;
        RECT -24.645 7.995 -24.315 8.325 ;
        RECT -24.645 6.635 -24.315 6.965 ;
        RECT -24.645 5.275 -24.315 5.605 ;
        RECT -24.645 3.915 -24.315 4.245 ;
        RECT -24.645 2.555 -24.315 2.885 ;
        RECT -24.645 1.195 -24.315 1.525 ;
        RECT -24.645 -0.165 -24.315 0.165 ;
        RECT -24.645 -1.525 -24.315 -1.195 ;
        RECT -24.645 -2.885 -24.315 -2.555 ;
        RECT -24.645 -6.965 -24.315 -6.635 ;
        RECT -24.645 -8.325 -24.315 -7.995 ;
        RECT -24.645 -9.48 -24.315 -9.15 ;
        RECT -24.645 -12.405 -24.315 -12.075 ;
        RECT -24.645 -15.125 -24.315 -14.795 ;
        RECT -24.645 -16.67 -24.315 -16.34 ;
        RECT -24.645 -17.845 -24.315 -17.515 ;
        RECT -24.645 -24.645 -24.315 -24.315 ;
        RECT -24.645 -30.66 -24.315 -30.33 ;
        RECT -24.645 -31.445 -24.315 -31.115 ;
        RECT -24.645 -32.805 -24.315 -32.475 ;
        RECT -24.645 -34.165 -24.315 -33.835 ;
        RECT -24.645 -36.885 -24.315 -36.555 ;
        RECT -24.645 -37.85 -24.315 -37.52 ;
        RECT -24.645 -40.965 -24.315 -40.635 ;
        RECT -24.645 -46.405 -24.315 -46.075 ;
        RECT -24.645 -49.125 -24.315 -48.795 ;
        RECT -24.645 -50.485 -24.315 -50.155 ;
        RECT -24.645 -53.205 -24.315 -52.875 ;
        RECT -24.645 -55.925 -24.315 -55.595 ;
        RECT -24.645 -61.365 -24.315 -61.035 ;
        RECT -24.645 -62.725 -24.315 -62.395 ;
        RECT -24.645 -64.085 -24.315 -63.755 ;
        RECT -24.645 -65.445 -24.315 -65.115 ;
        RECT -24.645 -68.165 -24.315 -67.835 ;
        RECT -24.645 -69.525 -24.315 -69.195 ;
        RECT -24.645 -70.79 -24.315 -70.46 ;
        RECT -24.645 -72.245 -24.315 -71.915 ;
        RECT -24.645 -73.605 -24.315 -73.275 ;
        RECT -24.645 -74.965 -24.315 -74.635 ;
        RECT -24.645 -76.325 -24.315 -75.995 ;
        RECT -24.645 -77.685 -24.315 -77.355 ;
        RECT -24.645 -79.045 -24.315 -78.715 ;
        RECT -24.645 -81.765 -24.315 -81.435 ;
        RECT -24.645 -83.125 -24.315 -82.795 ;
        RECT -24.645 -84.485 -24.315 -84.155 ;
        RECT -24.645 -85.845 -24.315 -85.515 ;
        RECT -24.645 -87.205 -24.315 -86.875 ;
        RECT -24.645 -88.565 -24.315 -88.235 ;
        RECT -24.645 -89.33 -24.315 -89 ;
        RECT -24.645 -91.285 -24.315 -90.955 ;
        RECT -24.645 -92.645 -24.315 -92.315 ;
        RECT -24.645 -94.005 -24.315 -93.675 ;
        RECT -24.645 -95.365 -24.315 -95.035 ;
        RECT -24.645 -96.725 -24.315 -96.395 ;
        RECT -24.645 -98.085 -24.315 -97.755 ;
        RECT -24.645 -100.805 -24.315 -100.475 ;
        RECT -24.645 -102.165 -24.315 -101.835 ;
        RECT -24.645 -103.525 -24.315 -103.195 ;
        RECT -24.645 -106.245 -24.315 -105.915 ;
        RECT -24.645 -107.605 -24.315 -107.275 ;
        RECT -24.645 -108.965 -24.315 -108.635 ;
        RECT -24.645 -110.325 -24.315 -109.995 ;
        RECT -24.645 -111.685 -24.315 -111.355 ;
        RECT -24.645 -113.045 -24.315 -112.715 ;
        RECT -24.645 -114.97 -24.315 -114.64 ;
        RECT -24.645 -115.765 -24.315 -115.435 ;
        RECT -24.645 -117.125 -24.315 -116.795 ;
        RECT -24.645 -118.485 -24.315 -118.155 ;
        RECT -24.645 -119.845 -24.315 -119.515 ;
        RECT -24.645 -121.205 -24.315 -120.875 ;
        RECT -24.645 -122.565 -24.315 -122.235 ;
        RECT -24.645 -129.365 -24.315 -129.035 ;
        RECT -24.645 -130.725 -24.315 -130.395 ;
        RECT -24.645 -132.085 -24.315 -131.755 ;
        RECT -24.645 -133.51 -24.315 -133.18 ;
        RECT -24.645 -136.165 -24.315 -135.835 ;
        RECT -24.645 -137.525 -24.315 -137.195 ;
        RECT -24.645 -138.885 -24.315 -138.555 ;
        RECT -24.645 -140.245 -24.315 -139.915 ;
        RECT -24.645 -141.605 -24.315 -141.275 ;
        RECT -24.645 -144.325 -24.315 -143.995 ;
        RECT -24.645 -145.685 -24.315 -145.355 ;
        RECT -24.645 -147.045 -24.315 -146.715 ;
        RECT -24.645 -152.485 -24.315 -152.155 ;
        RECT -24.645 -153.845 -24.315 -153.515 ;
        RECT -24.645 -155.205 -24.315 -154.875 ;
        RECT -24.645 -156.565 -24.315 -156.235 ;
        RECT -24.645 -157.925 -24.315 -157.595 ;
        RECT -24.645 -159.285 -24.315 -158.955 ;
        RECT -24.645 -162.005 -24.315 -161.675 ;
        RECT -24.645 -163.365 -24.315 -163.035 ;
        RECT -24.645 -164.725 -24.315 -164.395 ;
        RECT -24.645 -166.085 -24.315 -165.755 ;
        RECT -24.645 -167.445 -24.315 -167.115 ;
        RECT -24.645 -168.805 -24.315 -168.475 ;
        RECT -24.645 -170.165 -24.315 -169.835 ;
        RECT -24.645 -171.525 -24.315 -171.195 ;
        RECT -24.645 -172.885 -24.315 -172.555 ;
        RECT -24.645 -174.245 -24.315 -173.915 ;
        RECT -24.645 -175.605 -24.315 -175.275 ;
        RECT -24.645 -176.965 -24.315 -176.635 ;
        RECT -24.645 -178.325 -24.315 -177.995 ;
        RECT -24.645 -179.685 -24.315 -179.355 ;
        RECT -24.645 -181.045 -24.315 -180.715 ;
        RECT -24.645 -182.405 -24.315 -182.075 ;
        RECT -24.645 -185.125 -24.315 -184.795 ;
        RECT -24.645 -186.485 -24.315 -186.155 ;
        RECT -24.645 -191.925 -24.315 -191.595 ;
        RECT -24.645 -193.285 -24.315 -192.955 ;
        RECT -24.645 -194.645 -24.315 -194.315 ;
        RECT -24.645 -196.005 -24.315 -195.675 ;
        RECT -24.645 -198.725 -24.315 -198.395 ;
        RECT -24.645 -200.085 -24.315 -199.755 ;
        RECT -24.645 -201.445 -24.315 -201.115 ;
        RECT -24.645 -204.165 -24.315 -203.835 ;
        RECT -24.645 -205.525 -24.315 -205.195 ;
        RECT -24.645 -209.605 -24.315 -209.275 ;
        RECT -24.645 -215.045 -24.315 -214.715 ;
        RECT -24.645 -216.405 -24.315 -216.075 ;
        RECT -24.645 -217.765 -24.315 -217.435 ;
        RECT -24.645 -219.125 -24.315 -218.795 ;
        RECT -24.645 -220.485 -24.315 -220.155 ;
        RECT -24.645 -221.845 -24.315 -221.515 ;
        RECT -24.645 -223.205 -24.315 -222.875 ;
        RECT -24.645 -224.565 -24.315 -224.235 ;
        RECT -24.645 -226.155 -24.315 -225.825 ;
        RECT -24.645 -227.285 -24.315 -226.955 ;
        RECT -24.645 -230.005 -24.315 -229.675 ;
        RECT -24.645 -231.365 -24.315 -231.035 ;
        RECT -24.645 -234.085 -24.315 -233.755 ;
        RECT -24.645 -235.445 -24.315 -235.115 ;
        RECT -24.645 -236.805 -24.315 -236.475 ;
        RECT -24.645 -238.165 -24.315 -237.835 ;
        RECT -24.645 -243.81 -24.315 -242.68 ;
        RECT -24.64 -243.925 -24.32 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 246.76 -22.955 247.89 ;
        RECT -23.285 241.915 -22.955 242.245 ;
        RECT -23.285 240.555 -22.955 240.885 ;
        RECT -23.285 239.195 -22.955 239.525 ;
        RECT -23.285 237.835 -22.955 238.165 ;
        RECT -23.285 236.475 -22.955 236.805 ;
        RECT -23.285 235.115 -22.955 235.445 ;
        RECT -23.285 233.755 -22.955 234.085 ;
        RECT -23.285 232.395 -22.955 232.725 ;
        RECT -23.285 231.035 -22.955 231.365 ;
        RECT -23.285 229.675 -22.955 230.005 ;
        RECT -23.285 228.315 -22.955 228.645 ;
        RECT -23.285 226.955 -22.955 227.285 ;
        RECT -23.285 225.595 -22.955 225.925 ;
        RECT -23.285 224.235 -22.955 224.565 ;
        RECT -23.285 222.875 -22.955 223.205 ;
        RECT -23.285 221.515 -22.955 221.845 ;
        RECT -23.285 220.155 -22.955 220.485 ;
        RECT -23.285 218.795 -22.955 219.125 ;
        RECT -23.285 217.435 -22.955 217.765 ;
        RECT -23.285 216.075 -22.955 216.405 ;
        RECT -23.285 214.715 -22.955 215.045 ;
        RECT -23.285 213.355 -22.955 213.685 ;
        RECT -23.285 211.995 -22.955 212.325 ;
        RECT -23.285 210.635 -22.955 210.965 ;
        RECT -23.285 209.275 -22.955 209.605 ;
        RECT -23.285 207.915 -22.955 208.245 ;
        RECT -23.285 206.555 -22.955 206.885 ;
        RECT -23.285 205.195 -22.955 205.525 ;
        RECT -23.285 203.835 -22.955 204.165 ;
        RECT -23.285 202.475 -22.955 202.805 ;
        RECT -23.285 201.115 -22.955 201.445 ;
        RECT -23.285 199.755 -22.955 200.085 ;
        RECT -23.285 198.395 -22.955 198.725 ;
        RECT -23.285 197.035 -22.955 197.365 ;
        RECT -23.285 195.675 -22.955 196.005 ;
        RECT -23.285 194.315 -22.955 194.645 ;
        RECT -23.285 192.955 -22.955 193.285 ;
        RECT -23.285 191.595 -22.955 191.925 ;
        RECT -23.285 190.235 -22.955 190.565 ;
        RECT -23.285 188.875 -22.955 189.205 ;
        RECT -23.285 187.515 -22.955 187.845 ;
        RECT -23.285 186.155 -22.955 186.485 ;
        RECT -23.285 184.795 -22.955 185.125 ;
        RECT -23.285 183.435 -22.955 183.765 ;
        RECT -23.285 182.075 -22.955 182.405 ;
        RECT -23.285 180.715 -22.955 181.045 ;
        RECT -23.285 179.355 -22.955 179.685 ;
        RECT -23.285 177.995 -22.955 178.325 ;
        RECT -23.285 176.635 -22.955 176.965 ;
        RECT -23.285 175.275 -22.955 175.605 ;
        RECT -23.285 173.915 -22.955 174.245 ;
        RECT -23.285 172.555 -22.955 172.885 ;
        RECT -23.285 171.195 -22.955 171.525 ;
        RECT -23.285 169.835 -22.955 170.165 ;
        RECT -23.285 168.475 -22.955 168.805 ;
        RECT -23.285 167.115 -22.955 167.445 ;
        RECT -23.285 165.755 -22.955 166.085 ;
        RECT -23.285 164.395 -22.955 164.725 ;
        RECT -23.285 163.035 -22.955 163.365 ;
        RECT -23.285 161.675 -22.955 162.005 ;
        RECT -23.285 160.315 -22.955 160.645 ;
        RECT -23.285 158.955 -22.955 159.285 ;
        RECT -23.285 157.595 -22.955 157.925 ;
        RECT -23.285 156.235 -22.955 156.565 ;
        RECT -23.285 154.875 -22.955 155.205 ;
        RECT -23.285 153.515 -22.955 153.845 ;
        RECT -23.285 152.155 -22.955 152.485 ;
        RECT -23.285 150.795 -22.955 151.125 ;
        RECT -23.285 149.435 -22.955 149.765 ;
        RECT -23.285 148.075 -22.955 148.405 ;
        RECT -23.285 146.715 -22.955 147.045 ;
        RECT -23.285 145.355 -22.955 145.685 ;
        RECT -23.285 143.995 -22.955 144.325 ;
        RECT -23.285 142.635 -22.955 142.965 ;
        RECT -23.285 141.275 -22.955 141.605 ;
        RECT -23.285 139.915 -22.955 140.245 ;
        RECT -23.285 138.555 -22.955 138.885 ;
        RECT -23.285 137.195 -22.955 137.525 ;
        RECT -23.285 135.835 -22.955 136.165 ;
        RECT -23.285 134.475 -22.955 134.805 ;
        RECT -23.285 133.115 -22.955 133.445 ;
        RECT -23.285 131.755 -22.955 132.085 ;
        RECT -23.285 130.395 -22.955 130.725 ;
        RECT -23.285 129.035 -22.955 129.365 ;
        RECT -23.285 127.675 -22.955 128.005 ;
        RECT -23.285 126.315 -22.955 126.645 ;
        RECT -23.285 124.955 -22.955 125.285 ;
        RECT -23.285 123.595 -22.955 123.925 ;
        RECT -23.285 122.235 -22.955 122.565 ;
        RECT -23.285 120.875 -22.955 121.205 ;
        RECT -23.285 119.515 -22.955 119.845 ;
        RECT -23.285 118.155 -22.955 118.485 ;
        RECT -23.285 116.795 -22.955 117.125 ;
        RECT -23.285 115.435 -22.955 115.765 ;
        RECT -23.285 114.075 -22.955 114.405 ;
        RECT -23.285 112.715 -22.955 113.045 ;
        RECT -23.285 111.355 -22.955 111.685 ;
        RECT -23.285 109.995 -22.955 110.325 ;
        RECT -23.285 108.635 -22.955 108.965 ;
        RECT -23.285 107.275 -22.955 107.605 ;
        RECT -23.285 105.915 -22.955 106.245 ;
        RECT -23.285 104.555 -22.955 104.885 ;
        RECT -23.285 103.195 -22.955 103.525 ;
        RECT -23.285 101.835 -22.955 102.165 ;
        RECT -23.285 100.475 -22.955 100.805 ;
        RECT -23.285 99.115 -22.955 99.445 ;
        RECT -23.285 97.755 -22.955 98.085 ;
        RECT -23.285 96.395 -22.955 96.725 ;
        RECT -23.285 95.035 -22.955 95.365 ;
        RECT -23.285 93.675 -22.955 94.005 ;
        RECT -23.285 92.315 -22.955 92.645 ;
        RECT -23.285 90.955 -22.955 91.285 ;
        RECT -23.285 89.595 -22.955 89.925 ;
        RECT -23.285 88.235 -22.955 88.565 ;
        RECT -23.285 86.875 -22.955 87.205 ;
        RECT -23.285 85.515 -22.955 85.845 ;
        RECT -23.285 84.155 -22.955 84.485 ;
        RECT -23.285 82.795 -22.955 83.125 ;
        RECT -23.285 81.435 -22.955 81.765 ;
        RECT -23.285 80.075 -22.955 80.405 ;
        RECT -23.285 78.715 -22.955 79.045 ;
        RECT -23.285 77.355 -22.955 77.685 ;
        RECT -23.285 75.995 -22.955 76.325 ;
        RECT -23.285 74.635 -22.955 74.965 ;
        RECT -23.285 73.275 -22.955 73.605 ;
        RECT -23.285 71.915 -22.955 72.245 ;
        RECT -23.285 70.555 -22.955 70.885 ;
        RECT -23.285 69.195 -22.955 69.525 ;
        RECT -23.285 67.835 -22.955 68.165 ;
        RECT -23.285 66.475 -22.955 66.805 ;
        RECT -23.285 65.115 -22.955 65.445 ;
        RECT -23.285 63.755 -22.955 64.085 ;
        RECT -23.285 62.395 -22.955 62.725 ;
        RECT -23.285 61.035 -22.955 61.365 ;
        RECT -23.285 59.675 -22.955 60.005 ;
        RECT -23.285 58.315 -22.955 58.645 ;
        RECT -23.285 56.955 -22.955 57.285 ;
        RECT -23.285 55.595 -22.955 55.925 ;
        RECT -23.285 54.235 -22.955 54.565 ;
        RECT -23.285 52.875 -22.955 53.205 ;
        RECT -23.285 51.515 -22.955 51.845 ;
        RECT -23.285 50.155 -22.955 50.485 ;
        RECT -23.285 48.795 -22.955 49.125 ;
        RECT -23.285 47.435 -22.955 47.765 ;
        RECT -23.285 46.075 -22.955 46.405 ;
        RECT -23.285 44.715 -22.955 45.045 ;
        RECT -23.285 43.355 -22.955 43.685 ;
        RECT -23.285 41.995 -22.955 42.325 ;
        RECT -23.285 40.635 -22.955 40.965 ;
        RECT -23.285 39.275 -22.955 39.605 ;
        RECT -23.285 37.915 -22.955 38.245 ;
        RECT -23.285 36.555 -22.955 36.885 ;
        RECT -23.285 35.195 -22.955 35.525 ;
        RECT -23.285 33.835 -22.955 34.165 ;
        RECT -23.285 32.475 -22.955 32.805 ;
        RECT -23.285 31.115 -22.955 31.445 ;
        RECT -23.285 29.755 -22.955 30.085 ;
        RECT -23.285 28.395 -22.955 28.725 ;
        RECT -23.285 27.035 -22.955 27.365 ;
        RECT -23.285 25.675 -22.955 26.005 ;
        RECT -23.285 24.315 -22.955 24.645 ;
        RECT -23.285 22.955 -22.955 23.285 ;
        RECT -23.285 21.595 -22.955 21.925 ;
        RECT -23.285 20.235 -22.955 20.565 ;
        RECT -23.285 18.875 -22.955 19.205 ;
        RECT -23.285 17.515 -22.955 17.845 ;
        RECT -23.285 16.155 -22.955 16.485 ;
        RECT -23.285 14.795 -22.955 15.125 ;
        RECT -23.285 13.435 -22.955 13.765 ;
        RECT -23.285 12.075 -22.955 12.405 ;
        RECT -23.285 10.715 -22.955 11.045 ;
        RECT -23.285 9.355 -22.955 9.685 ;
        RECT -23.285 7.995 -22.955 8.325 ;
        RECT -23.285 6.635 -22.955 6.965 ;
        RECT -23.285 5.275 -22.955 5.605 ;
        RECT -23.285 3.915 -22.955 4.245 ;
        RECT -23.285 2.555 -22.955 2.885 ;
        RECT -23.285 1.195 -22.955 1.525 ;
        RECT -23.285 -0.165 -22.955 0.165 ;
        RECT -23.285 -1.525 -22.955 -1.195 ;
        RECT -23.285 -2.885 -22.955 -2.555 ;
        RECT -23.285 -6.965 -22.955 -6.635 ;
        RECT -23.285 -8.325 -22.955 -7.995 ;
        RECT -23.285 -9.48 -22.955 -9.15 ;
        RECT -23.285 -12.405 -22.955 -12.075 ;
        RECT -23.285 -15.125 -22.955 -14.795 ;
        RECT -23.285 -16.67 -22.955 -16.34 ;
        RECT -23.285 -17.845 -22.955 -17.515 ;
        RECT -23.285 -24.645 -22.955 -24.315 ;
        RECT -23.285 -30.66 -22.955 -30.33 ;
        RECT -23.285 -31.445 -22.955 -31.115 ;
        RECT -23.285 -32.805 -22.955 -32.475 ;
        RECT -23.285 -34.165 -22.955 -33.835 ;
        RECT -23.285 -36.885 -22.955 -36.555 ;
        RECT -23.285 -37.85 -22.955 -37.52 ;
        RECT -23.285 -40.965 -22.955 -40.635 ;
        RECT -23.285 -46.405 -22.955 -46.075 ;
        RECT -23.285 -47.765 -22.955 -47.435 ;
        RECT -23.285 -49.125 -22.955 -48.795 ;
        RECT -23.285 -50.485 -22.955 -50.155 ;
        RECT -23.285 -51.845 -22.955 -51.515 ;
        RECT -23.285 -53.205 -22.955 -52.875 ;
        RECT -23.285 -54.565 -22.955 -54.235 ;
        RECT -23.285 -55.925 -22.955 -55.595 ;
        RECT -23.285 -57.285 -22.955 -56.955 ;
        RECT -23.285 -58.645 -22.955 -58.315 ;
        RECT -23.285 -60.005 -22.955 -59.675 ;
        RECT -23.285 -61.365 -22.955 -61.035 ;
        RECT -23.285 -62.725 -22.955 -62.395 ;
        RECT -23.285 -64.085 -22.955 -63.755 ;
        RECT -23.285 -65.445 -22.955 -65.115 ;
        RECT -23.285 -68.165 -22.955 -67.835 ;
        RECT -23.285 -69.525 -22.955 -69.195 ;
        RECT -23.285 -70.79 -22.955 -70.46 ;
        RECT -23.285 -72.245 -22.955 -71.915 ;
        RECT -23.285 -73.605 -22.955 -73.275 ;
        RECT -23.285 -74.965 -22.955 -74.635 ;
        RECT -23.285 -76.325 -22.955 -75.995 ;
        RECT -23.285 -77.685 -22.955 -77.355 ;
        RECT -23.285 -79.045 -22.955 -78.715 ;
        RECT -23.285 -81.765 -22.955 -81.435 ;
        RECT -23.285 -83.125 -22.955 -82.795 ;
        RECT -23.285 -84.485 -22.955 -84.155 ;
        RECT -23.285 -85.845 -22.955 -85.515 ;
        RECT -23.285 -87.205 -22.955 -86.875 ;
        RECT -23.285 -88.565 -22.955 -88.235 ;
        RECT -23.285 -89.33 -22.955 -89 ;
        RECT -23.285 -91.285 -22.955 -90.955 ;
        RECT -23.285 -92.645 -22.955 -92.315 ;
        RECT -23.285 -94.005 -22.955 -93.675 ;
        RECT -23.285 -95.365 -22.955 -95.035 ;
        RECT -23.285 -96.725 -22.955 -96.395 ;
        RECT -23.285 -98.085 -22.955 -97.755 ;
        RECT -23.285 -100.805 -22.955 -100.475 ;
        RECT -23.285 -102.165 -22.955 -101.835 ;
        RECT -23.285 -103.525 -22.955 -103.195 ;
        RECT -23.285 -106.245 -22.955 -105.915 ;
        RECT -23.285 -107.605 -22.955 -107.275 ;
        RECT -23.285 -108.965 -22.955 -108.635 ;
        RECT -23.285 -110.325 -22.955 -109.995 ;
        RECT -23.285 -111.685 -22.955 -111.355 ;
        RECT -23.285 -113.045 -22.955 -112.715 ;
        RECT -23.285 -114.97 -22.955 -114.64 ;
        RECT -23.285 -115.765 -22.955 -115.435 ;
        RECT -23.285 -117.125 -22.955 -116.795 ;
        RECT -23.285 -118.485 -22.955 -118.155 ;
        RECT -23.285 -119.845 -22.955 -119.515 ;
        RECT -23.285 -121.205 -22.955 -120.875 ;
        RECT -23.285 -122.565 -22.955 -122.235 ;
        RECT -23.285 -129.365 -22.955 -129.035 ;
        RECT -23.285 -130.725 -22.955 -130.395 ;
        RECT -23.285 -132.085 -22.955 -131.755 ;
        RECT -23.285 -133.51 -22.955 -133.18 ;
        RECT -23.285 -137.525 -22.955 -137.195 ;
        RECT -23.285 -138.885 -22.955 -138.555 ;
        RECT -23.285 -140.245 -22.955 -139.915 ;
        RECT -23.285 -141.605 -22.955 -141.275 ;
        RECT -23.285 -144.325 -22.955 -143.995 ;
        RECT -23.285 -145.685 -22.955 -145.355 ;
        RECT -23.285 -147.045 -22.955 -146.715 ;
        RECT -23.285 -152.485 -22.955 -152.155 ;
        RECT -23.285 -153.845 -22.955 -153.515 ;
        RECT -23.285 -155.205 -22.955 -154.875 ;
        RECT -23.285 -156.565 -22.955 -156.235 ;
        RECT -23.285 -157.925 -22.955 -157.595 ;
        RECT -23.285 -159.285 -22.955 -158.955 ;
        RECT -23.285 -162.005 -22.955 -161.675 ;
        RECT -23.285 -163.365 -22.955 -163.035 ;
        RECT -23.285 -164.725 -22.955 -164.395 ;
        RECT -23.285 -166.085 -22.955 -165.755 ;
        RECT -23.285 -167.445 -22.955 -167.115 ;
        RECT -23.285 -168.805 -22.955 -168.475 ;
        RECT -23.285 -170.165 -22.955 -169.835 ;
        RECT -23.285 -171.525 -22.955 -171.195 ;
        RECT -23.285 -174.245 -22.955 -173.915 ;
        RECT -23.285 -175.605 -22.955 -175.275 ;
        RECT -23.285 -176.965 -22.955 -176.635 ;
        RECT -23.285 -178.325 -22.955 -177.995 ;
        RECT -23.285 -179.685 -22.955 -179.355 ;
        RECT -23.285 -181.045 -22.955 -180.715 ;
        RECT -23.285 -182.405 -22.955 -182.075 ;
        RECT -23.285 -185.125 -22.955 -184.795 ;
        RECT -23.285 -191.925 -22.955 -191.595 ;
        RECT -23.285 -193.285 -22.955 -192.955 ;
        RECT -23.285 -194.645 -22.955 -194.315 ;
        RECT -23.285 -196.005 -22.955 -195.675 ;
        RECT -23.285 -198.725 -22.955 -198.395 ;
        RECT -23.285 -200.085 -22.955 -199.755 ;
        RECT -23.285 -202.805 -22.955 -202.475 ;
        RECT -23.285 -204.165 -22.955 -203.835 ;
        RECT -23.285 -205.525 -22.955 -205.195 ;
        RECT -23.285 -209.605 -22.955 -209.275 ;
        RECT -23.285 -215.045 -22.955 -214.715 ;
        RECT -23.285 -216.405 -22.955 -216.075 ;
        RECT -23.285 -217.765 -22.955 -217.435 ;
        RECT -23.285 -219.125 -22.955 -218.795 ;
        RECT -23.285 -220.485 -22.955 -220.155 ;
        RECT -23.285 -221.845 -22.955 -221.515 ;
        RECT -23.285 -223.205 -22.955 -222.875 ;
        RECT -23.285 -224.565 -22.955 -224.235 ;
        RECT -23.285 -226.155 -22.955 -225.825 ;
        RECT -23.28 -226.6 -22.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 -234.085 -22.955 -233.755 ;
        RECT -23.285 -235.445 -22.955 -235.115 ;
        RECT -23.285 -236.805 -22.955 -236.475 ;
        RECT -23.285 -238.165 -22.955 -237.835 ;
        RECT -23.285 -243.81 -22.955 -242.68 ;
        RECT -23.28 -243.925 -22.96 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 13.435 -21.595 13.765 ;
        RECT -21.925 12.075 -21.595 12.405 ;
        RECT -21.925 10.715 -21.595 11.045 ;
        RECT -21.925 9.355 -21.595 9.685 ;
        RECT -21.925 7.995 -21.595 8.325 ;
        RECT -21.925 6.635 -21.595 6.965 ;
        RECT -21.925 5.275 -21.595 5.605 ;
        RECT -21.925 3.915 -21.595 4.245 ;
        RECT -21.925 2.555 -21.595 2.885 ;
        RECT -21.925 1.195 -21.595 1.525 ;
        RECT -21.925 -0.165 -21.595 0.165 ;
        RECT -21.925 -1.525 -21.595 -1.195 ;
        RECT -21.925 -2.885 -21.595 -2.555 ;
        RECT -21.925 -4.245 -21.595 -3.915 ;
        RECT -21.925 -6.965 -21.595 -6.635 ;
        RECT -21.925 -8.325 -21.595 -7.995 ;
        RECT -21.925 -9.48 -21.595 -9.15 ;
        RECT -21.925 -12.405 -21.595 -12.075 ;
        RECT -21.925 -15.125 -21.595 -14.795 ;
        RECT -21.925 -16.67 -21.595 -16.34 ;
        RECT -21.925 -17.845 -21.595 -17.515 ;
        RECT -21.92 -21.92 -21.6 248.005 ;
        RECT -21.925 246.76 -21.595 247.89 ;
        RECT -21.925 241.915 -21.595 242.245 ;
        RECT -21.925 240.555 -21.595 240.885 ;
        RECT -21.925 239.195 -21.595 239.525 ;
        RECT -21.925 237.835 -21.595 238.165 ;
        RECT -21.925 236.475 -21.595 236.805 ;
        RECT -21.925 235.115 -21.595 235.445 ;
        RECT -21.925 233.755 -21.595 234.085 ;
        RECT -21.925 232.395 -21.595 232.725 ;
        RECT -21.925 231.035 -21.595 231.365 ;
        RECT -21.925 229.675 -21.595 230.005 ;
        RECT -21.925 228.315 -21.595 228.645 ;
        RECT -21.925 226.955 -21.595 227.285 ;
        RECT -21.925 225.595 -21.595 225.925 ;
        RECT -21.925 224.235 -21.595 224.565 ;
        RECT -21.925 222.875 -21.595 223.205 ;
        RECT -21.925 221.515 -21.595 221.845 ;
        RECT -21.925 220.155 -21.595 220.485 ;
        RECT -21.925 218.795 -21.595 219.125 ;
        RECT -21.925 217.435 -21.595 217.765 ;
        RECT -21.925 216.075 -21.595 216.405 ;
        RECT -21.925 214.715 -21.595 215.045 ;
        RECT -21.925 213.355 -21.595 213.685 ;
        RECT -21.925 211.995 -21.595 212.325 ;
        RECT -21.925 210.635 -21.595 210.965 ;
        RECT -21.925 209.275 -21.595 209.605 ;
        RECT -21.925 207.915 -21.595 208.245 ;
        RECT -21.925 206.555 -21.595 206.885 ;
        RECT -21.925 205.195 -21.595 205.525 ;
        RECT -21.925 203.835 -21.595 204.165 ;
        RECT -21.925 202.475 -21.595 202.805 ;
        RECT -21.925 201.115 -21.595 201.445 ;
        RECT -21.925 199.755 -21.595 200.085 ;
        RECT -21.925 198.395 -21.595 198.725 ;
        RECT -21.925 197.035 -21.595 197.365 ;
        RECT -21.925 195.675 -21.595 196.005 ;
        RECT -21.925 194.315 -21.595 194.645 ;
        RECT -21.925 192.955 -21.595 193.285 ;
        RECT -21.925 191.595 -21.595 191.925 ;
        RECT -21.925 190.235 -21.595 190.565 ;
        RECT -21.925 188.875 -21.595 189.205 ;
        RECT -21.925 187.515 -21.595 187.845 ;
        RECT -21.925 186.155 -21.595 186.485 ;
        RECT -21.925 184.795 -21.595 185.125 ;
        RECT -21.925 183.435 -21.595 183.765 ;
        RECT -21.925 182.075 -21.595 182.405 ;
        RECT -21.925 180.715 -21.595 181.045 ;
        RECT -21.925 179.355 -21.595 179.685 ;
        RECT -21.925 177.995 -21.595 178.325 ;
        RECT -21.925 176.635 -21.595 176.965 ;
        RECT -21.925 175.275 -21.595 175.605 ;
        RECT -21.925 173.915 -21.595 174.245 ;
        RECT -21.925 172.555 -21.595 172.885 ;
        RECT -21.925 171.195 -21.595 171.525 ;
        RECT -21.925 169.835 -21.595 170.165 ;
        RECT -21.925 168.475 -21.595 168.805 ;
        RECT -21.925 167.115 -21.595 167.445 ;
        RECT -21.925 165.755 -21.595 166.085 ;
        RECT -21.925 164.395 -21.595 164.725 ;
        RECT -21.925 163.035 -21.595 163.365 ;
        RECT -21.925 161.675 -21.595 162.005 ;
        RECT -21.925 160.315 -21.595 160.645 ;
        RECT -21.925 158.955 -21.595 159.285 ;
        RECT -21.925 157.595 -21.595 157.925 ;
        RECT -21.925 156.235 -21.595 156.565 ;
        RECT -21.925 154.875 -21.595 155.205 ;
        RECT -21.925 153.515 -21.595 153.845 ;
        RECT -21.925 152.155 -21.595 152.485 ;
        RECT -21.925 150.795 -21.595 151.125 ;
        RECT -21.925 149.435 -21.595 149.765 ;
        RECT -21.925 148.075 -21.595 148.405 ;
        RECT -21.925 146.715 -21.595 147.045 ;
        RECT -21.925 145.355 -21.595 145.685 ;
        RECT -21.925 143.995 -21.595 144.325 ;
        RECT -21.925 142.635 -21.595 142.965 ;
        RECT -21.925 141.275 -21.595 141.605 ;
        RECT -21.925 139.915 -21.595 140.245 ;
        RECT -21.925 138.555 -21.595 138.885 ;
        RECT -21.925 137.195 -21.595 137.525 ;
        RECT -21.925 135.835 -21.595 136.165 ;
        RECT -21.925 134.475 -21.595 134.805 ;
        RECT -21.925 133.115 -21.595 133.445 ;
        RECT -21.925 131.755 -21.595 132.085 ;
        RECT -21.925 130.395 -21.595 130.725 ;
        RECT -21.925 129.035 -21.595 129.365 ;
        RECT -21.925 127.675 -21.595 128.005 ;
        RECT -21.925 126.315 -21.595 126.645 ;
        RECT -21.925 124.955 -21.595 125.285 ;
        RECT -21.925 123.595 -21.595 123.925 ;
        RECT -21.925 122.235 -21.595 122.565 ;
        RECT -21.925 120.875 -21.595 121.205 ;
        RECT -21.925 119.515 -21.595 119.845 ;
        RECT -21.925 118.155 -21.595 118.485 ;
        RECT -21.925 116.795 -21.595 117.125 ;
        RECT -21.925 115.435 -21.595 115.765 ;
        RECT -21.925 114.075 -21.595 114.405 ;
        RECT -21.925 112.715 -21.595 113.045 ;
        RECT -21.925 111.355 -21.595 111.685 ;
        RECT -21.925 109.995 -21.595 110.325 ;
        RECT -21.925 108.635 -21.595 108.965 ;
        RECT -21.925 107.275 -21.595 107.605 ;
        RECT -21.925 105.915 -21.595 106.245 ;
        RECT -21.925 104.555 -21.595 104.885 ;
        RECT -21.925 103.195 -21.595 103.525 ;
        RECT -21.925 101.835 -21.595 102.165 ;
        RECT -21.925 100.475 -21.595 100.805 ;
        RECT -21.925 99.115 -21.595 99.445 ;
        RECT -21.925 97.755 -21.595 98.085 ;
        RECT -21.925 96.395 -21.595 96.725 ;
        RECT -21.925 95.035 -21.595 95.365 ;
        RECT -21.925 93.675 -21.595 94.005 ;
        RECT -21.925 92.315 -21.595 92.645 ;
        RECT -21.925 90.955 -21.595 91.285 ;
        RECT -21.925 89.595 -21.595 89.925 ;
        RECT -21.925 88.235 -21.595 88.565 ;
        RECT -21.925 86.875 -21.595 87.205 ;
        RECT -21.925 85.515 -21.595 85.845 ;
        RECT -21.925 84.155 -21.595 84.485 ;
        RECT -21.925 82.795 -21.595 83.125 ;
        RECT -21.925 81.435 -21.595 81.765 ;
        RECT -21.925 80.075 -21.595 80.405 ;
        RECT -21.925 78.715 -21.595 79.045 ;
        RECT -21.925 77.355 -21.595 77.685 ;
        RECT -21.925 75.995 -21.595 76.325 ;
        RECT -21.925 74.635 -21.595 74.965 ;
        RECT -21.925 73.275 -21.595 73.605 ;
        RECT -21.925 71.915 -21.595 72.245 ;
        RECT -21.925 70.555 -21.595 70.885 ;
        RECT -21.925 69.195 -21.595 69.525 ;
        RECT -21.925 67.835 -21.595 68.165 ;
        RECT -21.925 66.475 -21.595 66.805 ;
        RECT -21.925 65.115 -21.595 65.445 ;
        RECT -21.925 63.755 -21.595 64.085 ;
        RECT -21.925 62.395 -21.595 62.725 ;
        RECT -21.925 61.035 -21.595 61.365 ;
        RECT -21.925 59.675 -21.595 60.005 ;
        RECT -21.925 58.315 -21.595 58.645 ;
        RECT -21.925 56.955 -21.595 57.285 ;
        RECT -21.925 55.595 -21.595 55.925 ;
        RECT -21.925 54.235 -21.595 54.565 ;
        RECT -21.925 52.875 -21.595 53.205 ;
        RECT -21.925 51.515 -21.595 51.845 ;
        RECT -21.925 50.155 -21.595 50.485 ;
        RECT -21.925 48.795 -21.595 49.125 ;
        RECT -21.925 47.435 -21.595 47.765 ;
        RECT -21.925 46.075 -21.595 46.405 ;
        RECT -21.925 44.715 -21.595 45.045 ;
        RECT -21.925 43.355 -21.595 43.685 ;
        RECT -21.925 41.995 -21.595 42.325 ;
        RECT -21.925 40.635 -21.595 40.965 ;
        RECT -21.925 39.275 -21.595 39.605 ;
        RECT -21.925 37.915 -21.595 38.245 ;
        RECT -21.925 36.555 -21.595 36.885 ;
        RECT -21.925 35.195 -21.595 35.525 ;
        RECT -21.925 33.835 -21.595 34.165 ;
        RECT -21.925 32.475 -21.595 32.805 ;
        RECT -21.925 31.115 -21.595 31.445 ;
        RECT -21.925 29.755 -21.595 30.085 ;
        RECT -21.925 28.395 -21.595 28.725 ;
        RECT -21.925 27.035 -21.595 27.365 ;
        RECT -21.925 25.675 -21.595 26.005 ;
        RECT -21.925 24.315 -21.595 24.645 ;
        RECT -21.925 22.955 -21.595 23.285 ;
        RECT -21.925 21.595 -21.595 21.925 ;
        RECT -21.925 20.235 -21.595 20.565 ;
        RECT -21.925 18.875 -21.595 19.205 ;
        RECT -21.925 17.515 -21.595 17.845 ;
        RECT -21.925 16.155 -21.595 16.485 ;
        RECT -21.925 14.795 -21.595 15.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 246.76 -29.755 247.89 ;
        RECT -30.085 241.915 -29.755 242.245 ;
        RECT -30.085 240.555 -29.755 240.885 ;
        RECT -30.085 239.195 -29.755 239.525 ;
        RECT -30.085 237.835 -29.755 238.165 ;
        RECT -30.085 236.475 -29.755 236.805 ;
        RECT -30.085 235.115 -29.755 235.445 ;
        RECT -30.085 233.755 -29.755 234.085 ;
        RECT -30.085 232.395 -29.755 232.725 ;
        RECT -30.085 231.035 -29.755 231.365 ;
        RECT -30.085 229.675 -29.755 230.005 ;
        RECT -30.085 228.315 -29.755 228.645 ;
        RECT -30.085 226.955 -29.755 227.285 ;
        RECT -30.085 225.595 -29.755 225.925 ;
        RECT -30.085 224.235 -29.755 224.565 ;
        RECT -30.085 222.875 -29.755 223.205 ;
        RECT -30.085 221.515 -29.755 221.845 ;
        RECT -30.085 220.155 -29.755 220.485 ;
        RECT -30.085 218.795 -29.755 219.125 ;
        RECT -30.085 217.435 -29.755 217.765 ;
        RECT -30.085 216.075 -29.755 216.405 ;
        RECT -30.085 214.715 -29.755 215.045 ;
        RECT -30.085 213.355 -29.755 213.685 ;
        RECT -30.085 211.995 -29.755 212.325 ;
        RECT -30.085 210.635 -29.755 210.965 ;
        RECT -30.085 209.275 -29.755 209.605 ;
        RECT -30.085 207.915 -29.755 208.245 ;
        RECT -30.085 206.555 -29.755 206.885 ;
        RECT -30.085 205.195 -29.755 205.525 ;
        RECT -30.085 203.835 -29.755 204.165 ;
        RECT -30.085 202.475 -29.755 202.805 ;
        RECT -30.085 201.115 -29.755 201.445 ;
        RECT -30.085 199.755 -29.755 200.085 ;
        RECT -30.085 198.395 -29.755 198.725 ;
        RECT -30.085 197.035 -29.755 197.365 ;
        RECT -30.085 195.675 -29.755 196.005 ;
        RECT -30.085 194.315 -29.755 194.645 ;
        RECT -30.085 192.955 -29.755 193.285 ;
        RECT -30.085 191.595 -29.755 191.925 ;
        RECT -30.085 190.235 -29.755 190.565 ;
        RECT -30.085 188.875 -29.755 189.205 ;
        RECT -30.085 187.515 -29.755 187.845 ;
        RECT -30.085 186.155 -29.755 186.485 ;
        RECT -30.085 184.795 -29.755 185.125 ;
        RECT -30.085 183.435 -29.755 183.765 ;
        RECT -30.085 182.075 -29.755 182.405 ;
        RECT -30.085 180.715 -29.755 181.045 ;
        RECT -30.085 179.355 -29.755 179.685 ;
        RECT -30.085 177.995 -29.755 178.325 ;
        RECT -30.085 176.635 -29.755 176.965 ;
        RECT -30.085 175.275 -29.755 175.605 ;
        RECT -30.085 173.915 -29.755 174.245 ;
        RECT -30.085 172.555 -29.755 172.885 ;
        RECT -30.085 171.195 -29.755 171.525 ;
        RECT -30.085 169.835 -29.755 170.165 ;
        RECT -30.085 168.475 -29.755 168.805 ;
        RECT -30.085 167.115 -29.755 167.445 ;
        RECT -30.085 165.755 -29.755 166.085 ;
        RECT -30.085 164.395 -29.755 164.725 ;
        RECT -30.085 163.035 -29.755 163.365 ;
        RECT -30.085 161.675 -29.755 162.005 ;
        RECT -30.085 160.315 -29.755 160.645 ;
        RECT -30.085 158.955 -29.755 159.285 ;
        RECT -30.085 157.595 -29.755 157.925 ;
        RECT -30.085 156.235 -29.755 156.565 ;
        RECT -30.085 154.875 -29.755 155.205 ;
        RECT -30.085 153.515 -29.755 153.845 ;
        RECT -30.085 152.155 -29.755 152.485 ;
        RECT -30.085 150.795 -29.755 151.125 ;
        RECT -30.085 149.435 -29.755 149.765 ;
        RECT -30.085 148.075 -29.755 148.405 ;
        RECT -30.085 146.715 -29.755 147.045 ;
        RECT -30.085 145.355 -29.755 145.685 ;
        RECT -30.085 143.995 -29.755 144.325 ;
        RECT -30.085 142.635 -29.755 142.965 ;
        RECT -30.085 141.275 -29.755 141.605 ;
        RECT -30.085 139.915 -29.755 140.245 ;
        RECT -30.085 138.555 -29.755 138.885 ;
        RECT -30.085 137.195 -29.755 137.525 ;
        RECT -30.085 135.835 -29.755 136.165 ;
        RECT -30.085 134.475 -29.755 134.805 ;
        RECT -30.085 133.115 -29.755 133.445 ;
        RECT -30.085 131.755 -29.755 132.085 ;
        RECT -30.085 130.395 -29.755 130.725 ;
        RECT -30.085 129.035 -29.755 129.365 ;
        RECT -30.085 127.675 -29.755 128.005 ;
        RECT -30.085 126.315 -29.755 126.645 ;
        RECT -30.085 124.955 -29.755 125.285 ;
        RECT -30.085 123.595 -29.755 123.925 ;
        RECT -30.085 122.235 -29.755 122.565 ;
        RECT -30.085 120.875 -29.755 121.205 ;
        RECT -30.085 119.515 -29.755 119.845 ;
        RECT -30.085 118.155 -29.755 118.485 ;
        RECT -30.085 116.795 -29.755 117.125 ;
        RECT -30.085 115.435 -29.755 115.765 ;
        RECT -30.085 114.075 -29.755 114.405 ;
        RECT -30.085 112.715 -29.755 113.045 ;
        RECT -30.085 111.355 -29.755 111.685 ;
        RECT -30.085 109.995 -29.755 110.325 ;
        RECT -30.085 108.635 -29.755 108.965 ;
        RECT -30.085 107.275 -29.755 107.605 ;
        RECT -30.085 105.915 -29.755 106.245 ;
        RECT -30.085 104.555 -29.755 104.885 ;
        RECT -30.085 103.195 -29.755 103.525 ;
        RECT -30.085 101.835 -29.755 102.165 ;
        RECT -30.085 100.475 -29.755 100.805 ;
        RECT -30.085 99.115 -29.755 99.445 ;
        RECT -30.085 97.755 -29.755 98.085 ;
        RECT -30.085 96.395 -29.755 96.725 ;
        RECT -30.085 95.035 -29.755 95.365 ;
        RECT -30.085 93.675 -29.755 94.005 ;
        RECT -30.085 92.315 -29.755 92.645 ;
        RECT -30.085 90.955 -29.755 91.285 ;
        RECT -30.085 89.595 -29.755 89.925 ;
        RECT -30.085 88.235 -29.755 88.565 ;
        RECT -30.085 86.875 -29.755 87.205 ;
        RECT -30.085 85.515 -29.755 85.845 ;
        RECT -30.085 84.155 -29.755 84.485 ;
        RECT -30.085 82.795 -29.755 83.125 ;
        RECT -30.085 81.435 -29.755 81.765 ;
        RECT -30.085 80.075 -29.755 80.405 ;
        RECT -30.085 78.715 -29.755 79.045 ;
        RECT -30.085 77.355 -29.755 77.685 ;
        RECT -30.085 75.995 -29.755 76.325 ;
        RECT -30.085 74.635 -29.755 74.965 ;
        RECT -30.085 73.275 -29.755 73.605 ;
        RECT -30.085 71.915 -29.755 72.245 ;
        RECT -30.085 70.555 -29.755 70.885 ;
        RECT -30.085 69.195 -29.755 69.525 ;
        RECT -30.085 67.835 -29.755 68.165 ;
        RECT -30.085 66.475 -29.755 66.805 ;
        RECT -30.085 65.115 -29.755 65.445 ;
        RECT -30.085 63.755 -29.755 64.085 ;
        RECT -30.085 62.395 -29.755 62.725 ;
        RECT -30.085 61.035 -29.755 61.365 ;
        RECT -30.085 59.675 -29.755 60.005 ;
        RECT -30.085 58.315 -29.755 58.645 ;
        RECT -30.085 56.955 -29.755 57.285 ;
        RECT -30.085 55.595 -29.755 55.925 ;
        RECT -30.085 54.235 -29.755 54.565 ;
        RECT -30.085 52.875 -29.755 53.205 ;
        RECT -30.085 51.515 -29.755 51.845 ;
        RECT -30.085 50.155 -29.755 50.485 ;
        RECT -30.085 48.795 -29.755 49.125 ;
        RECT -30.085 47.435 -29.755 47.765 ;
        RECT -30.085 46.075 -29.755 46.405 ;
        RECT -30.085 44.715 -29.755 45.045 ;
        RECT -30.085 43.355 -29.755 43.685 ;
        RECT -30.085 41.995 -29.755 42.325 ;
        RECT -30.085 40.635 -29.755 40.965 ;
        RECT -30.085 39.275 -29.755 39.605 ;
        RECT -30.085 37.915 -29.755 38.245 ;
        RECT -30.085 36.555 -29.755 36.885 ;
        RECT -30.085 35.195 -29.755 35.525 ;
        RECT -30.085 33.835 -29.755 34.165 ;
        RECT -30.085 32.475 -29.755 32.805 ;
        RECT -30.085 31.115 -29.755 31.445 ;
        RECT -30.085 29.755 -29.755 30.085 ;
        RECT -30.085 28.395 -29.755 28.725 ;
        RECT -30.085 27.035 -29.755 27.365 ;
        RECT -30.085 25.675 -29.755 26.005 ;
        RECT -30.085 24.315 -29.755 24.645 ;
        RECT -30.085 22.955 -29.755 23.285 ;
        RECT -30.085 21.595 -29.755 21.925 ;
        RECT -30.085 20.235 -29.755 20.565 ;
        RECT -30.085 18.875 -29.755 19.205 ;
        RECT -30.085 17.515 -29.755 17.845 ;
        RECT -30.085 16.155 -29.755 16.485 ;
        RECT -30.085 14.795 -29.755 15.125 ;
        RECT -30.085 13.435 -29.755 13.765 ;
        RECT -30.085 12.075 -29.755 12.405 ;
        RECT -30.085 10.715 -29.755 11.045 ;
        RECT -30.085 9.355 -29.755 9.685 ;
        RECT -30.085 7.995 -29.755 8.325 ;
        RECT -30.085 6.635 -29.755 6.965 ;
        RECT -30.085 5.275 -29.755 5.605 ;
        RECT -30.085 3.915 -29.755 4.245 ;
        RECT -30.085 2.555 -29.755 2.885 ;
        RECT -30.085 1.195 -29.755 1.525 ;
        RECT -30.085 -0.165 -29.755 0.165 ;
        RECT -30.085 -2.885 -29.755 -2.555 ;
        RECT -30.085 -6.965 -29.755 -6.635 ;
        RECT -30.085 -8.325 -29.755 -7.995 ;
        RECT -30.085 -9.48 -29.755 -9.15 ;
        RECT -30.085 -12.405 -29.755 -12.075 ;
        RECT -30.085 -15.125 -29.755 -14.795 ;
        RECT -30.085 -16.67 -29.755 -16.34 ;
        RECT -30.085 -17.845 -29.755 -17.515 ;
        RECT -30.085 -30.66 -29.755 -30.33 ;
        RECT -30.085 -31.445 -29.755 -31.115 ;
        RECT -30.085 -32.805 -29.755 -32.475 ;
        RECT -30.085 -34.165 -29.755 -33.835 ;
        RECT -30.085 -36.885 -29.755 -36.555 ;
        RECT -30.085 -37.85 -29.755 -37.52 ;
        RECT -30.085 -40.965 -29.755 -40.635 ;
        RECT -30.085 -46.405 -29.755 -46.075 ;
        RECT -30.085 -49.125 -29.755 -48.795 ;
        RECT -30.085 -50.485 -29.755 -50.155 ;
        RECT -30.085 -53.205 -29.755 -52.875 ;
        RECT -30.085 -55.925 -29.755 -55.595 ;
        RECT -30.08 -58.64 -29.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 -129.365 -29.755 -129.035 ;
        RECT -30.085 -130.725 -29.755 -130.395 ;
        RECT -30.085 -132.085 -29.755 -131.755 ;
        RECT -30.085 -133.51 -29.755 -133.18 ;
        RECT -30.085 -134.805 -29.755 -134.475 ;
        RECT -30.085 -136.165 -29.755 -135.835 ;
        RECT -30.085 -137.525 -29.755 -137.195 ;
        RECT -30.085 -138.885 -29.755 -138.555 ;
        RECT -30.085 -140.245 -29.755 -139.915 ;
        RECT -30.085 -141.605 -29.755 -141.275 ;
        RECT -30.085 -144.325 -29.755 -143.995 ;
        RECT -30.085 -145.685 -29.755 -145.355 ;
        RECT -30.085 -147.045 -29.755 -146.715 ;
        RECT -30.085 -152.485 -29.755 -152.155 ;
        RECT -30.085 -153.845 -29.755 -153.515 ;
        RECT -30.085 -155.205 -29.755 -154.875 ;
        RECT -30.085 -156.565 -29.755 -156.235 ;
        RECT -30.085 -157.925 -29.755 -157.595 ;
        RECT -30.085 -159.285 -29.755 -158.955 ;
        RECT -30.085 -162.005 -29.755 -161.675 ;
        RECT -30.085 -163.365 -29.755 -163.035 ;
        RECT -30.085 -164.725 -29.755 -164.395 ;
        RECT -30.085 -166.085 -29.755 -165.755 ;
        RECT -30.085 -167.445 -29.755 -167.115 ;
        RECT -30.085 -168.805 -29.755 -168.475 ;
        RECT -30.085 -170.165 -29.755 -169.835 ;
        RECT -30.085 -171.525 -29.755 -171.195 ;
        RECT -30.085 -172.885 -29.755 -172.555 ;
        RECT -30.085 -174.245 -29.755 -173.915 ;
        RECT -30.085 -175.605 -29.755 -175.275 ;
        RECT -30.085 -176.965 -29.755 -176.635 ;
        RECT -30.085 -178.325 -29.755 -177.995 ;
        RECT -30.085 -179.685 -29.755 -179.355 ;
        RECT -30.085 -181.045 -29.755 -180.715 ;
        RECT -30.085 -182.405 -29.755 -182.075 ;
        RECT -30.085 -183.765 -29.755 -183.435 ;
        RECT -30.085 -185.125 -29.755 -184.795 ;
        RECT -30.085 -186.485 -29.755 -186.155 ;
        RECT -30.085 -190.565 -29.755 -190.235 ;
        RECT -30.085 -191.925 -29.755 -191.595 ;
        RECT -30.085 -193.285 -29.755 -192.955 ;
        RECT -30.085 -194.645 -29.755 -194.315 ;
        RECT -30.085 -196.005 -29.755 -195.675 ;
        RECT -30.085 -197.365 -29.755 -197.035 ;
        RECT -30.085 -198.725 -29.755 -198.395 ;
        RECT -30.085 -200.085 -29.755 -199.755 ;
        RECT -30.085 -201.445 -29.755 -201.115 ;
        RECT -30.085 -202.805 -29.755 -202.475 ;
        RECT -30.085 -204.165 -29.755 -203.835 ;
        RECT -30.085 -205.525 -29.755 -205.195 ;
        RECT -30.085 -208.245 -29.755 -207.915 ;
        RECT -30.085 -209.605 -29.755 -209.275 ;
        RECT -30.085 -213.685 -29.755 -213.355 ;
        RECT -30.085 -215.045 -29.755 -214.715 ;
        RECT -30.085 -216.405 -29.755 -216.075 ;
        RECT -30.085 -217.765 -29.755 -217.435 ;
        RECT -30.085 -219.125 -29.755 -218.795 ;
        RECT -30.085 -220.485 -29.755 -220.155 ;
        RECT -30.085 -221.845 -29.755 -221.515 ;
        RECT -30.085 -223.205 -29.755 -222.875 ;
        RECT -30.085 -224.565 -29.755 -224.235 ;
        RECT -30.085 -226.155 -29.755 -225.825 ;
        RECT -30.085 -227.285 -29.755 -226.955 ;
        RECT -30.08 -227.285 -29.76 -121.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 -234.085 -29.755 -233.755 ;
        RECT -30.085 -235.445 -29.755 -235.115 ;
        RECT -30.085 -236.805 -29.755 -236.475 ;
        RECT -30.085 -238.165 -29.755 -237.835 ;
        RECT -30.085 -243.81 -29.755 -242.68 ;
        RECT -30.08 -243.925 -29.76 -231.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 246.76 -28.395 247.89 ;
        RECT -28.725 241.915 -28.395 242.245 ;
        RECT -28.725 240.555 -28.395 240.885 ;
        RECT -28.725 239.195 -28.395 239.525 ;
        RECT -28.725 237.835 -28.395 238.165 ;
        RECT -28.725 236.475 -28.395 236.805 ;
        RECT -28.725 235.115 -28.395 235.445 ;
        RECT -28.725 233.755 -28.395 234.085 ;
        RECT -28.725 232.395 -28.395 232.725 ;
        RECT -28.725 231.035 -28.395 231.365 ;
        RECT -28.725 229.675 -28.395 230.005 ;
        RECT -28.725 228.315 -28.395 228.645 ;
        RECT -28.725 226.955 -28.395 227.285 ;
        RECT -28.725 225.595 -28.395 225.925 ;
        RECT -28.725 224.235 -28.395 224.565 ;
        RECT -28.725 222.875 -28.395 223.205 ;
        RECT -28.725 221.515 -28.395 221.845 ;
        RECT -28.725 220.155 -28.395 220.485 ;
        RECT -28.725 218.795 -28.395 219.125 ;
        RECT -28.725 217.435 -28.395 217.765 ;
        RECT -28.725 216.075 -28.395 216.405 ;
        RECT -28.725 214.715 -28.395 215.045 ;
        RECT -28.725 213.355 -28.395 213.685 ;
        RECT -28.725 211.995 -28.395 212.325 ;
        RECT -28.725 210.635 -28.395 210.965 ;
        RECT -28.725 209.275 -28.395 209.605 ;
        RECT -28.725 207.915 -28.395 208.245 ;
        RECT -28.725 206.555 -28.395 206.885 ;
        RECT -28.725 205.195 -28.395 205.525 ;
        RECT -28.725 203.835 -28.395 204.165 ;
        RECT -28.725 202.475 -28.395 202.805 ;
        RECT -28.725 201.115 -28.395 201.445 ;
        RECT -28.725 199.755 -28.395 200.085 ;
        RECT -28.725 198.395 -28.395 198.725 ;
        RECT -28.725 197.035 -28.395 197.365 ;
        RECT -28.725 195.675 -28.395 196.005 ;
        RECT -28.725 194.315 -28.395 194.645 ;
        RECT -28.725 192.955 -28.395 193.285 ;
        RECT -28.725 191.595 -28.395 191.925 ;
        RECT -28.725 190.235 -28.395 190.565 ;
        RECT -28.725 188.875 -28.395 189.205 ;
        RECT -28.725 187.515 -28.395 187.845 ;
        RECT -28.725 186.155 -28.395 186.485 ;
        RECT -28.725 184.795 -28.395 185.125 ;
        RECT -28.725 183.435 -28.395 183.765 ;
        RECT -28.725 182.075 -28.395 182.405 ;
        RECT -28.725 180.715 -28.395 181.045 ;
        RECT -28.725 179.355 -28.395 179.685 ;
        RECT -28.725 177.995 -28.395 178.325 ;
        RECT -28.725 176.635 -28.395 176.965 ;
        RECT -28.725 175.275 -28.395 175.605 ;
        RECT -28.725 173.915 -28.395 174.245 ;
        RECT -28.725 172.555 -28.395 172.885 ;
        RECT -28.725 171.195 -28.395 171.525 ;
        RECT -28.725 169.835 -28.395 170.165 ;
        RECT -28.725 168.475 -28.395 168.805 ;
        RECT -28.725 167.115 -28.395 167.445 ;
        RECT -28.725 165.755 -28.395 166.085 ;
        RECT -28.725 164.395 -28.395 164.725 ;
        RECT -28.725 163.035 -28.395 163.365 ;
        RECT -28.725 161.675 -28.395 162.005 ;
        RECT -28.725 160.315 -28.395 160.645 ;
        RECT -28.725 158.955 -28.395 159.285 ;
        RECT -28.725 157.595 -28.395 157.925 ;
        RECT -28.725 156.235 -28.395 156.565 ;
        RECT -28.725 154.875 -28.395 155.205 ;
        RECT -28.725 153.515 -28.395 153.845 ;
        RECT -28.725 152.155 -28.395 152.485 ;
        RECT -28.725 150.795 -28.395 151.125 ;
        RECT -28.725 149.435 -28.395 149.765 ;
        RECT -28.725 148.075 -28.395 148.405 ;
        RECT -28.725 146.715 -28.395 147.045 ;
        RECT -28.725 145.355 -28.395 145.685 ;
        RECT -28.725 143.995 -28.395 144.325 ;
        RECT -28.725 142.635 -28.395 142.965 ;
        RECT -28.725 141.275 -28.395 141.605 ;
        RECT -28.725 139.915 -28.395 140.245 ;
        RECT -28.725 138.555 -28.395 138.885 ;
        RECT -28.725 137.195 -28.395 137.525 ;
        RECT -28.725 135.835 -28.395 136.165 ;
        RECT -28.725 134.475 -28.395 134.805 ;
        RECT -28.725 133.115 -28.395 133.445 ;
        RECT -28.725 131.755 -28.395 132.085 ;
        RECT -28.725 130.395 -28.395 130.725 ;
        RECT -28.725 129.035 -28.395 129.365 ;
        RECT -28.725 127.675 -28.395 128.005 ;
        RECT -28.725 126.315 -28.395 126.645 ;
        RECT -28.725 124.955 -28.395 125.285 ;
        RECT -28.725 123.595 -28.395 123.925 ;
        RECT -28.725 122.235 -28.395 122.565 ;
        RECT -28.725 120.875 -28.395 121.205 ;
        RECT -28.725 119.515 -28.395 119.845 ;
        RECT -28.725 118.155 -28.395 118.485 ;
        RECT -28.725 116.795 -28.395 117.125 ;
        RECT -28.725 115.435 -28.395 115.765 ;
        RECT -28.725 114.075 -28.395 114.405 ;
        RECT -28.725 112.715 -28.395 113.045 ;
        RECT -28.725 111.355 -28.395 111.685 ;
        RECT -28.725 109.995 -28.395 110.325 ;
        RECT -28.725 108.635 -28.395 108.965 ;
        RECT -28.725 107.275 -28.395 107.605 ;
        RECT -28.725 105.915 -28.395 106.245 ;
        RECT -28.725 104.555 -28.395 104.885 ;
        RECT -28.725 103.195 -28.395 103.525 ;
        RECT -28.725 101.835 -28.395 102.165 ;
        RECT -28.725 100.475 -28.395 100.805 ;
        RECT -28.725 99.115 -28.395 99.445 ;
        RECT -28.725 97.755 -28.395 98.085 ;
        RECT -28.725 96.395 -28.395 96.725 ;
        RECT -28.725 95.035 -28.395 95.365 ;
        RECT -28.725 93.675 -28.395 94.005 ;
        RECT -28.725 92.315 -28.395 92.645 ;
        RECT -28.725 90.955 -28.395 91.285 ;
        RECT -28.725 89.595 -28.395 89.925 ;
        RECT -28.725 88.235 -28.395 88.565 ;
        RECT -28.725 86.875 -28.395 87.205 ;
        RECT -28.725 85.515 -28.395 85.845 ;
        RECT -28.725 84.155 -28.395 84.485 ;
        RECT -28.725 82.795 -28.395 83.125 ;
        RECT -28.725 81.435 -28.395 81.765 ;
        RECT -28.725 80.075 -28.395 80.405 ;
        RECT -28.725 78.715 -28.395 79.045 ;
        RECT -28.725 77.355 -28.395 77.685 ;
        RECT -28.725 75.995 -28.395 76.325 ;
        RECT -28.725 74.635 -28.395 74.965 ;
        RECT -28.725 73.275 -28.395 73.605 ;
        RECT -28.725 71.915 -28.395 72.245 ;
        RECT -28.725 70.555 -28.395 70.885 ;
        RECT -28.725 69.195 -28.395 69.525 ;
        RECT -28.725 67.835 -28.395 68.165 ;
        RECT -28.725 66.475 -28.395 66.805 ;
        RECT -28.725 65.115 -28.395 65.445 ;
        RECT -28.725 63.755 -28.395 64.085 ;
        RECT -28.725 62.395 -28.395 62.725 ;
        RECT -28.725 61.035 -28.395 61.365 ;
        RECT -28.725 59.675 -28.395 60.005 ;
        RECT -28.725 58.315 -28.395 58.645 ;
        RECT -28.725 56.955 -28.395 57.285 ;
        RECT -28.725 55.595 -28.395 55.925 ;
        RECT -28.725 54.235 -28.395 54.565 ;
        RECT -28.725 52.875 -28.395 53.205 ;
        RECT -28.725 51.515 -28.395 51.845 ;
        RECT -28.725 50.155 -28.395 50.485 ;
        RECT -28.725 48.795 -28.395 49.125 ;
        RECT -28.725 47.435 -28.395 47.765 ;
        RECT -28.725 46.075 -28.395 46.405 ;
        RECT -28.725 44.715 -28.395 45.045 ;
        RECT -28.725 43.355 -28.395 43.685 ;
        RECT -28.725 41.995 -28.395 42.325 ;
        RECT -28.725 40.635 -28.395 40.965 ;
        RECT -28.725 39.275 -28.395 39.605 ;
        RECT -28.725 37.915 -28.395 38.245 ;
        RECT -28.725 36.555 -28.395 36.885 ;
        RECT -28.725 35.195 -28.395 35.525 ;
        RECT -28.725 33.835 -28.395 34.165 ;
        RECT -28.725 32.475 -28.395 32.805 ;
        RECT -28.725 31.115 -28.395 31.445 ;
        RECT -28.725 29.755 -28.395 30.085 ;
        RECT -28.725 28.395 -28.395 28.725 ;
        RECT -28.725 27.035 -28.395 27.365 ;
        RECT -28.725 25.675 -28.395 26.005 ;
        RECT -28.725 24.315 -28.395 24.645 ;
        RECT -28.725 22.955 -28.395 23.285 ;
        RECT -28.725 21.595 -28.395 21.925 ;
        RECT -28.725 20.235 -28.395 20.565 ;
        RECT -28.725 18.875 -28.395 19.205 ;
        RECT -28.725 17.515 -28.395 17.845 ;
        RECT -28.725 16.155 -28.395 16.485 ;
        RECT -28.725 14.795 -28.395 15.125 ;
        RECT -28.725 13.435 -28.395 13.765 ;
        RECT -28.725 12.075 -28.395 12.405 ;
        RECT -28.725 10.715 -28.395 11.045 ;
        RECT -28.725 9.355 -28.395 9.685 ;
        RECT -28.725 7.995 -28.395 8.325 ;
        RECT -28.725 6.635 -28.395 6.965 ;
        RECT -28.725 5.275 -28.395 5.605 ;
        RECT -28.725 3.915 -28.395 4.245 ;
        RECT -28.725 2.555 -28.395 2.885 ;
        RECT -28.725 1.195 -28.395 1.525 ;
        RECT -28.725 -0.165 -28.395 0.165 ;
        RECT -28.725 -2.885 -28.395 -2.555 ;
        RECT -28.725 -6.965 -28.395 -6.635 ;
        RECT -28.725 -8.325 -28.395 -7.995 ;
        RECT -28.725 -9.48 -28.395 -9.15 ;
        RECT -28.725 -12.405 -28.395 -12.075 ;
        RECT -28.725 -15.125 -28.395 -14.795 ;
        RECT -28.725 -16.67 -28.395 -16.34 ;
        RECT -28.725 -17.845 -28.395 -17.515 ;
        RECT -28.725 -30.66 -28.395 -30.33 ;
        RECT -28.725 -31.445 -28.395 -31.115 ;
        RECT -28.725 -32.805 -28.395 -32.475 ;
        RECT -28.725 -34.165 -28.395 -33.835 ;
        RECT -28.725 -36.885 -28.395 -36.555 ;
        RECT -28.725 -37.85 -28.395 -37.52 ;
        RECT -28.725 -40.965 -28.395 -40.635 ;
        RECT -28.725 -46.405 -28.395 -46.075 ;
        RECT -28.725 -49.125 -28.395 -48.795 ;
        RECT -28.725 -50.485 -28.395 -50.155 ;
        RECT -28.725 -53.205 -28.395 -52.875 ;
        RECT -28.725 -55.925 -28.395 -55.595 ;
        RECT -28.72 -57.96 -28.4 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 -122.565 -28.395 -122.235 ;
        RECT -28.725 -129.365 -28.395 -129.035 ;
        RECT -28.725 -130.725 -28.395 -130.395 ;
        RECT -28.725 -132.085 -28.395 -131.755 ;
        RECT -28.725 -133.51 -28.395 -133.18 ;
        RECT -28.725 -134.805 -28.395 -134.475 ;
        RECT -28.725 -136.165 -28.395 -135.835 ;
        RECT -28.725 -137.525 -28.395 -137.195 ;
        RECT -28.725 -138.885 -28.395 -138.555 ;
        RECT -28.725 -140.245 -28.395 -139.915 ;
        RECT -28.725 -141.605 -28.395 -141.275 ;
        RECT -28.725 -144.325 -28.395 -143.995 ;
        RECT -28.725 -145.685 -28.395 -145.355 ;
        RECT -28.725 -147.045 -28.395 -146.715 ;
        RECT -28.725 -152.485 -28.395 -152.155 ;
        RECT -28.725 -153.845 -28.395 -153.515 ;
        RECT -28.725 -155.205 -28.395 -154.875 ;
        RECT -28.725 -156.565 -28.395 -156.235 ;
        RECT -28.725 -157.925 -28.395 -157.595 ;
        RECT -28.725 -159.285 -28.395 -158.955 ;
        RECT -28.725 -162.005 -28.395 -161.675 ;
        RECT -28.725 -163.365 -28.395 -163.035 ;
        RECT -28.725 -164.725 -28.395 -164.395 ;
        RECT -28.725 -166.085 -28.395 -165.755 ;
        RECT -28.725 -167.445 -28.395 -167.115 ;
        RECT -28.725 -168.805 -28.395 -168.475 ;
        RECT -28.725 -170.165 -28.395 -169.835 ;
        RECT -28.725 -171.525 -28.395 -171.195 ;
        RECT -28.725 -172.885 -28.395 -172.555 ;
        RECT -28.725 -174.245 -28.395 -173.915 ;
        RECT -28.725 -175.605 -28.395 -175.275 ;
        RECT -28.725 -176.965 -28.395 -176.635 ;
        RECT -28.725 -178.325 -28.395 -177.995 ;
        RECT -28.725 -179.685 -28.395 -179.355 ;
        RECT -28.725 -181.045 -28.395 -180.715 ;
        RECT -28.725 -182.405 -28.395 -182.075 ;
        RECT -28.725 -183.765 -28.395 -183.435 ;
        RECT -28.725 -185.125 -28.395 -184.795 ;
        RECT -28.725 -186.485 -28.395 -186.155 ;
        RECT -28.725 -190.565 -28.395 -190.235 ;
        RECT -28.725 -191.925 -28.395 -191.595 ;
        RECT -28.725 -193.285 -28.395 -192.955 ;
        RECT -28.725 -194.645 -28.395 -194.315 ;
        RECT -28.725 -196.005 -28.395 -195.675 ;
        RECT -28.725 -198.725 -28.395 -198.395 ;
        RECT -28.725 -200.085 -28.395 -199.755 ;
        RECT -28.725 -201.445 -28.395 -201.115 ;
        RECT -28.725 -202.805 -28.395 -202.475 ;
        RECT -28.725 -204.165 -28.395 -203.835 ;
        RECT -28.725 -205.525 -28.395 -205.195 ;
        RECT -28.725 -208.245 -28.395 -207.915 ;
        RECT -28.725 -209.605 -28.395 -209.275 ;
        RECT -28.725 -215.045 -28.395 -214.715 ;
        RECT -28.725 -216.405 -28.395 -216.075 ;
        RECT -28.725 -217.765 -28.395 -217.435 ;
        RECT -28.725 -219.125 -28.395 -218.795 ;
        RECT -28.725 -220.485 -28.395 -220.155 ;
        RECT -28.725 -221.845 -28.395 -221.515 ;
        RECT -28.725 -223.205 -28.395 -222.875 ;
        RECT -28.725 -224.565 -28.395 -224.235 ;
        RECT -28.725 -227.285 -28.395 -226.955 ;
        RECT -28.725 -231.365 -28.395 -231.035 ;
        RECT -28.725 -234.085 -28.395 -233.755 ;
        RECT -28.725 -235.445 -28.395 -235.115 ;
        RECT -28.725 -236.805 -28.395 -236.475 ;
        RECT -28.725 -238.165 -28.395 -237.835 ;
        RECT -28.725 -243.81 -28.395 -242.68 ;
        RECT -28.72 -243.925 -28.4 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.365 171.195 -27.035 171.525 ;
        RECT -27.365 169.835 -27.035 170.165 ;
        RECT -27.365 168.475 -27.035 168.805 ;
        RECT -27.365 167.115 -27.035 167.445 ;
        RECT -27.365 165.755 -27.035 166.085 ;
        RECT -27.365 164.395 -27.035 164.725 ;
        RECT -27.365 163.035 -27.035 163.365 ;
        RECT -27.365 161.675 -27.035 162.005 ;
        RECT -27.365 160.315 -27.035 160.645 ;
        RECT -27.365 158.955 -27.035 159.285 ;
        RECT -27.365 157.595 -27.035 157.925 ;
        RECT -27.365 156.235 -27.035 156.565 ;
        RECT -27.365 154.875 -27.035 155.205 ;
        RECT -27.365 153.515 -27.035 153.845 ;
        RECT -27.365 152.155 -27.035 152.485 ;
        RECT -27.365 150.795 -27.035 151.125 ;
        RECT -27.365 149.435 -27.035 149.765 ;
        RECT -27.365 148.075 -27.035 148.405 ;
        RECT -27.365 146.715 -27.035 147.045 ;
        RECT -27.365 145.355 -27.035 145.685 ;
        RECT -27.365 143.995 -27.035 144.325 ;
        RECT -27.365 142.635 -27.035 142.965 ;
        RECT -27.365 141.275 -27.035 141.605 ;
        RECT -27.365 139.915 -27.035 140.245 ;
        RECT -27.365 138.555 -27.035 138.885 ;
        RECT -27.365 137.195 -27.035 137.525 ;
        RECT -27.365 135.835 -27.035 136.165 ;
        RECT -27.365 134.475 -27.035 134.805 ;
        RECT -27.365 133.115 -27.035 133.445 ;
        RECT -27.365 131.755 -27.035 132.085 ;
        RECT -27.365 130.395 -27.035 130.725 ;
        RECT -27.365 129.035 -27.035 129.365 ;
        RECT -27.365 127.675 -27.035 128.005 ;
        RECT -27.365 126.315 -27.035 126.645 ;
        RECT -27.365 124.955 -27.035 125.285 ;
        RECT -27.365 123.595 -27.035 123.925 ;
        RECT -27.365 122.235 -27.035 122.565 ;
        RECT -27.365 120.875 -27.035 121.205 ;
        RECT -27.365 119.515 -27.035 119.845 ;
        RECT -27.365 118.155 -27.035 118.485 ;
        RECT -27.365 116.795 -27.035 117.125 ;
        RECT -27.365 115.435 -27.035 115.765 ;
        RECT -27.365 114.075 -27.035 114.405 ;
        RECT -27.365 112.715 -27.035 113.045 ;
        RECT -27.365 111.355 -27.035 111.685 ;
        RECT -27.365 109.995 -27.035 110.325 ;
        RECT -27.365 108.635 -27.035 108.965 ;
        RECT -27.365 107.275 -27.035 107.605 ;
        RECT -27.365 105.915 -27.035 106.245 ;
        RECT -27.365 104.555 -27.035 104.885 ;
        RECT -27.365 103.195 -27.035 103.525 ;
        RECT -27.365 101.835 -27.035 102.165 ;
        RECT -27.365 100.475 -27.035 100.805 ;
        RECT -27.365 99.115 -27.035 99.445 ;
        RECT -27.365 97.755 -27.035 98.085 ;
        RECT -27.365 96.395 -27.035 96.725 ;
        RECT -27.365 95.035 -27.035 95.365 ;
        RECT -27.365 93.675 -27.035 94.005 ;
        RECT -27.365 92.315 -27.035 92.645 ;
        RECT -27.365 90.955 -27.035 91.285 ;
        RECT -27.365 89.595 -27.035 89.925 ;
        RECT -27.365 88.235 -27.035 88.565 ;
        RECT -27.365 86.875 -27.035 87.205 ;
        RECT -27.365 85.515 -27.035 85.845 ;
        RECT -27.365 84.155 -27.035 84.485 ;
        RECT -27.365 82.795 -27.035 83.125 ;
        RECT -27.365 81.435 -27.035 81.765 ;
        RECT -27.365 80.075 -27.035 80.405 ;
        RECT -27.365 78.715 -27.035 79.045 ;
        RECT -27.365 77.355 -27.035 77.685 ;
        RECT -27.365 75.995 -27.035 76.325 ;
        RECT -27.365 74.635 -27.035 74.965 ;
        RECT -27.365 73.275 -27.035 73.605 ;
        RECT -27.365 71.915 -27.035 72.245 ;
        RECT -27.365 70.555 -27.035 70.885 ;
        RECT -27.365 69.195 -27.035 69.525 ;
        RECT -27.365 67.835 -27.035 68.165 ;
        RECT -27.365 66.475 -27.035 66.805 ;
        RECT -27.365 65.115 -27.035 65.445 ;
        RECT -27.365 63.755 -27.035 64.085 ;
        RECT -27.365 62.395 -27.035 62.725 ;
        RECT -27.365 61.035 -27.035 61.365 ;
        RECT -27.365 59.675 -27.035 60.005 ;
        RECT -27.365 58.315 -27.035 58.645 ;
        RECT -27.365 56.955 -27.035 57.285 ;
        RECT -27.365 55.595 -27.035 55.925 ;
        RECT -27.365 54.235 -27.035 54.565 ;
        RECT -27.365 52.875 -27.035 53.205 ;
        RECT -27.365 51.515 -27.035 51.845 ;
        RECT -27.365 50.155 -27.035 50.485 ;
        RECT -27.365 48.795 -27.035 49.125 ;
        RECT -27.365 47.435 -27.035 47.765 ;
        RECT -27.365 46.075 -27.035 46.405 ;
        RECT -27.365 44.715 -27.035 45.045 ;
        RECT -27.365 43.355 -27.035 43.685 ;
        RECT -27.365 41.995 -27.035 42.325 ;
        RECT -27.365 40.635 -27.035 40.965 ;
        RECT -27.365 39.275 -27.035 39.605 ;
        RECT -27.365 37.915 -27.035 38.245 ;
        RECT -27.365 36.555 -27.035 36.885 ;
        RECT -27.365 35.195 -27.035 35.525 ;
        RECT -27.365 33.835 -27.035 34.165 ;
        RECT -27.365 32.475 -27.035 32.805 ;
        RECT -27.365 31.115 -27.035 31.445 ;
        RECT -27.365 29.755 -27.035 30.085 ;
        RECT -27.365 28.395 -27.035 28.725 ;
        RECT -27.365 27.035 -27.035 27.365 ;
        RECT -27.365 25.675 -27.035 26.005 ;
        RECT -27.365 24.315 -27.035 24.645 ;
        RECT -27.365 22.955 -27.035 23.285 ;
        RECT -27.365 21.595 -27.035 21.925 ;
        RECT -27.365 20.235 -27.035 20.565 ;
        RECT -27.365 18.875 -27.035 19.205 ;
        RECT -27.365 17.515 -27.035 17.845 ;
        RECT -27.365 16.155 -27.035 16.485 ;
        RECT -27.365 14.795 -27.035 15.125 ;
        RECT -27.365 13.435 -27.035 13.765 ;
        RECT -27.365 12.075 -27.035 12.405 ;
        RECT -27.365 10.715 -27.035 11.045 ;
        RECT -27.365 9.355 -27.035 9.685 ;
        RECT -27.365 7.995 -27.035 8.325 ;
        RECT -27.365 6.635 -27.035 6.965 ;
        RECT -27.365 5.275 -27.035 5.605 ;
        RECT -27.365 3.915 -27.035 4.245 ;
        RECT -27.365 2.555 -27.035 2.885 ;
        RECT -27.365 1.195 -27.035 1.525 ;
        RECT -27.365 -0.165 -27.035 0.165 ;
        RECT -27.365 -2.885 -27.035 -2.555 ;
        RECT -27.365 -6.965 -27.035 -6.635 ;
        RECT -27.365 -8.325 -27.035 -7.995 ;
        RECT -27.365 -9.48 -27.035 -9.15 ;
        RECT -27.365 -12.405 -27.035 -12.075 ;
        RECT -27.365 -15.125 -27.035 -14.795 ;
        RECT -27.365 -16.67 -27.035 -16.34 ;
        RECT -27.365 -17.845 -27.035 -17.515 ;
        RECT -27.365 -30.66 -27.035 -30.33 ;
        RECT -27.365 -31.445 -27.035 -31.115 ;
        RECT -27.365 -32.805 -27.035 -32.475 ;
        RECT -27.365 -34.165 -27.035 -33.835 ;
        RECT -27.365 -36.885 -27.035 -36.555 ;
        RECT -27.365 -37.85 -27.035 -37.52 ;
        RECT -27.365 -40.965 -27.035 -40.635 ;
        RECT -27.365 -46.405 -27.035 -46.075 ;
        RECT -27.365 -49.125 -27.035 -48.795 ;
        RECT -27.365 -50.485 -27.035 -50.155 ;
        RECT -27.365 -53.205 -27.035 -52.875 ;
        RECT -27.365 -55.925 -27.035 -55.595 ;
        RECT -27.365 -61.365 -27.035 -61.035 ;
        RECT -27.365 -62.725 -27.035 -62.395 ;
        RECT -27.365 -64.085 -27.035 -63.755 ;
        RECT -27.365 -65.445 -27.035 -65.115 ;
        RECT -27.365 -68.165 -27.035 -67.835 ;
        RECT -27.365 -69.525 -27.035 -69.195 ;
        RECT -27.365 -70.79 -27.035 -70.46 ;
        RECT -27.365 -72.245 -27.035 -71.915 ;
        RECT -27.365 -73.605 -27.035 -73.275 ;
        RECT -27.365 -74.965 -27.035 -74.635 ;
        RECT -27.365 -76.325 -27.035 -75.995 ;
        RECT -27.365 -77.685 -27.035 -77.355 ;
        RECT -27.365 -79.045 -27.035 -78.715 ;
        RECT -27.365 -81.765 -27.035 -81.435 ;
        RECT -27.365 -83.125 -27.035 -82.795 ;
        RECT -27.365 -84.485 -27.035 -84.155 ;
        RECT -27.365 -85.845 -27.035 -85.515 ;
        RECT -27.365 -87.205 -27.035 -86.875 ;
        RECT -27.365 -88.565 -27.035 -88.235 ;
        RECT -27.365 -89.33 -27.035 -89 ;
        RECT -27.365 -91.285 -27.035 -90.955 ;
        RECT -27.365 -92.645 -27.035 -92.315 ;
        RECT -27.365 -94.005 -27.035 -93.675 ;
        RECT -27.365 -95.365 -27.035 -95.035 ;
        RECT -27.365 -96.725 -27.035 -96.395 ;
        RECT -27.365 -98.085 -27.035 -97.755 ;
        RECT -27.365 -100.805 -27.035 -100.475 ;
        RECT -27.365 -102.165 -27.035 -101.835 ;
        RECT -27.365 -103.525 -27.035 -103.195 ;
        RECT -27.365 -106.245 -27.035 -105.915 ;
        RECT -27.365 -107.605 -27.035 -107.275 ;
        RECT -27.365 -108.965 -27.035 -108.635 ;
        RECT -27.365 -110.325 -27.035 -109.995 ;
        RECT -27.365 -111.685 -27.035 -111.355 ;
        RECT -27.365 -113.045 -27.035 -112.715 ;
        RECT -27.365 -114.97 -27.035 -114.64 ;
        RECT -27.365 -115.765 -27.035 -115.435 ;
        RECT -27.365 -117.125 -27.035 -116.795 ;
        RECT -27.365 -118.485 -27.035 -118.155 ;
        RECT -27.365 -119.845 -27.035 -119.515 ;
        RECT -27.365 -121.205 -27.035 -120.875 ;
        RECT -27.365 -122.565 -27.035 -122.235 ;
        RECT -27.365 -129.365 -27.035 -129.035 ;
        RECT -27.365 -130.725 -27.035 -130.395 ;
        RECT -27.365 -132.085 -27.035 -131.755 ;
        RECT -27.365 -133.51 -27.035 -133.18 ;
        RECT -27.365 -136.165 -27.035 -135.835 ;
        RECT -27.365 -137.525 -27.035 -137.195 ;
        RECT -27.365 -138.885 -27.035 -138.555 ;
        RECT -27.365 -140.245 -27.035 -139.915 ;
        RECT -27.365 -141.605 -27.035 -141.275 ;
        RECT -27.365 -144.325 -27.035 -143.995 ;
        RECT -27.365 -145.685 -27.035 -145.355 ;
        RECT -27.365 -147.045 -27.035 -146.715 ;
        RECT -27.365 -152.485 -27.035 -152.155 ;
        RECT -27.365 -153.845 -27.035 -153.515 ;
        RECT -27.365 -155.205 -27.035 -154.875 ;
        RECT -27.365 -156.565 -27.035 -156.235 ;
        RECT -27.365 -157.925 -27.035 -157.595 ;
        RECT -27.365 -159.285 -27.035 -158.955 ;
        RECT -27.365 -162.005 -27.035 -161.675 ;
        RECT -27.365 -163.365 -27.035 -163.035 ;
        RECT -27.365 -164.725 -27.035 -164.395 ;
        RECT -27.365 -166.085 -27.035 -165.755 ;
        RECT -27.365 -167.445 -27.035 -167.115 ;
        RECT -27.365 -168.805 -27.035 -168.475 ;
        RECT -27.365 -170.165 -27.035 -169.835 ;
        RECT -27.365 -171.525 -27.035 -171.195 ;
        RECT -27.365 -172.885 -27.035 -172.555 ;
        RECT -27.365 -174.245 -27.035 -173.915 ;
        RECT -27.365 -175.605 -27.035 -175.275 ;
        RECT -27.365 -176.965 -27.035 -176.635 ;
        RECT -27.365 -178.325 -27.035 -177.995 ;
        RECT -27.365 -179.685 -27.035 -179.355 ;
        RECT -27.365 -181.045 -27.035 -180.715 ;
        RECT -27.365 -182.405 -27.035 -182.075 ;
        RECT -27.365 -185.125 -27.035 -184.795 ;
        RECT -27.365 -186.485 -27.035 -186.155 ;
        RECT -27.365 -190.565 -27.035 -190.235 ;
        RECT -27.365 -191.925 -27.035 -191.595 ;
        RECT -27.365 -193.285 -27.035 -192.955 ;
        RECT -27.365 -194.645 -27.035 -194.315 ;
        RECT -27.365 -196.005 -27.035 -195.675 ;
        RECT -27.365 -198.725 -27.035 -198.395 ;
        RECT -27.365 -200.085 -27.035 -199.755 ;
        RECT -27.365 -201.445 -27.035 -201.115 ;
        RECT -27.365 -202.805 -27.035 -202.475 ;
        RECT -27.365 -204.165 -27.035 -203.835 ;
        RECT -27.365 -205.525 -27.035 -205.195 ;
        RECT -27.365 -208.245 -27.035 -207.915 ;
        RECT -27.365 -209.605 -27.035 -209.275 ;
        RECT -27.365 -215.045 -27.035 -214.715 ;
        RECT -27.365 -216.405 -27.035 -216.075 ;
        RECT -27.365 -217.765 -27.035 -217.435 ;
        RECT -27.365 -219.125 -27.035 -218.795 ;
        RECT -27.365 -220.485 -27.035 -220.155 ;
        RECT -27.365 -221.845 -27.035 -221.515 ;
        RECT -27.365 -223.205 -27.035 -222.875 ;
        RECT -27.365 -224.565 -27.035 -224.235 ;
        RECT -27.365 -226.155 -27.035 -225.825 ;
        RECT -27.365 -227.285 -27.035 -226.955 ;
        RECT -27.365 -231.365 -27.035 -231.035 ;
        RECT -27.365 -234.085 -27.035 -233.755 ;
        RECT -27.365 -235.445 -27.035 -235.115 ;
        RECT -27.365 -236.805 -27.035 -236.475 ;
        RECT -27.365 -238.165 -27.035 -237.835 ;
        RECT -27.365 -243.81 -27.035 -242.68 ;
        RECT -27.36 -243.925 -27.04 248.005 ;
        RECT -27.365 246.76 -27.035 247.89 ;
        RECT -27.365 241.915 -27.035 242.245 ;
        RECT -27.365 240.555 -27.035 240.885 ;
        RECT -27.365 239.195 -27.035 239.525 ;
        RECT -27.365 237.835 -27.035 238.165 ;
        RECT -27.365 236.475 -27.035 236.805 ;
        RECT -27.365 235.115 -27.035 235.445 ;
        RECT -27.365 233.755 -27.035 234.085 ;
        RECT -27.365 232.395 -27.035 232.725 ;
        RECT -27.365 231.035 -27.035 231.365 ;
        RECT -27.365 229.675 -27.035 230.005 ;
        RECT -27.365 228.315 -27.035 228.645 ;
        RECT -27.365 226.955 -27.035 227.285 ;
        RECT -27.365 225.595 -27.035 225.925 ;
        RECT -27.365 224.235 -27.035 224.565 ;
        RECT -27.365 222.875 -27.035 223.205 ;
        RECT -27.365 221.515 -27.035 221.845 ;
        RECT -27.365 220.155 -27.035 220.485 ;
        RECT -27.365 218.795 -27.035 219.125 ;
        RECT -27.365 217.435 -27.035 217.765 ;
        RECT -27.365 216.075 -27.035 216.405 ;
        RECT -27.365 214.715 -27.035 215.045 ;
        RECT -27.365 213.355 -27.035 213.685 ;
        RECT -27.365 211.995 -27.035 212.325 ;
        RECT -27.365 210.635 -27.035 210.965 ;
        RECT -27.365 209.275 -27.035 209.605 ;
        RECT -27.365 207.915 -27.035 208.245 ;
        RECT -27.365 206.555 -27.035 206.885 ;
        RECT -27.365 205.195 -27.035 205.525 ;
        RECT -27.365 203.835 -27.035 204.165 ;
        RECT -27.365 202.475 -27.035 202.805 ;
        RECT -27.365 201.115 -27.035 201.445 ;
        RECT -27.365 199.755 -27.035 200.085 ;
        RECT -27.365 198.395 -27.035 198.725 ;
        RECT -27.365 197.035 -27.035 197.365 ;
        RECT -27.365 195.675 -27.035 196.005 ;
        RECT -27.365 194.315 -27.035 194.645 ;
        RECT -27.365 192.955 -27.035 193.285 ;
        RECT -27.365 191.595 -27.035 191.925 ;
        RECT -27.365 190.235 -27.035 190.565 ;
        RECT -27.365 188.875 -27.035 189.205 ;
        RECT -27.365 187.515 -27.035 187.845 ;
        RECT -27.365 186.155 -27.035 186.485 ;
        RECT -27.365 184.795 -27.035 185.125 ;
        RECT -27.365 183.435 -27.035 183.765 ;
        RECT -27.365 182.075 -27.035 182.405 ;
        RECT -27.365 180.715 -27.035 181.045 ;
        RECT -27.365 179.355 -27.035 179.685 ;
        RECT -27.365 177.995 -27.035 178.325 ;
        RECT -27.365 176.635 -27.035 176.965 ;
        RECT -27.365 175.275 -27.035 175.605 ;
        RECT -27.365 173.915 -27.035 174.245 ;
        RECT -27.365 172.555 -27.035 172.885 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 -234.085 -35.195 -233.755 ;
        RECT -35.525 -235.445 -35.195 -235.115 ;
        RECT -35.525 -236.805 -35.195 -236.475 ;
        RECT -35.525 -238.165 -35.195 -237.835 ;
        RECT -35.525 -243.81 -35.195 -242.68 ;
        RECT -35.52 -243.925 -35.2 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.165 246.76 -33.835 247.89 ;
        RECT -34.165 241.915 -33.835 242.245 ;
        RECT -34.165 240.555 -33.835 240.885 ;
        RECT -34.165 239.195 -33.835 239.525 ;
        RECT -34.165 237.835 -33.835 238.165 ;
        RECT -34.165 236.475 -33.835 236.805 ;
        RECT -34.165 235.115 -33.835 235.445 ;
        RECT -34.165 233.755 -33.835 234.085 ;
        RECT -34.165 232.395 -33.835 232.725 ;
        RECT -34.165 231.035 -33.835 231.365 ;
        RECT -34.165 229.675 -33.835 230.005 ;
        RECT -34.165 228.315 -33.835 228.645 ;
        RECT -34.165 226.955 -33.835 227.285 ;
        RECT -34.165 225.595 -33.835 225.925 ;
        RECT -34.165 224.235 -33.835 224.565 ;
        RECT -34.165 222.875 -33.835 223.205 ;
        RECT -34.165 221.515 -33.835 221.845 ;
        RECT -34.165 220.155 -33.835 220.485 ;
        RECT -34.165 218.795 -33.835 219.125 ;
        RECT -34.165 217.435 -33.835 217.765 ;
        RECT -34.165 216.075 -33.835 216.405 ;
        RECT -34.165 214.715 -33.835 215.045 ;
        RECT -34.165 213.355 -33.835 213.685 ;
        RECT -34.165 211.995 -33.835 212.325 ;
        RECT -34.165 210.635 -33.835 210.965 ;
        RECT -34.165 209.275 -33.835 209.605 ;
        RECT -34.165 207.915 -33.835 208.245 ;
        RECT -34.165 206.555 -33.835 206.885 ;
        RECT -34.165 205.195 -33.835 205.525 ;
        RECT -34.165 203.835 -33.835 204.165 ;
        RECT -34.165 202.475 -33.835 202.805 ;
        RECT -34.165 201.115 -33.835 201.445 ;
        RECT -34.165 199.755 -33.835 200.085 ;
        RECT -34.165 198.395 -33.835 198.725 ;
        RECT -34.165 197.035 -33.835 197.365 ;
        RECT -34.165 195.675 -33.835 196.005 ;
        RECT -34.165 194.315 -33.835 194.645 ;
        RECT -34.165 192.955 -33.835 193.285 ;
        RECT -34.165 191.595 -33.835 191.925 ;
        RECT -34.165 190.235 -33.835 190.565 ;
        RECT -34.165 188.875 -33.835 189.205 ;
        RECT -34.165 187.515 -33.835 187.845 ;
        RECT -34.165 186.155 -33.835 186.485 ;
        RECT -34.165 184.795 -33.835 185.125 ;
        RECT -34.165 183.435 -33.835 183.765 ;
        RECT -34.165 182.075 -33.835 182.405 ;
        RECT -34.165 180.715 -33.835 181.045 ;
        RECT -34.165 179.355 -33.835 179.685 ;
        RECT -34.165 177.995 -33.835 178.325 ;
        RECT -34.165 176.635 -33.835 176.965 ;
        RECT -34.165 175.275 -33.835 175.605 ;
        RECT -34.165 173.915 -33.835 174.245 ;
        RECT -34.165 172.555 -33.835 172.885 ;
        RECT -34.165 171.195 -33.835 171.525 ;
        RECT -34.165 169.835 -33.835 170.165 ;
        RECT -34.165 168.475 -33.835 168.805 ;
        RECT -34.165 167.115 -33.835 167.445 ;
        RECT -34.165 165.755 -33.835 166.085 ;
        RECT -34.165 164.395 -33.835 164.725 ;
        RECT -34.165 163.035 -33.835 163.365 ;
        RECT -34.165 161.675 -33.835 162.005 ;
        RECT -34.165 160.315 -33.835 160.645 ;
        RECT -34.165 158.955 -33.835 159.285 ;
        RECT -34.165 157.595 -33.835 157.925 ;
        RECT -34.165 156.235 -33.835 156.565 ;
        RECT -34.165 154.875 -33.835 155.205 ;
        RECT -34.165 153.515 -33.835 153.845 ;
        RECT -34.165 152.155 -33.835 152.485 ;
        RECT -34.165 150.795 -33.835 151.125 ;
        RECT -34.165 149.435 -33.835 149.765 ;
        RECT -34.165 148.075 -33.835 148.405 ;
        RECT -34.165 146.715 -33.835 147.045 ;
        RECT -34.165 145.355 -33.835 145.685 ;
        RECT -34.165 143.995 -33.835 144.325 ;
        RECT -34.165 142.635 -33.835 142.965 ;
        RECT -34.165 141.275 -33.835 141.605 ;
        RECT -34.165 139.915 -33.835 140.245 ;
        RECT -34.165 138.555 -33.835 138.885 ;
        RECT -34.165 137.195 -33.835 137.525 ;
        RECT -34.165 135.835 -33.835 136.165 ;
        RECT -34.165 134.475 -33.835 134.805 ;
        RECT -34.165 133.115 -33.835 133.445 ;
        RECT -34.165 131.755 -33.835 132.085 ;
        RECT -34.165 130.395 -33.835 130.725 ;
        RECT -34.165 129.035 -33.835 129.365 ;
        RECT -34.165 127.675 -33.835 128.005 ;
        RECT -34.165 126.315 -33.835 126.645 ;
        RECT -34.165 124.955 -33.835 125.285 ;
        RECT -34.165 123.595 -33.835 123.925 ;
        RECT -34.165 122.235 -33.835 122.565 ;
        RECT -34.165 120.875 -33.835 121.205 ;
        RECT -34.165 119.515 -33.835 119.845 ;
        RECT -34.165 118.155 -33.835 118.485 ;
        RECT -34.165 116.795 -33.835 117.125 ;
        RECT -34.165 115.435 -33.835 115.765 ;
        RECT -34.165 114.075 -33.835 114.405 ;
        RECT -34.165 112.715 -33.835 113.045 ;
        RECT -34.165 111.355 -33.835 111.685 ;
        RECT -34.165 109.995 -33.835 110.325 ;
        RECT -34.165 108.635 -33.835 108.965 ;
        RECT -34.165 107.275 -33.835 107.605 ;
        RECT -34.165 105.915 -33.835 106.245 ;
        RECT -34.165 104.555 -33.835 104.885 ;
        RECT -34.165 103.195 -33.835 103.525 ;
        RECT -34.165 101.835 -33.835 102.165 ;
        RECT -34.165 100.475 -33.835 100.805 ;
        RECT -34.165 99.115 -33.835 99.445 ;
        RECT -34.165 97.755 -33.835 98.085 ;
        RECT -34.165 96.395 -33.835 96.725 ;
        RECT -34.165 95.035 -33.835 95.365 ;
        RECT -34.165 93.675 -33.835 94.005 ;
        RECT -34.165 92.315 -33.835 92.645 ;
        RECT -34.165 90.955 -33.835 91.285 ;
        RECT -34.165 89.595 -33.835 89.925 ;
        RECT -34.165 88.235 -33.835 88.565 ;
        RECT -34.165 86.875 -33.835 87.205 ;
        RECT -34.165 85.515 -33.835 85.845 ;
        RECT -34.165 84.155 -33.835 84.485 ;
        RECT -34.165 82.795 -33.835 83.125 ;
        RECT -34.165 81.435 -33.835 81.765 ;
        RECT -34.165 80.075 -33.835 80.405 ;
        RECT -34.165 78.715 -33.835 79.045 ;
        RECT -34.165 77.355 -33.835 77.685 ;
        RECT -34.165 75.995 -33.835 76.325 ;
        RECT -34.165 74.635 -33.835 74.965 ;
        RECT -34.165 73.275 -33.835 73.605 ;
        RECT -34.165 71.915 -33.835 72.245 ;
        RECT -34.165 70.555 -33.835 70.885 ;
        RECT -34.165 69.195 -33.835 69.525 ;
        RECT -34.165 67.835 -33.835 68.165 ;
        RECT -34.165 66.475 -33.835 66.805 ;
        RECT -34.165 65.115 -33.835 65.445 ;
        RECT -34.165 63.755 -33.835 64.085 ;
        RECT -34.165 62.395 -33.835 62.725 ;
        RECT -34.165 61.035 -33.835 61.365 ;
        RECT -34.165 59.675 -33.835 60.005 ;
        RECT -34.165 58.315 -33.835 58.645 ;
        RECT -34.165 56.955 -33.835 57.285 ;
        RECT -34.165 55.595 -33.835 55.925 ;
        RECT -34.165 54.235 -33.835 54.565 ;
        RECT -34.165 52.875 -33.835 53.205 ;
        RECT -34.165 51.515 -33.835 51.845 ;
        RECT -34.165 50.155 -33.835 50.485 ;
        RECT -34.165 48.795 -33.835 49.125 ;
        RECT -34.165 47.435 -33.835 47.765 ;
        RECT -34.165 46.075 -33.835 46.405 ;
        RECT -34.165 44.715 -33.835 45.045 ;
        RECT -34.165 43.355 -33.835 43.685 ;
        RECT -34.165 41.995 -33.835 42.325 ;
        RECT -34.165 40.635 -33.835 40.965 ;
        RECT -34.165 39.275 -33.835 39.605 ;
        RECT -34.165 37.915 -33.835 38.245 ;
        RECT -34.165 36.555 -33.835 36.885 ;
        RECT -34.165 35.195 -33.835 35.525 ;
        RECT -34.165 33.835 -33.835 34.165 ;
        RECT -34.165 32.475 -33.835 32.805 ;
        RECT -34.165 31.115 -33.835 31.445 ;
        RECT -34.165 29.755 -33.835 30.085 ;
        RECT -34.165 28.395 -33.835 28.725 ;
        RECT -34.165 27.035 -33.835 27.365 ;
        RECT -34.165 25.675 -33.835 26.005 ;
        RECT -34.165 24.315 -33.835 24.645 ;
        RECT -34.165 22.955 -33.835 23.285 ;
        RECT -34.165 21.595 -33.835 21.925 ;
        RECT -34.165 20.235 -33.835 20.565 ;
        RECT -34.165 18.875 -33.835 19.205 ;
        RECT -34.165 17.515 -33.835 17.845 ;
        RECT -34.165 16.155 -33.835 16.485 ;
        RECT -34.165 14.795 -33.835 15.125 ;
        RECT -34.165 13.435 -33.835 13.765 ;
        RECT -34.165 12.075 -33.835 12.405 ;
        RECT -34.165 10.715 -33.835 11.045 ;
        RECT -34.165 9.355 -33.835 9.685 ;
        RECT -34.165 7.995 -33.835 8.325 ;
        RECT -34.165 6.635 -33.835 6.965 ;
        RECT -34.165 5.275 -33.835 5.605 ;
        RECT -34.165 3.915 -33.835 4.245 ;
        RECT -34.165 2.555 -33.835 2.885 ;
        RECT -34.165 1.195 -33.835 1.525 ;
        RECT -34.165 -0.165 -33.835 0.165 ;
        RECT -34.165 -1.525 -33.835 -1.195 ;
        RECT -34.165 -8.325 -33.835 -7.995 ;
        RECT -34.165 -9.685 -33.835 -9.355 ;
        RECT -34.165 -12.405 -33.835 -12.075 ;
        RECT -34.165 -13.765 -33.835 -13.435 ;
        RECT -34.165 -15.125 -33.835 -14.795 ;
        RECT -34.165 -16.485 -33.835 -16.155 ;
        RECT -34.165 -17.845 -33.835 -17.515 ;
        RECT -34.165 -19.205 -33.835 -18.875 ;
        RECT -34.165 -20.565 -33.835 -20.235 ;
        RECT -34.165 -21.925 -33.835 -21.595 ;
        RECT -34.165 -23.285 -33.835 -22.955 ;
        RECT -34.165 -30.66 -33.835 -30.33 ;
        RECT -34.165 -31.445 -33.835 -31.115 ;
        RECT -34.165 -32.805 -33.835 -32.475 ;
        RECT -34.165 -34.165 -33.835 -33.835 ;
        RECT -34.165 -36.885 -33.835 -36.555 ;
        RECT -34.165 -37.85 -33.835 -37.52 ;
        RECT -34.165 -40.965 -33.835 -40.635 ;
        RECT -34.165 -46.405 -33.835 -46.075 ;
        RECT -34.165 -49.125 -33.835 -48.795 ;
        RECT -34.165 -50.485 -33.835 -50.155 ;
        RECT -34.165 -53.205 -33.835 -52.875 ;
        RECT -34.165 -55.925 -33.835 -55.595 ;
        RECT -34.165 -61.365 -33.835 -61.035 ;
        RECT -34.165 -62.725 -33.835 -62.395 ;
        RECT -34.165 -64.085 -33.835 -63.755 ;
        RECT -34.165 -65.445 -33.835 -65.115 ;
        RECT -34.165 -66.805 -33.835 -66.475 ;
        RECT -34.165 -68.165 -33.835 -67.835 ;
        RECT -34.165 -69.525 -33.835 -69.195 ;
        RECT -34.165 -70.885 -33.835 -70.555 ;
        RECT -34.165 -72.245 -33.835 -71.915 ;
        RECT -34.165 -73.605 -33.835 -73.275 ;
        RECT -34.165 -74.965 -33.835 -74.635 ;
        RECT -34.165 -76.325 -33.835 -75.995 ;
        RECT -34.165 -77.685 -33.835 -77.355 ;
        RECT -34.165 -79.045 -33.835 -78.715 ;
        RECT -34.165 -80.405 -33.835 -80.075 ;
        RECT -34.165 -81.765 -33.835 -81.435 ;
        RECT -34.165 -83.125 -33.835 -82.795 ;
        RECT -34.165 -84.485 -33.835 -84.155 ;
        RECT -34.165 -85.845 -33.835 -85.515 ;
        RECT -34.165 -87.205 -33.835 -86.875 ;
        RECT -34.165 -88.565 -33.835 -88.235 ;
        RECT -34.165 -89.925 -33.835 -89.595 ;
        RECT -34.165 -91.285 -33.835 -90.955 ;
        RECT -34.165 -92.645 -33.835 -92.315 ;
        RECT -34.165 -94.005 -33.835 -93.675 ;
        RECT -34.165 -95.365 -33.835 -95.035 ;
        RECT -34.165 -96.725 -33.835 -96.395 ;
        RECT -34.165 -98.085 -33.835 -97.755 ;
        RECT -34.165 -99.445 -33.835 -99.115 ;
        RECT -34.165 -100.805 -33.835 -100.475 ;
        RECT -34.165 -102.165 -33.835 -101.835 ;
        RECT -34.165 -103.525 -33.835 -103.195 ;
        RECT -34.165 -104.885 -33.835 -104.555 ;
        RECT -34.165 -106.245 -33.835 -105.915 ;
        RECT -34.165 -107.605 -33.835 -107.275 ;
        RECT -34.165 -108.965 -33.835 -108.635 ;
        RECT -34.165 -110.325 -33.835 -109.995 ;
        RECT -34.165 -111.685 -33.835 -111.355 ;
        RECT -34.165 -113.045 -33.835 -112.715 ;
        RECT -34.165 -114.405 -33.835 -114.075 ;
        RECT -34.165 -115.765 -33.835 -115.435 ;
        RECT -34.165 -117.125 -33.835 -116.795 ;
        RECT -34.165 -118.485 -33.835 -118.155 ;
        RECT -34.165 -119.845 -33.835 -119.515 ;
        RECT -34.165 -123.925 -33.835 -123.595 ;
        RECT -34.165 -129.365 -33.835 -129.035 ;
        RECT -34.165 -130.725 -33.835 -130.395 ;
        RECT -34.165 -132.085 -33.835 -131.755 ;
        RECT -34.165 -133.445 -33.835 -133.115 ;
        RECT -34.165 -134.805 -33.835 -134.475 ;
        RECT -34.165 -136.165 -33.835 -135.835 ;
        RECT -34.165 -137.525 -33.835 -137.195 ;
        RECT -34.165 -138.885 -33.835 -138.555 ;
        RECT -34.165 -140.245 -33.835 -139.915 ;
        RECT -34.165 -141.605 -33.835 -141.275 ;
        RECT -34.165 -142.965 -33.835 -142.635 ;
        RECT -34.165 -144.325 -33.835 -143.995 ;
        RECT -34.165 -145.685 -33.835 -145.355 ;
        RECT -34.165 -147.045 -33.835 -146.715 ;
        RECT -34.165 -148.405 -33.835 -148.075 ;
        RECT -34.165 -149.765 -33.835 -149.435 ;
        RECT -34.165 -151.125 -33.835 -150.795 ;
        RECT -34.165 -152.485 -33.835 -152.155 ;
        RECT -34.165 -153.845 -33.835 -153.515 ;
        RECT -34.165 -155.205 -33.835 -154.875 ;
        RECT -34.165 -156.565 -33.835 -156.235 ;
        RECT -34.165 -157.925 -33.835 -157.595 ;
        RECT -34.165 -159.285 -33.835 -158.955 ;
        RECT -34.165 -162.005 -33.835 -161.675 ;
        RECT -34.165 -163.365 -33.835 -163.035 ;
        RECT -34.165 -164.725 -33.835 -164.395 ;
        RECT -34.165 -166.085 -33.835 -165.755 ;
        RECT -34.165 -167.445 -33.835 -167.115 ;
        RECT -34.165 -168.805 -33.835 -168.475 ;
        RECT -34.165 -170.165 -33.835 -169.835 ;
        RECT -34.165 -171.525 -33.835 -171.195 ;
        RECT -34.165 -172.885 -33.835 -172.555 ;
        RECT -34.165 -174.245 -33.835 -173.915 ;
        RECT -34.165 -175.605 -33.835 -175.275 ;
        RECT -34.165 -176.965 -33.835 -176.635 ;
        RECT -34.165 -178.325 -33.835 -177.995 ;
        RECT -34.165 -179.685 -33.835 -179.355 ;
        RECT -34.165 -181.045 -33.835 -180.715 ;
        RECT -34.165 -182.405 -33.835 -182.075 ;
        RECT -34.165 -183.765 -33.835 -183.435 ;
        RECT -34.165 -185.125 -33.835 -184.795 ;
        RECT -34.165 -186.485 -33.835 -186.155 ;
        RECT -34.165 -187.845 -33.835 -187.515 ;
        RECT -34.165 -190.565 -33.835 -190.235 ;
        RECT -34.165 -191.925 -33.835 -191.595 ;
        RECT -34.165 -193.285 -33.835 -192.955 ;
        RECT -34.165 -194.645 -33.835 -194.315 ;
        RECT -34.165 -196.005 -33.835 -195.675 ;
        RECT -34.165 -197.365 -33.835 -197.035 ;
        RECT -34.165 -198.725 -33.835 -198.395 ;
        RECT -34.165 -200.085 -33.835 -199.755 ;
        RECT -34.165 -201.445 -33.835 -201.115 ;
        RECT -34.165 -202.805 -33.835 -202.475 ;
        RECT -34.165 -204.165 -33.835 -203.835 ;
        RECT -34.165 -205.525 -33.835 -205.195 ;
        RECT -34.165 -208.245 -33.835 -207.915 ;
        RECT -34.165 -209.605 -33.835 -209.275 ;
        RECT -34.165 -212.325 -33.835 -211.995 ;
        RECT -34.165 -215.045 -33.835 -214.715 ;
        RECT -34.165 -216.405 -33.835 -216.075 ;
        RECT -34.165 -217.765 -33.835 -217.435 ;
        RECT -34.165 -219.125 -33.835 -218.795 ;
        RECT -34.165 -220.485 -33.835 -220.155 ;
        RECT -34.165 -221.845 -33.835 -221.515 ;
        RECT -34.165 -223.205 -33.835 -222.875 ;
        RECT -34.165 -224.565 -33.835 -224.235 ;
        RECT -34.165 -226.155 -33.835 -225.825 ;
        RECT -34.165 -227.285 -33.835 -226.955 ;
        RECT -34.165 -228.645 -33.835 -228.315 ;
        RECT -34.16 -229.32 -33.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.805 246.76 -32.475 247.89 ;
        RECT -32.805 241.915 -32.475 242.245 ;
        RECT -32.805 240.555 -32.475 240.885 ;
        RECT -32.805 239.195 -32.475 239.525 ;
        RECT -32.805 237.835 -32.475 238.165 ;
        RECT -32.805 236.475 -32.475 236.805 ;
        RECT -32.805 235.115 -32.475 235.445 ;
        RECT -32.805 233.755 -32.475 234.085 ;
        RECT -32.805 232.395 -32.475 232.725 ;
        RECT -32.805 231.035 -32.475 231.365 ;
        RECT -32.805 229.675 -32.475 230.005 ;
        RECT -32.805 228.315 -32.475 228.645 ;
        RECT -32.805 226.955 -32.475 227.285 ;
        RECT -32.805 225.595 -32.475 225.925 ;
        RECT -32.805 224.235 -32.475 224.565 ;
        RECT -32.805 222.875 -32.475 223.205 ;
        RECT -32.805 221.515 -32.475 221.845 ;
        RECT -32.805 220.155 -32.475 220.485 ;
        RECT -32.805 218.795 -32.475 219.125 ;
        RECT -32.805 217.435 -32.475 217.765 ;
        RECT -32.805 216.075 -32.475 216.405 ;
        RECT -32.805 214.715 -32.475 215.045 ;
        RECT -32.805 213.355 -32.475 213.685 ;
        RECT -32.805 211.995 -32.475 212.325 ;
        RECT -32.805 210.635 -32.475 210.965 ;
        RECT -32.805 209.275 -32.475 209.605 ;
        RECT -32.805 207.915 -32.475 208.245 ;
        RECT -32.805 206.555 -32.475 206.885 ;
        RECT -32.805 205.195 -32.475 205.525 ;
        RECT -32.805 203.835 -32.475 204.165 ;
        RECT -32.805 202.475 -32.475 202.805 ;
        RECT -32.805 201.115 -32.475 201.445 ;
        RECT -32.805 199.755 -32.475 200.085 ;
        RECT -32.805 198.395 -32.475 198.725 ;
        RECT -32.805 197.035 -32.475 197.365 ;
        RECT -32.805 195.675 -32.475 196.005 ;
        RECT -32.805 194.315 -32.475 194.645 ;
        RECT -32.805 192.955 -32.475 193.285 ;
        RECT -32.805 191.595 -32.475 191.925 ;
        RECT -32.805 190.235 -32.475 190.565 ;
        RECT -32.805 188.875 -32.475 189.205 ;
        RECT -32.805 187.515 -32.475 187.845 ;
        RECT -32.805 186.155 -32.475 186.485 ;
        RECT -32.805 184.795 -32.475 185.125 ;
        RECT -32.805 183.435 -32.475 183.765 ;
        RECT -32.805 182.075 -32.475 182.405 ;
        RECT -32.805 180.715 -32.475 181.045 ;
        RECT -32.805 179.355 -32.475 179.685 ;
        RECT -32.805 177.995 -32.475 178.325 ;
        RECT -32.805 176.635 -32.475 176.965 ;
        RECT -32.805 175.275 -32.475 175.605 ;
        RECT -32.805 173.915 -32.475 174.245 ;
        RECT -32.805 172.555 -32.475 172.885 ;
        RECT -32.805 171.195 -32.475 171.525 ;
        RECT -32.805 169.835 -32.475 170.165 ;
        RECT -32.805 168.475 -32.475 168.805 ;
        RECT -32.805 167.115 -32.475 167.445 ;
        RECT -32.805 165.755 -32.475 166.085 ;
        RECT -32.805 164.395 -32.475 164.725 ;
        RECT -32.805 163.035 -32.475 163.365 ;
        RECT -32.805 161.675 -32.475 162.005 ;
        RECT -32.805 160.315 -32.475 160.645 ;
        RECT -32.805 158.955 -32.475 159.285 ;
        RECT -32.805 157.595 -32.475 157.925 ;
        RECT -32.805 156.235 -32.475 156.565 ;
        RECT -32.805 154.875 -32.475 155.205 ;
        RECT -32.805 153.515 -32.475 153.845 ;
        RECT -32.805 152.155 -32.475 152.485 ;
        RECT -32.805 150.795 -32.475 151.125 ;
        RECT -32.805 149.435 -32.475 149.765 ;
        RECT -32.805 148.075 -32.475 148.405 ;
        RECT -32.805 146.715 -32.475 147.045 ;
        RECT -32.805 145.355 -32.475 145.685 ;
        RECT -32.805 143.995 -32.475 144.325 ;
        RECT -32.805 142.635 -32.475 142.965 ;
        RECT -32.805 141.275 -32.475 141.605 ;
        RECT -32.805 139.915 -32.475 140.245 ;
        RECT -32.805 138.555 -32.475 138.885 ;
        RECT -32.805 137.195 -32.475 137.525 ;
        RECT -32.805 135.835 -32.475 136.165 ;
        RECT -32.805 134.475 -32.475 134.805 ;
        RECT -32.805 133.115 -32.475 133.445 ;
        RECT -32.805 131.755 -32.475 132.085 ;
        RECT -32.805 130.395 -32.475 130.725 ;
        RECT -32.805 129.035 -32.475 129.365 ;
        RECT -32.805 127.675 -32.475 128.005 ;
        RECT -32.805 126.315 -32.475 126.645 ;
        RECT -32.805 124.955 -32.475 125.285 ;
        RECT -32.805 123.595 -32.475 123.925 ;
        RECT -32.805 122.235 -32.475 122.565 ;
        RECT -32.805 120.875 -32.475 121.205 ;
        RECT -32.805 119.515 -32.475 119.845 ;
        RECT -32.805 118.155 -32.475 118.485 ;
        RECT -32.805 116.795 -32.475 117.125 ;
        RECT -32.805 115.435 -32.475 115.765 ;
        RECT -32.805 114.075 -32.475 114.405 ;
        RECT -32.805 112.715 -32.475 113.045 ;
        RECT -32.805 111.355 -32.475 111.685 ;
        RECT -32.805 109.995 -32.475 110.325 ;
        RECT -32.805 108.635 -32.475 108.965 ;
        RECT -32.805 107.275 -32.475 107.605 ;
        RECT -32.805 105.915 -32.475 106.245 ;
        RECT -32.805 104.555 -32.475 104.885 ;
        RECT -32.805 103.195 -32.475 103.525 ;
        RECT -32.805 101.835 -32.475 102.165 ;
        RECT -32.805 100.475 -32.475 100.805 ;
        RECT -32.805 99.115 -32.475 99.445 ;
        RECT -32.805 97.755 -32.475 98.085 ;
        RECT -32.805 96.395 -32.475 96.725 ;
        RECT -32.805 95.035 -32.475 95.365 ;
        RECT -32.805 93.675 -32.475 94.005 ;
        RECT -32.805 92.315 -32.475 92.645 ;
        RECT -32.805 90.955 -32.475 91.285 ;
        RECT -32.805 89.595 -32.475 89.925 ;
        RECT -32.805 88.235 -32.475 88.565 ;
        RECT -32.805 86.875 -32.475 87.205 ;
        RECT -32.805 85.515 -32.475 85.845 ;
        RECT -32.805 84.155 -32.475 84.485 ;
        RECT -32.805 82.795 -32.475 83.125 ;
        RECT -32.805 81.435 -32.475 81.765 ;
        RECT -32.805 80.075 -32.475 80.405 ;
        RECT -32.805 78.715 -32.475 79.045 ;
        RECT -32.805 77.355 -32.475 77.685 ;
        RECT -32.805 75.995 -32.475 76.325 ;
        RECT -32.805 74.635 -32.475 74.965 ;
        RECT -32.805 73.275 -32.475 73.605 ;
        RECT -32.805 71.915 -32.475 72.245 ;
        RECT -32.805 70.555 -32.475 70.885 ;
        RECT -32.805 69.195 -32.475 69.525 ;
        RECT -32.805 67.835 -32.475 68.165 ;
        RECT -32.805 66.475 -32.475 66.805 ;
        RECT -32.805 65.115 -32.475 65.445 ;
        RECT -32.805 63.755 -32.475 64.085 ;
        RECT -32.805 62.395 -32.475 62.725 ;
        RECT -32.805 61.035 -32.475 61.365 ;
        RECT -32.805 59.675 -32.475 60.005 ;
        RECT -32.805 58.315 -32.475 58.645 ;
        RECT -32.805 56.955 -32.475 57.285 ;
        RECT -32.805 55.595 -32.475 55.925 ;
        RECT -32.805 54.235 -32.475 54.565 ;
        RECT -32.805 52.875 -32.475 53.205 ;
        RECT -32.805 51.515 -32.475 51.845 ;
        RECT -32.805 50.155 -32.475 50.485 ;
        RECT -32.805 48.795 -32.475 49.125 ;
        RECT -32.805 47.435 -32.475 47.765 ;
        RECT -32.805 46.075 -32.475 46.405 ;
        RECT -32.805 44.715 -32.475 45.045 ;
        RECT -32.805 43.355 -32.475 43.685 ;
        RECT -32.805 41.995 -32.475 42.325 ;
        RECT -32.805 40.635 -32.475 40.965 ;
        RECT -32.805 39.275 -32.475 39.605 ;
        RECT -32.805 37.915 -32.475 38.245 ;
        RECT -32.805 36.555 -32.475 36.885 ;
        RECT -32.805 35.195 -32.475 35.525 ;
        RECT -32.805 33.835 -32.475 34.165 ;
        RECT -32.805 32.475 -32.475 32.805 ;
        RECT -32.805 31.115 -32.475 31.445 ;
        RECT -32.805 29.755 -32.475 30.085 ;
        RECT -32.805 28.395 -32.475 28.725 ;
        RECT -32.805 27.035 -32.475 27.365 ;
        RECT -32.805 25.675 -32.475 26.005 ;
        RECT -32.805 24.315 -32.475 24.645 ;
        RECT -32.805 22.955 -32.475 23.285 ;
        RECT -32.805 21.595 -32.475 21.925 ;
        RECT -32.805 20.235 -32.475 20.565 ;
        RECT -32.805 18.875 -32.475 19.205 ;
        RECT -32.805 17.515 -32.475 17.845 ;
        RECT -32.805 16.155 -32.475 16.485 ;
        RECT -32.805 14.795 -32.475 15.125 ;
        RECT -32.805 13.435 -32.475 13.765 ;
        RECT -32.805 12.075 -32.475 12.405 ;
        RECT -32.805 10.715 -32.475 11.045 ;
        RECT -32.805 9.355 -32.475 9.685 ;
        RECT -32.805 7.995 -32.475 8.325 ;
        RECT -32.805 6.635 -32.475 6.965 ;
        RECT -32.805 5.275 -32.475 5.605 ;
        RECT -32.805 3.915 -32.475 4.245 ;
        RECT -32.805 2.555 -32.475 2.885 ;
        RECT -32.805 1.195 -32.475 1.525 ;
        RECT -32.805 -0.165 -32.475 0.165 ;
        RECT -32.805 -8.325 -32.475 -7.995 ;
        RECT -32.805 -9.685 -32.475 -9.355 ;
        RECT -32.805 -12.405 -32.475 -12.075 ;
        RECT -32.805 -13.765 -32.475 -13.435 ;
        RECT -32.805 -15.125 -32.475 -14.795 ;
        RECT -32.805 -16.485 -32.475 -16.155 ;
        RECT -32.805 -17.845 -32.475 -17.515 ;
        RECT -32.805 -19.205 -32.475 -18.875 ;
        RECT -32.805 -20.565 -32.475 -20.235 ;
        RECT -32.805 -21.925 -32.475 -21.595 ;
        RECT -32.805 -23.285 -32.475 -22.955 ;
        RECT -32.805 -30.66 -32.475 -30.33 ;
        RECT -32.805 -31.445 -32.475 -31.115 ;
        RECT -32.805 -32.805 -32.475 -32.475 ;
        RECT -32.805 -34.165 -32.475 -33.835 ;
        RECT -32.805 -36.885 -32.475 -36.555 ;
        RECT -32.805 -37.85 -32.475 -37.52 ;
        RECT -32.805 -40.965 -32.475 -40.635 ;
        RECT -32.805 -46.405 -32.475 -46.075 ;
        RECT -32.805 -49.125 -32.475 -48.795 ;
        RECT -32.805 -50.485 -32.475 -50.155 ;
        RECT -32.805 -53.205 -32.475 -52.875 ;
        RECT -32.805 -55.925 -32.475 -55.595 ;
        RECT -32.805 -61.365 -32.475 -61.035 ;
        RECT -32.805 -62.725 -32.475 -62.395 ;
        RECT -32.805 -64.085 -32.475 -63.755 ;
        RECT -32.805 -65.445 -32.475 -65.115 ;
        RECT -32.805 -66.805 -32.475 -66.475 ;
        RECT -32.805 -68.165 -32.475 -67.835 ;
        RECT -32.805 -69.525 -32.475 -69.195 ;
        RECT -32.805 -70.885 -32.475 -70.555 ;
        RECT -32.805 -72.245 -32.475 -71.915 ;
        RECT -32.805 -73.605 -32.475 -73.275 ;
        RECT -32.805 -74.965 -32.475 -74.635 ;
        RECT -32.805 -76.325 -32.475 -75.995 ;
        RECT -32.805 -77.685 -32.475 -77.355 ;
        RECT -32.805 -79.045 -32.475 -78.715 ;
        RECT -32.805 -80.405 -32.475 -80.075 ;
        RECT -32.805 -81.765 -32.475 -81.435 ;
        RECT -32.805 -83.125 -32.475 -82.795 ;
        RECT -32.805 -84.485 -32.475 -84.155 ;
        RECT -32.805 -85.845 -32.475 -85.515 ;
        RECT -32.805 -87.205 -32.475 -86.875 ;
        RECT -32.805 -88.565 -32.475 -88.235 ;
        RECT -32.805 -89.925 -32.475 -89.595 ;
        RECT -32.805 -91.285 -32.475 -90.955 ;
        RECT -32.805 -92.645 -32.475 -92.315 ;
        RECT -32.805 -94.005 -32.475 -93.675 ;
        RECT -32.805 -95.365 -32.475 -95.035 ;
        RECT -32.805 -96.725 -32.475 -96.395 ;
        RECT -32.805 -98.085 -32.475 -97.755 ;
        RECT -32.805 -99.445 -32.475 -99.115 ;
        RECT -32.805 -100.805 -32.475 -100.475 ;
        RECT -32.805 -102.165 -32.475 -101.835 ;
        RECT -32.805 -103.525 -32.475 -103.195 ;
        RECT -32.805 -104.885 -32.475 -104.555 ;
        RECT -32.805 -106.245 -32.475 -105.915 ;
        RECT -32.805 -107.605 -32.475 -107.275 ;
        RECT -32.805 -108.965 -32.475 -108.635 ;
        RECT -32.805 -110.325 -32.475 -109.995 ;
        RECT -32.805 -111.685 -32.475 -111.355 ;
        RECT -32.805 -113.045 -32.475 -112.715 ;
        RECT -32.805 -114.405 -32.475 -114.075 ;
        RECT -32.805 -115.765 -32.475 -115.435 ;
        RECT -32.805 -117.125 -32.475 -116.795 ;
        RECT -32.805 -118.485 -32.475 -118.155 ;
        RECT -32.805 -119.845 -32.475 -119.515 ;
        RECT -32.805 -123.925 -32.475 -123.595 ;
        RECT -32.805 -129.365 -32.475 -129.035 ;
        RECT -32.805 -130.725 -32.475 -130.395 ;
        RECT -32.805 -132.085 -32.475 -131.755 ;
        RECT -32.805 -133.445 -32.475 -133.115 ;
        RECT -32.805 -134.805 -32.475 -134.475 ;
        RECT -32.805 -136.165 -32.475 -135.835 ;
        RECT -32.805 -137.525 -32.475 -137.195 ;
        RECT -32.805 -138.885 -32.475 -138.555 ;
        RECT -32.805 -140.245 -32.475 -139.915 ;
        RECT -32.805 -141.605 -32.475 -141.275 ;
        RECT -32.805 -142.965 -32.475 -142.635 ;
        RECT -32.805 -144.325 -32.475 -143.995 ;
        RECT -32.805 -145.685 -32.475 -145.355 ;
        RECT -32.805 -147.045 -32.475 -146.715 ;
        RECT -32.805 -148.405 -32.475 -148.075 ;
        RECT -32.805 -149.765 -32.475 -149.435 ;
        RECT -32.805 -151.125 -32.475 -150.795 ;
        RECT -32.805 -152.485 -32.475 -152.155 ;
        RECT -32.805 -153.845 -32.475 -153.515 ;
        RECT -32.805 -155.205 -32.475 -154.875 ;
        RECT -32.805 -156.565 -32.475 -156.235 ;
        RECT -32.805 -157.925 -32.475 -157.595 ;
        RECT -32.805 -159.285 -32.475 -158.955 ;
        RECT -32.805 -162.005 -32.475 -161.675 ;
        RECT -32.805 -163.365 -32.475 -163.035 ;
        RECT -32.805 -164.725 -32.475 -164.395 ;
        RECT -32.805 -166.085 -32.475 -165.755 ;
        RECT -32.805 -167.445 -32.475 -167.115 ;
        RECT -32.805 -168.805 -32.475 -168.475 ;
        RECT -32.805 -170.165 -32.475 -169.835 ;
        RECT -32.805 -171.525 -32.475 -171.195 ;
        RECT -32.805 -172.885 -32.475 -172.555 ;
        RECT -32.805 -174.245 -32.475 -173.915 ;
        RECT -32.805 -175.605 -32.475 -175.275 ;
        RECT -32.805 -176.965 -32.475 -176.635 ;
        RECT -32.805 -178.325 -32.475 -177.995 ;
        RECT -32.805 -179.685 -32.475 -179.355 ;
        RECT -32.805 -181.045 -32.475 -180.715 ;
        RECT -32.805 -182.405 -32.475 -182.075 ;
        RECT -32.805 -183.765 -32.475 -183.435 ;
        RECT -32.805 -185.125 -32.475 -184.795 ;
        RECT -32.805 -186.485 -32.475 -186.155 ;
        RECT -32.805 -190.565 -32.475 -190.235 ;
        RECT -32.805 -191.925 -32.475 -191.595 ;
        RECT -32.805 -193.285 -32.475 -192.955 ;
        RECT -32.805 -194.645 -32.475 -194.315 ;
        RECT -32.805 -196.005 -32.475 -195.675 ;
        RECT -32.805 -197.365 -32.475 -197.035 ;
        RECT -32.805 -198.725 -32.475 -198.395 ;
        RECT -32.805 -200.085 -32.475 -199.755 ;
        RECT -32.805 -201.445 -32.475 -201.115 ;
        RECT -32.805 -202.805 -32.475 -202.475 ;
        RECT -32.805 -204.165 -32.475 -203.835 ;
        RECT -32.805 -205.525 -32.475 -205.195 ;
        RECT -32.805 -208.245 -32.475 -207.915 ;
        RECT -32.805 -209.605 -32.475 -209.275 ;
        RECT -32.805 -212.325 -32.475 -211.995 ;
        RECT -32.805 -213.685 -32.475 -213.355 ;
        RECT -32.805 -215.045 -32.475 -214.715 ;
        RECT -32.805 -216.405 -32.475 -216.075 ;
        RECT -32.805 -217.765 -32.475 -217.435 ;
        RECT -32.805 -219.125 -32.475 -218.795 ;
        RECT -32.805 -220.485 -32.475 -220.155 ;
        RECT -32.805 -221.845 -32.475 -221.515 ;
        RECT -32.805 -223.205 -32.475 -222.875 ;
        RECT -32.805 -224.565 -32.475 -224.235 ;
        RECT -32.805 -226.155 -32.475 -225.825 ;
        RECT -32.805 -227.285 -32.475 -226.955 ;
        RECT -32.805 -228.645 -32.475 -228.315 ;
        RECT -32.805 -231.365 -32.475 -231.035 ;
        RECT -32.805 -234.085 -32.475 -233.755 ;
        RECT -32.805 -235.445 -32.475 -235.115 ;
        RECT -32.805 -236.805 -32.475 -236.475 ;
        RECT -32.805 -238.165 -32.475 -237.835 ;
        RECT -32.805 -243.81 -32.475 -242.68 ;
        RECT -32.8 -243.925 -32.48 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.445 -61.365 -31.115 -61.035 ;
        RECT -31.445 -62.725 -31.115 -62.395 ;
        RECT -31.445 -64.085 -31.115 -63.755 ;
        RECT -31.445 -65.445 -31.115 -65.115 ;
        RECT -31.445 -66.805 -31.115 -66.475 ;
        RECT -31.445 -68.165 -31.115 -67.835 ;
        RECT -31.445 -69.525 -31.115 -69.195 ;
        RECT -31.445 -70.885 -31.115 -70.555 ;
        RECT -31.445 -72.245 -31.115 -71.915 ;
        RECT -31.445 -73.605 -31.115 -73.275 ;
        RECT -31.445 -74.965 -31.115 -74.635 ;
        RECT -31.445 -76.325 -31.115 -75.995 ;
        RECT -31.445 -77.685 -31.115 -77.355 ;
        RECT -31.445 -79.045 -31.115 -78.715 ;
        RECT -31.445 -80.405 -31.115 -80.075 ;
        RECT -31.445 -81.765 -31.115 -81.435 ;
        RECT -31.445 -83.125 -31.115 -82.795 ;
        RECT -31.445 -84.485 -31.115 -84.155 ;
        RECT -31.445 -85.845 -31.115 -85.515 ;
        RECT -31.445 -87.205 -31.115 -86.875 ;
        RECT -31.445 -88.565 -31.115 -88.235 ;
        RECT -31.445 -89.925 -31.115 -89.595 ;
        RECT -31.445 -91.285 -31.115 -90.955 ;
        RECT -31.445 -92.645 -31.115 -92.315 ;
        RECT -31.445 -94.005 -31.115 -93.675 ;
        RECT -31.445 -95.365 -31.115 -95.035 ;
        RECT -31.445 -96.725 -31.115 -96.395 ;
        RECT -31.445 -98.085 -31.115 -97.755 ;
        RECT -31.445 -99.445 -31.115 -99.115 ;
        RECT -31.445 -100.805 -31.115 -100.475 ;
        RECT -31.445 -102.165 -31.115 -101.835 ;
        RECT -31.445 -103.525 -31.115 -103.195 ;
        RECT -31.445 -104.885 -31.115 -104.555 ;
        RECT -31.445 -106.245 -31.115 -105.915 ;
        RECT -31.445 -107.605 -31.115 -107.275 ;
        RECT -31.445 -108.965 -31.115 -108.635 ;
        RECT -31.445 -110.325 -31.115 -109.995 ;
        RECT -31.445 -111.685 -31.115 -111.355 ;
        RECT -31.445 -113.045 -31.115 -112.715 ;
        RECT -31.445 -114.405 -31.115 -114.075 ;
        RECT -31.445 -115.765 -31.115 -115.435 ;
        RECT -31.445 -117.125 -31.115 -116.795 ;
        RECT -31.445 -118.485 -31.115 -118.155 ;
        RECT -31.445 -119.845 -31.115 -119.515 ;
        RECT -31.445 -123.925 -31.115 -123.595 ;
        RECT -31.445 -129.365 -31.115 -129.035 ;
        RECT -31.445 -130.725 -31.115 -130.395 ;
        RECT -31.445 -132.085 -31.115 -131.755 ;
        RECT -31.445 -133.445 -31.115 -133.115 ;
        RECT -31.445 -134.805 -31.115 -134.475 ;
        RECT -31.445 -136.165 -31.115 -135.835 ;
        RECT -31.445 -137.525 -31.115 -137.195 ;
        RECT -31.445 -138.885 -31.115 -138.555 ;
        RECT -31.445 -140.245 -31.115 -139.915 ;
        RECT -31.445 -141.605 -31.115 -141.275 ;
        RECT -31.445 -142.965 -31.115 -142.635 ;
        RECT -31.445 -144.325 -31.115 -143.995 ;
        RECT -31.445 -145.685 -31.115 -145.355 ;
        RECT -31.445 -147.045 -31.115 -146.715 ;
        RECT -31.445 -148.405 -31.115 -148.075 ;
        RECT -31.445 -149.765 -31.115 -149.435 ;
        RECT -31.445 -151.125 -31.115 -150.795 ;
        RECT -31.445 -152.485 -31.115 -152.155 ;
        RECT -31.445 -153.845 -31.115 -153.515 ;
        RECT -31.445 -155.205 -31.115 -154.875 ;
        RECT -31.445 -156.565 -31.115 -156.235 ;
        RECT -31.445 -157.925 -31.115 -157.595 ;
        RECT -31.445 -159.285 -31.115 -158.955 ;
        RECT -31.445 -162.005 -31.115 -161.675 ;
        RECT -31.445 -163.365 -31.115 -163.035 ;
        RECT -31.445 -164.725 -31.115 -164.395 ;
        RECT -31.445 -166.085 -31.115 -165.755 ;
        RECT -31.445 -167.445 -31.115 -167.115 ;
        RECT -31.445 -168.805 -31.115 -168.475 ;
        RECT -31.445 -170.165 -31.115 -169.835 ;
        RECT -31.445 -171.525 -31.115 -171.195 ;
        RECT -31.445 -172.885 -31.115 -172.555 ;
        RECT -31.445 -174.245 -31.115 -173.915 ;
        RECT -31.445 -175.605 -31.115 -175.275 ;
        RECT -31.445 -176.965 -31.115 -176.635 ;
        RECT -31.445 -178.325 -31.115 -177.995 ;
        RECT -31.445 -179.685 -31.115 -179.355 ;
        RECT -31.445 -181.045 -31.115 -180.715 ;
        RECT -31.445 -182.405 -31.115 -182.075 ;
        RECT -31.445 -183.765 -31.115 -183.435 ;
        RECT -31.445 -185.125 -31.115 -184.795 ;
        RECT -31.445 -186.485 -31.115 -186.155 ;
        RECT -31.445 -190.565 -31.115 -190.235 ;
        RECT -31.445 -191.925 -31.115 -191.595 ;
        RECT -31.445 -193.285 -31.115 -192.955 ;
        RECT -31.445 -194.645 -31.115 -194.315 ;
        RECT -31.445 -196.005 -31.115 -195.675 ;
        RECT -31.445 -197.365 -31.115 -197.035 ;
        RECT -31.445 -198.725 -31.115 -198.395 ;
        RECT -31.445 -200.085 -31.115 -199.755 ;
        RECT -31.445 -201.445 -31.115 -201.115 ;
        RECT -31.445 -202.805 -31.115 -202.475 ;
        RECT -31.445 -204.165 -31.115 -203.835 ;
        RECT -31.445 -205.525 -31.115 -205.195 ;
        RECT -31.445 -208.245 -31.115 -207.915 ;
        RECT -31.445 -209.605 -31.115 -209.275 ;
        RECT -31.445 -213.685 -31.115 -213.355 ;
        RECT -31.445 -215.045 -31.115 -214.715 ;
        RECT -31.445 -216.405 -31.115 -216.075 ;
        RECT -31.445 -217.765 -31.115 -217.435 ;
        RECT -31.445 -219.125 -31.115 -218.795 ;
        RECT -31.445 -220.485 -31.115 -220.155 ;
        RECT -31.445 -221.845 -31.115 -221.515 ;
        RECT -31.445 -223.205 -31.115 -222.875 ;
        RECT -31.445 -224.565 -31.115 -224.235 ;
        RECT -31.445 -226.155 -31.115 -225.825 ;
        RECT -31.445 -227.285 -31.115 -226.955 ;
        RECT -31.445 -228.645 -31.115 -228.315 ;
        RECT -31.445 -230.005 -31.115 -229.675 ;
        RECT -31.445 -231.365 -31.115 -231.035 ;
        RECT -31.445 -234.085 -31.115 -233.755 ;
        RECT -31.445 -235.445 -31.115 -235.115 ;
        RECT -31.445 -236.805 -31.115 -236.475 ;
        RECT -31.445 -238.165 -31.115 -237.835 ;
        RECT -31.445 -243.81 -31.115 -242.68 ;
        RECT -31.44 -243.925 -31.12 248.005 ;
        RECT -31.445 246.76 -31.115 247.89 ;
        RECT -31.445 241.915 -31.115 242.245 ;
        RECT -31.445 240.555 -31.115 240.885 ;
        RECT -31.445 239.195 -31.115 239.525 ;
        RECT -31.445 237.835 -31.115 238.165 ;
        RECT -31.445 236.475 -31.115 236.805 ;
        RECT -31.445 235.115 -31.115 235.445 ;
        RECT -31.445 233.755 -31.115 234.085 ;
        RECT -31.445 232.395 -31.115 232.725 ;
        RECT -31.445 231.035 -31.115 231.365 ;
        RECT -31.445 229.675 -31.115 230.005 ;
        RECT -31.445 228.315 -31.115 228.645 ;
        RECT -31.445 226.955 -31.115 227.285 ;
        RECT -31.445 225.595 -31.115 225.925 ;
        RECT -31.445 224.235 -31.115 224.565 ;
        RECT -31.445 222.875 -31.115 223.205 ;
        RECT -31.445 221.515 -31.115 221.845 ;
        RECT -31.445 220.155 -31.115 220.485 ;
        RECT -31.445 218.795 -31.115 219.125 ;
        RECT -31.445 217.435 -31.115 217.765 ;
        RECT -31.445 216.075 -31.115 216.405 ;
        RECT -31.445 214.715 -31.115 215.045 ;
        RECT -31.445 213.355 -31.115 213.685 ;
        RECT -31.445 211.995 -31.115 212.325 ;
        RECT -31.445 210.635 -31.115 210.965 ;
        RECT -31.445 209.275 -31.115 209.605 ;
        RECT -31.445 207.915 -31.115 208.245 ;
        RECT -31.445 206.555 -31.115 206.885 ;
        RECT -31.445 205.195 -31.115 205.525 ;
        RECT -31.445 203.835 -31.115 204.165 ;
        RECT -31.445 202.475 -31.115 202.805 ;
        RECT -31.445 201.115 -31.115 201.445 ;
        RECT -31.445 199.755 -31.115 200.085 ;
        RECT -31.445 198.395 -31.115 198.725 ;
        RECT -31.445 197.035 -31.115 197.365 ;
        RECT -31.445 195.675 -31.115 196.005 ;
        RECT -31.445 194.315 -31.115 194.645 ;
        RECT -31.445 192.955 -31.115 193.285 ;
        RECT -31.445 191.595 -31.115 191.925 ;
        RECT -31.445 190.235 -31.115 190.565 ;
        RECT -31.445 188.875 -31.115 189.205 ;
        RECT -31.445 187.515 -31.115 187.845 ;
        RECT -31.445 186.155 -31.115 186.485 ;
        RECT -31.445 184.795 -31.115 185.125 ;
        RECT -31.445 183.435 -31.115 183.765 ;
        RECT -31.445 182.075 -31.115 182.405 ;
        RECT -31.445 180.715 -31.115 181.045 ;
        RECT -31.445 179.355 -31.115 179.685 ;
        RECT -31.445 177.995 -31.115 178.325 ;
        RECT -31.445 176.635 -31.115 176.965 ;
        RECT -31.445 175.275 -31.115 175.605 ;
        RECT -31.445 173.915 -31.115 174.245 ;
        RECT -31.445 172.555 -31.115 172.885 ;
        RECT -31.445 171.195 -31.115 171.525 ;
        RECT -31.445 169.835 -31.115 170.165 ;
        RECT -31.445 168.475 -31.115 168.805 ;
        RECT -31.445 167.115 -31.115 167.445 ;
        RECT -31.445 165.755 -31.115 166.085 ;
        RECT -31.445 164.395 -31.115 164.725 ;
        RECT -31.445 163.035 -31.115 163.365 ;
        RECT -31.445 161.675 -31.115 162.005 ;
        RECT -31.445 160.315 -31.115 160.645 ;
        RECT -31.445 158.955 -31.115 159.285 ;
        RECT -31.445 157.595 -31.115 157.925 ;
        RECT -31.445 156.235 -31.115 156.565 ;
        RECT -31.445 154.875 -31.115 155.205 ;
        RECT -31.445 153.515 -31.115 153.845 ;
        RECT -31.445 152.155 -31.115 152.485 ;
        RECT -31.445 150.795 -31.115 151.125 ;
        RECT -31.445 149.435 -31.115 149.765 ;
        RECT -31.445 148.075 -31.115 148.405 ;
        RECT -31.445 146.715 -31.115 147.045 ;
        RECT -31.445 145.355 -31.115 145.685 ;
        RECT -31.445 143.995 -31.115 144.325 ;
        RECT -31.445 142.635 -31.115 142.965 ;
        RECT -31.445 141.275 -31.115 141.605 ;
        RECT -31.445 139.915 -31.115 140.245 ;
        RECT -31.445 138.555 -31.115 138.885 ;
        RECT -31.445 137.195 -31.115 137.525 ;
        RECT -31.445 135.835 -31.115 136.165 ;
        RECT -31.445 134.475 -31.115 134.805 ;
        RECT -31.445 133.115 -31.115 133.445 ;
        RECT -31.445 131.755 -31.115 132.085 ;
        RECT -31.445 130.395 -31.115 130.725 ;
        RECT -31.445 129.035 -31.115 129.365 ;
        RECT -31.445 127.675 -31.115 128.005 ;
        RECT -31.445 126.315 -31.115 126.645 ;
        RECT -31.445 124.955 -31.115 125.285 ;
        RECT -31.445 123.595 -31.115 123.925 ;
        RECT -31.445 122.235 -31.115 122.565 ;
        RECT -31.445 120.875 -31.115 121.205 ;
        RECT -31.445 119.515 -31.115 119.845 ;
        RECT -31.445 118.155 -31.115 118.485 ;
        RECT -31.445 116.795 -31.115 117.125 ;
        RECT -31.445 115.435 -31.115 115.765 ;
        RECT -31.445 114.075 -31.115 114.405 ;
        RECT -31.445 112.715 -31.115 113.045 ;
        RECT -31.445 111.355 -31.115 111.685 ;
        RECT -31.445 109.995 -31.115 110.325 ;
        RECT -31.445 108.635 -31.115 108.965 ;
        RECT -31.445 107.275 -31.115 107.605 ;
        RECT -31.445 105.915 -31.115 106.245 ;
        RECT -31.445 104.555 -31.115 104.885 ;
        RECT -31.445 103.195 -31.115 103.525 ;
        RECT -31.445 101.835 -31.115 102.165 ;
        RECT -31.445 100.475 -31.115 100.805 ;
        RECT -31.445 99.115 -31.115 99.445 ;
        RECT -31.445 97.755 -31.115 98.085 ;
        RECT -31.445 96.395 -31.115 96.725 ;
        RECT -31.445 95.035 -31.115 95.365 ;
        RECT -31.445 93.675 -31.115 94.005 ;
        RECT -31.445 92.315 -31.115 92.645 ;
        RECT -31.445 90.955 -31.115 91.285 ;
        RECT -31.445 89.595 -31.115 89.925 ;
        RECT -31.445 88.235 -31.115 88.565 ;
        RECT -31.445 86.875 -31.115 87.205 ;
        RECT -31.445 85.515 -31.115 85.845 ;
        RECT -31.445 84.155 -31.115 84.485 ;
        RECT -31.445 82.795 -31.115 83.125 ;
        RECT -31.445 81.435 -31.115 81.765 ;
        RECT -31.445 80.075 -31.115 80.405 ;
        RECT -31.445 78.715 -31.115 79.045 ;
        RECT -31.445 77.355 -31.115 77.685 ;
        RECT -31.445 75.995 -31.115 76.325 ;
        RECT -31.445 74.635 -31.115 74.965 ;
        RECT -31.445 73.275 -31.115 73.605 ;
        RECT -31.445 71.915 -31.115 72.245 ;
        RECT -31.445 70.555 -31.115 70.885 ;
        RECT -31.445 69.195 -31.115 69.525 ;
        RECT -31.445 67.835 -31.115 68.165 ;
        RECT -31.445 66.475 -31.115 66.805 ;
        RECT -31.445 65.115 -31.115 65.445 ;
        RECT -31.445 63.755 -31.115 64.085 ;
        RECT -31.445 62.395 -31.115 62.725 ;
        RECT -31.445 61.035 -31.115 61.365 ;
        RECT -31.445 59.675 -31.115 60.005 ;
        RECT -31.445 58.315 -31.115 58.645 ;
        RECT -31.445 56.955 -31.115 57.285 ;
        RECT -31.445 55.595 -31.115 55.925 ;
        RECT -31.445 54.235 -31.115 54.565 ;
        RECT -31.445 52.875 -31.115 53.205 ;
        RECT -31.445 51.515 -31.115 51.845 ;
        RECT -31.445 50.155 -31.115 50.485 ;
        RECT -31.445 48.795 -31.115 49.125 ;
        RECT -31.445 47.435 -31.115 47.765 ;
        RECT -31.445 46.075 -31.115 46.405 ;
        RECT -31.445 44.715 -31.115 45.045 ;
        RECT -31.445 43.355 -31.115 43.685 ;
        RECT -31.445 41.995 -31.115 42.325 ;
        RECT -31.445 40.635 -31.115 40.965 ;
        RECT -31.445 39.275 -31.115 39.605 ;
        RECT -31.445 37.915 -31.115 38.245 ;
        RECT -31.445 36.555 -31.115 36.885 ;
        RECT -31.445 35.195 -31.115 35.525 ;
        RECT -31.445 33.835 -31.115 34.165 ;
        RECT -31.445 32.475 -31.115 32.805 ;
        RECT -31.445 31.115 -31.115 31.445 ;
        RECT -31.445 29.755 -31.115 30.085 ;
        RECT -31.445 28.395 -31.115 28.725 ;
        RECT -31.445 27.035 -31.115 27.365 ;
        RECT -31.445 25.675 -31.115 26.005 ;
        RECT -31.445 24.315 -31.115 24.645 ;
        RECT -31.445 22.955 -31.115 23.285 ;
        RECT -31.445 21.595 -31.115 21.925 ;
        RECT -31.445 20.235 -31.115 20.565 ;
        RECT -31.445 18.875 -31.115 19.205 ;
        RECT -31.445 17.515 -31.115 17.845 ;
        RECT -31.445 16.155 -31.115 16.485 ;
        RECT -31.445 14.795 -31.115 15.125 ;
        RECT -31.445 13.435 -31.115 13.765 ;
        RECT -31.445 12.075 -31.115 12.405 ;
        RECT -31.445 10.715 -31.115 11.045 ;
        RECT -31.445 9.355 -31.115 9.685 ;
        RECT -31.445 7.995 -31.115 8.325 ;
        RECT -31.445 6.635 -31.115 6.965 ;
        RECT -31.445 5.275 -31.115 5.605 ;
        RECT -31.445 3.915 -31.115 4.245 ;
        RECT -31.445 2.555 -31.115 2.885 ;
        RECT -31.445 1.195 -31.115 1.525 ;
        RECT -31.445 -0.165 -31.115 0.165 ;
        RECT -31.445 -2.885 -31.115 -2.555 ;
        RECT -31.445 -6.965 -31.115 -6.635 ;
        RECT -31.445 -8.325 -31.115 -7.995 ;
        RECT -31.445 -9.685 -31.115 -9.355 ;
        RECT -31.445 -12.405 -31.115 -12.075 ;
        RECT -31.445 -13.765 -31.115 -13.435 ;
        RECT -31.445 -15.125 -31.115 -14.795 ;
        RECT -31.445 -16.485 -31.115 -16.155 ;
        RECT -31.445 -17.845 -31.115 -17.515 ;
        RECT -31.445 -19.205 -31.115 -18.875 ;
        RECT -31.445 -20.565 -31.115 -20.235 ;
        RECT -31.445 -21.925 -31.115 -21.595 ;
        RECT -31.445 -23.285 -31.115 -22.955 ;
        RECT -31.445 -30.66 -31.115 -30.33 ;
        RECT -31.445 -31.445 -31.115 -31.115 ;
        RECT -31.445 -32.805 -31.115 -32.475 ;
        RECT -31.445 -34.165 -31.115 -33.835 ;
        RECT -31.445 -36.885 -31.115 -36.555 ;
        RECT -31.445 -37.85 -31.115 -37.52 ;
        RECT -31.445 -40.965 -31.115 -40.635 ;
        RECT -31.445 -46.405 -31.115 -46.075 ;
        RECT -31.445 -49.125 -31.115 -48.795 ;
        RECT -31.445 -50.485 -31.115 -50.155 ;
        RECT -31.445 -53.205 -31.115 -52.875 ;
        RECT -31.445 -55.925 -31.115 -55.595 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.245 246.76 -37.915 247.89 ;
        RECT -38.245 241.915 -37.915 242.245 ;
        RECT -38.245 240.555 -37.915 240.885 ;
        RECT -38.245 239.195 -37.915 239.525 ;
        RECT -38.245 237.835 -37.915 238.165 ;
        RECT -38.245 236.475 -37.915 236.805 ;
        RECT -38.245 235.115 -37.915 235.445 ;
        RECT -38.245 233.755 -37.915 234.085 ;
        RECT -38.245 232.395 -37.915 232.725 ;
        RECT -38.245 231.035 -37.915 231.365 ;
        RECT -38.245 229.675 -37.915 230.005 ;
        RECT -38.245 228.315 -37.915 228.645 ;
        RECT -38.245 226.955 -37.915 227.285 ;
        RECT -38.245 225.595 -37.915 225.925 ;
        RECT -38.245 224.235 -37.915 224.565 ;
        RECT -38.245 222.875 -37.915 223.205 ;
        RECT -38.245 221.515 -37.915 221.845 ;
        RECT -38.245 220.155 -37.915 220.485 ;
        RECT -38.245 218.795 -37.915 219.125 ;
        RECT -38.245 217.435 -37.915 217.765 ;
        RECT -38.245 216.075 -37.915 216.405 ;
        RECT -38.245 214.715 -37.915 215.045 ;
        RECT -38.245 213.355 -37.915 213.685 ;
        RECT -38.245 211.995 -37.915 212.325 ;
        RECT -38.245 210.635 -37.915 210.965 ;
        RECT -38.245 209.275 -37.915 209.605 ;
        RECT -38.245 207.915 -37.915 208.245 ;
        RECT -38.245 206.555 -37.915 206.885 ;
        RECT -38.245 205.195 -37.915 205.525 ;
        RECT -38.245 203.835 -37.915 204.165 ;
        RECT -38.245 202.475 -37.915 202.805 ;
        RECT -38.245 201.115 -37.915 201.445 ;
        RECT -38.245 199.755 -37.915 200.085 ;
        RECT -38.245 198.395 -37.915 198.725 ;
        RECT -38.245 197.035 -37.915 197.365 ;
        RECT -38.245 195.675 -37.915 196.005 ;
        RECT -38.245 194.315 -37.915 194.645 ;
        RECT -38.245 192.955 -37.915 193.285 ;
        RECT -38.245 191.595 -37.915 191.925 ;
        RECT -38.245 190.235 -37.915 190.565 ;
        RECT -38.245 188.875 -37.915 189.205 ;
        RECT -38.245 187.515 -37.915 187.845 ;
        RECT -38.245 186.155 -37.915 186.485 ;
        RECT -38.245 184.795 -37.915 185.125 ;
        RECT -38.245 183.435 -37.915 183.765 ;
        RECT -38.245 182.075 -37.915 182.405 ;
        RECT -38.245 180.715 -37.915 181.045 ;
        RECT -38.245 179.355 -37.915 179.685 ;
        RECT -38.245 177.995 -37.915 178.325 ;
        RECT -38.245 176.635 -37.915 176.965 ;
        RECT -38.245 175.275 -37.915 175.605 ;
        RECT -38.245 173.915 -37.915 174.245 ;
        RECT -38.245 172.555 -37.915 172.885 ;
        RECT -38.245 171.195 -37.915 171.525 ;
        RECT -38.245 169.835 -37.915 170.165 ;
        RECT -38.245 168.475 -37.915 168.805 ;
        RECT -38.245 167.115 -37.915 167.445 ;
        RECT -38.245 165.755 -37.915 166.085 ;
        RECT -38.245 164.395 -37.915 164.725 ;
        RECT -38.245 163.035 -37.915 163.365 ;
        RECT -38.245 161.675 -37.915 162.005 ;
        RECT -38.245 160.315 -37.915 160.645 ;
        RECT -38.245 158.955 -37.915 159.285 ;
        RECT -38.245 157.595 -37.915 157.925 ;
        RECT -38.245 156.235 -37.915 156.565 ;
        RECT -38.245 154.875 -37.915 155.205 ;
        RECT -38.245 153.515 -37.915 153.845 ;
        RECT -38.245 152.155 -37.915 152.485 ;
        RECT -38.245 150.795 -37.915 151.125 ;
        RECT -38.245 149.435 -37.915 149.765 ;
        RECT -38.245 148.075 -37.915 148.405 ;
        RECT -38.245 146.715 -37.915 147.045 ;
        RECT -38.245 145.355 -37.915 145.685 ;
        RECT -38.245 143.995 -37.915 144.325 ;
        RECT -38.245 142.635 -37.915 142.965 ;
        RECT -38.245 141.275 -37.915 141.605 ;
        RECT -38.245 139.915 -37.915 140.245 ;
        RECT -38.245 138.555 -37.915 138.885 ;
        RECT -38.245 137.195 -37.915 137.525 ;
        RECT -38.245 135.835 -37.915 136.165 ;
        RECT -38.245 134.475 -37.915 134.805 ;
        RECT -38.245 133.115 -37.915 133.445 ;
        RECT -38.245 131.755 -37.915 132.085 ;
        RECT -38.245 130.395 -37.915 130.725 ;
        RECT -38.245 129.035 -37.915 129.365 ;
        RECT -38.245 127.675 -37.915 128.005 ;
        RECT -38.245 126.315 -37.915 126.645 ;
        RECT -38.245 124.955 -37.915 125.285 ;
        RECT -38.245 123.595 -37.915 123.925 ;
        RECT -38.245 122.235 -37.915 122.565 ;
        RECT -38.245 120.875 -37.915 121.205 ;
        RECT -38.245 119.515 -37.915 119.845 ;
        RECT -38.245 118.155 -37.915 118.485 ;
        RECT -38.245 116.795 -37.915 117.125 ;
        RECT -38.245 115.435 -37.915 115.765 ;
        RECT -38.245 114.075 -37.915 114.405 ;
        RECT -38.245 112.715 -37.915 113.045 ;
        RECT -38.245 111.355 -37.915 111.685 ;
        RECT -38.245 109.995 -37.915 110.325 ;
        RECT -38.245 108.635 -37.915 108.965 ;
        RECT -38.245 107.275 -37.915 107.605 ;
        RECT -38.245 105.915 -37.915 106.245 ;
        RECT -38.245 104.555 -37.915 104.885 ;
        RECT -38.245 103.195 -37.915 103.525 ;
        RECT -38.245 101.835 -37.915 102.165 ;
        RECT -38.245 100.475 -37.915 100.805 ;
        RECT -38.245 99.115 -37.915 99.445 ;
        RECT -38.245 97.755 -37.915 98.085 ;
        RECT -38.245 96.395 -37.915 96.725 ;
        RECT -38.245 95.035 -37.915 95.365 ;
        RECT -38.245 93.675 -37.915 94.005 ;
        RECT -38.245 92.315 -37.915 92.645 ;
        RECT -38.245 90.955 -37.915 91.285 ;
        RECT -38.245 89.595 -37.915 89.925 ;
        RECT -38.245 88.235 -37.915 88.565 ;
        RECT -38.245 86.875 -37.915 87.205 ;
        RECT -38.245 85.515 -37.915 85.845 ;
        RECT -38.245 84.155 -37.915 84.485 ;
        RECT -38.245 82.795 -37.915 83.125 ;
        RECT -38.245 81.435 -37.915 81.765 ;
        RECT -38.245 80.075 -37.915 80.405 ;
        RECT -38.245 78.715 -37.915 79.045 ;
        RECT -38.245 77.355 -37.915 77.685 ;
        RECT -38.245 75.995 -37.915 76.325 ;
        RECT -38.245 74.635 -37.915 74.965 ;
        RECT -38.245 73.275 -37.915 73.605 ;
        RECT -38.245 71.915 -37.915 72.245 ;
        RECT -38.245 70.555 -37.915 70.885 ;
        RECT -38.245 69.195 -37.915 69.525 ;
        RECT -38.245 67.835 -37.915 68.165 ;
        RECT -38.245 66.475 -37.915 66.805 ;
        RECT -38.245 65.115 -37.915 65.445 ;
        RECT -38.245 63.755 -37.915 64.085 ;
        RECT -38.245 62.395 -37.915 62.725 ;
        RECT -38.245 61.035 -37.915 61.365 ;
        RECT -38.245 59.675 -37.915 60.005 ;
        RECT -38.245 58.315 -37.915 58.645 ;
        RECT -38.245 56.955 -37.915 57.285 ;
        RECT -38.245 55.595 -37.915 55.925 ;
        RECT -38.245 54.235 -37.915 54.565 ;
        RECT -38.245 52.875 -37.915 53.205 ;
        RECT -38.245 51.515 -37.915 51.845 ;
        RECT -38.245 50.155 -37.915 50.485 ;
        RECT -38.245 48.795 -37.915 49.125 ;
        RECT -38.245 47.435 -37.915 47.765 ;
        RECT -38.245 46.075 -37.915 46.405 ;
        RECT -38.245 44.715 -37.915 45.045 ;
        RECT -38.245 43.355 -37.915 43.685 ;
        RECT -38.245 41.995 -37.915 42.325 ;
        RECT -38.245 40.635 -37.915 40.965 ;
        RECT -38.245 39.275 -37.915 39.605 ;
        RECT -38.245 37.915 -37.915 38.245 ;
        RECT -38.245 36.555 -37.915 36.885 ;
        RECT -38.245 35.195 -37.915 35.525 ;
        RECT -38.245 33.835 -37.915 34.165 ;
        RECT -38.245 32.475 -37.915 32.805 ;
        RECT -38.245 31.115 -37.915 31.445 ;
        RECT -38.245 29.755 -37.915 30.085 ;
        RECT -38.245 28.395 -37.915 28.725 ;
        RECT -38.245 27.035 -37.915 27.365 ;
        RECT -38.245 25.675 -37.915 26.005 ;
        RECT -38.245 24.315 -37.915 24.645 ;
        RECT -38.245 22.955 -37.915 23.285 ;
        RECT -38.245 21.595 -37.915 21.925 ;
        RECT -38.245 20.235 -37.915 20.565 ;
        RECT -38.245 18.875 -37.915 19.205 ;
        RECT -38.245 17.515 -37.915 17.845 ;
        RECT -38.245 16.155 -37.915 16.485 ;
        RECT -38.245 14.795 -37.915 15.125 ;
        RECT -38.245 13.435 -37.915 13.765 ;
        RECT -38.245 12.075 -37.915 12.405 ;
        RECT -38.245 10.715 -37.915 11.045 ;
        RECT -38.245 9.355 -37.915 9.685 ;
        RECT -38.245 7.995 -37.915 8.325 ;
        RECT -38.245 6.635 -37.915 6.965 ;
        RECT -38.245 5.275 -37.915 5.605 ;
        RECT -38.245 3.915 -37.915 4.245 ;
        RECT -38.245 2.555 -37.915 2.885 ;
        RECT -38.245 1.195 -37.915 1.525 ;
        RECT -38.245 -0.165 -37.915 0.165 ;
        RECT -38.245 -1.525 -37.915 -1.195 ;
        RECT -38.245 -4.245 -37.915 -3.915 ;
        RECT -38.245 -8.325 -37.915 -7.995 ;
        RECT -38.245 -9.685 -37.915 -9.355 ;
        RECT -38.245 -12.405 -37.915 -12.075 ;
        RECT -38.245 -13.765 -37.915 -13.435 ;
        RECT -38.245 -15.125 -37.915 -14.795 ;
        RECT -38.245 -16.485 -37.915 -16.155 ;
        RECT -38.245 -17.845 -37.915 -17.515 ;
        RECT -38.245 -19.205 -37.915 -18.875 ;
        RECT -38.245 -20.565 -37.915 -20.235 ;
        RECT -38.245 -21.925 -37.915 -21.595 ;
        RECT -38.245 -23.285 -37.915 -22.955 ;
        RECT -38.245 -30.66 -37.915 -30.33 ;
        RECT -38.245 -31.445 -37.915 -31.115 ;
        RECT -38.245 -32.805 -37.915 -32.475 ;
        RECT -38.245 -34.165 -37.915 -33.835 ;
        RECT -38.245 -36.885 -37.915 -36.555 ;
        RECT -38.245 -37.85 -37.915 -37.52 ;
        RECT -38.245 -40.965 -37.915 -40.635 ;
        RECT -38.245 -46.405 -37.915 -46.075 ;
        RECT -38.245 -47.765 -37.915 -47.435 ;
        RECT -38.245 -49.125 -37.915 -48.795 ;
        RECT -38.245 -50.485 -37.915 -50.155 ;
        RECT -38.245 -51.845 -37.915 -51.515 ;
        RECT -38.245 -53.205 -37.915 -52.875 ;
        RECT -38.245 -54.565 -37.915 -54.235 ;
        RECT -38.245 -55.925 -37.915 -55.595 ;
        RECT -38.245 -57.285 -37.915 -56.955 ;
        RECT -38.245 -58.645 -37.915 -58.315 ;
        RECT -38.245 -60.005 -37.915 -59.675 ;
        RECT -38.245 -61.365 -37.915 -61.035 ;
        RECT -38.245 -62.725 -37.915 -62.395 ;
        RECT -38.245 -64.085 -37.915 -63.755 ;
        RECT -38.245 -65.445 -37.915 -65.115 ;
        RECT -38.245 -66.805 -37.915 -66.475 ;
        RECT -38.245 -68.165 -37.915 -67.835 ;
        RECT -38.245 -69.525 -37.915 -69.195 ;
        RECT -38.245 -70.885 -37.915 -70.555 ;
        RECT -38.245 -72.245 -37.915 -71.915 ;
        RECT -38.245 -73.605 -37.915 -73.275 ;
        RECT -38.245 -74.965 -37.915 -74.635 ;
        RECT -38.245 -76.325 -37.915 -75.995 ;
        RECT -38.245 -77.685 -37.915 -77.355 ;
        RECT -38.245 -79.045 -37.915 -78.715 ;
        RECT -38.245 -80.405 -37.915 -80.075 ;
        RECT -38.245 -81.765 -37.915 -81.435 ;
        RECT -38.245 -83.125 -37.915 -82.795 ;
        RECT -38.245 -84.485 -37.915 -84.155 ;
        RECT -38.245 -85.845 -37.915 -85.515 ;
        RECT -38.245 -87.205 -37.915 -86.875 ;
        RECT -38.245 -88.565 -37.915 -88.235 ;
        RECT -38.245 -89.925 -37.915 -89.595 ;
        RECT -38.245 -91.285 -37.915 -90.955 ;
        RECT -38.245 -92.645 -37.915 -92.315 ;
        RECT -38.245 -94.005 -37.915 -93.675 ;
        RECT -38.245 -95.365 -37.915 -95.035 ;
        RECT -38.245 -96.725 -37.915 -96.395 ;
        RECT -38.245 -98.085 -37.915 -97.755 ;
        RECT -38.245 -99.445 -37.915 -99.115 ;
        RECT -38.245 -100.805 -37.915 -100.475 ;
        RECT -38.245 -102.165 -37.915 -101.835 ;
        RECT -38.245 -103.525 -37.915 -103.195 ;
        RECT -38.245 -104.885 -37.915 -104.555 ;
        RECT -38.245 -106.245 -37.915 -105.915 ;
        RECT -38.245 -107.605 -37.915 -107.275 ;
        RECT -38.245 -108.965 -37.915 -108.635 ;
        RECT -38.245 -110.325 -37.915 -109.995 ;
        RECT -38.245 -111.685 -37.915 -111.355 ;
        RECT -38.245 -113.045 -37.915 -112.715 ;
        RECT -38.245 -114.405 -37.915 -114.075 ;
        RECT -38.245 -115.765 -37.915 -115.435 ;
        RECT -38.245 -117.125 -37.915 -116.795 ;
        RECT -38.245 -118.485 -37.915 -118.155 ;
        RECT -38.245 -119.845 -37.915 -119.515 ;
        RECT -38.245 -123.925 -37.915 -123.595 ;
        RECT -38.245 -129.365 -37.915 -129.035 ;
        RECT -38.245 -130.725 -37.915 -130.395 ;
        RECT -38.245 -131.47 -37.915 -131.14 ;
        RECT -38.245 -133.445 -37.915 -133.115 ;
        RECT -38.245 -134.805 -37.915 -134.475 ;
        RECT -38.245 -136.165 -37.915 -135.835 ;
        RECT -38.245 -137.525 -37.915 -137.195 ;
        RECT -38.245 -140.245 -37.915 -139.915 ;
        RECT -38.245 -141.605 -37.915 -141.275 ;
        RECT -38.245 -142.965 -37.915 -142.635 ;
        RECT -38.245 -144.31 -37.915 -143.98 ;
        RECT -38.245 -145.685 -37.915 -145.355 ;
        RECT -38.245 -147.045 -37.915 -146.715 ;
        RECT -38.245 -149.765 -37.915 -149.435 ;
        RECT -38.245 -153.845 -37.915 -153.515 ;
        RECT -38.245 -155.205 -37.915 -154.875 ;
        RECT -38.245 -156.565 -37.915 -156.235 ;
        RECT -38.245 -157.925 -37.915 -157.595 ;
        RECT -38.245 -159.285 -37.915 -158.955 ;
        RECT -38.245 -162.005 -37.915 -161.675 ;
        RECT -38.245 -163.365 -37.915 -163.035 ;
        RECT -38.245 -164.725 -37.915 -164.395 ;
        RECT -38.245 -166.085 -37.915 -165.755 ;
        RECT -38.245 -167.445 -37.915 -167.115 ;
        RECT -38.245 -168.805 -37.915 -168.475 ;
        RECT -38.245 -170.165 -37.915 -169.835 ;
        RECT -38.245 -171.525 -37.915 -171.195 ;
        RECT -38.245 -172.885 -37.915 -172.555 ;
        RECT -38.245 -174.245 -37.915 -173.915 ;
        RECT -38.245 -175.605 -37.915 -175.275 ;
        RECT -38.245 -176.965 -37.915 -176.635 ;
        RECT -38.245 -178.325 -37.915 -177.995 ;
        RECT -38.245 -179.685 -37.915 -179.355 ;
        RECT -38.245 -181.045 -37.915 -180.715 ;
        RECT -38.245 -182.405 -37.915 -182.075 ;
        RECT -38.245 -183.765 -37.915 -183.435 ;
        RECT -38.245 -185.125 -37.915 -184.795 ;
        RECT -38.245 -186.485 -37.915 -186.155 ;
        RECT -38.245 -187.845 -37.915 -187.515 ;
        RECT -38.245 -189.205 -37.915 -188.875 ;
        RECT -38.245 -190.565 -37.915 -190.235 ;
        RECT -38.245 -191.925 -37.915 -191.595 ;
        RECT -38.245 -193.285 -37.915 -192.955 ;
        RECT -38.245 -194.645 -37.915 -194.315 ;
        RECT -38.245 -196.005 -37.915 -195.675 ;
        RECT -38.245 -197.365 -37.915 -197.035 ;
        RECT -38.245 -198.725 -37.915 -198.395 ;
        RECT -38.245 -200.085 -37.915 -199.755 ;
        RECT -38.245 -201.445 -37.915 -201.115 ;
        RECT -38.245 -202.805 -37.915 -202.475 ;
        RECT -38.245 -204.165 -37.915 -203.835 ;
        RECT -38.245 -205.525 -37.915 -205.195 ;
        RECT -38.245 -206.885 -37.915 -206.555 ;
        RECT -38.245 -208.245 -37.915 -207.915 ;
        RECT -38.245 -209.605 -37.915 -209.275 ;
        RECT -38.245 -210.965 -37.915 -210.635 ;
        RECT -38.245 -212.325 -37.915 -211.995 ;
        RECT -38.245 -213.685 -37.915 -213.355 ;
        RECT -38.245 -215.045 -37.915 -214.715 ;
        RECT -38.245 -216.405 -37.915 -216.075 ;
        RECT -38.245 -217.765 -37.915 -217.435 ;
        RECT -38.245 -219.125 -37.915 -218.795 ;
        RECT -38.245 -220.485 -37.915 -220.155 ;
        RECT -38.245 -221.845 -37.915 -221.515 ;
        RECT -38.245 -223.205 -37.915 -222.875 ;
        RECT -38.245 -224.565 -37.915 -224.235 ;
        RECT -38.245 -226.155 -37.915 -225.825 ;
        RECT -38.245 -227.285 -37.915 -226.955 ;
        RECT -38.245 -228.645 -37.915 -228.315 ;
        RECT -38.245 -230.005 -37.915 -229.675 ;
        RECT -38.245 -234.085 -37.915 -233.755 ;
        RECT -38.245 -235.445 -37.915 -235.115 ;
        RECT -38.245 -236.805 -37.915 -236.475 ;
        RECT -38.245 -238.165 -37.915 -237.835 ;
        RECT -38.245 -243.81 -37.915 -242.68 ;
        RECT -38.24 -243.925 -37.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.885 246.76 -36.555 247.89 ;
        RECT -36.885 241.915 -36.555 242.245 ;
        RECT -36.885 240.555 -36.555 240.885 ;
        RECT -36.885 239.195 -36.555 239.525 ;
        RECT -36.885 237.835 -36.555 238.165 ;
        RECT -36.885 236.475 -36.555 236.805 ;
        RECT -36.885 235.115 -36.555 235.445 ;
        RECT -36.885 233.755 -36.555 234.085 ;
        RECT -36.885 232.395 -36.555 232.725 ;
        RECT -36.885 231.035 -36.555 231.365 ;
        RECT -36.885 229.675 -36.555 230.005 ;
        RECT -36.885 228.315 -36.555 228.645 ;
        RECT -36.885 226.955 -36.555 227.285 ;
        RECT -36.885 225.595 -36.555 225.925 ;
        RECT -36.885 224.235 -36.555 224.565 ;
        RECT -36.885 222.875 -36.555 223.205 ;
        RECT -36.885 221.515 -36.555 221.845 ;
        RECT -36.885 220.155 -36.555 220.485 ;
        RECT -36.885 218.795 -36.555 219.125 ;
        RECT -36.885 217.435 -36.555 217.765 ;
        RECT -36.885 216.075 -36.555 216.405 ;
        RECT -36.885 214.715 -36.555 215.045 ;
        RECT -36.885 213.355 -36.555 213.685 ;
        RECT -36.885 211.995 -36.555 212.325 ;
        RECT -36.885 210.635 -36.555 210.965 ;
        RECT -36.885 209.275 -36.555 209.605 ;
        RECT -36.885 207.915 -36.555 208.245 ;
        RECT -36.885 206.555 -36.555 206.885 ;
        RECT -36.885 205.195 -36.555 205.525 ;
        RECT -36.885 203.835 -36.555 204.165 ;
        RECT -36.885 202.475 -36.555 202.805 ;
        RECT -36.885 201.115 -36.555 201.445 ;
        RECT -36.885 199.755 -36.555 200.085 ;
        RECT -36.885 198.395 -36.555 198.725 ;
        RECT -36.885 197.035 -36.555 197.365 ;
        RECT -36.885 195.675 -36.555 196.005 ;
        RECT -36.885 194.315 -36.555 194.645 ;
        RECT -36.885 192.955 -36.555 193.285 ;
        RECT -36.885 191.595 -36.555 191.925 ;
        RECT -36.885 190.235 -36.555 190.565 ;
        RECT -36.885 188.875 -36.555 189.205 ;
        RECT -36.885 187.515 -36.555 187.845 ;
        RECT -36.885 186.155 -36.555 186.485 ;
        RECT -36.885 184.795 -36.555 185.125 ;
        RECT -36.885 183.435 -36.555 183.765 ;
        RECT -36.885 182.075 -36.555 182.405 ;
        RECT -36.885 180.715 -36.555 181.045 ;
        RECT -36.885 179.355 -36.555 179.685 ;
        RECT -36.885 177.995 -36.555 178.325 ;
        RECT -36.885 176.635 -36.555 176.965 ;
        RECT -36.885 175.275 -36.555 175.605 ;
        RECT -36.885 173.915 -36.555 174.245 ;
        RECT -36.885 172.555 -36.555 172.885 ;
        RECT -36.885 171.195 -36.555 171.525 ;
        RECT -36.885 169.835 -36.555 170.165 ;
        RECT -36.885 168.475 -36.555 168.805 ;
        RECT -36.885 167.115 -36.555 167.445 ;
        RECT -36.885 165.755 -36.555 166.085 ;
        RECT -36.885 164.395 -36.555 164.725 ;
        RECT -36.885 163.035 -36.555 163.365 ;
        RECT -36.885 161.675 -36.555 162.005 ;
        RECT -36.885 160.315 -36.555 160.645 ;
        RECT -36.885 158.955 -36.555 159.285 ;
        RECT -36.885 157.595 -36.555 157.925 ;
        RECT -36.885 156.235 -36.555 156.565 ;
        RECT -36.885 154.875 -36.555 155.205 ;
        RECT -36.885 153.515 -36.555 153.845 ;
        RECT -36.885 152.155 -36.555 152.485 ;
        RECT -36.885 150.795 -36.555 151.125 ;
        RECT -36.885 149.435 -36.555 149.765 ;
        RECT -36.885 148.075 -36.555 148.405 ;
        RECT -36.885 146.715 -36.555 147.045 ;
        RECT -36.885 145.355 -36.555 145.685 ;
        RECT -36.885 143.995 -36.555 144.325 ;
        RECT -36.885 142.635 -36.555 142.965 ;
        RECT -36.885 141.275 -36.555 141.605 ;
        RECT -36.885 139.915 -36.555 140.245 ;
        RECT -36.885 138.555 -36.555 138.885 ;
        RECT -36.885 137.195 -36.555 137.525 ;
        RECT -36.885 135.835 -36.555 136.165 ;
        RECT -36.885 134.475 -36.555 134.805 ;
        RECT -36.885 133.115 -36.555 133.445 ;
        RECT -36.885 131.755 -36.555 132.085 ;
        RECT -36.885 130.395 -36.555 130.725 ;
        RECT -36.885 129.035 -36.555 129.365 ;
        RECT -36.885 127.675 -36.555 128.005 ;
        RECT -36.885 126.315 -36.555 126.645 ;
        RECT -36.885 124.955 -36.555 125.285 ;
        RECT -36.885 123.595 -36.555 123.925 ;
        RECT -36.885 122.235 -36.555 122.565 ;
        RECT -36.885 120.875 -36.555 121.205 ;
        RECT -36.885 119.515 -36.555 119.845 ;
        RECT -36.885 118.155 -36.555 118.485 ;
        RECT -36.885 116.795 -36.555 117.125 ;
        RECT -36.885 115.435 -36.555 115.765 ;
        RECT -36.885 114.075 -36.555 114.405 ;
        RECT -36.885 112.715 -36.555 113.045 ;
        RECT -36.885 111.355 -36.555 111.685 ;
        RECT -36.885 109.995 -36.555 110.325 ;
        RECT -36.885 108.635 -36.555 108.965 ;
        RECT -36.885 107.275 -36.555 107.605 ;
        RECT -36.885 105.915 -36.555 106.245 ;
        RECT -36.885 104.555 -36.555 104.885 ;
        RECT -36.885 103.195 -36.555 103.525 ;
        RECT -36.885 101.835 -36.555 102.165 ;
        RECT -36.885 100.475 -36.555 100.805 ;
        RECT -36.885 99.115 -36.555 99.445 ;
        RECT -36.885 97.755 -36.555 98.085 ;
        RECT -36.885 96.395 -36.555 96.725 ;
        RECT -36.885 95.035 -36.555 95.365 ;
        RECT -36.885 93.675 -36.555 94.005 ;
        RECT -36.885 92.315 -36.555 92.645 ;
        RECT -36.885 90.955 -36.555 91.285 ;
        RECT -36.885 89.595 -36.555 89.925 ;
        RECT -36.885 88.235 -36.555 88.565 ;
        RECT -36.885 86.875 -36.555 87.205 ;
        RECT -36.885 85.515 -36.555 85.845 ;
        RECT -36.885 84.155 -36.555 84.485 ;
        RECT -36.885 82.795 -36.555 83.125 ;
        RECT -36.885 81.435 -36.555 81.765 ;
        RECT -36.885 80.075 -36.555 80.405 ;
        RECT -36.885 78.715 -36.555 79.045 ;
        RECT -36.885 77.355 -36.555 77.685 ;
        RECT -36.885 75.995 -36.555 76.325 ;
        RECT -36.885 74.635 -36.555 74.965 ;
        RECT -36.885 73.275 -36.555 73.605 ;
        RECT -36.885 71.915 -36.555 72.245 ;
        RECT -36.885 70.555 -36.555 70.885 ;
        RECT -36.885 69.195 -36.555 69.525 ;
        RECT -36.885 67.835 -36.555 68.165 ;
        RECT -36.885 66.475 -36.555 66.805 ;
        RECT -36.885 65.115 -36.555 65.445 ;
        RECT -36.885 63.755 -36.555 64.085 ;
        RECT -36.885 62.395 -36.555 62.725 ;
        RECT -36.885 61.035 -36.555 61.365 ;
        RECT -36.885 59.675 -36.555 60.005 ;
        RECT -36.885 58.315 -36.555 58.645 ;
        RECT -36.885 56.955 -36.555 57.285 ;
        RECT -36.885 55.595 -36.555 55.925 ;
        RECT -36.885 54.235 -36.555 54.565 ;
        RECT -36.885 52.875 -36.555 53.205 ;
        RECT -36.885 51.515 -36.555 51.845 ;
        RECT -36.885 50.155 -36.555 50.485 ;
        RECT -36.885 48.795 -36.555 49.125 ;
        RECT -36.885 47.435 -36.555 47.765 ;
        RECT -36.885 46.075 -36.555 46.405 ;
        RECT -36.885 44.715 -36.555 45.045 ;
        RECT -36.885 43.355 -36.555 43.685 ;
        RECT -36.885 41.995 -36.555 42.325 ;
        RECT -36.885 40.635 -36.555 40.965 ;
        RECT -36.885 39.275 -36.555 39.605 ;
        RECT -36.885 37.915 -36.555 38.245 ;
        RECT -36.885 36.555 -36.555 36.885 ;
        RECT -36.885 35.195 -36.555 35.525 ;
        RECT -36.885 33.835 -36.555 34.165 ;
        RECT -36.885 32.475 -36.555 32.805 ;
        RECT -36.885 31.115 -36.555 31.445 ;
        RECT -36.885 29.755 -36.555 30.085 ;
        RECT -36.885 28.395 -36.555 28.725 ;
        RECT -36.885 27.035 -36.555 27.365 ;
        RECT -36.885 25.675 -36.555 26.005 ;
        RECT -36.885 24.315 -36.555 24.645 ;
        RECT -36.885 22.955 -36.555 23.285 ;
        RECT -36.885 21.595 -36.555 21.925 ;
        RECT -36.885 20.235 -36.555 20.565 ;
        RECT -36.885 18.875 -36.555 19.205 ;
        RECT -36.885 17.515 -36.555 17.845 ;
        RECT -36.885 16.155 -36.555 16.485 ;
        RECT -36.885 14.795 -36.555 15.125 ;
        RECT -36.885 13.435 -36.555 13.765 ;
        RECT -36.885 12.075 -36.555 12.405 ;
        RECT -36.885 10.715 -36.555 11.045 ;
        RECT -36.885 9.355 -36.555 9.685 ;
        RECT -36.885 7.995 -36.555 8.325 ;
        RECT -36.885 6.635 -36.555 6.965 ;
        RECT -36.885 5.275 -36.555 5.605 ;
        RECT -36.885 3.915 -36.555 4.245 ;
        RECT -36.885 2.555 -36.555 2.885 ;
        RECT -36.885 1.195 -36.555 1.525 ;
        RECT -36.885 -0.165 -36.555 0.165 ;
        RECT -36.885 -1.525 -36.555 -1.195 ;
        RECT -36.88 -1.525 -36.56 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.885 -4.245 -36.555 -3.915 ;
        RECT -36.885 -5.605 -36.555 -5.275 ;
        RECT -36.885 -8.325 -36.555 -7.995 ;
        RECT -36.885 -9.685 -36.555 -9.355 ;
        RECT -36.885 -12.405 -36.555 -12.075 ;
        RECT -36.885 -13.765 -36.555 -13.435 ;
        RECT -36.885 -15.125 -36.555 -14.795 ;
        RECT -36.885 -16.485 -36.555 -16.155 ;
        RECT -36.885 -17.845 -36.555 -17.515 ;
        RECT -36.885 -19.205 -36.555 -18.875 ;
        RECT -36.885 -20.565 -36.555 -20.235 ;
        RECT -36.885 -21.925 -36.555 -21.595 ;
        RECT -36.885 -23.285 -36.555 -22.955 ;
        RECT -36.885 -30.66 -36.555 -30.33 ;
        RECT -36.885 -31.445 -36.555 -31.115 ;
        RECT -36.885 -32.805 -36.555 -32.475 ;
        RECT -36.885 -34.165 -36.555 -33.835 ;
        RECT -36.885 -36.885 -36.555 -36.555 ;
        RECT -36.885 -37.85 -36.555 -37.52 ;
        RECT -36.885 -40.965 -36.555 -40.635 ;
        RECT -36.885 -46.405 -36.555 -46.075 ;
        RECT -36.885 -47.765 -36.555 -47.435 ;
        RECT -36.885 -49.125 -36.555 -48.795 ;
        RECT -36.885 -50.485 -36.555 -50.155 ;
        RECT -36.885 -51.845 -36.555 -51.515 ;
        RECT -36.885 -53.205 -36.555 -52.875 ;
        RECT -36.885 -54.565 -36.555 -54.235 ;
        RECT -36.885 -55.925 -36.555 -55.595 ;
        RECT -36.885 -57.285 -36.555 -56.955 ;
        RECT -36.885 -58.645 -36.555 -58.315 ;
        RECT -36.885 -60.005 -36.555 -59.675 ;
        RECT -36.885 -61.365 -36.555 -61.035 ;
        RECT -36.885 -62.725 -36.555 -62.395 ;
        RECT -36.885 -64.085 -36.555 -63.755 ;
        RECT -36.885 -65.445 -36.555 -65.115 ;
        RECT -36.885 -66.805 -36.555 -66.475 ;
        RECT -36.885 -68.165 -36.555 -67.835 ;
        RECT -36.885 -69.525 -36.555 -69.195 ;
        RECT -36.885 -70.885 -36.555 -70.555 ;
        RECT -36.885 -72.245 -36.555 -71.915 ;
        RECT -36.885 -73.605 -36.555 -73.275 ;
        RECT -36.885 -74.965 -36.555 -74.635 ;
        RECT -36.885 -76.325 -36.555 -75.995 ;
        RECT -36.885 -77.685 -36.555 -77.355 ;
        RECT -36.885 -79.045 -36.555 -78.715 ;
        RECT -36.885 -80.405 -36.555 -80.075 ;
        RECT -36.885 -81.765 -36.555 -81.435 ;
        RECT -36.885 -83.125 -36.555 -82.795 ;
        RECT -36.885 -84.485 -36.555 -84.155 ;
        RECT -36.885 -85.845 -36.555 -85.515 ;
        RECT -36.885 -87.205 -36.555 -86.875 ;
        RECT -36.885 -88.565 -36.555 -88.235 ;
        RECT -36.885 -89.925 -36.555 -89.595 ;
        RECT -36.885 -91.285 -36.555 -90.955 ;
        RECT -36.885 -92.645 -36.555 -92.315 ;
        RECT -36.885 -94.005 -36.555 -93.675 ;
        RECT -36.885 -95.365 -36.555 -95.035 ;
        RECT -36.885 -96.725 -36.555 -96.395 ;
        RECT -36.885 -98.085 -36.555 -97.755 ;
        RECT -36.885 -99.445 -36.555 -99.115 ;
        RECT -36.885 -100.805 -36.555 -100.475 ;
        RECT -36.885 -102.165 -36.555 -101.835 ;
        RECT -36.885 -103.525 -36.555 -103.195 ;
        RECT -36.885 -104.885 -36.555 -104.555 ;
        RECT -36.885 -106.245 -36.555 -105.915 ;
        RECT -36.885 -107.605 -36.555 -107.275 ;
        RECT -36.885 -108.965 -36.555 -108.635 ;
        RECT -36.885 -110.325 -36.555 -109.995 ;
        RECT -36.885 -111.685 -36.555 -111.355 ;
        RECT -36.885 -113.045 -36.555 -112.715 ;
        RECT -36.885 -114.405 -36.555 -114.075 ;
        RECT -36.885 -115.765 -36.555 -115.435 ;
        RECT -36.885 -117.125 -36.555 -116.795 ;
        RECT -36.885 -118.485 -36.555 -118.155 ;
        RECT -36.885 -119.845 -36.555 -119.515 ;
        RECT -36.885 -123.925 -36.555 -123.595 ;
        RECT -36.885 -129.365 -36.555 -129.035 ;
        RECT -36.885 -130.725 -36.555 -130.395 ;
        RECT -36.885 -131.47 -36.555 -131.14 ;
        RECT -36.885 -133.445 -36.555 -133.115 ;
        RECT -36.885 -134.805 -36.555 -134.475 ;
        RECT -36.885 -136.165 -36.555 -135.835 ;
        RECT -36.885 -137.525 -36.555 -137.195 ;
        RECT -36.885 -140.245 -36.555 -139.915 ;
        RECT -36.885 -141.605 -36.555 -141.275 ;
        RECT -36.885 -142.965 -36.555 -142.635 ;
        RECT -36.885 -144.31 -36.555 -143.98 ;
        RECT -36.885 -145.685 -36.555 -145.355 ;
        RECT -36.885 -147.045 -36.555 -146.715 ;
        RECT -36.885 -149.765 -36.555 -149.435 ;
        RECT -36.885 -153.845 -36.555 -153.515 ;
        RECT -36.885 -155.205 -36.555 -154.875 ;
        RECT -36.885 -156.565 -36.555 -156.235 ;
        RECT -36.885 -157.925 -36.555 -157.595 ;
        RECT -36.885 -159.285 -36.555 -158.955 ;
        RECT -36.885 -162.005 -36.555 -161.675 ;
        RECT -36.885 -163.365 -36.555 -163.035 ;
        RECT -36.885 -164.725 -36.555 -164.395 ;
        RECT -36.885 -166.085 -36.555 -165.755 ;
        RECT -36.885 -167.445 -36.555 -167.115 ;
        RECT -36.885 -168.805 -36.555 -168.475 ;
        RECT -36.885 -170.165 -36.555 -169.835 ;
        RECT -36.885 -171.525 -36.555 -171.195 ;
        RECT -36.885 -172.885 -36.555 -172.555 ;
        RECT -36.885 -174.245 -36.555 -173.915 ;
        RECT -36.885 -175.605 -36.555 -175.275 ;
        RECT -36.885 -176.965 -36.555 -176.635 ;
        RECT -36.885 -178.325 -36.555 -177.995 ;
        RECT -36.885 -179.685 -36.555 -179.355 ;
        RECT -36.885 -181.045 -36.555 -180.715 ;
        RECT -36.885 -182.405 -36.555 -182.075 ;
        RECT -36.885 -183.765 -36.555 -183.435 ;
        RECT -36.885 -185.125 -36.555 -184.795 ;
        RECT -36.885 -186.485 -36.555 -186.155 ;
        RECT -36.885 -187.845 -36.555 -187.515 ;
        RECT -36.885 -189.205 -36.555 -188.875 ;
        RECT -36.885 -190.565 -36.555 -190.235 ;
        RECT -36.885 -191.925 -36.555 -191.595 ;
        RECT -36.885 -193.285 -36.555 -192.955 ;
        RECT -36.885 -194.645 -36.555 -194.315 ;
        RECT -36.885 -196.005 -36.555 -195.675 ;
        RECT -36.885 -197.365 -36.555 -197.035 ;
        RECT -36.885 -198.725 -36.555 -198.395 ;
        RECT -36.885 -200.085 -36.555 -199.755 ;
        RECT -36.885 -201.445 -36.555 -201.115 ;
        RECT -36.885 -202.805 -36.555 -202.475 ;
        RECT -36.885 -204.165 -36.555 -203.835 ;
        RECT -36.885 -205.525 -36.555 -205.195 ;
        RECT -36.885 -206.885 -36.555 -206.555 ;
        RECT -36.885 -208.245 -36.555 -207.915 ;
        RECT -36.885 -209.605 -36.555 -209.275 ;
        RECT -36.885 -210.965 -36.555 -210.635 ;
        RECT -36.885 -212.325 -36.555 -211.995 ;
        RECT -36.885 -213.685 -36.555 -213.355 ;
        RECT -36.885 -215.045 -36.555 -214.715 ;
        RECT -36.885 -216.405 -36.555 -216.075 ;
        RECT -36.885 -217.765 -36.555 -217.435 ;
        RECT -36.885 -219.125 -36.555 -218.795 ;
        RECT -36.885 -220.485 -36.555 -220.155 ;
        RECT -36.885 -221.845 -36.555 -221.515 ;
        RECT -36.885 -223.205 -36.555 -222.875 ;
        RECT -36.885 -224.565 -36.555 -224.235 ;
        RECT -36.885 -226.155 -36.555 -225.825 ;
        RECT -36.885 -227.285 -36.555 -226.955 ;
        RECT -36.885 -228.645 -36.555 -228.315 ;
        RECT -36.885 -230.005 -36.555 -229.675 ;
        RECT -36.885 -234.085 -36.555 -233.755 ;
        RECT -36.885 -235.445 -36.555 -235.115 ;
        RECT -36.885 -236.805 -36.555 -236.475 ;
        RECT -36.885 -238.165 -36.555 -237.835 ;
        RECT -36.885 -243.81 -36.555 -242.68 ;
        RECT -36.88 -243.925 -36.56 -3.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 -95.365 -35.195 -95.035 ;
        RECT -35.525 -96.725 -35.195 -96.395 ;
        RECT -35.525 -98.085 -35.195 -97.755 ;
        RECT -35.525 -99.445 -35.195 -99.115 ;
        RECT -35.525 -100.805 -35.195 -100.475 ;
        RECT -35.525 -102.165 -35.195 -101.835 ;
        RECT -35.525 -103.525 -35.195 -103.195 ;
        RECT -35.525 -104.885 -35.195 -104.555 ;
        RECT -35.525 -106.245 -35.195 -105.915 ;
        RECT -35.525 -107.605 -35.195 -107.275 ;
        RECT -35.525 -108.965 -35.195 -108.635 ;
        RECT -35.525 -110.325 -35.195 -109.995 ;
        RECT -35.525 -111.685 -35.195 -111.355 ;
        RECT -35.525 -113.045 -35.195 -112.715 ;
        RECT -35.525 -114.405 -35.195 -114.075 ;
        RECT -35.525 -115.765 -35.195 -115.435 ;
        RECT -35.525 -117.125 -35.195 -116.795 ;
        RECT -35.525 -118.485 -35.195 -118.155 ;
        RECT -35.525 -119.845 -35.195 -119.515 ;
        RECT -35.525 -123.925 -35.195 -123.595 ;
        RECT -35.525 -129.365 -35.195 -129.035 ;
        RECT -35.525 -130.725 -35.195 -130.395 ;
        RECT -35.525 -132.085 -35.195 -131.755 ;
        RECT -35.525 -133.445 -35.195 -133.115 ;
        RECT -35.525 -134.805 -35.195 -134.475 ;
        RECT -35.525 -136.165 -35.195 -135.835 ;
        RECT -35.525 -137.525 -35.195 -137.195 ;
        RECT -35.525 -138.885 -35.195 -138.555 ;
        RECT -35.525 -140.245 -35.195 -139.915 ;
        RECT -35.525 -141.605 -35.195 -141.275 ;
        RECT -35.525 -142.965 -35.195 -142.635 ;
        RECT -35.525 -144.325 -35.195 -143.995 ;
        RECT -35.525 -145.685 -35.195 -145.355 ;
        RECT -35.525 -147.045 -35.195 -146.715 ;
        RECT -35.525 -148.405 -35.195 -148.075 ;
        RECT -35.525 -149.765 -35.195 -149.435 ;
        RECT -35.525 -151.125 -35.195 -150.795 ;
        RECT -35.52 -151.8 -35.2 248.005 ;
        RECT -35.525 246.76 -35.195 247.89 ;
        RECT -35.525 241.915 -35.195 242.245 ;
        RECT -35.525 240.555 -35.195 240.885 ;
        RECT -35.525 239.195 -35.195 239.525 ;
        RECT -35.525 237.835 -35.195 238.165 ;
        RECT -35.525 236.475 -35.195 236.805 ;
        RECT -35.525 235.115 -35.195 235.445 ;
        RECT -35.525 233.755 -35.195 234.085 ;
        RECT -35.525 232.395 -35.195 232.725 ;
        RECT -35.525 231.035 -35.195 231.365 ;
        RECT -35.525 229.675 -35.195 230.005 ;
        RECT -35.525 228.315 -35.195 228.645 ;
        RECT -35.525 226.955 -35.195 227.285 ;
        RECT -35.525 225.595 -35.195 225.925 ;
        RECT -35.525 224.235 -35.195 224.565 ;
        RECT -35.525 222.875 -35.195 223.205 ;
        RECT -35.525 221.515 -35.195 221.845 ;
        RECT -35.525 220.155 -35.195 220.485 ;
        RECT -35.525 218.795 -35.195 219.125 ;
        RECT -35.525 217.435 -35.195 217.765 ;
        RECT -35.525 216.075 -35.195 216.405 ;
        RECT -35.525 214.715 -35.195 215.045 ;
        RECT -35.525 213.355 -35.195 213.685 ;
        RECT -35.525 211.995 -35.195 212.325 ;
        RECT -35.525 210.635 -35.195 210.965 ;
        RECT -35.525 209.275 -35.195 209.605 ;
        RECT -35.525 207.915 -35.195 208.245 ;
        RECT -35.525 206.555 -35.195 206.885 ;
        RECT -35.525 205.195 -35.195 205.525 ;
        RECT -35.525 203.835 -35.195 204.165 ;
        RECT -35.525 202.475 -35.195 202.805 ;
        RECT -35.525 201.115 -35.195 201.445 ;
        RECT -35.525 199.755 -35.195 200.085 ;
        RECT -35.525 198.395 -35.195 198.725 ;
        RECT -35.525 197.035 -35.195 197.365 ;
        RECT -35.525 195.675 -35.195 196.005 ;
        RECT -35.525 194.315 -35.195 194.645 ;
        RECT -35.525 192.955 -35.195 193.285 ;
        RECT -35.525 191.595 -35.195 191.925 ;
        RECT -35.525 190.235 -35.195 190.565 ;
        RECT -35.525 188.875 -35.195 189.205 ;
        RECT -35.525 187.515 -35.195 187.845 ;
        RECT -35.525 186.155 -35.195 186.485 ;
        RECT -35.525 184.795 -35.195 185.125 ;
        RECT -35.525 183.435 -35.195 183.765 ;
        RECT -35.525 182.075 -35.195 182.405 ;
        RECT -35.525 180.715 -35.195 181.045 ;
        RECT -35.525 179.355 -35.195 179.685 ;
        RECT -35.525 177.995 -35.195 178.325 ;
        RECT -35.525 176.635 -35.195 176.965 ;
        RECT -35.525 175.275 -35.195 175.605 ;
        RECT -35.525 173.915 -35.195 174.245 ;
        RECT -35.525 172.555 -35.195 172.885 ;
        RECT -35.525 171.195 -35.195 171.525 ;
        RECT -35.525 169.835 -35.195 170.165 ;
        RECT -35.525 168.475 -35.195 168.805 ;
        RECT -35.525 167.115 -35.195 167.445 ;
        RECT -35.525 165.755 -35.195 166.085 ;
        RECT -35.525 164.395 -35.195 164.725 ;
        RECT -35.525 163.035 -35.195 163.365 ;
        RECT -35.525 161.675 -35.195 162.005 ;
        RECT -35.525 160.315 -35.195 160.645 ;
        RECT -35.525 158.955 -35.195 159.285 ;
        RECT -35.525 157.595 -35.195 157.925 ;
        RECT -35.525 156.235 -35.195 156.565 ;
        RECT -35.525 154.875 -35.195 155.205 ;
        RECT -35.525 153.515 -35.195 153.845 ;
        RECT -35.525 152.155 -35.195 152.485 ;
        RECT -35.525 150.795 -35.195 151.125 ;
        RECT -35.525 149.435 -35.195 149.765 ;
        RECT -35.525 148.075 -35.195 148.405 ;
        RECT -35.525 146.715 -35.195 147.045 ;
        RECT -35.525 145.355 -35.195 145.685 ;
        RECT -35.525 143.995 -35.195 144.325 ;
        RECT -35.525 142.635 -35.195 142.965 ;
        RECT -35.525 141.275 -35.195 141.605 ;
        RECT -35.525 139.915 -35.195 140.245 ;
        RECT -35.525 138.555 -35.195 138.885 ;
        RECT -35.525 137.195 -35.195 137.525 ;
        RECT -35.525 135.835 -35.195 136.165 ;
        RECT -35.525 134.475 -35.195 134.805 ;
        RECT -35.525 133.115 -35.195 133.445 ;
        RECT -35.525 131.755 -35.195 132.085 ;
        RECT -35.525 130.395 -35.195 130.725 ;
        RECT -35.525 129.035 -35.195 129.365 ;
        RECT -35.525 127.675 -35.195 128.005 ;
        RECT -35.525 126.315 -35.195 126.645 ;
        RECT -35.525 124.955 -35.195 125.285 ;
        RECT -35.525 123.595 -35.195 123.925 ;
        RECT -35.525 122.235 -35.195 122.565 ;
        RECT -35.525 120.875 -35.195 121.205 ;
        RECT -35.525 119.515 -35.195 119.845 ;
        RECT -35.525 118.155 -35.195 118.485 ;
        RECT -35.525 116.795 -35.195 117.125 ;
        RECT -35.525 115.435 -35.195 115.765 ;
        RECT -35.525 114.075 -35.195 114.405 ;
        RECT -35.525 112.715 -35.195 113.045 ;
        RECT -35.525 111.355 -35.195 111.685 ;
        RECT -35.525 109.995 -35.195 110.325 ;
        RECT -35.525 108.635 -35.195 108.965 ;
        RECT -35.525 107.275 -35.195 107.605 ;
        RECT -35.525 105.915 -35.195 106.245 ;
        RECT -35.525 104.555 -35.195 104.885 ;
        RECT -35.525 103.195 -35.195 103.525 ;
        RECT -35.525 101.835 -35.195 102.165 ;
        RECT -35.525 100.475 -35.195 100.805 ;
        RECT -35.525 99.115 -35.195 99.445 ;
        RECT -35.525 97.755 -35.195 98.085 ;
        RECT -35.525 96.395 -35.195 96.725 ;
        RECT -35.525 95.035 -35.195 95.365 ;
        RECT -35.525 93.675 -35.195 94.005 ;
        RECT -35.525 92.315 -35.195 92.645 ;
        RECT -35.525 90.955 -35.195 91.285 ;
        RECT -35.525 89.595 -35.195 89.925 ;
        RECT -35.525 88.235 -35.195 88.565 ;
        RECT -35.525 86.875 -35.195 87.205 ;
        RECT -35.525 85.515 -35.195 85.845 ;
        RECT -35.525 84.155 -35.195 84.485 ;
        RECT -35.525 82.795 -35.195 83.125 ;
        RECT -35.525 81.435 -35.195 81.765 ;
        RECT -35.525 80.075 -35.195 80.405 ;
        RECT -35.525 78.715 -35.195 79.045 ;
        RECT -35.525 77.355 -35.195 77.685 ;
        RECT -35.525 75.995 -35.195 76.325 ;
        RECT -35.525 74.635 -35.195 74.965 ;
        RECT -35.525 73.275 -35.195 73.605 ;
        RECT -35.525 71.915 -35.195 72.245 ;
        RECT -35.525 70.555 -35.195 70.885 ;
        RECT -35.525 69.195 -35.195 69.525 ;
        RECT -35.525 67.835 -35.195 68.165 ;
        RECT -35.525 66.475 -35.195 66.805 ;
        RECT -35.525 65.115 -35.195 65.445 ;
        RECT -35.525 63.755 -35.195 64.085 ;
        RECT -35.525 62.395 -35.195 62.725 ;
        RECT -35.525 61.035 -35.195 61.365 ;
        RECT -35.525 59.675 -35.195 60.005 ;
        RECT -35.525 58.315 -35.195 58.645 ;
        RECT -35.525 56.955 -35.195 57.285 ;
        RECT -35.525 55.595 -35.195 55.925 ;
        RECT -35.525 54.235 -35.195 54.565 ;
        RECT -35.525 52.875 -35.195 53.205 ;
        RECT -35.525 51.515 -35.195 51.845 ;
        RECT -35.525 50.155 -35.195 50.485 ;
        RECT -35.525 48.795 -35.195 49.125 ;
        RECT -35.525 47.435 -35.195 47.765 ;
        RECT -35.525 46.075 -35.195 46.405 ;
        RECT -35.525 44.715 -35.195 45.045 ;
        RECT -35.525 43.355 -35.195 43.685 ;
        RECT -35.525 41.995 -35.195 42.325 ;
        RECT -35.525 40.635 -35.195 40.965 ;
        RECT -35.525 39.275 -35.195 39.605 ;
        RECT -35.525 37.915 -35.195 38.245 ;
        RECT -35.525 36.555 -35.195 36.885 ;
        RECT -35.525 35.195 -35.195 35.525 ;
        RECT -35.525 33.835 -35.195 34.165 ;
        RECT -35.525 32.475 -35.195 32.805 ;
        RECT -35.525 31.115 -35.195 31.445 ;
        RECT -35.525 29.755 -35.195 30.085 ;
        RECT -35.525 28.395 -35.195 28.725 ;
        RECT -35.525 27.035 -35.195 27.365 ;
        RECT -35.525 25.675 -35.195 26.005 ;
        RECT -35.525 24.315 -35.195 24.645 ;
        RECT -35.525 22.955 -35.195 23.285 ;
        RECT -35.525 21.595 -35.195 21.925 ;
        RECT -35.525 20.235 -35.195 20.565 ;
        RECT -35.525 18.875 -35.195 19.205 ;
        RECT -35.525 17.515 -35.195 17.845 ;
        RECT -35.525 16.155 -35.195 16.485 ;
        RECT -35.525 14.795 -35.195 15.125 ;
        RECT -35.525 13.435 -35.195 13.765 ;
        RECT -35.525 12.075 -35.195 12.405 ;
        RECT -35.525 10.715 -35.195 11.045 ;
        RECT -35.525 9.355 -35.195 9.685 ;
        RECT -35.525 7.995 -35.195 8.325 ;
        RECT -35.525 6.635 -35.195 6.965 ;
        RECT -35.525 5.275 -35.195 5.605 ;
        RECT -35.525 3.915 -35.195 4.245 ;
        RECT -35.525 2.555 -35.195 2.885 ;
        RECT -35.525 1.195 -35.195 1.525 ;
        RECT -35.525 -0.165 -35.195 0.165 ;
        RECT -35.525 -1.525 -35.195 -1.195 ;
        RECT -35.525 -4.245 -35.195 -3.915 ;
        RECT -35.525 -8.325 -35.195 -7.995 ;
        RECT -35.525 -9.685 -35.195 -9.355 ;
        RECT -35.525 -12.405 -35.195 -12.075 ;
        RECT -35.525 -13.765 -35.195 -13.435 ;
        RECT -35.525 -15.125 -35.195 -14.795 ;
        RECT -35.525 -16.485 -35.195 -16.155 ;
        RECT -35.525 -17.845 -35.195 -17.515 ;
        RECT -35.525 -19.205 -35.195 -18.875 ;
        RECT -35.525 -20.565 -35.195 -20.235 ;
        RECT -35.525 -21.925 -35.195 -21.595 ;
        RECT -35.525 -23.285 -35.195 -22.955 ;
        RECT -35.525 -30.66 -35.195 -30.33 ;
        RECT -35.525 -31.445 -35.195 -31.115 ;
        RECT -35.525 -32.805 -35.195 -32.475 ;
        RECT -35.525 -34.165 -35.195 -33.835 ;
        RECT -35.525 -36.885 -35.195 -36.555 ;
        RECT -35.525 -37.85 -35.195 -37.52 ;
        RECT -35.525 -40.965 -35.195 -40.635 ;
        RECT -35.525 -46.405 -35.195 -46.075 ;
        RECT -35.525 -49.125 -35.195 -48.795 ;
        RECT -35.525 -50.485 -35.195 -50.155 ;
        RECT -35.525 -53.205 -35.195 -52.875 ;
        RECT -35.525 -55.925 -35.195 -55.595 ;
        RECT -35.525 -61.365 -35.195 -61.035 ;
        RECT -35.525 -62.725 -35.195 -62.395 ;
        RECT -35.525 -64.085 -35.195 -63.755 ;
        RECT -35.525 -65.445 -35.195 -65.115 ;
        RECT -35.525 -66.805 -35.195 -66.475 ;
        RECT -35.525 -68.165 -35.195 -67.835 ;
        RECT -35.525 -69.525 -35.195 -69.195 ;
        RECT -35.525 -70.885 -35.195 -70.555 ;
        RECT -35.525 -72.245 -35.195 -71.915 ;
        RECT -35.525 -73.605 -35.195 -73.275 ;
        RECT -35.525 -74.965 -35.195 -74.635 ;
        RECT -35.525 -76.325 -35.195 -75.995 ;
        RECT -35.525 -77.685 -35.195 -77.355 ;
        RECT -35.525 -79.045 -35.195 -78.715 ;
        RECT -35.525 -80.405 -35.195 -80.075 ;
        RECT -35.525 -81.765 -35.195 -81.435 ;
        RECT -35.525 -83.125 -35.195 -82.795 ;
        RECT -35.525 -84.485 -35.195 -84.155 ;
        RECT -35.525 -85.845 -35.195 -85.515 ;
        RECT -35.525 -87.205 -35.195 -86.875 ;
        RECT -35.525 -88.565 -35.195 -88.235 ;
        RECT -35.525 -89.925 -35.195 -89.595 ;
        RECT -35.525 -91.285 -35.195 -90.955 ;
        RECT -35.525 -92.645 -35.195 -92.315 ;
        RECT -35.525 -94.005 -35.195 -93.675 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 -129.365 -44.715 -129.035 ;
        RECT -45.045 -130.725 -44.715 -130.395 ;
        RECT -45.045 -131.47 -44.715 -131.14 ;
        RECT -45.045 -133.445 -44.715 -133.115 ;
        RECT -45.045 -134.805 -44.715 -134.475 ;
        RECT -45.045 -136.165 -44.715 -135.835 ;
        RECT -45.045 -137.525 -44.715 -137.195 ;
        RECT -45.045 -140.245 -44.715 -139.915 ;
        RECT -45.045 -141.605 -44.715 -141.275 ;
        RECT -45.045 -142.965 -44.715 -142.635 ;
        RECT -45.045 -144.31 -44.715 -143.98 ;
        RECT -45.045 -145.685 -44.715 -145.355 ;
        RECT -45.045 -147.045 -44.715 -146.715 ;
        RECT -45.045 -149.765 -44.715 -149.435 ;
        RECT -45.045 -152.485 -44.715 -152.155 ;
        RECT -45.045 -153.845 -44.715 -153.515 ;
        RECT -45.045 -155.205 -44.715 -154.875 ;
        RECT -45.045 -156.565 -44.715 -156.235 ;
        RECT -45.045 -157.925 -44.715 -157.595 ;
        RECT -45.045 -159.285 -44.715 -158.955 ;
        RECT -45.045 -162.005 -44.715 -161.675 ;
        RECT -45.045 -163.365 -44.715 -163.035 ;
        RECT -45.045 -164.725 -44.715 -164.395 ;
        RECT -45.045 -166.085 -44.715 -165.755 ;
        RECT -45.045 -167.445 -44.715 -167.115 ;
        RECT -45.045 -168.805 -44.715 -168.475 ;
        RECT -45.045 -170.165 -44.715 -169.835 ;
        RECT -45.045 -171.525 -44.715 -171.195 ;
        RECT -45.045 -172.885 -44.715 -172.555 ;
        RECT -45.045 -174.245 -44.715 -173.915 ;
        RECT -45.045 -175.605 -44.715 -175.275 ;
        RECT -45.045 -176.965 -44.715 -176.635 ;
        RECT -45.045 -178.325 -44.715 -177.995 ;
        RECT -45.045 -179.685 -44.715 -179.355 ;
        RECT -45.045 -181.045 -44.715 -180.715 ;
        RECT -45.045 -182.405 -44.715 -182.075 ;
        RECT -45.045 -183.765 -44.715 -183.435 ;
        RECT -45.045 -185.125 -44.715 -184.795 ;
        RECT -45.045 -186.485 -44.715 -186.155 ;
        RECT -45.045 -187.845 -44.715 -187.515 ;
        RECT -45.045 -189.205 -44.715 -188.875 ;
        RECT -45.045 -190.565 -44.715 -190.235 ;
        RECT -45.045 -191.925 -44.715 -191.595 ;
        RECT -45.045 -193.285 -44.715 -192.955 ;
        RECT -45.045 -194.645 -44.715 -194.315 ;
        RECT -45.045 -196.005 -44.715 -195.675 ;
        RECT -45.045 -197.365 -44.715 -197.035 ;
        RECT -45.045 -198.725 -44.715 -198.395 ;
        RECT -45.045 -200.085 -44.715 -199.755 ;
        RECT -45.045 -201.445 -44.715 -201.115 ;
        RECT -45.045 -202.805 -44.715 -202.475 ;
        RECT -45.045 -204.165 -44.715 -203.835 ;
        RECT -45.045 -205.525 -44.715 -205.195 ;
        RECT -45.045 -206.885 -44.715 -206.555 ;
        RECT -45.045 -208.245 -44.715 -207.915 ;
        RECT -45.045 -209.605 -44.715 -209.275 ;
        RECT -45.045 -210.965 -44.715 -210.635 ;
        RECT -45.045 -212.325 -44.715 -211.995 ;
        RECT -45.045 -213.685 -44.715 -213.355 ;
        RECT -45.045 -215.045 -44.715 -214.715 ;
        RECT -45.045 -216.405 -44.715 -216.075 ;
        RECT -45.045 -217.765 -44.715 -217.435 ;
        RECT -45.045 -219.125 -44.715 -218.795 ;
        RECT -45.045 -220.485 -44.715 -220.155 ;
        RECT -45.045 -221.845 -44.715 -221.515 ;
        RECT -45.045 -223.205 -44.715 -222.875 ;
        RECT -45.045 -224.565 -44.715 -224.235 ;
        RECT -45.045 -226.155 -44.715 -225.825 ;
        RECT -45.045 -227.285 -44.715 -226.955 ;
        RECT -45.045 -228.645 -44.715 -228.315 ;
        RECT -45.045 -231.365 -44.715 -231.035 ;
        RECT -45.045 -234.085 -44.715 -233.755 ;
        RECT -45.045 -235.445 -44.715 -235.115 ;
        RECT -45.045 -236.805 -44.715 -236.475 ;
        RECT -45.045 -238.165 -44.715 -237.835 ;
        RECT -45.045 -243.81 -44.715 -242.68 ;
        RECT -45.04 -243.925 -44.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 246.76 -43.355 247.89 ;
        RECT -43.685 241.915 -43.355 242.245 ;
        RECT -43.685 240.555 -43.355 240.885 ;
        RECT -43.685 239.195 -43.355 239.525 ;
        RECT -43.685 237.835 -43.355 238.165 ;
        RECT -43.685 236.475 -43.355 236.805 ;
        RECT -43.685 235.115 -43.355 235.445 ;
        RECT -43.685 233.755 -43.355 234.085 ;
        RECT -43.685 232.395 -43.355 232.725 ;
        RECT -43.685 231.035 -43.355 231.365 ;
        RECT -43.685 229.675 -43.355 230.005 ;
        RECT -43.685 228.315 -43.355 228.645 ;
        RECT -43.685 226.955 -43.355 227.285 ;
        RECT -43.685 225.595 -43.355 225.925 ;
        RECT -43.685 224.235 -43.355 224.565 ;
        RECT -43.685 222.875 -43.355 223.205 ;
        RECT -43.685 221.515 -43.355 221.845 ;
        RECT -43.685 220.155 -43.355 220.485 ;
        RECT -43.685 218.795 -43.355 219.125 ;
        RECT -43.685 217.435 -43.355 217.765 ;
        RECT -43.685 216.075 -43.355 216.405 ;
        RECT -43.685 214.715 -43.355 215.045 ;
        RECT -43.685 213.355 -43.355 213.685 ;
        RECT -43.685 211.995 -43.355 212.325 ;
        RECT -43.685 210.635 -43.355 210.965 ;
        RECT -43.685 209.275 -43.355 209.605 ;
        RECT -43.685 207.915 -43.355 208.245 ;
        RECT -43.685 206.555 -43.355 206.885 ;
        RECT -43.685 205.195 -43.355 205.525 ;
        RECT -43.685 203.835 -43.355 204.165 ;
        RECT -43.685 202.475 -43.355 202.805 ;
        RECT -43.685 201.115 -43.355 201.445 ;
        RECT -43.685 199.755 -43.355 200.085 ;
        RECT -43.685 198.395 -43.355 198.725 ;
        RECT -43.685 197.035 -43.355 197.365 ;
        RECT -43.685 195.675 -43.355 196.005 ;
        RECT -43.685 194.315 -43.355 194.645 ;
        RECT -43.685 192.955 -43.355 193.285 ;
        RECT -43.685 191.595 -43.355 191.925 ;
        RECT -43.685 190.235 -43.355 190.565 ;
        RECT -43.685 188.875 -43.355 189.205 ;
        RECT -43.685 187.515 -43.355 187.845 ;
        RECT -43.685 186.155 -43.355 186.485 ;
        RECT -43.685 184.795 -43.355 185.125 ;
        RECT -43.685 183.435 -43.355 183.765 ;
        RECT -43.685 182.075 -43.355 182.405 ;
        RECT -43.685 180.715 -43.355 181.045 ;
        RECT -43.685 179.355 -43.355 179.685 ;
        RECT -43.685 177.995 -43.355 178.325 ;
        RECT -43.685 176.635 -43.355 176.965 ;
        RECT -43.685 175.275 -43.355 175.605 ;
        RECT -43.685 173.915 -43.355 174.245 ;
        RECT -43.685 172.555 -43.355 172.885 ;
        RECT -43.685 171.195 -43.355 171.525 ;
        RECT -43.685 169.835 -43.355 170.165 ;
        RECT -43.685 168.475 -43.355 168.805 ;
        RECT -43.685 167.115 -43.355 167.445 ;
        RECT -43.685 165.755 -43.355 166.085 ;
        RECT -43.685 164.395 -43.355 164.725 ;
        RECT -43.685 163.035 -43.355 163.365 ;
        RECT -43.685 161.675 -43.355 162.005 ;
        RECT -43.685 160.315 -43.355 160.645 ;
        RECT -43.685 158.955 -43.355 159.285 ;
        RECT -43.685 157.595 -43.355 157.925 ;
        RECT -43.685 156.235 -43.355 156.565 ;
        RECT -43.685 154.875 -43.355 155.205 ;
        RECT -43.685 153.515 -43.355 153.845 ;
        RECT -43.685 152.155 -43.355 152.485 ;
        RECT -43.685 150.795 -43.355 151.125 ;
        RECT -43.685 149.435 -43.355 149.765 ;
        RECT -43.685 148.075 -43.355 148.405 ;
        RECT -43.685 146.715 -43.355 147.045 ;
        RECT -43.685 145.355 -43.355 145.685 ;
        RECT -43.685 143.995 -43.355 144.325 ;
        RECT -43.685 142.635 -43.355 142.965 ;
        RECT -43.685 141.275 -43.355 141.605 ;
        RECT -43.685 139.915 -43.355 140.245 ;
        RECT -43.685 138.555 -43.355 138.885 ;
        RECT -43.685 137.195 -43.355 137.525 ;
        RECT -43.685 135.835 -43.355 136.165 ;
        RECT -43.685 134.475 -43.355 134.805 ;
        RECT -43.685 133.115 -43.355 133.445 ;
        RECT -43.685 131.755 -43.355 132.085 ;
        RECT -43.685 130.395 -43.355 130.725 ;
        RECT -43.685 129.035 -43.355 129.365 ;
        RECT -43.685 127.675 -43.355 128.005 ;
        RECT -43.685 126.315 -43.355 126.645 ;
        RECT -43.685 124.955 -43.355 125.285 ;
        RECT -43.685 123.595 -43.355 123.925 ;
        RECT -43.685 122.235 -43.355 122.565 ;
        RECT -43.685 120.875 -43.355 121.205 ;
        RECT -43.685 119.515 -43.355 119.845 ;
        RECT -43.685 118.155 -43.355 118.485 ;
        RECT -43.685 116.795 -43.355 117.125 ;
        RECT -43.685 115.435 -43.355 115.765 ;
        RECT -43.685 114.075 -43.355 114.405 ;
        RECT -43.685 112.715 -43.355 113.045 ;
        RECT -43.685 111.355 -43.355 111.685 ;
        RECT -43.685 109.995 -43.355 110.325 ;
        RECT -43.685 108.635 -43.355 108.965 ;
        RECT -43.685 107.275 -43.355 107.605 ;
        RECT -43.685 105.915 -43.355 106.245 ;
        RECT -43.685 104.555 -43.355 104.885 ;
        RECT -43.685 103.195 -43.355 103.525 ;
        RECT -43.685 101.835 -43.355 102.165 ;
        RECT -43.685 100.475 -43.355 100.805 ;
        RECT -43.685 99.115 -43.355 99.445 ;
        RECT -43.685 97.755 -43.355 98.085 ;
        RECT -43.685 96.395 -43.355 96.725 ;
        RECT -43.685 95.035 -43.355 95.365 ;
        RECT -43.685 93.675 -43.355 94.005 ;
        RECT -43.685 92.315 -43.355 92.645 ;
        RECT -43.685 90.955 -43.355 91.285 ;
        RECT -43.685 89.595 -43.355 89.925 ;
        RECT -43.685 88.235 -43.355 88.565 ;
        RECT -43.685 86.875 -43.355 87.205 ;
        RECT -43.685 85.515 -43.355 85.845 ;
        RECT -43.685 84.155 -43.355 84.485 ;
        RECT -43.685 82.795 -43.355 83.125 ;
        RECT -43.685 81.435 -43.355 81.765 ;
        RECT -43.685 80.075 -43.355 80.405 ;
        RECT -43.685 78.715 -43.355 79.045 ;
        RECT -43.685 77.355 -43.355 77.685 ;
        RECT -43.685 75.995 -43.355 76.325 ;
        RECT -43.685 74.635 -43.355 74.965 ;
        RECT -43.685 73.275 -43.355 73.605 ;
        RECT -43.685 71.915 -43.355 72.245 ;
        RECT -43.685 70.555 -43.355 70.885 ;
        RECT -43.685 69.195 -43.355 69.525 ;
        RECT -43.685 67.835 -43.355 68.165 ;
        RECT -43.685 66.475 -43.355 66.805 ;
        RECT -43.685 65.115 -43.355 65.445 ;
        RECT -43.685 63.755 -43.355 64.085 ;
        RECT -43.685 62.395 -43.355 62.725 ;
        RECT -43.685 61.035 -43.355 61.365 ;
        RECT -43.685 59.675 -43.355 60.005 ;
        RECT -43.685 58.315 -43.355 58.645 ;
        RECT -43.685 56.955 -43.355 57.285 ;
        RECT -43.685 55.595 -43.355 55.925 ;
        RECT -43.685 54.235 -43.355 54.565 ;
        RECT -43.685 52.875 -43.355 53.205 ;
        RECT -43.685 51.515 -43.355 51.845 ;
        RECT -43.685 50.155 -43.355 50.485 ;
        RECT -43.685 48.795 -43.355 49.125 ;
        RECT -43.685 47.435 -43.355 47.765 ;
        RECT -43.685 46.075 -43.355 46.405 ;
        RECT -43.685 44.715 -43.355 45.045 ;
        RECT -43.685 43.355 -43.355 43.685 ;
        RECT -43.685 41.995 -43.355 42.325 ;
        RECT -43.685 40.635 -43.355 40.965 ;
        RECT -43.685 39.275 -43.355 39.605 ;
        RECT -43.685 37.915 -43.355 38.245 ;
        RECT -43.685 36.555 -43.355 36.885 ;
        RECT -43.685 35.195 -43.355 35.525 ;
        RECT -43.685 33.835 -43.355 34.165 ;
        RECT -43.685 32.475 -43.355 32.805 ;
        RECT -43.685 31.115 -43.355 31.445 ;
        RECT -43.685 29.755 -43.355 30.085 ;
        RECT -43.685 28.395 -43.355 28.725 ;
        RECT -43.685 27.035 -43.355 27.365 ;
        RECT -43.685 25.675 -43.355 26.005 ;
        RECT -43.685 24.315 -43.355 24.645 ;
        RECT -43.685 22.955 -43.355 23.285 ;
        RECT -43.685 21.595 -43.355 21.925 ;
        RECT -43.685 20.235 -43.355 20.565 ;
        RECT -43.685 18.875 -43.355 19.205 ;
        RECT -43.685 17.515 -43.355 17.845 ;
        RECT -43.685 16.155 -43.355 16.485 ;
        RECT -43.685 14.795 -43.355 15.125 ;
        RECT -43.685 13.435 -43.355 13.765 ;
        RECT -43.685 12.075 -43.355 12.405 ;
        RECT -43.685 10.715 -43.355 11.045 ;
        RECT -43.685 9.355 -43.355 9.685 ;
        RECT -43.685 7.995 -43.355 8.325 ;
        RECT -43.685 6.635 -43.355 6.965 ;
        RECT -43.685 5.275 -43.355 5.605 ;
        RECT -43.685 3.915 -43.355 4.245 ;
        RECT -43.685 2.555 -43.355 2.885 ;
        RECT -43.685 1.195 -43.355 1.525 ;
        RECT -43.685 -0.165 -43.355 0.165 ;
        RECT -43.685 -1.525 -43.355 -1.195 ;
        RECT -43.685 -4.245 -43.355 -3.915 ;
        RECT -43.685 -5.605 -43.355 -5.275 ;
        RECT -43.685 -6.965 -43.355 -6.635 ;
        RECT -43.685 -8.325 -43.355 -7.995 ;
        RECT -43.685 -9.685 -43.355 -9.355 ;
        RECT -43.685 -12.405 -43.355 -12.075 ;
        RECT -43.685 -13.765 -43.355 -13.435 ;
        RECT -43.685 -15.125 -43.355 -14.795 ;
        RECT -43.685 -16.485 -43.355 -16.155 ;
        RECT -43.685 -17.845 -43.355 -17.515 ;
        RECT -43.685 -19.205 -43.355 -18.875 ;
        RECT -43.685 -20.565 -43.355 -20.235 ;
        RECT -43.685 -21.925 -43.355 -21.595 ;
        RECT -43.685 -23.285 -43.355 -22.955 ;
        RECT -43.685 -30.66 -43.355 -30.33 ;
        RECT -43.685 -31.445 -43.355 -31.115 ;
        RECT -43.685 -32.805 -43.355 -32.475 ;
        RECT -43.685 -34.165 -43.355 -33.835 ;
        RECT -43.685 -36.885 -43.355 -36.555 ;
        RECT -43.685 -37.85 -43.355 -37.52 ;
        RECT -43.685 -40.965 -43.355 -40.635 ;
        RECT -43.685 -46.405 -43.355 -46.075 ;
        RECT -43.685 -49.125 -43.355 -48.795 ;
        RECT -43.685 -50.485 -43.355 -50.155 ;
        RECT -43.685 -53.205 -43.355 -52.875 ;
        RECT -43.685 -55.925 -43.355 -55.595 ;
        RECT -43.68 -58.64 -43.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 -129.365 -43.355 -129.035 ;
        RECT -43.685 -130.725 -43.355 -130.395 ;
        RECT -43.685 -131.47 -43.355 -131.14 ;
        RECT -43.685 -133.445 -43.355 -133.115 ;
        RECT -43.685 -134.805 -43.355 -134.475 ;
        RECT -43.685 -136.165 -43.355 -135.835 ;
        RECT -43.685 -137.525 -43.355 -137.195 ;
        RECT -43.685 -140.245 -43.355 -139.915 ;
        RECT -43.685 -141.605 -43.355 -141.275 ;
        RECT -43.685 -142.965 -43.355 -142.635 ;
        RECT -43.685 -144.31 -43.355 -143.98 ;
        RECT -43.685 -145.685 -43.355 -145.355 ;
        RECT -43.685 -147.045 -43.355 -146.715 ;
        RECT -43.685 -149.765 -43.355 -149.435 ;
        RECT -43.68 -152.48 -43.36 -124.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 -234.085 -43.355 -233.755 ;
        RECT -43.685 -235.445 -43.355 -235.115 ;
        RECT -43.685 -236.805 -43.355 -236.475 ;
        RECT -43.685 -238.165 -43.355 -237.835 ;
        RECT -43.685 -243.81 -43.355 -242.68 ;
        RECT -43.68 -243.925 -43.36 -231.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 246.76 -41.995 247.89 ;
        RECT -42.325 241.915 -41.995 242.245 ;
        RECT -42.325 240.555 -41.995 240.885 ;
        RECT -42.325 239.195 -41.995 239.525 ;
        RECT -42.325 237.835 -41.995 238.165 ;
        RECT -42.325 236.475 -41.995 236.805 ;
        RECT -42.325 235.115 -41.995 235.445 ;
        RECT -42.325 233.755 -41.995 234.085 ;
        RECT -42.325 232.395 -41.995 232.725 ;
        RECT -42.325 231.035 -41.995 231.365 ;
        RECT -42.325 229.675 -41.995 230.005 ;
        RECT -42.325 228.315 -41.995 228.645 ;
        RECT -42.325 226.955 -41.995 227.285 ;
        RECT -42.325 225.595 -41.995 225.925 ;
        RECT -42.325 224.235 -41.995 224.565 ;
        RECT -42.325 222.875 -41.995 223.205 ;
        RECT -42.325 221.515 -41.995 221.845 ;
        RECT -42.325 220.155 -41.995 220.485 ;
        RECT -42.325 218.795 -41.995 219.125 ;
        RECT -42.325 217.435 -41.995 217.765 ;
        RECT -42.325 216.075 -41.995 216.405 ;
        RECT -42.325 214.715 -41.995 215.045 ;
        RECT -42.325 213.355 -41.995 213.685 ;
        RECT -42.325 211.995 -41.995 212.325 ;
        RECT -42.325 210.635 -41.995 210.965 ;
        RECT -42.325 209.275 -41.995 209.605 ;
        RECT -42.325 207.915 -41.995 208.245 ;
        RECT -42.325 206.555 -41.995 206.885 ;
        RECT -42.325 205.195 -41.995 205.525 ;
        RECT -42.325 203.835 -41.995 204.165 ;
        RECT -42.325 202.475 -41.995 202.805 ;
        RECT -42.325 201.115 -41.995 201.445 ;
        RECT -42.325 199.755 -41.995 200.085 ;
        RECT -42.325 198.395 -41.995 198.725 ;
        RECT -42.325 197.035 -41.995 197.365 ;
        RECT -42.325 195.675 -41.995 196.005 ;
        RECT -42.325 194.315 -41.995 194.645 ;
        RECT -42.325 192.955 -41.995 193.285 ;
        RECT -42.325 191.595 -41.995 191.925 ;
        RECT -42.325 190.235 -41.995 190.565 ;
        RECT -42.325 188.875 -41.995 189.205 ;
        RECT -42.325 187.515 -41.995 187.845 ;
        RECT -42.325 186.155 -41.995 186.485 ;
        RECT -42.325 184.795 -41.995 185.125 ;
        RECT -42.325 183.435 -41.995 183.765 ;
        RECT -42.325 182.075 -41.995 182.405 ;
        RECT -42.325 180.715 -41.995 181.045 ;
        RECT -42.325 179.355 -41.995 179.685 ;
        RECT -42.325 177.995 -41.995 178.325 ;
        RECT -42.325 176.635 -41.995 176.965 ;
        RECT -42.325 175.275 -41.995 175.605 ;
        RECT -42.325 173.915 -41.995 174.245 ;
        RECT -42.325 172.555 -41.995 172.885 ;
        RECT -42.325 171.195 -41.995 171.525 ;
        RECT -42.325 169.835 -41.995 170.165 ;
        RECT -42.325 168.475 -41.995 168.805 ;
        RECT -42.325 167.115 -41.995 167.445 ;
        RECT -42.325 165.755 -41.995 166.085 ;
        RECT -42.325 164.395 -41.995 164.725 ;
        RECT -42.325 163.035 -41.995 163.365 ;
        RECT -42.325 161.675 -41.995 162.005 ;
        RECT -42.325 160.315 -41.995 160.645 ;
        RECT -42.325 158.955 -41.995 159.285 ;
        RECT -42.325 157.595 -41.995 157.925 ;
        RECT -42.325 156.235 -41.995 156.565 ;
        RECT -42.325 154.875 -41.995 155.205 ;
        RECT -42.325 153.515 -41.995 153.845 ;
        RECT -42.325 152.155 -41.995 152.485 ;
        RECT -42.325 150.795 -41.995 151.125 ;
        RECT -42.325 149.435 -41.995 149.765 ;
        RECT -42.325 148.075 -41.995 148.405 ;
        RECT -42.325 146.715 -41.995 147.045 ;
        RECT -42.325 145.355 -41.995 145.685 ;
        RECT -42.325 143.995 -41.995 144.325 ;
        RECT -42.325 142.635 -41.995 142.965 ;
        RECT -42.325 141.275 -41.995 141.605 ;
        RECT -42.325 139.915 -41.995 140.245 ;
        RECT -42.325 138.555 -41.995 138.885 ;
        RECT -42.325 137.195 -41.995 137.525 ;
        RECT -42.325 135.835 -41.995 136.165 ;
        RECT -42.325 134.475 -41.995 134.805 ;
        RECT -42.325 133.115 -41.995 133.445 ;
        RECT -42.325 131.755 -41.995 132.085 ;
        RECT -42.325 130.395 -41.995 130.725 ;
        RECT -42.325 129.035 -41.995 129.365 ;
        RECT -42.325 127.675 -41.995 128.005 ;
        RECT -42.325 126.315 -41.995 126.645 ;
        RECT -42.325 124.955 -41.995 125.285 ;
        RECT -42.325 123.595 -41.995 123.925 ;
        RECT -42.325 122.235 -41.995 122.565 ;
        RECT -42.325 120.875 -41.995 121.205 ;
        RECT -42.325 119.515 -41.995 119.845 ;
        RECT -42.325 118.155 -41.995 118.485 ;
        RECT -42.325 116.795 -41.995 117.125 ;
        RECT -42.325 115.435 -41.995 115.765 ;
        RECT -42.325 114.075 -41.995 114.405 ;
        RECT -42.325 112.715 -41.995 113.045 ;
        RECT -42.325 111.355 -41.995 111.685 ;
        RECT -42.325 109.995 -41.995 110.325 ;
        RECT -42.325 108.635 -41.995 108.965 ;
        RECT -42.325 107.275 -41.995 107.605 ;
        RECT -42.325 105.915 -41.995 106.245 ;
        RECT -42.325 104.555 -41.995 104.885 ;
        RECT -42.325 103.195 -41.995 103.525 ;
        RECT -42.325 101.835 -41.995 102.165 ;
        RECT -42.325 100.475 -41.995 100.805 ;
        RECT -42.325 99.115 -41.995 99.445 ;
        RECT -42.325 97.755 -41.995 98.085 ;
        RECT -42.325 96.395 -41.995 96.725 ;
        RECT -42.325 95.035 -41.995 95.365 ;
        RECT -42.325 93.675 -41.995 94.005 ;
        RECT -42.325 92.315 -41.995 92.645 ;
        RECT -42.325 90.955 -41.995 91.285 ;
        RECT -42.325 89.595 -41.995 89.925 ;
        RECT -42.325 88.235 -41.995 88.565 ;
        RECT -42.325 86.875 -41.995 87.205 ;
        RECT -42.325 85.515 -41.995 85.845 ;
        RECT -42.325 84.155 -41.995 84.485 ;
        RECT -42.325 82.795 -41.995 83.125 ;
        RECT -42.325 81.435 -41.995 81.765 ;
        RECT -42.325 80.075 -41.995 80.405 ;
        RECT -42.325 78.715 -41.995 79.045 ;
        RECT -42.325 77.355 -41.995 77.685 ;
        RECT -42.325 75.995 -41.995 76.325 ;
        RECT -42.325 74.635 -41.995 74.965 ;
        RECT -42.325 73.275 -41.995 73.605 ;
        RECT -42.325 71.915 -41.995 72.245 ;
        RECT -42.325 70.555 -41.995 70.885 ;
        RECT -42.325 69.195 -41.995 69.525 ;
        RECT -42.325 67.835 -41.995 68.165 ;
        RECT -42.325 66.475 -41.995 66.805 ;
        RECT -42.325 65.115 -41.995 65.445 ;
        RECT -42.325 63.755 -41.995 64.085 ;
        RECT -42.325 62.395 -41.995 62.725 ;
        RECT -42.325 61.035 -41.995 61.365 ;
        RECT -42.325 59.675 -41.995 60.005 ;
        RECT -42.325 58.315 -41.995 58.645 ;
        RECT -42.325 56.955 -41.995 57.285 ;
        RECT -42.325 55.595 -41.995 55.925 ;
        RECT -42.325 54.235 -41.995 54.565 ;
        RECT -42.325 52.875 -41.995 53.205 ;
        RECT -42.325 51.515 -41.995 51.845 ;
        RECT -42.325 50.155 -41.995 50.485 ;
        RECT -42.325 48.795 -41.995 49.125 ;
        RECT -42.325 47.435 -41.995 47.765 ;
        RECT -42.325 46.075 -41.995 46.405 ;
        RECT -42.325 44.715 -41.995 45.045 ;
        RECT -42.325 43.355 -41.995 43.685 ;
        RECT -42.325 41.995 -41.995 42.325 ;
        RECT -42.325 40.635 -41.995 40.965 ;
        RECT -42.325 39.275 -41.995 39.605 ;
        RECT -42.325 37.915 -41.995 38.245 ;
        RECT -42.325 36.555 -41.995 36.885 ;
        RECT -42.325 35.195 -41.995 35.525 ;
        RECT -42.325 33.835 -41.995 34.165 ;
        RECT -42.325 32.475 -41.995 32.805 ;
        RECT -42.325 31.115 -41.995 31.445 ;
        RECT -42.325 29.755 -41.995 30.085 ;
        RECT -42.325 28.395 -41.995 28.725 ;
        RECT -42.325 27.035 -41.995 27.365 ;
        RECT -42.325 25.675 -41.995 26.005 ;
        RECT -42.325 24.315 -41.995 24.645 ;
        RECT -42.325 22.955 -41.995 23.285 ;
        RECT -42.325 21.595 -41.995 21.925 ;
        RECT -42.325 20.235 -41.995 20.565 ;
        RECT -42.325 18.875 -41.995 19.205 ;
        RECT -42.325 17.515 -41.995 17.845 ;
        RECT -42.325 16.155 -41.995 16.485 ;
        RECT -42.325 14.795 -41.995 15.125 ;
        RECT -42.325 13.435 -41.995 13.765 ;
        RECT -42.325 12.075 -41.995 12.405 ;
        RECT -42.325 10.715 -41.995 11.045 ;
        RECT -42.325 9.355 -41.995 9.685 ;
        RECT -42.325 7.995 -41.995 8.325 ;
        RECT -42.325 6.635 -41.995 6.965 ;
        RECT -42.325 5.275 -41.995 5.605 ;
        RECT -42.325 3.915 -41.995 4.245 ;
        RECT -42.325 2.555 -41.995 2.885 ;
        RECT -42.325 1.195 -41.995 1.525 ;
        RECT -42.325 -0.165 -41.995 0.165 ;
        RECT -42.325 -1.525 -41.995 -1.195 ;
        RECT -42.32 -1.525 -42 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 -8.325 -41.995 -7.995 ;
        RECT -42.325 -9.685 -41.995 -9.355 ;
        RECT -42.325 -12.405 -41.995 -12.075 ;
        RECT -42.325 -13.765 -41.995 -13.435 ;
        RECT -42.325 -15.125 -41.995 -14.795 ;
        RECT -42.325 -16.485 -41.995 -16.155 ;
        RECT -42.325 -17.845 -41.995 -17.515 ;
        RECT -42.325 -19.205 -41.995 -18.875 ;
        RECT -42.325 -20.565 -41.995 -20.235 ;
        RECT -42.325 -21.925 -41.995 -21.595 ;
        RECT -42.325 -23.285 -41.995 -22.955 ;
        RECT -42.325 -30.66 -41.995 -30.33 ;
        RECT -42.325 -31.445 -41.995 -31.115 ;
        RECT -42.325 -32.805 -41.995 -32.475 ;
        RECT -42.325 -34.165 -41.995 -33.835 ;
        RECT -42.325 -36.885 -41.995 -36.555 ;
        RECT -42.325 -37.85 -41.995 -37.52 ;
        RECT -42.325 -40.965 -41.995 -40.635 ;
        RECT -42.325 -46.405 -41.995 -46.075 ;
        RECT -42.325 -49.125 -41.995 -48.795 ;
        RECT -42.325 -50.485 -41.995 -50.155 ;
        RECT -42.325 -53.205 -41.995 -52.875 ;
        RECT -42.325 -55.925 -41.995 -55.595 ;
        RECT -42.325 -61.365 -41.995 -61.035 ;
        RECT -42.325 -62.725 -41.995 -62.395 ;
        RECT -42.325 -64.085 -41.995 -63.755 ;
        RECT -42.325 -65.445 -41.995 -65.115 ;
        RECT -42.325 -66.805 -41.995 -66.475 ;
        RECT -42.325 -68.165 -41.995 -67.835 ;
        RECT -42.325 -69.525 -41.995 -69.195 ;
        RECT -42.325 -70.885 -41.995 -70.555 ;
        RECT -42.325 -72.245 -41.995 -71.915 ;
        RECT -42.325 -73.605 -41.995 -73.275 ;
        RECT -42.325 -74.965 -41.995 -74.635 ;
        RECT -42.325 -76.325 -41.995 -75.995 ;
        RECT -42.325 -77.685 -41.995 -77.355 ;
        RECT -42.325 -79.045 -41.995 -78.715 ;
        RECT -42.325 -80.405 -41.995 -80.075 ;
        RECT -42.325 -81.765 -41.995 -81.435 ;
        RECT -42.325 -83.125 -41.995 -82.795 ;
        RECT -42.325 -84.485 -41.995 -84.155 ;
        RECT -42.325 -85.845 -41.995 -85.515 ;
        RECT -42.325 -87.205 -41.995 -86.875 ;
        RECT -42.325 -88.565 -41.995 -88.235 ;
        RECT -42.325 -89.925 -41.995 -89.595 ;
        RECT -42.325 -91.285 -41.995 -90.955 ;
        RECT -42.325 -92.645 -41.995 -92.315 ;
        RECT -42.325 -94.005 -41.995 -93.675 ;
        RECT -42.325 -95.365 -41.995 -95.035 ;
        RECT -42.325 -96.725 -41.995 -96.395 ;
        RECT -42.325 -98.085 -41.995 -97.755 ;
        RECT -42.325 -99.445 -41.995 -99.115 ;
        RECT -42.325 -100.805 -41.995 -100.475 ;
        RECT -42.325 -102.165 -41.995 -101.835 ;
        RECT -42.325 -103.525 -41.995 -103.195 ;
        RECT -42.325 -104.885 -41.995 -104.555 ;
        RECT -42.325 -106.245 -41.995 -105.915 ;
        RECT -42.325 -107.605 -41.995 -107.275 ;
        RECT -42.325 -108.965 -41.995 -108.635 ;
        RECT -42.325 -110.325 -41.995 -109.995 ;
        RECT -42.325 -111.685 -41.995 -111.355 ;
        RECT -42.325 -113.045 -41.995 -112.715 ;
        RECT -42.325 -114.405 -41.995 -114.075 ;
        RECT -42.325 -115.765 -41.995 -115.435 ;
        RECT -42.325 -117.125 -41.995 -116.795 ;
        RECT -42.325 -118.485 -41.995 -118.155 ;
        RECT -42.325 -119.845 -41.995 -119.515 ;
        RECT -42.325 -121.205 -41.995 -120.875 ;
        RECT -42.325 -123.925 -41.995 -123.595 ;
        RECT -42.325 -129.365 -41.995 -129.035 ;
        RECT -42.325 -130.725 -41.995 -130.395 ;
        RECT -42.325 -131.47 -41.995 -131.14 ;
        RECT -42.325 -133.445 -41.995 -133.115 ;
        RECT -42.325 -134.805 -41.995 -134.475 ;
        RECT -42.325 -136.165 -41.995 -135.835 ;
        RECT -42.325 -137.525 -41.995 -137.195 ;
        RECT -42.325 -140.245 -41.995 -139.915 ;
        RECT -42.325 -141.605 -41.995 -141.275 ;
        RECT -42.325 -142.965 -41.995 -142.635 ;
        RECT -42.325 -144.31 -41.995 -143.98 ;
        RECT -42.325 -145.685 -41.995 -145.355 ;
        RECT -42.325 -147.045 -41.995 -146.715 ;
        RECT -42.325 -149.765 -41.995 -149.435 ;
        RECT -42.325 -153.845 -41.995 -153.515 ;
        RECT -42.325 -155.205 -41.995 -154.875 ;
        RECT -42.325 -156.565 -41.995 -156.235 ;
        RECT -42.325 -157.925 -41.995 -157.595 ;
        RECT -42.325 -159.285 -41.995 -158.955 ;
        RECT -42.325 -162.005 -41.995 -161.675 ;
        RECT -42.325 -163.365 -41.995 -163.035 ;
        RECT -42.325 -164.725 -41.995 -164.395 ;
        RECT -42.325 -166.085 -41.995 -165.755 ;
        RECT -42.325 -167.445 -41.995 -167.115 ;
        RECT -42.325 -168.805 -41.995 -168.475 ;
        RECT -42.325 -170.165 -41.995 -169.835 ;
        RECT -42.325 -171.525 -41.995 -171.195 ;
        RECT -42.325 -172.885 -41.995 -172.555 ;
        RECT -42.325 -174.245 -41.995 -173.915 ;
        RECT -42.325 -175.605 -41.995 -175.275 ;
        RECT -42.325 -176.965 -41.995 -176.635 ;
        RECT -42.325 -178.325 -41.995 -177.995 ;
        RECT -42.325 -179.685 -41.995 -179.355 ;
        RECT -42.325 -181.045 -41.995 -180.715 ;
        RECT -42.325 -182.405 -41.995 -182.075 ;
        RECT -42.325 -183.765 -41.995 -183.435 ;
        RECT -42.325 -185.125 -41.995 -184.795 ;
        RECT -42.325 -186.485 -41.995 -186.155 ;
        RECT -42.325 -187.845 -41.995 -187.515 ;
        RECT -42.325 -189.205 -41.995 -188.875 ;
        RECT -42.325 -190.565 -41.995 -190.235 ;
        RECT -42.325 -191.925 -41.995 -191.595 ;
        RECT -42.325 -193.285 -41.995 -192.955 ;
        RECT -42.325 -194.645 -41.995 -194.315 ;
        RECT -42.325 -196.005 -41.995 -195.675 ;
        RECT -42.325 -197.365 -41.995 -197.035 ;
        RECT -42.325 -198.725 -41.995 -198.395 ;
        RECT -42.325 -200.085 -41.995 -199.755 ;
        RECT -42.325 -201.445 -41.995 -201.115 ;
        RECT -42.325 -202.805 -41.995 -202.475 ;
        RECT -42.325 -204.165 -41.995 -203.835 ;
        RECT -42.325 -205.525 -41.995 -205.195 ;
        RECT -42.325 -206.885 -41.995 -206.555 ;
        RECT -42.325 -208.245 -41.995 -207.915 ;
        RECT -42.325 -209.605 -41.995 -209.275 ;
        RECT -42.325 -210.965 -41.995 -210.635 ;
        RECT -42.325 -212.325 -41.995 -211.995 ;
        RECT -42.325 -213.685 -41.995 -213.355 ;
        RECT -42.325 -215.045 -41.995 -214.715 ;
        RECT -42.325 -216.405 -41.995 -216.075 ;
        RECT -42.325 -217.765 -41.995 -217.435 ;
        RECT -42.325 -219.125 -41.995 -218.795 ;
        RECT -42.325 -220.485 -41.995 -220.155 ;
        RECT -42.325 -221.845 -41.995 -221.515 ;
        RECT -42.325 -223.205 -41.995 -222.875 ;
        RECT -42.325 -224.565 -41.995 -224.235 ;
        RECT -42.325 -226.155 -41.995 -225.825 ;
        RECT -42.325 -227.285 -41.995 -226.955 ;
        RECT -42.325 -228.645 -41.995 -228.315 ;
        RECT -42.325 -234.085 -41.995 -233.755 ;
        RECT -42.325 -235.445 -41.995 -235.115 ;
        RECT -42.325 -236.805 -41.995 -236.475 ;
        RECT -42.325 -238.165 -41.995 -237.835 ;
        RECT -42.325 -243.81 -41.995 -242.68 ;
        RECT -42.32 -243.925 -42 -7.32 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.965 246.76 -40.635 247.89 ;
        RECT -40.965 241.915 -40.635 242.245 ;
        RECT -40.965 240.555 -40.635 240.885 ;
        RECT -40.965 239.195 -40.635 239.525 ;
        RECT -40.965 237.835 -40.635 238.165 ;
        RECT -40.965 236.475 -40.635 236.805 ;
        RECT -40.965 235.115 -40.635 235.445 ;
        RECT -40.965 233.755 -40.635 234.085 ;
        RECT -40.965 232.395 -40.635 232.725 ;
        RECT -40.965 231.035 -40.635 231.365 ;
        RECT -40.965 229.675 -40.635 230.005 ;
        RECT -40.965 228.315 -40.635 228.645 ;
        RECT -40.965 226.955 -40.635 227.285 ;
        RECT -40.965 225.595 -40.635 225.925 ;
        RECT -40.965 224.235 -40.635 224.565 ;
        RECT -40.965 222.875 -40.635 223.205 ;
        RECT -40.965 221.515 -40.635 221.845 ;
        RECT -40.965 220.155 -40.635 220.485 ;
        RECT -40.965 218.795 -40.635 219.125 ;
        RECT -40.965 217.435 -40.635 217.765 ;
        RECT -40.965 216.075 -40.635 216.405 ;
        RECT -40.965 214.715 -40.635 215.045 ;
        RECT -40.965 213.355 -40.635 213.685 ;
        RECT -40.965 211.995 -40.635 212.325 ;
        RECT -40.965 210.635 -40.635 210.965 ;
        RECT -40.965 209.275 -40.635 209.605 ;
        RECT -40.965 207.915 -40.635 208.245 ;
        RECT -40.965 206.555 -40.635 206.885 ;
        RECT -40.965 205.195 -40.635 205.525 ;
        RECT -40.965 203.835 -40.635 204.165 ;
        RECT -40.965 202.475 -40.635 202.805 ;
        RECT -40.965 201.115 -40.635 201.445 ;
        RECT -40.965 199.755 -40.635 200.085 ;
        RECT -40.965 198.395 -40.635 198.725 ;
        RECT -40.965 197.035 -40.635 197.365 ;
        RECT -40.965 195.675 -40.635 196.005 ;
        RECT -40.965 194.315 -40.635 194.645 ;
        RECT -40.965 192.955 -40.635 193.285 ;
        RECT -40.965 191.595 -40.635 191.925 ;
        RECT -40.965 190.235 -40.635 190.565 ;
        RECT -40.965 188.875 -40.635 189.205 ;
        RECT -40.965 187.515 -40.635 187.845 ;
        RECT -40.965 186.155 -40.635 186.485 ;
        RECT -40.965 184.795 -40.635 185.125 ;
        RECT -40.965 183.435 -40.635 183.765 ;
        RECT -40.965 182.075 -40.635 182.405 ;
        RECT -40.965 180.715 -40.635 181.045 ;
        RECT -40.965 179.355 -40.635 179.685 ;
        RECT -40.965 177.995 -40.635 178.325 ;
        RECT -40.965 176.635 -40.635 176.965 ;
        RECT -40.965 175.275 -40.635 175.605 ;
        RECT -40.965 173.915 -40.635 174.245 ;
        RECT -40.965 172.555 -40.635 172.885 ;
        RECT -40.965 171.195 -40.635 171.525 ;
        RECT -40.965 169.835 -40.635 170.165 ;
        RECT -40.965 168.475 -40.635 168.805 ;
        RECT -40.965 167.115 -40.635 167.445 ;
        RECT -40.965 165.755 -40.635 166.085 ;
        RECT -40.965 164.395 -40.635 164.725 ;
        RECT -40.965 163.035 -40.635 163.365 ;
        RECT -40.965 161.675 -40.635 162.005 ;
        RECT -40.965 160.315 -40.635 160.645 ;
        RECT -40.965 158.955 -40.635 159.285 ;
        RECT -40.965 157.595 -40.635 157.925 ;
        RECT -40.965 156.235 -40.635 156.565 ;
        RECT -40.965 154.875 -40.635 155.205 ;
        RECT -40.965 153.515 -40.635 153.845 ;
        RECT -40.965 152.155 -40.635 152.485 ;
        RECT -40.965 150.795 -40.635 151.125 ;
        RECT -40.965 149.435 -40.635 149.765 ;
        RECT -40.965 148.075 -40.635 148.405 ;
        RECT -40.965 146.715 -40.635 147.045 ;
        RECT -40.965 145.355 -40.635 145.685 ;
        RECT -40.965 143.995 -40.635 144.325 ;
        RECT -40.965 142.635 -40.635 142.965 ;
        RECT -40.965 141.275 -40.635 141.605 ;
        RECT -40.965 139.915 -40.635 140.245 ;
        RECT -40.965 138.555 -40.635 138.885 ;
        RECT -40.965 137.195 -40.635 137.525 ;
        RECT -40.965 135.835 -40.635 136.165 ;
        RECT -40.965 134.475 -40.635 134.805 ;
        RECT -40.965 133.115 -40.635 133.445 ;
        RECT -40.965 131.755 -40.635 132.085 ;
        RECT -40.965 130.395 -40.635 130.725 ;
        RECT -40.965 129.035 -40.635 129.365 ;
        RECT -40.965 127.675 -40.635 128.005 ;
        RECT -40.965 126.315 -40.635 126.645 ;
        RECT -40.965 124.955 -40.635 125.285 ;
        RECT -40.965 123.595 -40.635 123.925 ;
        RECT -40.965 122.235 -40.635 122.565 ;
        RECT -40.965 120.875 -40.635 121.205 ;
        RECT -40.965 119.515 -40.635 119.845 ;
        RECT -40.965 118.155 -40.635 118.485 ;
        RECT -40.965 116.795 -40.635 117.125 ;
        RECT -40.965 115.435 -40.635 115.765 ;
        RECT -40.965 114.075 -40.635 114.405 ;
        RECT -40.965 112.715 -40.635 113.045 ;
        RECT -40.965 111.355 -40.635 111.685 ;
        RECT -40.965 109.995 -40.635 110.325 ;
        RECT -40.965 108.635 -40.635 108.965 ;
        RECT -40.965 107.275 -40.635 107.605 ;
        RECT -40.965 105.915 -40.635 106.245 ;
        RECT -40.965 104.555 -40.635 104.885 ;
        RECT -40.965 103.195 -40.635 103.525 ;
        RECT -40.965 101.835 -40.635 102.165 ;
        RECT -40.965 100.475 -40.635 100.805 ;
        RECT -40.965 99.115 -40.635 99.445 ;
        RECT -40.965 97.755 -40.635 98.085 ;
        RECT -40.965 96.395 -40.635 96.725 ;
        RECT -40.965 95.035 -40.635 95.365 ;
        RECT -40.965 93.675 -40.635 94.005 ;
        RECT -40.965 92.315 -40.635 92.645 ;
        RECT -40.965 90.955 -40.635 91.285 ;
        RECT -40.965 89.595 -40.635 89.925 ;
        RECT -40.965 88.235 -40.635 88.565 ;
        RECT -40.965 86.875 -40.635 87.205 ;
        RECT -40.965 85.515 -40.635 85.845 ;
        RECT -40.965 84.155 -40.635 84.485 ;
        RECT -40.965 82.795 -40.635 83.125 ;
        RECT -40.965 81.435 -40.635 81.765 ;
        RECT -40.965 80.075 -40.635 80.405 ;
        RECT -40.965 78.715 -40.635 79.045 ;
        RECT -40.965 77.355 -40.635 77.685 ;
        RECT -40.965 75.995 -40.635 76.325 ;
        RECT -40.965 74.635 -40.635 74.965 ;
        RECT -40.965 73.275 -40.635 73.605 ;
        RECT -40.965 71.915 -40.635 72.245 ;
        RECT -40.965 70.555 -40.635 70.885 ;
        RECT -40.965 69.195 -40.635 69.525 ;
        RECT -40.965 67.835 -40.635 68.165 ;
        RECT -40.965 66.475 -40.635 66.805 ;
        RECT -40.965 65.115 -40.635 65.445 ;
        RECT -40.965 63.755 -40.635 64.085 ;
        RECT -40.965 62.395 -40.635 62.725 ;
        RECT -40.965 61.035 -40.635 61.365 ;
        RECT -40.965 59.675 -40.635 60.005 ;
        RECT -40.965 58.315 -40.635 58.645 ;
        RECT -40.965 56.955 -40.635 57.285 ;
        RECT -40.965 55.595 -40.635 55.925 ;
        RECT -40.965 54.235 -40.635 54.565 ;
        RECT -40.965 52.875 -40.635 53.205 ;
        RECT -40.965 51.515 -40.635 51.845 ;
        RECT -40.965 50.155 -40.635 50.485 ;
        RECT -40.965 48.795 -40.635 49.125 ;
        RECT -40.965 47.435 -40.635 47.765 ;
        RECT -40.965 46.075 -40.635 46.405 ;
        RECT -40.965 44.715 -40.635 45.045 ;
        RECT -40.965 43.355 -40.635 43.685 ;
        RECT -40.965 41.995 -40.635 42.325 ;
        RECT -40.965 40.635 -40.635 40.965 ;
        RECT -40.965 39.275 -40.635 39.605 ;
        RECT -40.965 37.915 -40.635 38.245 ;
        RECT -40.965 36.555 -40.635 36.885 ;
        RECT -40.965 35.195 -40.635 35.525 ;
        RECT -40.965 33.835 -40.635 34.165 ;
        RECT -40.965 32.475 -40.635 32.805 ;
        RECT -40.965 31.115 -40.635 31.445 ;
        RECT -40.965 29.755 -40.635 30.085 ;
        RECT -40.965 28.395 -40.635 28.725 ;
        RECT -40.965 27.035 -40.635 27.365 ;
        RECT -40.965 25.675 -40.635 26.005 ;
        RECT -40.965 24.315 -40.635 24.645 ;
        RECT -40.965 22.955 -40.635 23.285 ;
        RECT -40.965 21.595 -40.635 21.925 ;
        RECT -40.965 20.235 -40.635 20.565 ;
        RECT -40.965 18.875 -40.635 19.205 ;
        RECT -40.965 17.515 -40.635 17.845 ;
        RECT -40.965 16.155 -40.635 16.485 ;
        RECT -40.965 14.795 -40.635 15.125 ;
        RECT -40.965 13.435 -40.635 13.765 ;
        RECT -40.965 12.075 -40.635 12.405 ;
        RECT -40.965 10.715 -40.635 11.045 ;
        RECT -40.965 9.355 -40.635 9.685 ;
        RECT -40.965 7.995 -40.635 8.325 ;
        RECT -40.965 6.635 -40.635 6.965 ;
        RECT -40.965 5.275 -40.635 5.605 ;
        RECT -40.965 3.915 -40.635 4.245 ;
        RECT -40.965 2.555 -40.635 2.885 ;
        RECT -40.965 1.195 -40.635 1.525 ;
        RECT -40.965 -0.165 -40.635 0.165 ;
        RECT -40.965 -1.525 -40.635 -1.195 ;
        RECT -40.965 -5.605 -40.635 -5.275 ;
        RECT -40.965 -8.325 -40.635 -7.995 ;
        RECT -40.965 -9.685 -40.635 -9.355 ;
        RECT -40.965 -12.405 -40.635 -12.075 ;
        RECT -40.965 -13.765 -40.635 -13.435 ;
        RECT -40.965 -15.125 -40.635 -14.795 ;
        RECT -40.965 -16.485 -40.635 -16.155 ;
        RECT -40.965 -17.845 -40.635 -17.515 ;
        RECT -40.965 -19.205 -40.635 -18.875 ;
        RECT -40.965 -20.565 -40.635 -20.235 ;
        RECT -40.965 -21.925 -40.635 -21.595 ;
        RECT -40.965 -23.285 -40.635 -22.955 ;
        RECT -40.965 -30.66 -40.635 -30.33 ;
        RECT -40.965 -31.445 -40.635 -31.115 ;
        RECT -40.965 -32.805 -40.635 -32.475 ;
        RECT -40.965 -34.165 -40.635 -33.835 ;
        RECT -40.965 -36.885 -40.635 -36.555 ;
        RECT -40.965 -37.85 -40.635 -37.52 ;
        RECT -40.965 -40.965 -40.635 -40.635 ;
        RECT -40.965 -46.405 -40.635 -46.075 ;
        RECT -40.965 -49.125 -40.635 -48.795 ;
        RECT -40.965 -50.485 -40.635 -50.155 ;
        RECT -40.965 -53.205 -40.635 -52.875 ;
        RECT -40.965 -55.925 -40.635 -55.595 ;
        RECT -40.965 -61.365 -40.635 -61.035 ;
        RECT -40.965 -62.725 -40.635 -62.395 ;
        RECT -40.965 -64.085 -40.635 -63.755 ;
        RECT -40.965 -65.445 -40.635 -65.115 ;
        RECT -40.965 -66.805 -40.635 -66.475 ;
        RECT -40.965 -68.165 -40.635 -67.835 ;
        RECT -40.965 -69.525 -40.635 -69.195 ;
        RECT -40.965 -70.885 -40.635 -70.555 ;
        RECT -40.965 -72.245 -40.635 -71.915 ;
        RECT -40.965 -73.605 -40.635 -73.275 ;
        RECT -40.965 -74.965 -40.635 -74.635 ;
        RECT -40.965 -76.325 -40.635 -75.995 ;
        RECT -40.965 -77.685 -40.635 -77.355 ;
        RECT -40.965 -79.045 -40.635 -78.715 ;
        RECT -40.965 -80.405 -40.635 -80.075 ;
        RECT -40.965 -81.765 -40.635 -81.435 ;
        RECT -40.965 -83.125 -40.635 -82.795 ;
        RECT -40.965 -84.485 -40.635 -84.155 ;
        RECT -40.965 -85.845 -40.635 -85.515 ;
        RECT -40.965 -87.205 -40.635 -86.875 ;
        RECT -40.965 -88.565 -40.635 -88.235 ;
        RECT -40.965 -89.925 -40.635 -89.595 ;
        RECT -40.965 -91.285 -40.635 -90.955 ;
        RECT -40.965 -92.645 -40.635 -92.315 ;
        RECT -40.965 -94.005 -40.635 -93.675 ;
        RECT -40.965 -95.365 -40.635 -95.035 ;
        RECT -40.965 -96.725 -40.635 -96.395 ;
        RECT -40.965 -98.085 -40.635 -97.755 ;
        RECT -40.965 -99.445 -40.635 -99.115 ;
        RECT -40.965 -100.805 -40.635 -100.475 ;
        RECT -40.965 -102.165 -40.635 -101.835 ;
        RECT -40.965 -103.525 -40.635 -103.195 ;
        RECT -40.965 -104.885 -40.635 -104.555 ;
        RECT -40.965 -106.245 -40.635 -105.915 ;
        RECT -40.965 -107.605 -40.635 -107.275 ;
        RECT -40.965 -108.965 -40.635 -108.635 ;
        RECT -40.965 -110.325 -40.635 -109.995 ;
        RECT -40.965 -111.685 -40.635 -111.355 ;
        RECT -40.965 -113.045 -40.635 -112.715 ;
        RECT -40.965 -114.405 -40.635 -114.075 ;
        RECT -40.965 -115.765 -40.635 -115.435 ;
        RECT -40.965 -117.125 -40.635 -116.795 ;
        RECT -40.965 -118.485 -40.635 -118.155 ;
        RECT -40.965 -119.845 -40.635 -119.515 ;
        RECT -40.965 -121.205 -40.635 -120.875 ;
        RECT -40.965 -123.925 -40.635 -123.595 ;
        RECT -40.965 -129.365 -40.635 -129.035 ;
        RECT -40.965 -130.725 -40.635 -130.395 ;
        RECT -40.965 -131.47 -40.635 -131.14 ;
        RECT -40.965 -133.445 -40.635 -133.115 ;
        RECT -40.965 -134.805 -40.635 -134.475 ;
        RECT -40.965 -136.165 -40.635 -135.835 ;
        RECT -40.965 -137.525 -40.635 -137.195 ;
        RECT -40.965 -140.245 -40.635 -139.915 ;
        RECT -40.965 -141.605 -40.635 -141.275 ;
        RECT -40.965 -142.965 -40.635 -142.635 ;
        RECT -40.965 -144.31 -40.635 -143.98 ;
        RECT -40.965 -145.685 -40.635 -145.355 ;
        RECT -40.965 -147.045 -40.635 -146.715 ;
        RECT -40.965 -149.765 -40.635 -149.435 ;
        RECT -40.965 -152.485 -40.635 -152.155 ;
        RECT -40.965 -153.845 -40.635 -153.515 ;
        RECT -40.965 -155.205 -40.635 -154.875 ;
        RECT -40.965 -156.565 -40.635 -156.235 ;
        RECT -40.965 -157.925 -40.635 -157.595 ;
        RECT -40.965 -159.285 -40.635 -158.955 ;
        RECT -40.965 -162.005 -40.635 -161.675 ;
        RECT -40.965 -163.365 -40.635 -163.035 ;
        RECT -40.965 -164.725 -40.635 -164.395 ;
        RECT -40.965 -166.085 -40.635 -165.755 ;
        RECT -40.965 -167.445 -40.635 -167.115 ;
        RECT -40.965 -168.805 -40.635 -168.475 ;
        RECT -40.965 -170.165 -40.635 -169.835 ;
        RECT -40.965 -171.525 -40.635 -171.195 ;
        RECT -40.965 -172.885 -40.635 -172.555 ;
        RECT -40.965 -174.245 -40.635 -173.915 ;
        RECT -40.965 -175.605 -40.635 -175.275 ;
        RECT -40.965 -176.965 -40.635 -176.635 ;
        RECT -40.965 -178.325 -40.635 -177.995 ;
        RECT -40.965 -179.685 -40.635 -179.355 ;
        RECT -40.965 -181.045 -40.635 -180.715 ;
        RECT -40.965 -182.405 -40.635 -182.075 ;
        RECT -40.965 -183.765 -40.635 -183.435 ;
        RECT -40.965 -185.125 -40.635 -184.795 ;
        RECT -40.965 -186.485 -40.635 -186.155 ;
        RECT -40.965 -187.845 -40.635 -187.515 ;
        RECT -40.965 -189.205 -40.635 -188.875 ;
        RECT -40.965 -190.565 -40.635 -190.235 ;
        RECT -40.965 -191.925 -40.635 -191.595 ;
        RECT -40.965 -193.285 -40.635 -192.955 ;
        RECT -40.965 -194.645 -40.635 -194.315 ;
        RECT -40.965 -196.005 -40.635 -195.675 ;
        RECT -40.965 -197.365 -40.635 -197.035 ;
        RECT -40.965 -198.725 -40.635 -198.395 ;
        RECT -40.965 -200.085 -40.635 -199.755 ;
        RECT -40.965 -201.445 -40.635 -201.115 ;
        RECT -40.965 -202.805 -40.635 -202.475 ;
        RECT -40.965 -204.165 -40.635 -203.835 ;
        RECT -40.965 -205.525 -40.635 -205.195 ;
        RECT -40.965 -206.885 -40.635 -206.555 ;
        RECT -40.965 -208.245 -40.635 -207.915 ;
        RECT -40.965 -209.605 -40.635 -209.275 ;
        RECT -40.965 -210.965 -40.635 -210.635 ;
        RECT -40.965 -212.325 -40.635 -211.995 ;
        RECT -40.965 -213.685 -40.635 -213.355 ;
        RECT -40.965 -215.045 -40.635 -214.715 ;
        RECT -40.965 -216.405 -40.635 -216.075 ;
        RECT -40.965 -217.765 -40.635 -217.435 ;
        RECT -40.965 -219.125 -40.635 -218.795 ;
        RECT -40.965 -220.485 -40.635 -220.155 ;
        RECT -40.965 -221.845 -40.635 -221.515 ;
        RECT -40.965 -223.205 -40.635 -222.875 ;
        RECT -40.965 -224.565 -40.635 -224.235 ;
        RECT -40.965 -226.155 -40.635 -225.825 ;
        RECT -40.965 -227.285 -40.635 -226.955 ;
        RECT -40.965 -228.645 -40.635 -228.315 ;
        RECT -40.965 -231.365 -40.635 -231.035 ;
        RECT -40.965 -234.085 -40.635 -233.755 ;
        RECT -40.965 -235.445 -40.635 -235.115 ;
        RECT -40.965 -236.805 -40.635 -236.475 ;
        RECT -40.965 -238.165 -40.635 -237.835 ;
        RECT -40.965 -243.81 -40.635 -242.68 ;
        RECT -40.96 -243.925 -40.64 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.605 -200.085 -39.275 -199.755 ;
        RECT -39.605 -201.445 -39.275 -201.115 ;
        RECT -39.605 -202.805 -39.275 -202.475 ;
        RECT -39.605 -204.165 -39.275 -203.835 ;
        RECT -39.605 -205.525 -39.275 -205.195 ;
        RECT -39.605 -206.885 -39.275 -206.555 ;
        RECT -39.605 -208.245 -39.275 -207.915 ;
        RECT -39.605 -209.605 -39.275 -209.275 ;
        RECT -39.605 -210.965 -39.275 -210.635 ;
        RECT -39.605 -212.325 -39.275 -211.995 ;
        RECT -39.605 -213.685 -39.275 -213.355 ;
        RECT -39.605 -215.045 -39.275 -214.715 ;
        RECT -39.605 -216.405 -39.275 -216.075 ;
        RECT -39.605 -217.765 -39.275 -217.435 ;
        RECT -39.605 -219.125 -39.275 -218.795 ;
        RECT -39.605 -220.485 -39.275 -220.155 ;
        RECT -39.605 -221.845 -39.275 -221.515 ;
        RECT -39.605 -223.205 -39.275 -222.875 ;
        RECT -39.605 -224.565 -39.275 -224.235 ;
        RECT -39.605 -226.155 -39.275 -225.825 ;
        RECT -39.605 -227.285 -39.275 -226.955 ;
        RECT -39.605 -228.645 -39.275 -228.315 ;
        RECT -39.605 -231.365 -39.275 -231.035 ;
        RECT -39.605 -234.085 -39.275 -233.755 ;
        RECT -39.605 -235.445 -39.275 -235.115 ;
        RECT -39.605 -236.805 -39.275 -236.475 ;
        RECT -39.605 -238.165 -39.275 -237.835 ;
        RECT -39.605 -243.81 -39.275 -242.68 ;
        RECT -39.6 -243.925 -39.28 248.005 ;
        RECT -39.605 246.76 -39.275 247.89 ;
        RECT -39.605 241.915 -39.275 242.245 ;
        RECT -39.605 240.555 -39.275 240.885 ;
        RECT -39.605 239.195 -39.275 239.525 ;
        RECT -39.605 237.835 -39.275 238.165 ;
        RECT -39.605 236.475 -39.275 236.805 ;
        RECT -39.605 235.115 -39.275 235.445 ;
        RECT -39.605 233.755 -39.275 234.085 ;
        RECT -39.605 232.395 -39.275 232.725 ;
        RECT -39.605 231.035 -39.275 231.365 ;
        RECT -39.605 229.675 -39.275 230.005 ;
        RECT -39.605 228.315 -39.275 228.645 ;
        RECT -39.605 226.955 -39.275 227.285 ;
        RECT -39.605 225.595 -39.275 225.925 ;
        RECT -39.605 224.235 -39.275 224.565 ;
        RECT -39.605 222.875 -39.275 223.205 ;
        RECT -39.605 221.515 -39.275 221.845 ;
        RECT -39.605 220.155 -39.275 220.485 ;
        RECT -39.605 218.795 -39.275 219.125 ;
        RECT -39.605 217.435 -39.275 217.765 ;
        RECT -39.605 216.075 -39.275 216.405 ;
        RECT -39.605 214.715 -39.275 215.045 ;
        RECT -39.605 213.355 -39.275 213.685 ;
        RECT -39.605 211.995 -39.275 212.325 ;
        RECT -39.605 210.635 -39.275 210.965 ;
        RECT -39.605 209.275 -39.275 209.605 ;
        RECT -39.605 207.915 -39.275 208.245 ;
        RECT -39.605 206.555 -39.275 206.885 ;
        RECT -39.605 205.195 -39.275 205.525 ;
        RECT -39.605 203.835 -39.275 204.165 ;
        RECT -39.605 202.475 -39.275 202.805 ;
        RECT -39.605 201.115 -39.275 201.445 ;
        RECT -39.605 199.755 -39.275 200.085 ;
        RECT -39.605 198.395 -39.275 198.725 ;
        RECT -39.605 197.035 -39.275 197.365 ;
        RECT -39.605 195.675 -39.275 196.005 ;
        RECT -39.605 194.315 -39.275 194.645 ;
        RECT -39.605 192.955 -39.275 193.285 ;
        RECT -39.605 191.595 -39.275 191.925 ;
        RECT -39.605 190.235 -39.275 190.565 ;
        RECT -39.605 188.875 -39.275 189.205 ;
        RECT -39.605 187.515 -39.275 187.845 ;
        RECT -39.605 186.155 -39.275 186.485 ;
        RECT -39.605 184.795 -39.275 185.125 ;
        RECT -39.605 183.435 -39.275 183.765 ;
        RECT -39.605 182.075 -39.275 182.405 ;
        RECT -39.605 180.715 -39.275 181.045 ;
        RECT -39.605 179.355 -39.275 179.685 ;
        RECT -39.605 177.995 -39.275 178.325 ;
        RECT -39.605 176.635 -39.275 176.965 ;
        RECT -39.605 175.275 -39.275 175.605 ;
        RECT -39.605 173.915 -39.275 174.245 ;
        RECT -39.605 172.555 -39.275 172.885 ;
        RECT -39.605 171.195 -39.275 171.525 ;
        RECT -39.605 169.835 -39.275 170.165 ;
        RECT -39.605 168.475 -39.275 168.805 ;
        RECT -39.605 167.115 -39.275 167.445 ;
        RECT -39.605 165.755 -39.275 166.085 ;
        RECT -39.605 164.395 -39.275 164.725 ;
        RECT -39.605 163.035 -39.275 163.365 ;
        RECT -39.605 161.675 -39.275 162.005 ;
        RECT -39.605 160.315 -39.275 160.645 ;
        RECT -39.605 158.955 -39.275 159.285 ;
        RECT -39.605 157.595 -39.275 157.925 ;
        RECT -39.605 156.235 -39.275 156.565 ;
        RECT -39.605 154.875 -39.275 155.205 ;
        RECT -39.605 153.515 -39.275 153.845 ;
        RECT -39.605 152.155 -39.275 152.485 ;
        RECT -39.605 150.795 -39.275 151.125 ;
        RECT -39.605 149.435 -39.275 149.765 ;
        RECT -39.605 148.075 -39.275 148.405 ;
        RECT -39.605 146.715 -39.275 147.045 ;
        RECT -39.605 145.355 -39.275 145.685 ;
        RECT -39.605 143.995 -39.275 144.325 ;
        RECT -39.605 142.635 -39.275 142.965 ;
        RECT -39.605 141.275 -39.275 141.605 ;
        RECT -39.605 139.915 -39.275 140.245 ;
        RECT -39.605 138.555 -39.275 138.885 ;
        RECT -39.605 137.195 -39.275 137.525 ;
        RECT -39.605 135.835 -39.275 136.165 ;
        RECT -39.605 134.475 -39.275 134.805 ;
        RECT -39.605 133.115 -39.275 133.445 ;
        RECT -39.605 131.755 -39.275 132.085 ;
        RECT -39.605 130.395 -39.275 130.725 ;
        RECT -39.605 129.035 -39.275 129.365 ;
        RECT -39.605 127.675 -39.275 128.005 ;
        RECT -39.605 126.315 -39.275 126.645 ;
        RECT -39.605 124.955 -39.275 125.285 ;
        RECT -39.605 123.595 -39.275 123.925 ;
        RECT -39.605 122.235 -39.275 122.565 ;
        RECT -39.605 120.875 -39.275 121.205 ;
        RECT -39.605 119.515 -39.275 119.845 ;
        RECT -39.605 118.155 -39.275 118.485 ;
        RECT -39.605 116.795 -39.275 117.125 ;
        RECT -39.605 115.435 -39.275 115.765 ;
        RECT -39.605 114.075 -39.275 114.405 ;
        RECT -39.605 112.715 -39.275 113.045 ;
        RECT -39.605 111.355 -39.275 111.685 ;
        RECT -39.605 109.995 -39.275 110.325 ;
        RECT -39.605 108.635 -39.275 108.965 ;
        RECT -39.605 107.275 -39.275 107.605 ;
        RECT -39.605 105.915 -39.275 106.245 ;
        RECT -39.605 104.555 -39.275 104.885 ;
        RECT -39.605 103.195 -39.275 103.525 ;
        RECT -39.605 101.835 -39.275 102.165 ;
        RECT -39.605 100.475 -39.275 100.805 ;
        RECT -39.605 99.115 -39.275 99.445 ;
        RECT -39.605 97.755 -39.275 98.085 ;
        RECT -39.605 96.395 -39.275 96.725 ;
        RECT -39.605 95.035 -39.275 95.365 ;
        RECT -39.605 93.675 -39.275 94.005 ;
        RECT -39.605 92.315 -39.275 92.645 ;
        RECT -39.605 90.955 -39.275 91.285 ;
        RECT -39.605 89.595 -39.275 89.925 ;
        RECT -39.605 88.235 -39.275 88.565 ;
        RECT -39.605 86.875 -39.275 87.205 ;
        RECT -39.605 85.515 -39.275 85.845 ;
        RECT -39.605 84.155 -39.275 84.485 ;
        RECT -39.605 82.795 -39.275 83.125 ;
        RECT -39.605 81.435 -39.275 81.765 ;
        RECT -39.605 80.075 -39.275 80.405 ;
        RECT -39.605 78.715 -39.275 79.045 ;
        RECT -39.605 77.355 -39.275 77.685 ;
        RECT -39.605 75.995 -39.275 76.325 ;
        RECT -39.605 74.635 -39.275 74.965 ;
        RECT -39.605 73.275 -39.275 73.605 ;
        RECT -39.605 71.915 -39.275 72.245 ;
        RECT -39.605 70.555 -39.275 70.885 ;
        RECT -39.605 69.195 -39.275 69.525 ;
        RECT -39.605 67.835 -39.275 68.165 ;
        RECT -39.605 66.475 -39.275 66.805 ;
        RECT -39.605 65.115 -39.275 65.445 ;
        RECT -39.605 63.755 -39.275 64.085 ;
        RECT -39.605 62.395 -39.275 62.725 ;
        RECT -39.605 61.035 -39.275 61.365 ;
        RECT -39.605 59.675 -39.275 60.005 ;
        RECT -39.605 58.315 -39.275 58.645 ;
        RECT -39.605 56.955 -39.275 57.285 ;
        RECT -39.605 55.595 -39.275 55.925 ;
        RECT -39.605 54.235 -39.275 54.565 ;
        RECT -39.605 52.875 -39.275 53.205 ;
        RECT -39.605 51.515 -39.275 51.845 ;
        RECT -39.605 50.155 -39.275 50.485 ;
        RECT -39.605 48.795 -39.275 49.125 ;
        RECT -39.605 47.435 -39.275 47.765 ;
        RECT -39.605 46.075 -39.275 46.405 ;
        RECT -39.605 44.715 -39.275 45.045 ;
        RECT -39.605 43.355 -39.275 43.685 ;
        RECT -39.605 41.995 -39.275 42.325 ;
        RECT -39.605 40.635 -39.275 40.965 ;
        RECT -39.605 39.275 -39.275 39.605 ;
        RECT -39.605 37.915 -39.275 38.245 ;
        RECT -39.605 36.555 -39.275 36.885 ;
        RECT -39.605 35.195 -39.275 35.525 ;
        RECT -39.605 33.835 -39.275 34.165 ;
        RECT -39.605 32.475 -39.275 32.805 ;
        RECT -39.605 31.115 -39.275 31.445 ;
        RECT -39.605 29.755 -39.275 30.085 ;
        RECT -39.605 28.395 -39.275 28.725 ;
        RECT -39.605 27.035 -39.275 27.365 ;
        RECT -39.605 25.675 -39.275 26.005 ;
        RECT -39.605 24.315 -39.275 24.645 ;
        RECT -39.605 22.955 -39.275 23.285 ;
        RECT -39.605 21.595 -39.275 21.925 ;
        RECT -39.605 20.235 -39.275 20.565 ;
        RECT -39.605 18.875 -39.275 19.205 ;
        RECT -39.605 17.515 -39.275 17.845 ;
        RECT -39.605 16.155 -39.275 16.485 ;
        RECT -39.605 14.795 -39.275 15.125 ;
        RECT -39.605 13.435 -39.275 13.765 ;
        RECT -39.605 12.075 -39.275 12.405 ;
        RECT -39.605 10.715 -39.275 11.045 ;
        RECT -39.605 9.355 -39.275 9.685 ;
        RECT -39.605 7.995 -39.275 8.325 ;
        RECT -39.605 6.635 -39.275 6.965 ;
        RECT -39.605 5.275 -39.275 5.605 ;
        RECT -39.605 3.915 -39.275 4.245 ;
        RECT -39.605 2.555 -39.275 2.885 ;
        RECT -39.605 1.195 -39.275 1.525 ;
        RECT -39.605 -0.165 -39.275 0.165 ;
        RECT -39.605 -1.525 -39.275 -1.195 ;
        RECT -39.605 -8.325 -39.275 -7.995 ;
        RECT -39.605 -9.685 -39.275 -9.355 ;
        RECT -39.605 -12.405 -39.275 -12.075 ;
        RECT -39.605 -13.765 -39.275 -13.435 ;
        RECT -39.605 -15.125 -39.275 -14.795 ;
        RECT -39.605 -16.485 -39.275 -16.155 ;
        RECT -39.605 -17.845 -39.275 -17.515 ;
        RECT -39.605 -19.205 -39.275 -18.875 ;
        RECT -39.605 -20.565 -39.275 -20.235 ;
        RECT -39.605 -21.925 -39.275 -21.595 ;
        RECT -39.605 -23.285 -39.275 -22.955 ;
        RECT -39.605 -30.66 -39.275 -30.33 ;
        RECT -39.605 -31.445 -39.275 -31.115 ;
        RECT -39.605 -32.805 -39.275 -32.475 ;
        RECT -39.605 -34.165 -39.275 -33.835 ;
        RECT -39.605 -36.885 -39.275 -36.555 ;
        RECT -39.605 -37.85 -39.275 -37.52 ;
        RECT -39.605 -40.965 -39.275 -40.635 ;
        RECT -39.605 -46.405 -39.275 -46.075 ;
        RECT -39.605 -49.125 -39.275 -48.795 ;
        RECT -39.605 -50.485 -39.275 -50.155 ;
        RECT -39.605 -53.205 -39.275 -52.875 ;
        RECT -39.605 -55.925 -39.275 -55.595 ;
        RECT -39.605 -61.365 -39.275 -61.035 ;
        RECT -39.605 -62.725 -39.275 -62.395 ;
        RECT -39.605 -64.085 -39.275 -63.755 ;
        RECT -39.605 -65.445 -39.275 -65.115 ;
        RECT -39.605 -66.805 -39.275 -66.475 ;
        RECT -39.605 -68.165 -39.275 -67.835 ;
        RECT -39.605 -69.525 -39.275 -69.195 ;
        RECT -39.605 -70.885 -39.275 -70.555 ;
        RECT -39.605 -72.245 -39.275 -71.915 ;
        RECT -39.605 -73.605 -39.275 -73.275 ;
        RECT -39.605 -74.965 -39.275 -74.635 ;
        RECT -39.605 -76.325 -39.275 -75.995 ;
        RECT -39.605 -77.685 -39.275 -77.355 ;
        RECT -39.605 -79.045 -39.275 -78.715 ;
        RECT -39.605 -80.405 -39.275 -80.075 ;
        RECT -39.605 -81.765 -39.275 -81.435 ;
        RECT -39.605 -83.125 -39.275 -82.795 ;
        RECT -39.605 -84.485 -39.275 -84.155 ;
        RECT -39.605 -85.845 -39.275 -85.515 ;
        RECT -39.605 -87.205 -39.275 -86.875 ;
        RECT -39.605 -88.565 -39.275 -88.235 ;
        RECT -39.605 -89.925 -39.275 -89.595 ;
        RECT -39.605 -91.285 -39.275 -90.955 ;
        RECT -39.605 -92.645 -39.275 -92.315 ;
        RECT -39.605 -94.005 -39.275 -93.675 ;
        RECT -39.605 -95.365 -39.275 -95.035 ;
        RECT -39.605 -96.725 -39.275 -96.395 ;
        RECT -39.605 -98.085 -39.275 -97.755 ;
        RECT -39.605 -99.445 -39.275 -99.115 ;
        RECT -39.605 -100.805 -39.275 -100.475 ;
        RECT -39.605 -102.165 -39.275 -101.835 ;
        RECT -39.605 -103.525 -39.275 -103.195 ;
        RECT -39.605 -104.885 -39.275 -104.555 ;
        RECT -39.605 -106.245 -39.275 -105.915 ;
        RECT -39.605 -107.605 -39.275 -107.275 ;
        RECT -39.605 -108.965 -39.275 -108.635 ;
        RECT -39.605 -110.325 -39.275 -109.995 ;
        RECT -39.605 -111.685 -39.275 -111.355 ;
        RECT -39.605 -113.045 -39.275 -112.715 ;
        RECT -39.605 -114.405 -39.275 -114.075 ;
        RECT -39.605 -115.765 -39.275 -115.435 ;
        RECT -39.605 -117.125 -39.275 -116.795 ;
        RECT -39.605 -118.485 -39.275 -118.155 ;
        RECT -39.605 -119.845 -39.275 -119.515 ;
        RECT -39.605 -123.925 -39.275 -123.595 ;
        RECT -39.605 -129.365 -39.275 -129.035 ;
        RECT -39.605 -130.725 -39.275 -130.395 ;
        RECT -39.605 -131.47 -39.275 -131.14 ;
        RECT -39.605 -133.445 -39.275 -133.115 ;
        RECT -39.605 -134.805 -39.275 -134.475 ;
        RECT -39.605 -136.165 -39.275 -135.835 ;
        RECT -39.605 -137.525 -39.275 -137.195 ;
        RECT -39.605 -140.245 -39.275 -139.915 ;
        RECT -39.605 -141.605 -39.275 -141.275 ;
        RECT -39.605 -142.965 -39.275 -142.635 ;
        RECT -39.605 -144.31 -39.275 -143.98 ;
        RECT -39.605 -145.685 -39.275 -145.355 ;
        RECT -39.605 -147.045 -39.275 -146.715 ;
        RECT -39.605 -149.765 -39.275 -149.435 ;
        RECT -39.605 -153.845 -39.275 -153.515 ;
        RECT -39.605 -155.205 -39.275 -154.875 ;
        RECT -39.605 -156.565 -39.275 -156.235 ;
        RECT -39.605 -157.925 -39.275 -157.595 ;
        RECT -39.605 -159.285 -39.275 -158.955 ;
        RECT -39.605 -162.005 -39.275 -161.675 ;
        RECT -39.605 -163.365 -39.275 -163.035 ;
        RECT -39.605 -164.725 -39.275 -164.395 ;
        RECT -39.605 -166.085 -39.275 -165.755 ;
        RECT -39.605 -167.445 -39.275 -167.115 ;
        RECT -39.605 -168.805 -39.275 -168.475 ;
        RECT -39.605 -170.165 -39.275 -169.835 ;
        RECT -39.605 -171.525 -39.275 -171.195 ;
        RECT -39.605 -172.885 -39.275 -172.555 ;
        RECT -39.605 -174.245 -39.275 -173.915 ;
        RECT -39.605 -175.605 -39.275 -175.275 ;
        RECT -39.605 -176.965 -39.275 -176.635 ;
        RECT -39.605 -178.325 -39.275 -177.995 ;
        RECT -39.605 -179.685 -39.275 -179.355 ;
        RECT -39.605 -181.045 -39.275 -180.715 ;
        RECT -39.605 -182.405 -39.275 -182.075 ;
        RECT -39.605 -183.765 -39.275 -183.435 ;
        RECT -39.605 -185.125 -39.275 -184.795 ;
        RECT -39.605 -186.485 -39.275 -186.155 ;
        RECT -39.605 -187.845 -39.275 -187.515 ;
        RECT -39.605 -189.205 -39.275 -188.875 ;
        RECT -39.605 -190.565 -39.275 -190.235 ;
        RECT -39.605 -191.925 -39.275 -191.595 ;
        RECT -39.605 -193.285 -39.275 -192.955 ;
        RECT -39.605 -194.645 -39.275 -194.315 ;
        RECT -39.605 -196.005 -39.275 -195.675 ;
        RECT -39.605 -197.365 -39.275 -197.035 ;
        RECT -39.605 -198.725 -39.275 -198.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 246.76 -48.795 247.89 ;
        RECT -49.125 241.915 -48.795 242.245 ;
        RECT -49.125 240.555 -48.795 240.885 ;
        RECT -49.125 239.195 -48.795 239.525 ;
        RECT -49.125 237.835 -48.795 238.165 ;
        RECT -49.125 236.475 -48.795 236.805 ;
        RECT -49.125 235.115 -48.795 235.445 ;
        RECT -49.125 233.755 -48.795 234.085 ;
        RECT -49.125 232.395 -48.795 232.725 ;
        RECT -49.125 231.035 -48.795 231.365 ;
        RECT -49.125 229.675 -48.795 230.005 ;
        RECT -49.125 228.315 -48.795 228.645 ;
        RECT -49.125 226.955 -48.795 227.285 ;
        RECT -49.125 225.595 -48.795 225.925 ;
        RECT -49.125 224.235 -48.795 224.565 ;
        RECT -49.125 222.875 -48.795 223.205 ;
        RECT -49.125 221.515 -48.795 221.845 ;
        RECT -49.125 220.155 -48.795 220.485 ;
        RECT -49.125 218.795 -48.795 219.125 ;
        RECT -49.125 217.435 -48.795 217.765 ;
        RECT -49.125 216.075 -48.795 216.405 ;
        RECT -49.125 214.715 -48.795 215.045 ;
        RECT -49.125 213.355 -48.795 213.685 ;
        RECT -49.125 211.995 -48.795 212.325 ;
        RECT -49.125 210.635 -48.795 210.965 ;
        RECT -49.125 209.275 -48.795 209.605 ;
        RECT -49.125 207.915 -48.795 208.245 ;
        RECT -49.125 206.555 -48.795 206.885 ;
        RECT -49.125 205.195 -48.795 205.525 ;
        RECT -49.125 203.835 -48.795 204.165 ;
        RECT -49.125 202.475 -48.795 202.805 ;
        RECT -49.125 201.115 -48.795 201.445 ;
        RECT -49.125 199.755 -48.795 200.085 ;
        RECT -49.125 198.395 -48.795 198.725 ;
        RECT -49.125 197.035 -48.795 197.365 ;
        RECT -49.125 195.675 -48.795 196.005 ;
        RECT -49.125 194.315 -48.795 194.645 ;
        RECT -49.125 192.955 -48.795 193.285 ;
        RECT -49.125 191.595 -48.795 191.925 ;
        RECT -49.125 190.235 -48.795 190.565 ;
        RECT -49.125 188.875 -48.795 189.205 ;
        RECT -49.125 187.515 -48.795 187.845 ;
        RECT -49.125 186.155 -48.795 186.485 ;
        RECT -49.125 184.795 -48.795 185.125 ;
        RECT -49.125 183.435 -48.795 183.765 ;
        RECT -49.125 182.075 -48.795 182.405 ;
        RECT -49.125 180.715 -48.795 181.045 ;
        RECT -49.125 179.355 -48.795 179.685 ;
        RECT -49.125 177.995 -48.795 178.325 ;
        RECT -49.125 176.635 -48.795 176.965 ;
        RECT -49.125 175.275 -48.795 175.605 ;
        RECT -49.125 173.915 -48.795 174.245 ;
        RECT -49.125 172.555 -48.795 172.885 ;
        RECT -49.125 171.195 -48.795 171.525 ;
        RECT -49.125 169.835 -48.795 170.165 ;
        RECT -49.125 168.475 -48.795 168.805 ;
        RECT -49.125 167.115 -48.795 167.445 ;
        RECT -49.125 165.755 -48.795 166.085 ;
        RECT -49.125 164.395 -48.795 164.725 ;
        RECT -49.125 163.035 -48.795 163.365 ;
        RECT -49.125 161.675 -48.795 162.005 ;
        RECT -49.125 160.315 -48.795 160.645 ;
        RECT -49.125 158.955 -48.795 159.285 ;
        RECT -49.125 157.595 -48.795 157.925 ;
        RECT -49.125 156.235 -48.795 156.565 ;
        RECT -49.125 154.875 -48.795 155.205 ;
        RECT -49.125 153.515 -48.795 153.845 ;
        RECT -49.125 152.155 -48.795 152.485 ;
        RECT -49.125 150.795 -48.795 151.125 ;
        RECT -49.125 149.435 -48.795 149.765 ;
        RECT -49.125 148.075 -48.795 148.405 ;
        RECT -49.125 146.715 -48.795 147.045 ;
        RECT -49.125 145.355 -48.795 145.685 ;
        RECT -49.125 143.995 -48.795 144.325 ;
        RECT -49.125 142.635 -48.795 142.965 ;
        RECT -49.125 141.275 -48.795 141.605 ;
        RECT -49.125 139.915 -48.795 140.245 ;
        RECT -49.125 138.555 -48.795 138.885 ;
        RECT -49.125 136.42 -48.795 136.75 ;
        RECT -49.125 134.245 -48.795 134.575 ;
        RECT -49.125 133.395 -48.795 133.725 ;
        RECT -49.125 131.085 -48.795 131.415 ;
        RECT -49.125 130.235 -48.795 130.565 ;
        RECT -49.125 127.925 -48.795 128.255 ;
        RECT -49.125 127.075 -48.795 127.405 ;
        RECT -49.125 124.765 -48.795 125.095 ;
        RECT -49.125 123.915 -48.795 124.245 ;
        RECT -49.125 121.605 -48.795 121.935 ;
        RECT -49.125 120.755 -48.795 121.085 ;
        RECT -49.125 118.445 -48.795 118.775 ;
        RECT -49.125 117.595 -48.795 117.925 ;
        RECT -49.12 117.48 -48.8 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 -159.285 -48.795 -158.955 ;
        RECT -49.125 -162.005 -48.795 -161.675 ;
        RECT -49.125 -163.365 -48.795 -163.035 ;
        RECT -49.125 -164.725 -48.795 -164.395 ;
        RECT -49.125 -166.085 -48.795 -165.755 ;
        RECT -49.125 -167.445 -48.795 -167.115 ;
        RECT -49.125 -168.805 -48.795 -168.475 ;
        RECT -49.125 -170.165 -48.795 -169.835 ;
        RECT -49.125 -171.525 -48.795 -171.195 ;
        RECT -49.125 -172.885 -48.795 -172.555 ;
        RECT -49.125 -174.245 -48.795 -173.915 ;
        RECT -49.125 -175.605 -48.795 -175.275 ;
        RECT -49.125 -176.965 -48.795 -176.635 ;
        RECT -49.125 -178.325 -48.795 -177.995 ;
        RECT -49.125 -179.685 -48.795 -179.355 ;
        RECT -49.125 -181.045 -48.795 -180.715 ;
        RECT -49.125 -182.405 -48.795 -182.075 ;
        RECT -49.125 -183.765 -48.795 -183.435 ;
        RECT -49.125 -185.125 -48.795 -184.795 ;
        RECT -49.125 -186.485 -48.795 -186.155 ;
        RECT -49.125 -187.845 -48.795 -187.515 ;
        RECT -49.125 -189.205 -48.795 -188.875 ;
        RECT -49.125 -190.565 -48.795 -190.235 ;
        RECT -49.125 -191.925 -48.795 -191.595 ;
        RECT -49.125 -193.285 -48.795 -192.955 ;
        RECT -49.125 -194.645 -48.795 -194.315 ;
        RECT -49.125 -196.005 -48.795 -195.675 ;
        RECT -49.125 -197.365 -48.795 -197.035 ;
        RECT -49.125 -198.725 -48.795 -198.395 ;
        RECT -49.125 -200.085 -48.795 -199.755 ;
        RECT -49.125 -201.445 -48.795 -201.115 ;
        RECT -49.125 -202.805 -48.795 -202.475 ;
        RECT -49.125 -204.165 -48.795 -203.835 ;
        RECT -49.125 -205.525 -48.795 -205.195 ;
        RECT -49.125 -206.885 -48.795 -206.555 ;
        RECT -49.125 -208.245 -48.795 -207.915 ;
        RECT -49.125 -209.605 -48.795 -209.275 ;
        RECT -49.125 -210.965 -48.795 -210.635 ;
        RECT -49.125 -212.325 -48.795 -211.995 ;
        RECT -49.125 -213.685 -48.795 -213.355 ;
        RECT -49.125 -215.045 -48.795 -214.715 ;
        RECT -49.125 -216.405 -48.795 -216.075 ;
        RECT -49.125 -217.765 -48.795 -217.435 ;
        RECT -49.125 -219.125 -48.795 -218.795 ;
        RECT -49.125 -220.485 -48.795 -220.155 ;
        RECT -49.125 -221.845 -48.795 -221.515 ;
        RECT -49.125 -223.205 -48.795 -222.875 ;
        RECT -49.125 -224.565 -48.795 -224.235 ;
        RECT -49.125 -226.155 -48.795 -225.825 ;
        RECT -49.125 -227.285 -48.795 -226.955 ;
        RECT -49.125 -228.645 -48.795 -228.315 ;
        RECT -49.125 -230.005 -48.795 -229.675 ;
        RECT -49.125 -231.365 -48.795 -231.035 ;
        RECT -49.125 -234.085 -48.795 -233.755 ;
        RECT -49.125 -235.445 -48.795 -235.115 ;
        RECT -49.125 -236.805 -48.795 -236.475 ;
        RECT -49.125 -238.165 -48.795 -237.835 ;
        RECT -49.125 -243.81 -48.795 -242.68 ;
        RECT -49.12 -243.925 -48.8 -158.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 246.76 -47.435 247.89 ;
        RECT -47.765 241.915 -47.435 242.245 ;
        RECT -47.765 240.555 -47.435 240.885 ;
        RECT -47.765 239.195 -47.435 239.525 ;
        RECT -47.765 237.835 -47.435 238.165 ;
        RECT -47.765 236.475 -47.435 236.805 ;
        RECT -47.765 235.115 -47.435 235.445 ;
        RECT -47.765 233.755 -47.435 234.085 ;
        RECT -47.765 232.395 -47.435 232.725 ;
        RECT -47.765 231.035 -47.435 231.365 ;
        RECT -47.765 229.675 -47.435 230.005 ;
        RECT -47.765 228.315 -47.435 228.645 ;
        RECT -47.765 226.955 -47.435 227.285 ;
        RECT -47.765 225.595 -47.435 225.925 ;
        RECT -47.765 224.235 -47.435 224.565 ;
        RECT -47.765 222.875 -47.435 223.205 ;
        RECT -47.765 221.515 -47.435 221.845 ;
        RECT -47.765 220.155 -47.435 220.485 ;
        RECT -47.765 218.795 -47.435 219.125 ;
        RECT -47.765 217.435 -47.435 217.765 ;
        RECT -47.765 216.075 -47.435 216.405 ;
        RECT -47.765 214.715 -47.435 215.045 ;
        RECT -47.765 213.355 -47.435 213.685 ;
        RECT -47.765 211.995 -47.435 212.325 ;
        RECT -47.765 210.635 -47.435 210.965 ;
        RECT -47.765 209.275 -47.435 209.605 ;
        RECT -47.765 207.915 -47.435 208.245 ;
        RECT -47.765 206.555 -47.435 206.885 ;
        RECT -47.765 205.195 -47.435 205.525 ;
        RECT -47.765 203.835 -47.435 204.165 ;
        RECT -47.765 202.475 -47.435 202.805 ;
        RECT -47.765 201.115 -47.435 201.445 ;
        RECT -47.765 199.755 -47.435 200.085 ;
        RECT -47.765 198.395 -47.435 198.725 ;
        RECT -47.765 197.035 -47.435 197.365 ;
        RECT -47.765 195.675 -47.435 196.005 ;
        RECT -47.765 194.315 -47.435 194.645 ;
        RECT -47.765 192.955 -47.435 193.285 ;
        RECT -47.765 191.595 -47.435 191.925 ;
        RECT -47.765 190.235 -47.435 190.565 ;
        RECT -47.765 188.875 -47.435 189.205 ;
        RECT -47.765 187.515 -47.435 187.845 ;
        RECT -47.765 186.155 -47.435 186.485 ;
        RECT -47.765 184.795 -47.435 185.125 ;
        RECT -47.765 183.435 -47.435 183.765 ;
        RECT -47.765 182.075 -47.435 182.405 ;
        RECT -47.765 180.715 -47.435 181.045 ;
        RECT -47.765 179.355 -47.435 179.685 ;
        RECT -47.765 177.995 -47.435 178.325 ;
        RECT -47.765 176.635 -47.435 176.965 ;
        RECT -47.765 175.275 -47.435 175.605 ;
        RECT -47.765 173.915 -47.435 174.245 ;
        RECT -47.765 172.555 -47.435 172.885 ;
        RECT -47.765 171.195 -47.435 171.525 ;
        RECT -47.765 169.835 -47.435 170.165 ;
        RECT -47.765 168.475 -47.435 168.805 ;
        RECT -47.765 167.115 -47.435 167.445 ;
        RECT -47.765 165.755 -47.435 166.085 ;
        RECT -47.765 164.395 -47.435 164.725 ;
        RECT -47.765 163.035 -47.435 163.365 ;
        RECT -47.765 161.675 -47.435 162.005 ;
        RECT -47.765 160.315 -47.435 160.645 ;
        RECT -47.765 158.955 -47.435 159.285 ;
        RECT -47.765 157.595 -47.435 157.925 ;
        RECT -47.765 156.235 -47.435 156.565 ;
        RECT -47.765 154.875 -47.435 155.205 ;
        RECT -47.765 153.515 -47.435 153.845 ;
        RECT -47.765 152.155 -47.435 152.485 ;
        RECT -47.765 150.795 -47.435 151.125 ;
        RECT -47.765 149.435 -47.435 149.765 ;
        RECT -47.765 148.075 -47.435 148.405 ;
        RECT -47.765 146.715 -47.435 147.045 ;
        RECT -47.765 145.355 -47.435 145.685 ;
        RECT -47.765 143.995 -47.435 144.325 ;
        RECT -47.765 142.635 -47.435 142.965 ;
        RECT -47.765 141.275 -47.435 141.605 ;
        RECT -47.765 139.915 -47.435 140.245 ;
        RECT -47.765 138.555 -47.435 138.885 ;
        RECT -47.765 136.42 -47.435 136.75 ;
        RECT -47.765 134.245 -47.435 134.575 ;
        RECT -47.765 133.395 -47.435 133.725 ;
        RECT -47.765 131.085 -47.435 131.415 ;
        RECT -47.765 130.235 -47.435 130.565 ;
        RECT -47.765 127.925 -47.435 128.255 ;
        RECT -47.765 127.075 -47.435 127.405 ;
        RECT -47.765 124.765 -47.435 125.095 ;
        RECT -47.765 123.915 -47.435 124.245 ;
        RECT -47.765 121.605 -47.435 121.935 ;
        RECT -47.765 120.755 -47.435 121.085 ;
        RECT -47.765 118.445 -47.435 118.775 ;
        RECT -47.765 117.595 -47.435 117.925 ;
        RECT -47.765 115.285 -47.435 115.615 ;
        RECT -47.765 114.435 -47.435 114.765 ;
        RECT -47.765 112.125 -47.435 112.455 ;
        RECT -47.765 111.275 -47.435 111.605 ;
        RECT -47.765 108.965 -47.435 109.295 ;
        RECT -47.765 108.115 -47.435 108.445 ;
        RECT -47.765 105.805 -47.435 106.135 ;
        RECT -47.765 104.955 -47.435 105.285 ;
        RECT -47.765 102.645 -47.435 102.975 ;
        RECT -47.765 101.795 -47.435 102.125 ;
        RECT -47.765 99.62 -47.435 99.95 ;
        RECT -47.765 97.755 -47.435 98.085 ;
        RECT -47.765 96.395 -47.435 96.725 ;
        RECT -47.765 95.035 -47.435 95.365 ;
        RECT -47.765 93.675 -47.435 94.005 ;
        RECT -47.765 92.315 -47.435 92.645 ;
        RECT -47.765 90.955 -47.435 91.285 ;
        RECT -47.765 89.595 -47.435 89.925 ;
        RECT -47.765 88.235 -47.435 88.565 ;
        RECT -47.765 86.875 -47.435 87.205 ;
        RECT -47.765 85.515 -47.435 85.845 ;
        RECT -47.765 84.155 -47.435 84.485 ;
        RECT -47.765 82.795 -47.435 83.125 ;
        RECT -47.765 81.435 -47.435 81.765 ;
        RECT -47.765 80.075 -47.435 80.405 ;
        RECT -47.765 78.715 -47.435 79.045 ;
        RECT -47.765 77.355 -47.435 77.685 ;
        RECT -47.765 75.995 -47.435 76.325 ;
        RECT -47.765 74.635 -47.435 74.965 ;
        RECT -47.765 73.275 -47.435 73.605 ;
        RECT -47.765 71.915 -47.435 72.245 ;
        RECT -47.765 70.555 -47.435 70.885 ;
        RECT -47.765 69.195 -47.435 69.525 ;
        RECT -47.765 67.835 -47.435 68.165 ;
        RECT -47.765 66.475 -47.435 66.805 ;
        RECT -47.765 65.115 -47.435 65.445 ;
        RECT -47.765 63.755 -47.435 64.085 ;
        RECT -47.765 62.395 -47.435 62.725 ;
        RECT -47.765 61.035 -47.435 61.365 ;
        RECT -47.765 59.675 -47.435 60.005 ;
        RECT -47.765 58.315 -47.435 58.645 ;
        RECT -47.765 56.955 -47.435 57.285 ;
        RECT -47.765 55.595 -47.435 55.925 ;
        RECT -47.765 54.235 -47.435 54.565 ;
        RECT -47.765 52.875 -47.435 53.205 ;
        RECT -47.765 51.515 -47.435 51.845 ;
        RECT -47.765 50.155 -47.435 50.485 ;
        RECT -47.765 48.795 -47.435 49.125 ;
        RECT -47.765 47.435 -47.435 47.765 ;
        RECT -47.765 46.075 -47.435 46.405 ;
        RECT -47.765 44.715 -47.435 45.045 ;
        RECT -47.765 43.355 -47.435 43.685 ;
        RECT -47.765 41.995 -47.435 42.325 ;
        RECT -47.765 40.635 -47.435 40.965 ;
        RECT -47.765 39.275 -47.435 39.605 ;
        RECT -47.765 37.915 -47.435 38.245 ;
        RECT -47.765 36.555 -47.435 36.885 ;
        RECT -47.765 35.195 -47.435 35.525 ;
        RECT -47.765 33.835 -47.435 34.165 ;
        RECT -47.765 32.475 -47.435 32.805 ;
        RECT -47.765 31.115 -47.435 31.445 ;
        RECT -47.765 29.755 -47.435 30.085 ;
        RECT -47.765 28.395 -47.435 28.725 ;
        RECT -47.765 27.035 -47.435 27.365 ;
        RECT -47.765 25.675 -47.435 26.005 ;
        RECT -47.765 24.315 -47.435 24.645 ;
        RECT -47.765 22.955 -47.435 23.285 ;
        RECT -47.765 21.595 -47.435 21.925 ;
        RECT -47.765 20.235 -47.435 20.565 ;
        RECT -47.765 18.875 -47.435 19.205 ;
        RECT -47.765 17.515 -47.435 17.845 ;
        RECT -47.765 16.155 -47.435 16.485 ;
        RECT -47.765 14.795 -47.435 15.125 ;
        RECT -47.765 13.435 -47.435 13.765 ;
        RECT -47.765 12.075 -47.435 12.405 ;
        RECT -47.765 10.715 -47.435 11.045 ;
        RECT -47.765 9.355 -47.435 9.685 ;
        RECT -47.765 7.995 -47.435 8.325 ;
        RECT -47.765 6.635 -47.435 6.965 ;
        RECT -47.765 5.275 -47.435 5.605 ;
        RECT -47.765 3.915 -47.435 4.245 ;
        RECT -47.765 2.555 -47.435 2.885 ;
        RECT -47.765 1.195 -47.435 1.525 ;
        RECT -47.765 -0.165 -47.435 0.165 ;
        RECT -47.765 -1.525 -47.435 -1.195 ;
        RECT -47.765 -2.885 -47.435 -2.555 ;
        RECT -47.765 -4.245 -47.435 -3.915 ;
        RECT -47.765 -5.605 -47.435 -5.275 ;
        RECT -47.765 -6.965 -47.435 -6.635 ;
        RECT -47.765 -8.325 -47.435 -7.995 ;
        RECT -47.765 -9.685 -47.435 -9.355 ;
        RECT -47.765 -12.405 -47.435 -12.075 ;
        RECT -47.765 -13.765 -47.435 -13.435 ;
        RECT -47.765 -15.125 -47.435 -14.795 ;
        RECT -47.765 -16.485 -47.435 -16.155 ;
        RECT -47.765 -17.845 -47.435 -17.515 ;
        RECT -47.765 -19.205 -47.435 -18.875 ;
        RECT -47.765 -20.565 -47.435 -20.235 ;
        RECT -47.765 -21.925 -47.435 -21.595 ;
        RECT -47.765 -23.285 -47.435 -22.955 ;
        RECT -47.765 -24.645 -47.435 -24.315 ;
        RECT -47.765 -26.005 -47.435 -25.675 ;
        RECT -47.765 -27.365 -47.435 -27.035 ;
        RECT -47.765 -30.66 -47.435 -30.33 ;
        RECT -47.765 -31.445 -47.435 -31.115 ;
        RECT -47.765 -32.805 -47.435 -32.475 ;
        RECT -47.765 -34.165 -47.435 -33.835 ;
        RECT -47.765 -36.885 -47.435 -36.555 ;
        RECT -47.765 -37.85 -47.435 -37.52 ;
        RECT -47.765 -40.965 -47.435 -40.635 ;
        RECT -47.765 -46.405 -47.435 -46.075 ;
        RECT -47.765 -49.125 -47.435 -48.795 ;
        RECT -47.765 -50.485 -47.435 -50.155 ;
        RECT -47.765 -53.205 -47.435 -52.875 ;
        RECT -47.765 -55.925 -47.435 -55.595 ;
        RECT -47.765 -61.365 -47.435 -61.035 ;
        RECT -47.765 -62.725 -47.435 -62.395 ;
        RECT -47.765 -64.085 -47.435 -63.755 ;
        RECT -47.765 -65.445 -47.435 -65.115 ;
        RECT -47.765 -66.805 -47.435 -66.475 ;
        RECT -47.765 -68.165 -47.435 -67.835 ;
        RECT -47.765 -69.525 -47.435 -69.195 ;
        RECT -47.765 -70.885 -47.435 -70.555 ;
        RECT -47.765 -72.245 -47.435 -71.915 ;
        RECT -47.765 -73.605 -47.435 -73.275 ;
        RECT -47.765 -74.965 -47.435 -74.635 ;
        RECT -47.765 -76.325 -47.435 -75.995 ;
        RECT -47.765 -77.685 -47.435 -77.355 ;
        RECT -47.765 -79.045 -47.435 -78.715 ;
        RECT -47.765 -80.405 -47.435 -80.075 ;
        RECT -47.765 -81.765 -47.435 -81.435 ;
        RECT -47.765 -83.125 -47.435 -82.795 ;
        RECT -47.765 -84.485 -47.435 -84.155 ;
        RECT -47.765 -85.845 -47.435 -85.515 ;
        RECT -47.765 -87.205 -47.435 -86.875 ;
        RECT -47.765 -88.565 -47.435 -88.235 ;
        RECT -47.765 -89.925 -47.435 -89.595 ;
        RECT -47.765 -91.285 -47.435 -90.955 ;
        RECT -47.765 -92.645 -47.435 -92.315 ;
        RECT -47.765 -94.005 -47.435 -93.675 ;
        RECT -47.765 -95.365 -47.435 -95.035 ;
        RECT -47.765 -96.725 -47.435 -96.395 ;
        RECT -47.765 -98.085 -47.435 -97.755 ;
        RECT -47.765 -99.445 -47.435 -99.115 ;
        RECT -47.765 -100.805 -47.435 -100.475 ;
        RECT -47.765 -102.165 -47.435 -101.835 ;
        RECT -47.765 -103.525 -47.435 -103.195 ;
        RECT -47.765 -104.885 -47.435 -104.555 ;
        RECT -47.765 -106.245 -47.435 -105.915 ;
        RECT -47.765 -107.605 -47.435 -107.275 ;
        RECT -47.765 -108.965 -47.435 -108.635 ;
        RECT -47.765 -110.325 -47.435 -109.995 ;
        RECT -47.765 -111.685 -47.435 -111.355 ;
        RECT -47.765 -113.045 -47.435 -112.715 ;
        RECT -47.765 -114.405 -47.435 -114.075 ;
        RECT -47.765 -115.765 -47.435 -115.435 ;
        RECT -47.765 -117.125 -47.435 -116.795 ;
        RECT -47.765 -118.485 -47.435 -118.155 ;
        RECT -47.765 -119.845 -47.435 -119.515 ;
        RECT -47.765 -121.205 -47.435 -120.875 ;
        RECT -47.765 -129.365 -47.435 -129.035 ;
        RECT -47.765 -130.725 -47.435 -130.395 ;
        RECT -47.765 -131.47 -47.435 -131.14 ;
        RECT -47.765 -133.445 -47.435 -133.115 ;
        RECT -47.765 -134.805 -47.435 -134.475 ;
        RECT -47.765 -136.165 -47.435 -135.835 ;
        RECT -47.765 -137.525 -47.435 -137.195 ;
        RECT -47.765 -140.245 -47.435 -139.915 ;
        RECT -47.765 -141.605 -47.435 -141.275 ;
        RECT -47.765 -142.965 -47.435 -142.635 ;
        RECT -47.765 -144.31 -47.435 -143.98 ;
        RECT -47.765 -145.685 -47.435 -145.355 ;
        RECT -47.765 -147.045 -47.435 -146.715 ;
        RECT -47.765 -149.765 -47.435 -149.435 ;
        RECT -47.76 -151.8 -47.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 -234.085 -47.435 -233.755 ;
        RECT -47.765 -235.445 -47.435 -235.115 ;
        RECT -47.765 -236.805 -47.435 -236.475 ;
        RECT -47.765 -238.165 -47.435 -237.835 ;
        RECT -47.765 -243.81 -47.435 -242.68 ;
        RECT -47.76 -243.925 -47.44 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 246.76 -46.075 247.89 ;
        RECT -46.405 241.915 -46.075 242.245 ;
        RECT -46.405 240.555 -46.075 240.885 ;
        RECT -46.405 239.195 -46.075 239.525 ;
        RECT -46.405 237.835 -46.075 238.165 ;
        RECT -46.405 236.475 -46.075 236.805 ;
        RECT -46.405 235.115 -46.075 235.445 ;
        RECT -46.405 233.755 -46.075 234.085 ;
        RECT -46.405 232.395 -46.075 232.725 ;
        RECT -46.405 231.035 -46.075 231.365 ;
        RECT -46.405 229.675 -46.075 230.005 ;
        RECT -46.405 228.315 -46.075 228.645 ;
        RECT -46.405 226.955 -46.075 227.285 ;
        RECT -46.405 225.595 -46.075 225.925 ;
        RECT -46.405 224.235 -46.075 224.565 ;
        RECT -46.405 222.875 -46.075 223.205 ;
        RECT -46.405 221.515 -46.075 221.845 ;
        RECT -46.405 220.155 -46.075 220.485 ;
        RECT -46.405 218.795 -46.075 219.125 ;
        RECT -46.405 217.435 -46.075 217.765 ;
        RECT -46.405 216.075 -46.075 216.405 ;
        RECT -46.405 214.715 -46.075 215.045 ;
        RECT -46.405 213.355 -46.075 213.685 ;
        RECT -46.405 211.995 -46.075 212.325 ;
        RECT -46.405 210.635 -46.075 210.965 ;
        RECT -46.405 209.275 -46.075 209.605 ;
        RECT -46.405 207.915 -46.075 208.245 ;
        RECT -46.405 206.555 -46.075 206.885 ;
        RECT -46.405 205.195 -46.075 205.525 ;
        RECT -46.405 203.835 -46.075 204.165 ;
        RECT -46.405 202.475 -46.075 202.805 ;
        RECT -46.405 201.115 -46.075 201.445 ;
        RECT -46.405 199.755 -46.075 200.085 ;
        RECT -46.405 198.395 -46.075 198.725 ;
        RECT -46.405 197.035 -46.075 197.365 ;
        RECT -46.405 195.675 -46.075 196.005 ;
        RECT -46.405 194.315 -46.075 194.645 ;
        RECT -46.405 192.955 -46.075 193.285 ;
        RECT -46.405 191.595 -46.075 191.925 ;
        RECT -46.405 190.235 -46.075 190.565 ;
        RECT -46.405 188.875 -46.075 189.205 ;
        RECT -46.405 187.515 -46.075 187.845 ;
        RECT -46.405 186.155 -46.075 186.485 ;
        RECT -46.405 184.795 -46.075 185.125 ;
        RECT -46.405 183.435 -46.075 183.765 ;
        RECT -46.405 182.075 -46.075 182.405 ;
        RECT -46.405 180.715 -46.075 181.045 ;
        RECT -46.405 179.355 -46.075 179.685 ;
        RECT -46.405 177.995 -46.075 178.325 ;
        RECT -46.405 176.635 -46.075 176.965 ;
        RECT -46.405 175.275 -46.075 175.605 ;
        RECT -46.405 173.915 -46.075 174.245 ;
        RECT -46.405 172.555 -46.075 172.885 ;
        RECT -46.405 171.195 -46.075 171.525 ;
        RECT -46.405 169.835 -46.075 170.165 ;
        RECT -46.405 168.475 -46.075 168.805 ;
        RECT -46.405 167.115 -46.075 167.445 ;
        RECT -46.405 165.755 -46.075 166.085 ;
        RECT -46.405 164.395 -46.075 164.725 ;
        RECT -46.405 163.035 -46.075 163.365 ;
        RECT -46.405 161.675 -46.075 162.005 ;
        RECT -46.405 160.315 -46.075 160.645 ;
        RECT -46.405 158.955 -46.075 159.285 ;
        RECT -46.405 157.595 -46.075 157.925 ;
        RECT -46.405 156.235 -46.075 156.565 ;
        RECT -46.405 154.875 -46.075 155.205 ;
        RECT -46.405 153.515 -46.075 153.845 ;
        RECT -46.405 152.155 -46.075 152.485 ;
        RECT -46.405 150.795 -46.075 151.125 ;
        RECT -46.405 149.435 -46.075 149.765 ;
        RECT -46.405 148.075 -46.075 148.405 ;
        RECT -46.405 146.715 -46.075 147.045 ;
        RECT -46.405 145.355 -46.075 145.685 ;
        RECT -46.405 143.995 -46.075 144.325 ;
        RECT -46.405 142.635 -46.075 142.965 ;
        RECT -46.405 141.275 -46.075 141.605 ;
        RECT -46.405 139.915 -46.075 140.245 ;
        RECT -46.405 138.555 -46.075 138.885 ;
        RECT -46.405 136.42 -46.075 136.75 ;
        RECT -46.405 134.245 -46.075 134.575 ;
        RECT -46.405 133.395 -46.075 133.725 ;
        RECT -46.405 131.085 -46.075 131.415 ;
        RECT -46.405 130.235 -46.075 130.565 ;
        RECT -46.405 127.925 -46.075 128.255 ;
        RECT -46.405 127.075 -46.075 127.405 ;
        RECT -46.405 124.765 -46.075 125.095 ;
        RECT -46.405 123.915 -46.075 124.245 ;
        RECT -46.405 121.605 -46.075 121.935 ;
        RECT -46.405 120.755 -46.075 121.085 ;
        RECT -46.405 118.445 -46.075 118.775 ;
        RECT -46.405 117.595 -46.075 117.925 ;
        RECT -46.405 115.285 -46.075 115.615 ;
        RECT -46.405 114.435 -46.075 114.765 ;
        RECT -46.405 112.125 -46.075 112.455 ;
        RECT -46.405 111.275 -46.075 111.605 ;
        RECT -46.405 108.965 -46.075 109.295 ;
        RECT -46.405 108.115 -46.075 108.445 ;
        RECT -46.405 105.805 -46.075 106.135 ;
        RECT -46.405 104.955 -46.075 105.285 ;
        RECT -46.405 102.645 -46.075 102.975 ;
        RECT -46.405 101.795 -46.075 102.125 ;
        RECT -46.405 99.62 -46.075 99.95 ;
        RECT -46.405 97.755 -46.075 98.085 ;
        RECT -46.405 96.395 -46.075 96.725 ;
        RECT -46.405 95.035 -46.075 95.365 ;
        RECT -46.405 93.675 -46.075 94.005 ;
        RECT -46.405 92.315 -46.075 92.645 ;
        RECT -46.405 90.955 -46.075 91.285 ;
        RECT -46.405 89.595 -46.075 89.925 ;
        RECT -46.405 88.235 -46.075 88.565 ;
        RECT -46.405 86.875 -46.075 87.205 ;
        RECT -46.405 85.515 -46.075 85.845 ;
        RECT -46.405 84.155 -46.075 84.485 ;
        RECT -46.405 82.795 -46.075 83.125 ;
        RECT -46.405 81.435 -46.075 81.765 ;
        RECT -46.405 80.075 -46.075 80.405 ;
        RECT -46.405 78.715 -46.075 79.045 ;
        RECT -46.405 77.355 -46.075 77.685 ;
        RECT -46.405 75.995 -46.075 76.325 ;
        RECT -46.405 74.635 -46.075 74.965 ;
        RECT -46.405 73.275 -46.075 73.605 ;
        RECT -46.405 71.915 -46.075 72.245 ;
        RECT -46.405 70.555 -46.075 70.885 ;
        RECT -46.405 69.195 -46.075 69.525 ;
        RECT -46.405 67.835 -46.075 68.165 ;
        RECT -46.405 66.475 -46.075 66.805 ;
        RECT -46.405 65.115 -46.075 65.445 ;
        RECT -46.405 63.755 -46.075 64.085 ;
        RECT -46.405 62.395 -46.075 62.725 ;
        RECT -46.405 61.035 -46.075 61.365 ;
        RECT -46.405 59.675 -46.075 60.005 ;
        RECT -46.405 58.315 -46.075 58.645 ;
        RECT -46.405 56.955 -46.075 57.285 ;
        RECT -46.405 55.595 -46.075 55.925 ;
        RECT -46.405 54.235 -46.075 54.565 ;
        RECT -46.405 52.875 -46.075 53.205 ;
        RECT -46.405 51.515 -46.075 51.845 ;
        RECT -46.405 50.155 -46.075 50.485 ;
        RECT -46.405 48.795 -46.075 49.125 ;
        RECT -46.405 47.435 -46.075 47.765 ;
        RECT -46.405 46.075 -46.075 46.405 ;
        RECT -46.405 44.715 -46.075 45.045 ;
        RECT -46.405 43.355 -46.075 43.685 ;
        RECT -46.405 41.995 -46.075 42.325 ;
        RECT -46.405 40.635 -46.075 40.965 ;
        RECT -46.405 39.275 -46.075 39.605 ;
        RECT -46.405 37.915 -46.075 38.245 ;
        RECT -46.405 36.555 -46.075 36.885 ;
        RECT -46.405 35.195 -46.075 35.525 ;
        RECT -46.405 33.835 -46.075 34.165 ;
        RECT -46.405 32.475 -46.075 32.805 ;
        RECT -46.405 31.115 -46.075 31.445 ;
        RECT -46.405 29.755 -46.075 30.085 ;
        RECT -46.405 28.395 -46.075 28.725 ;
        RECT -46.405 27.035 -46.075 27.365 ;
        RECT -46.405 25.675 -46.075 26.005 ;
        RECT -46.405 24.315 -46.075 24.645 ;
        RECT -46.405 22.955 -46.075 23.285 ;
        RECT -46.405 21.595 -46.075 21.925 ;
        RECT -46.405 20.235 -46.075 20.565 ;
        RECT -46.405 18.875 -46.075 19.205 ;
        RECT -46.405 17.515 -46.075 17.845 ;
        RECT -46.405 16.155 -46.075 16.485 ;
        RECT -46.405 14.795 -46.075 15.125 ;
        RECT -46.405 13.435 -46.075 13.765 ;
        RECT -46.405 12.075 -46.075 12.405 ;
        RECT -46.405 10.715 -46.075 11.045 ;
        RECT -46.405 9.355 -46.075 9.685 ;
        RECT -46.405 7.995 -46.075 8.325 ;
        RECT -46.405 6.635 -46.075 6.965 ;
        RECT -46.405 5.275 -46.075 5.605 ;
        RECT -46.405 3.915 -46.075 4.245 ;
        RECT -46.405 2.555 -46.075 2.885 ;
        RECT -46.405 1.195 -46.075 1.525 ;
        RECT -46.405 -0.165 -46.075 0.165 ;
        RECT -46.405 -1.525 -46.075 -1.195 ;
        RECT -46.4 -1.525 -46.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 -30.66 -46.075 -30.33 ;
        RECT -46.405 -31.445 -46.075 -31.115 ;
        RECT -46.405 -32.805 -46.075 -32.475 ;
        RECT -46.405 -34.165 -46.075 -33.835 ;
        RECT -46.405 -36.885 -46.075 -36.555 ;
        RECT -46.405 -37.85 -46.075 -37.52 ;
        RECT -46.405 -40.965 -46.075 -40.635 ;
        RECT -46.405 -46.405 -46.075 -46.075 ;
        RECT -46.405 -49.125 -46.075 -48.795 ;
        RECT -46.405 -50.485 -46.075 -50.155 ;
        RECT -46.405 -53.205 -46.075 -52.875 ;
        RECT -46.405 -55.925 -46.075 -55.595 ;
        RECT -46.405 -61.365 -46.075 -61.035 ;
        RECT -46.405 -62.725 -46.075 -62.395 ;
        RECT -46.405 -64.085 -46.075 -63.755 ;
        RECT -46.405 -65.445 -46.075 -65.115 ;
        RECT -46.405 -66.805 -46.075 -66.475 ;
        RECT -46.405 -68.165 -46.075 -67.835 ;
        RECT -46.405 -69.525 -46.075 -69.195 ;
        RECT -46.405 -70.885 -46.075 -70.555 ;
        RECT -46.405 -72.245 -46.075 -71.915 ;
        RECT -46.405 -73.605 -46.075 -73.275 ;
        RECT -46.405 -74.965 -46.075 -74.635 ;
        RECT -46.405 -76.325 -46.075 -75.995 ;
        RECT -46.405 -77.685 -46.075 -77.355 ;
        RECT -46.405 -79.045 -46.075 -78.715 ;
        RECT -46.405 -80.405 -46.075 -80.075 ;
        RECT -46.405 -81.765 -46.075 -81.435 ;
        RECT -46.405 -83.125 -46.075 -82.795 ;
        RECT -46.405 -84.485 -46.075 -84.155 ;
        RECT -46.405 -85.845 -46.075 -85.515 ;
        RECT -46.405 -87.205 -46.075 -86.875 ;
        RECT -46.405 -88.565 -46.075 -88.235 ;
        RECT -46.405 -89.925 -46.075 -89.595 ;
        RECT -46.405 -91.285 -46.075 -90.955 ;
        RECT -46.405 -92.645 -46.075 -92.315 ;
        RECT -46.405 -94.005 -46.075 -93.675 ;
        RECT -46.405 -95.365 -46.075 -95.035 ;
        RECT -46.405 -96.725 -46.075 -96.395 ;
        RECT -46.405 -98.085 -46.075 -97.755 ;
        RECT -46.405 -99.445 -46.075 -99.115 ;
        RECT -46.405 -100.805 -46.075 -100.475 ;
        RECT -46.405 -102.165 -46.075 -101.835 ;
        RECT -46.405 -103.525 -46.075 -103.195 ;
        RECT -46.405 -104.885 -46.075 -104.555 ;
        RECT -46.405 -106.245 -46.075 -105.915 ;
        RECT -46.405 -107.605 -46.075 -107.275 ;
        RECT -46.405 -108.965 -46.075 -108.635 ;
        RECT -46.405 -110.325 -46.075 -109.995 ;
        RECT -46.405 -111.685 -46.075 -111.355 ;
        RECT -46.405 -113.045 -46.075 -112.715 ;
        RECT -46.405 -114.405 -46.075 -114.075 ;
        RECT -46.405 -115.765 -46.075 -115.435 ;
        RECT -46.405 -117.125 -46.075 -116.795 ;
        RECT -46.405 -118.485 -46.075 -118.155 ;
        RECT -46.405 -119.845 -46.075 -119.515 ;
        RECT -46.405 -121.205 -46.075 -120.875 ;
        RECT -46.405 -129.365 -46.075 -129.035 ;
        RECT -46.405 -130.725 -46.075 -130.395 ;
        RECT -46.405 -131.47 -46.075 -131.14 ;
        RECT -46.405 -133.445 -46.075 -133.115 ;
        RECT -46.405 -134.805 -46.075 -134.475 ;
        RECT -46.405 -136.165 -46.075 -135.835 ;
        RECT -46.405 -137.525 -46.075 -137.195 ;
        RECT -46.405 -140.245 -46.075 -139.915 ;
        RECT -46.405 -141.605 -46.075 -141.275 ;
        RECT -46.405 -142.965 -46.075 -142.635 ;
        RECT -46.405 -144.31 -46.075 -143.98 ;
        RECT -46.405 -145.685 -46.075 -145.355 ;
        RECT -46.405 -147.045 -46.075 -146.715 ;
        RECT -46.405 -149.765 -46.075 -149.435 ;
        RECT -46.405 -152.485 -46.075 -152.155 ;
        RECT -46.405 -153.845 -46.075 -153.515 ;
        RECT -46.405 -155.205 -46.075 -154.875 ;
        RECT -46.405 -156.565 -46.075 -156.235 ;
        RECT -46.405 -157.925 -46.075 -157.595 ;
        RECT -46.405 -159.285 -46.075 -158.955 ;
        RECT -46.405 -162.005 -46.075 -161.675 ;
        RECT -46.405 -163.365 -46.075 -163.035 ;
        RECT -46.405 -164.725 -46.075 -164.395 ;
        RECT -46.405 -166.085 -46.075 -165.755 ;
        RECT -46.405 -167.445 -46.075 -167.115 ;
        RECT -46.405 -168.805 -46.075 -168.475 ;
        RECT -46.405 -170.165 -46.075 -169.835 ;
        RECT -46.405 -171.525 -46.075 -171.195 ;
        RECT -46.405 -172.885 -46.075 -172.555 ;
        RECT -46.405 -174.245 -46.075 -173.915 ;
        RECT -46.405 -175.605 -46.075 -175.275 ;
        RECT -46.405 -176.965 -46.075 -176.635 ;
        RECT -46.405 -178.325 -46.075 -177.995 ;
        RECT -46.405 -179.685 -46.075 -179.355 ;
        RECT -46.405 -181.045 -46.075 -180.715 ;
        RECT -46.405 -182.405 -46.075 -182.075 ;
        RECT -46.405 -183.765 -46.075 -183.435 ;
        RECT -46.405 -185.125 -46.075 -184.795 ;
        RECT -46.405 -186.485 -46.075 -186.155 ;
        RECT -46.405 -187.845 -46.075 -187.515 ;
        RECT -46.405 -189.205 -46.075 -188.875 ;
        RECT -46.405 -190.565 -46.075 -190.235 ;
        RECT -46.405 -191.925 -46.075 -191.595 ;
        RECT -46.405 -193.285 -46.075 -192.955 ;
        RECT -46.405 -194.645 -46.075 -194.315 ;
        RECT -46.405 -196.005 -46.075 -195.675 ;
        RECT -46.405 -197.365 -46.075 -197.035 ;
        RECT -46.405 -198.725 -46.075 -198.395 ;
        RECT -46.405 -200.085 -46.075 -199.755 ;
        RECT -46.405 -201.445 -46.075 -201.115 ;
        RECT -46.405 -202.805 -46.075 -202.475 ;
        RECT -46.405 -204.165 -46.075 -203.835 ;
        RECT -46.405 -205.525 -46.075 -205.195 ;
        RECT -46.405 -206.885 -46.075 -206.555 ;
        RECT -46.405 -208.245 -46.075 -207.915 ;
        RECT -46.405 -209.605 -46.075 -209.275 ;
        RECT -46.405 -210.965 -46.075 -210.635 ;
        RECT -46.405 -212.325 -46.075 -211.995 ;
        RECT -46.405 -213.685 -46.075 -213.355 ;
        RECT -46.405 -215.045 -46.075 -214.715 ;
        RECT -46.405 -216.405 -46.075 -216.075 ;
        RECT -46.405 -217.765 -46.075 -217.435 ;
        RECT -46.405 -219.125 -46.075 -218.795 ;
        RECT -46.405 -220.485 -46.075 -220.155 ;
        RECT -46.405 -221.845 -46.075 -221.515 ;
        RECT -46.405 -223.205 -46.075 -222.875 ;
        RECT -46.405 -224.565 -46.075 -224.235 ;
        RECT -46.405 -226.155 -46.075 -225.825 ;
        RECT -46.405 -227.285 -46.075 -226.955 ;
        RECT -46.405 -228.645 -46.075 -228.315 ;
        RECT -46.4 -229.32 -46.08 -27.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 228.315 -44.715 228.645 ;
        RECT -45.045 226.955 -44.715 227.285 ;
        RECT -45.045 225.595 -44.715 225.925 ;
        RECT -45.045 224.235 -44.715 224.565 ;
        RECT -45.045 222.875 -44.715 223.205 ;
        RECT -45.045 221.515 -44.715 221.845 ;
        RECT -45.045 220.155 -44.715 220.485 ;
        RECT -45.045 218.795 -44.715 219.125 ;
        RECT -45.045 217.435 -44.715 217.765 ;
        RECT -45.045 216.075 -44.715 216.405 ;
        RECT -45.045 214.715 -44.715 215.045 ;
        RECT -45.045 213.355 -44.715 213.685 ;
        RECT -45.045 211.995 -44.715 212.325 ;
        RECT -45.045 210.635 -44.715 210.965 ;
        RECT -45.045 209.275 -44.715 209.605 ;
        RECT -45.045 207.915 -44.715 208.245 ;
        RECT -45.045 206.555 -44.715 206.885 ;
        RECT -45.045 205.195 -44.715 205.525 ;
        RECT -45.045 203.835 -44.715 204.165 ;
        RECT -45.045 202.475 -44.715 202.805 ;
        RECT -45.045 201.115 -44.715 201.445 ;
        RECT -45.045 199.755 -44.715 200.085 ;
        RECT -45.045 198.395 -44.715 198.725 ;
        RECT -45.045 197.035 -44.715 197.365 ;
        RECT -45.045 195.675 -44.715 196.005 ;
        RECT -45.045 194.315 -44.715 194.645 ;
        RECT -45.045 192.955 -44.715 193.285 ;
        RECT -45.045 191.595 -44.715 191.925 ;
        RECT -45.045 190.235 -44.715 190.565 ;
        RECT -45.045 188.875 -44.715 189.205 ;
        RECT -45.045 187.515 -44.715 187.845 ;
        RECT -45.045 186.155 -44.715 186.485 ;
        RECT -45.045 184.795 -44.715 185.125 ;
        RECT -45.045 183.435 -44.715 183.765 ;
        RECT -45.045 182.075 -44.715 182.405 ;
        RECT -45.045 180.715 -44.715 181.045 ;
        RECT -45.045 179.355 -44.715 179.685 ;
        RECT -45.045 177.995 -44.715 178.325 ;
        RECT -45.045 176.635 -44.715 176.965 ;
        RECT -45.045 175.275 -44.715 175.605 ;
        RECT -45.045 173.915 -44.715 174.245 ;
        RECT -45.045 172.555 -44.715 172.885 ;
        RECT -45.045 171.195 -44.715 171.525 ;
        RECT -45.045 169.835 -44.715 170.165 ;
        RECT -45.045 168.475 -44.715 168.805 ;
        RECT -45.045 167.115 -44.715 167.445 ;
        RECT -45.045 165.755 -44.715 166.085 ;
        RECT -45.045 164.395 -44.715 164.725 ;
        RECT -45.045 163.035 -44.715 163.365 ;
        RECT -45.045 161.675 -44.715 162.005 ;
        RECT -45.045 160.315 -44.715 160.645 ;
        RECT -45.045 158.955 -44.715 159.285 ;
        RECT -45.045 157.595 -44.715 157.925 ;
        RECT -45.045 156.235 -44.715 156.565 ;
        RECT -45.045 154.875 -44.715 155.205 ;
        RECT -45.045 153.515 -44.715 153.845 ;
        RECT -45.045 152.155 -44.715 152.485 ;
        RECT -45.045 150.795 -44.715 151.125 ;
        RECT -45.045 149.435 -44.715 149.765 ;
        RECT -45.045 148.075 -44.715 148.405 ;
        RECT -45.045 146.715 -44.715 147.045 ;
        RECT -45.045 145.355 -44.715 145.685 ;
        RECT -45.045 143.995 -44.715 144.325 ;
        RECT -45.045 142.635 -44.715 142.965 ;
        RECT -45.045 141.275 -44.715 141.605 ;
        RECT -45.045 139.915 -44.715 140.245 ;
        RECT -45.045 138.555 -44.715 138.885 ;
        RECT -45.045 136.42 -44.715 136.75 ;
        RECT -45.045 134.245 -44.715 134.575 ;
        RECT -45.045 133.395 -44.715 133.725 ;
        RECT -45.045 131.085 -44.715 131.415 ;
        RECT -45.045 130.235 -44.715 130.565 ;
        RECT -45.045 127.925 -44.715 128.255 ;
        RECT -45.045 127.075 -44.715 127.405 ;
        RECT -45.045 124.765 -44.715 125.095 ;
        RECT -45.045 123.915 -44.715 124.245 ;
        RECT -45.045 121.605 -44.715 121.935 ;
        RECT -45.045 120.755 -44.715 121.085 ;
        RECT -45.045 118.445 -44.715 118.775 ;
        RECT -45.045 117.595 -44.715 117.925 ;
        RECT -45.045 115.285 -44.715 115.615 ;
        RECT -45.045 114.435 -44.715 114.765 ;
        RECT -45.045 112.125 -44.715 112.455 ;
        RECT -45.045 111.275 -44.715 111.605 ;
        RECT -45.045 108.965 -44.715 109.295 ;
        RECT -45.045 108.115 -44.715 108.445 ;
        RECT -45.045 105.805 -44.715 106.135 ;
        RECT -45.045 104.955 -44.715 105.285 ;
        RECT -45.045 102.645 -44.715 102.975 ;
        RECT -45.045 101.795 -44.715 102.125 ;
        RECT -45.045 99.62 -44.715 99.95 ;
        RECT -45.045 97.755 -44.715 98.085 ;
        RECT -45.045 96.395 -44.715 96.725 ;
        RECT -45.045 95.035 -44.715 95.365 ;
        RECT -45.045 93.675 -44.715 94.005 ;
        RECT -45.045 92.315 -44.715 92.645 ;
        RECT -45.045 90.955 -44.715 91.285 ;
        RECT -45.045 89.595 -44.715 89.925 ;
        RECT -45.045 88.235 -44.715 88.565 ;
        RECT -45.045 86.875 -44.715 87.205 ;
        RECT -45.045 85.515 -44.715 85.845 ;
        RECT -45.045 84.155 -44.715 84.485 ;
        RECT -45.045 82.795 -44.715 83.125 ;
        RECT -45.045 81.435 -44.715 81.765 ;
        RECT -45.045 80.075 -44.715 80.405 ;
        RECT -45.045 78.715 -44.715 79.045 ;
        RECT -45.045 77.355 -44.715 77.685 ;
        RECT -45.045 75.995 -44.715 76.325 ;
        RECT -45.045 74.635 -44.715 74.965 ;
        RECT -45.045 73.275 -44.715 73.605 ;
        RECT -45.045 71.915 -44.715 72.245 ;
        RECT -45.045 70.555 -44.715 70.885 ;
        RECT -45.045 69.195 -44.715 69.525 ;
        RECT -45.045 67.835 -44.715 68.165 ;
        RECT -45.045 66.475 -44.715 66.805 ;
        RECT -45.045 65.115 -44.715 65.445 ;
        RECT -45.045 63.755 -44.715 64.085 ;
        RECT -45.045 62.395 -44.715 62.725 ;
        RECT -45.045 61.035 -44.715 61.365 ;
        RECT -45.045 59.675 -44.715 60.005 ;
        RECT -45.045 58.315 -44.715 58.645 ;
        RECT -45.045 56.955 -44.715 57.285 ;
        RECT -45.045 55.595 -44.715 55.925 ;
        RECT -45.045 54.235 -44.715 54.565 ;
        RECT -45.045 52.875 -44.715 53.205 ;
        RECT -45.045 51.515 -44.715 51.845 ;
        RECT -45.045 50.155 -44.715 50.485 ;
        RECT -45.045 48.795 -44.715 49.125 ;
        RECT -45.045 47.435 -44.715 47.765 ;
        RECT -45.045 46.075 -44.715 46.405 ;
        RECT -45.045 44.715 -44.715 45.045 ;
        RECT -45.045 43.355 -44.715 43.685 ;
        RECT -45.045 41.995 -44.715 42.325 ;
        RECT -45.045 40.635 -44.715 40.965 ;
        RECT -45.045 39.275 -44.715 39.605 ;
        RECT -45.045 37.915 -44.715 38.245 ;
        RECT -45.045 36.555 -44.715 36.885 ;
        RECT -45.045 35.195 -44.715 35.525 ;
        RECT -45.045 33.835 -44.715 34.165 ;
        RECT -45.045 32.475 -44.715 32.805 ;
        RECT -45.045 31.115 -44.715 31.445 ;
        RECT -45.045 29.755 -44.715 30.085 ;
        RECT -45.045 28.395 -44.715 28.725 ;
        RECT -45.045 27.035 -44.715 27.365 ;
        RECT -45.045 25.675 -44.715 26.005 ;
        RECT -45.045 24.315 -44.715 24.645 ;
        RECT -45.045 22.955 -44.715 23.285 ;
        RECT -45.045 21.595 -44.715 21.925 ;
        RECT -45.045 20.235 -44.715 20.565 ;
        RECT -45.045 18.875 -44.715 19.205 ;
        RECT -45.045 17.515 -44.715 17.845 ;
        RECT -45.045 16.155 -44.715 16.485 ;
        RECT -45.045 14.795 -44.715 15.125 ;
        RECT -45.045 13.435 -44.715 13.765 ;
        RECT -45.045 12.075 -44.715 12.405 ;
        RECT -45.045 10.715 -44.715 11.045 ;
        RECT -45.045 9.355 -44.715 9.685 ;
        RECT -45.045 7.995 -44.715 8.325 ;
        RECT -45.045 6.635 -44.715 6.965 ;
        RECT -45.045 5.275 -44.715 5.605 ;
        RECT -45.045 3.915 -44.715 4.245 ;
        RECT -45.045 2.555 -44.715 2.885 ;
        RECT -45.045 1.195 -44.715 1.525 ;
        RECT -45.045 -0.165 -44.715 0.165 ;
        RECT -45.045 -1.525 -44.715 -1.195 ;
        RECT -45.045 -4.245 -44.715 -3.915 ;
        RECT -45.045 -5.605 -44.715 -5.275 ;
        RECT -45.045 -6.965 -44.715 -6.635 ;
        RECT -45.045 -8.325 -44.715 -7.995 ;
        RECT -45.045 -9.685 -44.715 -9.355 ;
        RECT -45.045 -12.405 -44.715 -12.075 ;
        RECT -45.045 -13.765 -44.715 -13.435 ;
        RECT -45.045 -15.125 -44.715 -14.795 ;
        RECT -45.045 -16.485 -44.715 -16.155 ;
        RECT -45.045 -17.845 -44.715 -17.515 ;
        RECT -45.045 -19.205 -44.715 -18.875 ;
        RECT -45.045 -20.565 -44.715 -20.235 ;
        RECT -45.045 -21.925 -44.715 -21.595 ;
        RECT -45.045 -23.285 -44.715 -22.955 ;
        RECT -45.045 -24.645 -44.715 -24.315 ;
        RECT -45.045 -30.66 -44.715 -30.33 ;
        RECT -45.045 -31.445 -44.715 -31.115 ;
        RECT -45.045 -32.805 -44.715 -32.475 ;
        RECT -45.045 -34.165 -44.715 -33.835 ;
        RECT -45.045 -36.885 -44.715 -36.555 ;
        RECT -45.045 -37.85 -44.715 -37.52 ;
        RECT -45.045 -40.965 -44.715 -40.635 ;
        RECT -45.045 -46.405 -44.715 -46.075 ;
        RECT -45.045 -49.125 -44.715 -48.795 ;
        RECT -45.045 -50.485 -44.715 -50.155 ;
        RECT -45.045 -53.205 -44.715 -52.875 ;
        RECT -45.045 -55.925 -44.715 -55.595 ;
        RECT -45.04 -59.32 -44.72 248.005 ;
        RECT -45.045 246.76 -44.715 247.89 ;
        RECT -45.045 241.915 -44.715 242.245 ;
        RECT -45.045 240.555 -44.715 240.885 ;
        RECT -45.045 239.195 -44.715 239.525 ;
        RECT -45.045 237.835 -44.715 238.165 ;
        RECT -45.045 236.475 -44.715 236.805 ;
        RECT -45.045 235.115 -44.715 235.445 ;
        RECT -45.045 233.755 -44.715 234.085 ;
        RECT -45.045 232.395 -44.715 232.725 ;
        RECT -45.045 231.035 -44.715 231.365 ;
        RECT -45.045 229.675 -44.715 230.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 97.755 -54.235 98.085 ;
        RECT -54.565 96.395 -54.235 96.725 ;
        RECT -54.565 95.035 -54.235 95.365 ;
        RECT -54.565 93.675 -54.235 94.005 ;
        RECT -54.565 92.315 -54.235 92.645 ;
        RECT -54.565 89.595 -54.235 89.925 ;
        RECT -54.565 88.235 -54.235 88.565 ;
        RECT -54.565 84.155 -54.235 84.485 ;
        RECT -54.565 82.795 -54.235 83.125 ;
        RECT -54.565 81.435 -54.235 81.765 ;
        RECT -54.565 80.075 -54.235 80.405 ;
        RECT -54.565 78.715 -54.235 79.045 ;
        RECT -54.565 77.355 -54.235 77.685 ;
        RECT -54.565 75.995 -54.235 76.325 ;
        RECT -54.565 74.635 -54.235 74.965 ;
        RECT -54.565 73.275 -54.235 73.605 ;
        RECT -54.565 71.915 -54.235 72.245 ;
        RECT -54.565 70.555 -54.235 70.885 ;
        RECT -54.565 69.195 -54.235 69.525 ;
        RECT -54.565 67.835 -54.235 68.165 ;
        RECT -54.565 66.475 -54.235 66.805 ;
        RECT -54.565 65.115 -54.235 65.445 ;
        RECT -54.565 63.755 -54.235 64.085 ;
        RECT -54.565 62.395 -54.235 62.725 ;
        RECT -54.565 61.035 -54.235 61.365 ;
        RECT -54.565 59.675 -54.235 60.005 ;
        RECT -54.565 58.315 -54.235 58.645 ;
        RECT -54.565 56.955 -54.235 57.285 ;
        RECT -54.565 55.595 -54.235 55.925 ;
        RECT -54.565 54.235 -54.235 54.565 ;
        RECT -54.565 52.875 -54.235 53.205 ;
        RECT -54.565 51.515 -54.235 51.845 ;
        RECT -54.565 50.155 -54.235 50.485 ;
        RECT -54.565 48.795 -54.235 49.125 ;
        RECT -54.565 47.435 -54.235 47.765 ;
        RECT -54.565 46.075 -54.235 46.405 ;
        RECT -54.565 44.715 -54.235 45.045 ;
        RECT -54.565 43.355 -54.235 43.685 ;
        RECT -54.565 41.995 -54.235 42.325 ;
        RECT -54.565 40.635 -54.235 40.965 ;
        RECT -54.565 39.275 -54.235 39.605 ;
        RECT -54.565 37.915 -54.235 38.245 ;
        RECT -54.565 36.555 -54.235 36.885 ;
        RECT -54.565 35.195 -54.235 35.525 ;
        RECT -54.565 33.835 -54.235 34.165 ;
        RECT -54.565 32.475 -54.235 32.805 ;
        RECT -54.565 31.115 -54.235 31.445 ;
        RECT -54.565 29.755 -54.235 30.085 ;
        RECT -54.565 28.395 -54.235 28.725 ;
        RECT -54.565 27.035 -54.235 27.365 ;
        RECT -54.565 25.675 -54.235 26.005 ;
        RECT -54.565 24.315 -54.235 24.645 ;
        RECT -54.565 22.955 -54.235 23.285 ;
        RECT -54.565 21.595 -54.235 21.925 ;
        RECT -54.565 20.235 -54.235 20.565 ;
        RECT -54.565 18.875 -54.235 19.205 ;
        RECT -54.565 17.515 -54.235 17.845 ;
        RECT -54.565 16.155 -54.235 16.485 ;
        RECT -54.565 14.795 -54.235 15.125 ;
        RECT -54.565 13.435 -54.235 13.765 ;
        RECT -54.565 12.075 -54.235 12.405 ;
        RECT -54.565 10.715 -54.235 11.045 ;
        RECT -54.565 9.355 -54.235 9.685 ;
        RECT -54.565 7.995 -54.235 8.325 ;
        RECT -54.565 6.635 -54.235 6.965 ;
        RECT -54.565 5.275 -54.235 5.605 ;
        RECT -54.565 3.915 -54.235 4.245 ;
        RECT -54.565 2.555 -54.235 2.885 ;
        RECT -54.565 1.195 -54.235 1.525 ;
        RECT -54.565 -0.165 -54.235 0.165 ;
        RECT -54.565 -1.525 -54.235 -1.195 ;
        RECT -54.565 -2.885 -54.235 -2.555 ;
        RECT -54.565 -4.245 -54.235 -3.915 ;
        RECT -54.565 -5.605 -54.235 -5.275 ;
        RECT -54.565 -6.965 -54.235 -6.635 ;
        RECT -54.565 -8.325 -54.235 -7.995 ;
        RECT -54.565 -9.685 -54.235 -9.355 ;
        RECT -54.565 -12.405 -54.235 -12.075 ;
        RECT -54.565 -13.765 -54.235 -13.435 ;
        RECT -54.565 -15.125 -54.235 -14.795 ;
        RECT -54.565 -16.485 -54.235 -16.155 ;
        RECT -54.565 -17.845 -54.235 -17.515 ;
        RECT -54.565 -19.205 -54.235 -18.875 ;
        RECT -54.565 -20.565 -54.235 -20.235 ;
        RECT -54.565 -21.925 -54.235 -21.595 ;
        RECT -54.565 -23.285 -54.235 -22.955 ;
        RECT -54.565 -24.645 -54.235 -24.315 ;
        RECT -54.565 -26.005 -54.235 -25.675 ;
        RECT -54.565 -27.365 -54.235 -27.035 ;
        RECT -54.565 -28.725 -54.235 -28.395 ;
        RECT -54.565 -30.085 -54.235 -29.755 ;
        RECT -54.565 -31.445 -54.235 -31.115 ;
        RECT -54.565 -32.805 -54.235 -32.475 ;
        RECT -54.565 -34.165 -54.235 -33.835 ;
        RECT -54.565 -35.525 -54.235 -35.195 ;
        RECT -54.565 -36.885 -54.235 -36.555 ;
        RECT -54.565 -38.245 -54.235 -37.915 ;
        RECT -54.565 -39.605 -54.235 -39.275 ;
        RECT -54.565 -40.965 -54.235 -40.635 ;
        RECT -54.565 -42.325 -54.235 -41.995 ;
        RECT -54.565 -43.685 -54.235 -43.355 ;
        RECT -54.565 -45.045 -54.235 -44.715 ;
        RECT -54.565 -46.405 -54.235 -46.075 ;
        RECT -54.565 -47.765 -54.235 -47.435 ;
        RECT -54.565 -49.125 -54.235 -48.795 ;
        RECT -54.565 -50.485 -54.235 -50.155 ;
        RECT -54.565 -51.845 -54.235 -51.515 ;
        RECT -54.565 -53.205 -54.235 -52.875 ;
        RECT -54.565 -54.565 -54.235 -54.235 ;
        RECT -54.565 -55.925 -54.235 -55.595 ;
        RECT -54.565 -57.285 -54.235 -56.955 ;
        RECT -54.565 -58.645 -54.235 -58.315 ;
        RECT -54.565 -60.005 -54.235 -59.675 ;
        RECT -54.565 -61.365 -54.235 -61.035 ;
        RECT -54.565 -62.725 -54.235 -62.395 ;
        RECT -54.565 -64.085 -54.235 -63.755 ;
        RECT -54.565 -65.445 -54.235 -65.115 ;
        RECT -54.565 -66.805 -54.235 -66.475 ;
        RECT -54.565 -68.165 -54.235 -67.835 ;
        RECT -54.565 -69.525 -54.235 -69.195 ;
        RECT -54.565 -70.885 -54.235 -70.555 ;
        RECT -54.565 -72.245 -54.235 -71.915 ;
        RECT -54.565 -73.605 -54.235 -73.275 ;
        RECT -54.565 -74.965 -54.235 -74.635 ;
        RECT -54.565 -76.325 -54.235 -75.995 ;
        RECT -54.565 -77.685 -54.235 -77.355 ;
        RECT -54.565 -79.045 -54.235 -78.715 ;
        RECT -54.565 -80.405 -54.235 -80.075 ;
        RECT -54.565 -81.765 -54.235 -81.435 ;
        RECT -54.565 -83.125 -54.235 -82.795 ;
        RECT -54.565 -84.485 -54.235 -84.155 ;
        RECT -54.565 -85.845 -54.235 -85.515 ;
        RECT -54.565 -87.205 -54.235 -86.875 ;
        RECT -54.565 -88.565 -54.235 -88.235 ;
        RECT -54.565 -89.925 -54.235 -89.595 ;
        RECT -54.565 -91.285 -54.235 -90.955 ;
        RECT -54.565 -92.645 -54.235 -92.315 ;
        RECT -54.565 -94.005 -54.235 -93.675 ;
        RECT -54.565 -95.365 -54.235 -95.035 ;
        RECT -54.565 -96.725 -54.235 -96.395 ;
        RECT -54.565 -98.085 -54.235 -97.755 ;
        RECT -54.565 -99.445 -54.235 -99.115 ;
        RECT -54.565 -100.805 -54.235 -100.475 ;
        RECT -54.565 -102.165 -54.235 -101.835 ;
        RECT -54.565 -103.525 -54.235 -103.195 ;
        RECT -54.565 -104.885 -54.235 -104.555 ;
        RECT -54.565 -106.245 -54.235 -105.915 ;
        RECT -54.565 -107.605 -54.235 -107.275 ;
        RECT -54.565 -108.965 -54.235 -108.635 ;
        RECT -54.565 -110.325 -54.235 -109.995 ;
        RECT -54.565 -111.685 -54.235 -111.355 ;
        RECT -54.565 -113.045 -54.235 -112.715 ;
        RECT -54.565 -114.405 -54.235 -114.075 ;
        RECT -54.565 -115.765 -54.235 -115.435 ;
        RECT -54.565 -117.125 -54.235 -116.795 ;
        RECT -54.565 -118.485 -54.235 -118.155 ;
        RECT -54.565 -119.845 -54.235 -119.515 ;
        RECT -54.565 -121.205 -54.235 -120.875 ;
        RECT -54.565 -122.565 -54.235 -122.235 ;
        RECT -54.565 -123.925 -54.235 -123.595 ;
        RECT -54.565 -129.365 -54.235 -129.035 ;
        RECT -54.565 -130.725 -54.235 -130.395 ;
        RECT -54.565 -131.47 -54.235 -131.14 ;
        RECT -54.565 -133.445 -54.235 -133.115 ;
        RECT -54.565 -134.805 -54.235 -134.475 ;
        RECT -54.565 -136.165 -54.235 -135.835 ;
        RECT -54.565 -137.525 -54.235 -137.195 ;
        RECT -54.565 -140.245 -54.235 -139.915 ;
        RECT -54.565 -141.605 -54.235 -141.275 ;
        RECT -54.565 -142.965 -54.235 -142.635 ;
        RECT -54.565 -144.31 -54.235 -143.98 ;
        RECT -54.565 -145.685 -54.235 -145.355 ;
        RECT -54.565 -147.045 -54.235 -146.715 ;
        RECT -54.565 -149.765 -54.235 -149.435 ;
        RECT -54.56 -151.8 -54.24 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 -234.085 -54.235 -233.755 ;
        RECT -54.565 -235.445 -54.235 -235.115 ;
        RECT -54.565 -236.805 -54.235 -236.475 ;
        RECT -54.565 -238.165 -54.235 -237.835 ;
        RECT -54.565 -243.81 -54.235 -242.68 ;
        RECT -54.56 -243.925 -54.24 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 246.76 -52.875 247.89 ;
        RECT -53.205 241.915 -52.875 242.245 ;
        RECT -53.205 240.555 -52.875 240.885 ;
        RECT -53.205 239.195 -52.875 239.525 ;
        RECT -53.205 237.835 -52.875 238.165 ;
        RECT -53.205 236.475 -52.875 236.805 ;
        RECT -53.205 235.115 -52.875 235.445 ;
        RECT -53.205 233.755 -52.875 234.085 ;
        RECT -53.205 232.395 -52.875 232.725 ;
        RECT -53.205 231.035 -52.875 231.365 ;
        RECT -53.205 229.675 -52.875 230.005 ;
        RECT -53.205 228.315 -52.875 228.645 ;
        RECT -53.205 226.955 -52.875 227.285 ;
        RECT -53.205 225.595 -52.875 225.925 ;
        RECT -53.205 224.235 -52.875 224.565 ;
        RECT -53.205 222.875 -52.875 223.205 ;
        RECT -53.205 221.515 -52.875 221.845 ;
        RECT -53.205 220.155 -52.875 220.485 ;
        RECT -53.205 218.795 -52.875 219.125 ;
        RECT -53.205 217.435 -52.875 217.765 ;
        RECT -53.205 216.075 -52.875 216.405 ;
        RECT -53.205 214.715 -52.875 215.045 ;
        RECT -53.205 213.355 -52.875 213.685 ;
        RECT -53.205 211.995 -52.875 212.325 ;
        RECT -53.205 210.635 -52.875 210.965 ;
        RECT -53.205 209.275 -52.875 209.605 ;
        RECT -53.205 207.915 -52.875 208.245 ;
        RECT -53.205 206.555 -52.875 206.885 ;
        RECT -53.205 205.195 -52.875 205.525 ;
        RECT -53.205 203.835 -52.875 204.165 ;
        RECT -53.205 202.475 -52.875 202.805 ;
        RECT -53.205 201.115 -52.875 201.445 ;
        RECT -53.205 199.755 -52.875 200.085 ;
        RECT -53.205 198.395 -52.875 198.725 ;
        RECT -53.205 197.035 -52.875 197.365 ;
        RECT -53.205 195.675 -52.875 196.005 ;
        RECT -53.205 194.315 -52.875 194.645 ;
        RECT -53.205 192.955 -52.875 193.285 ;
        RECT -53.205 191.595 -52.875 191.925 ;
        RECT -53.205 190.235 -52.875 190.565 ;
        RECT -53.205 188.875 -52.875 189.205 ;
        RECT -53.205 187.515 -52.875 187.845 ;
        RECT -53.205 186.155 -52.875 186.485 ;
        RECT -53.205 184.795 -52.875 185.125 ;
        RECT -53.205 183.435 -52.875 183.765 ;
        RECT -53.205 182.075 -52.875 182.405 ;
        RECT -53.205 180.715 -52.875 181.045 ;
        RECT -53.205 179.355 -52.875 179.685 ;
        RECT -53.205 177.995 -52.875 178.325 ;
        RECT -53.205 176.635 -52.875 176.965 ;
        RECT -53.205 175.275 -52.875 175.605 ;
        RECT -53.205 173.915 -52.875 174.245 ;
        RECT -53.205 172.555 -52.875 172.885 ;
        RECT -53.205 171.195 -52.875 171.525 ;
        RECT -53.205 169.835 -52.875 170.165 ;
        RECT -53.205 168.475 -52.875 168.805 ;
        RECT -53.205 167.115 -52.875 167.445 ;
        RECT -53.205 165.755 -52.875 166.085 ;
        RECT -53.205 164.395 -52.875 164.725 ;
        RECT -53.205 163.035 -52.875 163.365 ;
        RECT -53.205 161.675 -52.875 162.005 ;
        RECT -53.205 160.315 -52.875 160.645 ;
        RECT -53.205 158.955 -52.875 159.285 ;
        RECT -53.205 157.595 -52.875 157.925 ;
        RECT -53.205 156.235 -52.875 156.565 ;
        RECT -53.205 154.875 -52.875 155.205 ;
        RECT -53.205 153.515 -52.875 153.845 ;
        RECT -53.205 152.155 -52.875 152.485 ;
        RECT -53.205 150.795 -52.875 151.125 ;
        RECT -53.205 149.435 -52.875 149.765 ;
        RECT -53.205 148.075 -52.875 148.405 ;
        RECT -53.205 146.715 -52.875 147.045 ;
        RECT -53.205 145.355 -52.875 145.685 ;
        RECT -53.205 143.995 -52.875 144.325 ;
        RECT -53.205 142.635 -52.875 142.965 ;
        RECT -53.205 141.275 -52.875 141.605 ;
        RECT -53.205 139.915 -52.875 140.245 ;
        RECT -53.205 138.555 -52.875 138.885 ;
        RECT -53.2 138.555 -52.88 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 97.755 -52.875 98.085 ;
        RECT -53.205 96.395 -52.875 96.725 ;
        RECT -53.205 95.035 -52.875 95.365 ;
        RECT -53.205 93.675 -52.875 94.005 ;
        RECT -53.205 92.315 -52.875 92.645 ;
        RECT -53.205 89.595 -52.875 89.925 ;
        RECT -53.205 88.235 -52.875 88.565 ;
        RECT -53.205 84.155 -52.875 84.485 ;
        RECT -53.205 82.795 -52.875 83.125 ;
        RECT -53.205 81.435 -52.875 81.765 ;
        RECT -53.205 80.075 -52.875 80.405 ;
        RECT -53.205 78.715 -52.875 79.045 ;
        RECT -53.205 77.355 -52.875 77.685 ;
        RECT -53.205 75.995 -52.875 76.325 ;
        RECT -53.205 74.635 -52.875 74.965 ;
        RECT -53.205 73.275 -52.875 73.605 ;
        RECT -53.205 71.915 -52.875 72.245 ;
        RECT -53.205 70.555 -52.875 70.885 ;
        RECT -53.205 69.195 -52.875 69.525 ;
        RECT -53.205 67.835 -52.875 68.165 ;
        RECT -53.205 66.475 -52.875 66.805 ;
        RECT -53.205 65.115 -52.875 65.445 ;
        RECT -53.205 63.755 -52.875 64.085 ;
        RECT -53.205 62.395 -52.875 62.725 ;
        RECT -53.205 61.035 -52.875 61.365 ;
        RECT -53.205 59.675 -52.875 60.005 ;
        RECT -53.205 58.315 -52.875 58.645 ;
        RECT -53.205 56.955 -52.875 57.285 ;
        RECT -53.205 55.595 -52.875 55.925 ;
        RECT -53.205 54.235 -52.875 54.565 ;
        RECT -53.205 52.875 -52.875 53.205 ;
        RECT -53.205 51.515 -52.875 51.845 ;
        RECT -53.205 50.155 -52.875 50.485 ;
        RECT -53.205 48.795 -52.875 49.125 ;
        RECT -53.205 47.435 -52.875 47.765 ;
        RECT -53.205 46.075 -52.875 46.405 ;
        RECT -53.205 44.715 -52.875 45.045 ;
        RECT -53.205 43.355 -52.875 43.685 ;
        RECT -53.205 41.995 -52.875 42.325 ;
        RECT -53.205 40.635 -52.875 40.965 ;
        RECT -53.205 39.275 -52.875 39.605 ;
        RECT -53.205 37.915 -52.875 38.245 ;
        RECT -53.205 36.555 -52.875 36.885 ;
        RECT -53.205 35.195 -52.875 35.525 ;
        RECT -53.205 33.835 -52.875 34.165 ;
        RECT -53.205 32.475 -52.875 32.805 ;
        RECT -53.205 31.115 -52.875 31.445 ;
        RECT -53.205 29.755 -52.875 30.085 ;
        RECT -53.205 28.395 -52.875 28.725 ;
        RECT -53.205 27.035 -52.875 27.365 ;
        RECT -53.205 25.675 -52.875 26.005 ;
        RECT -53.205 24.315 -52.875 24.645 ;
        RECT -53.205 22.955 -52.875 23.285 ;
        RECT -53.205 21.595 -52.875 21.925 ;
        RECT -53.205 20.235 -52.875 20.565 ;
        RECT -53.205 18.875 -52.875 19.205 ;
        RECT -53.205 17.515 -52.875 17.845 ;
        RECT -53.205 16.155 -52.875 16.485 ;
        RECT -53.205 14.795 -52.875 15.125 ;
        RECT -53.205 13.435 -52.875 13.765 ;
        RECT -53.205 12.075 -52.875 12.405 ;
        RECT -53.205 10.715 -52.875 11.045 ;
        RECT -53.205 9.355 -52.875 9.685 ;
        RECT -53.205 7.995 -52.875 8.325 ;
        RECT -53.205 6.635 -52.875 6.965 ;
        RECT -53.205 5.275 -52.875 5.605 ;
        RECT -53.205 3.915 -52.875 4.245 ;
        RECT -53.205 2.555 -52.875 2.885 ;
        RECT -53.205 1.195 -52.875 1.525 ;
        RECT -53.205 -0.165 -52.875 0.165 ;
        RECT -53.205 -1.525 -52.875 -1.195 ;
        RECT -53.205 -2.885 -52.875 -2.555 ;
        RECT -53.205 -4.245 -52.875 -3.915 ;
        RECT -53.205 -5.605 -52.875 -5.275 ;
        RECT -53.205 -6.965 -52.875 -6.635 ;
        RECT -53.205 -8.325 -52.875 -7.995 ;
        RECT -53.205 -9.685 -52.875 -9.355 ;
        RECT -53.205 -12.405 -52.875 -12.075 ;
        RECT -53.205 -13.765 -52.875 -13.435 ;
        RECT -53.205 -15.125 -52.875 -14.795 ;
        RECT -53.205 -16.485 -52.875 -16.155 ;
        RECT -53.205 -17.845 -52.875 -17.515 ;
        RECT -53.205 -19.205 -52.875 -18.875 ;
        RECT -53.205 -20.565 -52.875 -20.235 ;
        RECT -53.205 -21.925 -52.875 -21.595 ;
        RECT -53.205 -23.285 -52.875 -22.955 ;
        RECT -53.205 -24.645 -52.875 -24.315 ;
        RECT -53.205 -26.005 -52.875 -25.675 ;
        RECT -53.205 -27.365 -52.875 -27.035 ;
        RECT -53.205 -28.725 -52.875 -28.395 ;
        RECT -53.205 -30.085 -52.875 -29.755 ;
        RECT -53.205 -31.445 -52.875 -31.115 ;
        RECT -53.205 -32.805 -52.875 -32.475 ;
        RECT -53.205 -34.165 -52.875 -33.835 ;
        RECT -53.205 -35.525 -52.875 -35.195 ;
        RECT -53.205 -36.885 -52.875 -36.555 ;
        RECT -53.205 -38.245 -52.875 -37.915 ;
        RECT -53.205 -39.605 -52.875 -39.275 ;
        RECT -53.205 -40.965 -52.875 -40.635 ;
        RECT -53.205 -42.325 -52.875 -41.995 ;
        RECT -53.205 -43.685 -52.875 -43.355 ;
        RECT -53.205 -45.045 -52.875 -44.715 ;
        RECT -53.205 -46.405 -52.875 -46.075 ;
        RECT -53.205 -47.765 -52.875 -47.435 ;
        RECT -53.205 -49.125 -52.875 -48.795 ;
        RECT -53.205 -50.485 -52.875 -50.155 ;
        RECT -53.205 -51.845 -52.875 -51.515 ;
        RECT -53.205 -53.205 -52.875 -52.875 ;
        RECT -53.205 -54.565 -52.875 -54.235 ;
        RECT -53.205 -55.925 -52.875 -55.595 ;
        RECT -53.205 -57.285 -52.875 -56.955 ;
        RECT -53.205 -58.645 -52.875 -58.315 ;
        RECT -53.205 -60.005 -52.875 -59.675 ;
        RECT -53.205 -61.365 -52.875 -61.035 ;
        RECT -53.205 -62.725 -52.875 -62.395 ;
        RECT -53.205 -64.085 -52.875 -63.755 ;
        RECT -53.205 -65.445 -52.875 -65.115 ;
        RECT -53.205 -66.805 -52.875 -66.475 ;
        RECT -53.205 -68.165 -52.875 -67.835 ;
        RECT -53.205 -69.525 -52.875 -69.195 ;
        RECT -53.205 -70.885 -52.875 -70.555 ;
        RECT -53.205 -72.245 -52.875 -71.915 ;
        RECT -53.205 -73.605 -52.875 -73.275 ;
        RECT -53.205 -74.965 -52.875 -74.635 ;
        RECT -53.205 -76.325 -52.875 -75.995 ;
        RECT -53.205 -77.685 -52.875 -77.355 ;
        RECT -53.205 -79.045 -52.875 -78.715 ;
        RECT -53.205 -80.405 -52.875 -80.075 ;
        RECT -53.205 -81.765 -52.875 -81.435 ;
        RECT -53.205 -83.125 -52.875 -82.795 ;
        RECT -53.205 -84.485 -52.875 -84.155 ;
        RECT -53.205 -85.845 -52.875 -85.515 ;
        RECT -53.205 -87.205 -52.875 -86.875 ;
        RECT -53.205 -88.565 -52.875 -88.235 ;
        RECT -53.205 -89.925 -52.875 -89.595 ;
        RECT -53.205 -91.285 -52.875 -90.955 ;
        RECT -53.205 -92.645 -52.875 -92.315 ;
        RECT -53.205 -94.005 -52.875 -93.675 ;
        RECT -53.205 -95.365 -52.875 -95.035 ;
        RECT -53.205 -96.725 -52.875 -96.395 ;
        RECT -53.205 -98.085 -52.875 -97.755 ;
        RECT -53.205 -99.445 -52.875 -99.115 ;
        RECT -53.205 -100.805 -52.875 -100.475 ;
        RECT -53.205 -102.165 -52.875 -101.835 ;
        RECT -53.205 -103.525 -52.875 -103.195 ;
        RECT -53.205 -104.885 -52.875 -104.555 ;
        RECT -53.205 -106.245 -52.875 -105.915 ;
        RECT -53.205 -107.605 -52.875 -107.275 ;
        RECT -53.205 -108.965 -52.875 -108.635 ;
        RECT -53.205 -110.325 -52.875 -109.995 ;
        RECT -53.205 -111.685 -52.875 -111.355 ;
        RECT -53.205 -113.045 -52.875 -112.715 ;
        RECT -53.205 -114.405 -52.875 -114.075 ;
        RECT -53.205 -115.765 -52.875 -115.435 ;
        RECT -53.205 -117.125 -52.875 -116.795 ;
        RECT -53.205 -118.485 -52.875 -118.155 ;
        RECT -53.205 -119.845 -52.875 -119.515 ;
        RECT -53.205 -121.205 -52.875 -120.875 ;
        RECT -53.205 -122.565 -52.875 -122.235 ;
        RECT -53.205 -129.365 -52.875 -129.035 ;
        RECT -53.205 -130.725 -52.875 -130.395 ;
        RECT -53.205 -131.47 -52.875 -131.14 ;
        RECT -53.205 -133.445 -52.875 -133.115 ;
        RECT -53.205 -134.805 -52.875 -134.475 ;
        RECT -53.205 -136.165 -52.875 -135.835 ;
        RECT -53.205 -137.525 -52.875 -137.195 ;
        RECT -53.205 -140.245 -52.875 -139.915 ;
        RECT -53.205 -141.605 -52.875 -141.275 ;
        RECT -53.205 -142.965 -52.875 -142.635 ;
        RECT -53.205 -144.31 -52.875 -143.98 ;
        RECT -53.205 -145.685 -52.875 -145.355 ;
        RECT -53.205 -147.045 -52.875 -146.715 ;
        RECT -53.205 -149.765 -52.875 -149.435 ;
        RECT -53.2 -149.765 -52.88 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 -234.085 -52.875 -233.755 ;
        RECT -53.205 -235.445 -52.875 -235.115 ;
        RECT -53.205 -236.805 -52.875 -236.475 ;
        RECT -53.205 -238.165 -52.875 -237.835 ;
        RECT -53.205 -243.81 -52.875 -242.68 ;
        RECT -53.2 -243.925 -52.88 -231.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 246.76 -51.515 247.89 ;
        RECT -51.845 241.915 -51.515 242.245 ;
        RECT -51.845 240.555 -51.515 240.885 ;
        RECT -51.845 239.195 -51.515 239.525 ;
        RECT -51.845 237.835 -51.515 238.165 ;
        RECT -51.845 236.475 -51.515 236.805 ;
        RECT -51.845 235.115 -51.515 235.445 ;
        RECT -51.845 233.755 -51.515 234.085 ;
        RECT -51.845 232.395 -51.515 232.725 ;
        RECT -51.845 231.035 -51.515 231.365 ;
        RECT -51.845 229.675 -51.515 230.005 ;
        RECT -51.845 228.315 -51.515 228.645 ;
        RECT -51.845 226.955 -51.515 227.285 ;
        RECT -51.845 225.595 -51.515 225.925 ;
        RECT -51.845 224.235 -51.515 224.565 ;
        RECT -51.845 222.875 -51.515 223.205 ;
        RECT -51.845 221.515 -51.515 221.845 ;
        RECT -51.845 220.155 -51.515 220.485 ;
        RECT -51.845 218.795 -51.515 219.125 ;
        RECT -51.845 217.435 -51.515 217.765 ;
        RECT -51.845 216.075 -51.515 216.405 ;
        RECT -51.845 214.715 -51.515 215.045 ;
        RECT -51.845 213.355 -51.515 213.685 ;
        RECT -51.845 211.995 -51.515 212.325 ;
        RECT -51.845 210.635 -51.515 210.965 ;
        RECT -51.845 209.275 -51.515 209.605 ;
        RECT -51.845 207.915 -51.515 208.245 ;
        RECT -51.845 206.555 -51.515 206.885 ;
        RECT -51.845 205.195 -51.515 205.525 ;
        RECT -51.845 203.835 -51.515 204.165 ;
        RECT -51.845 202.475 -51.515 202.805 ;
        RECT -51.845 201.115 -51.515 201.445 ;
        RECT -51.845 199.755 -51.515 200.085 ;
        RECT -51.845 198.395 -51.515 198.725 ;
        RECT -51.845 197.035 -51.515 197.365 ;
        RECT -51.845 195.675 -51.515 196.005 ;
        RECT -51.845 194.315 -51.515 194.645 ;
        RECT -51.845 192.955 -51.515 193.285 ;
        RECT -51.845 191.595 -51.515 191.925 ;
        RECT -51.845 190.235 -51.515 190.565 ;
        RECT -51.845 188.875 -51.515 189.205 ;
        RECT -51.845 187.515 -51.515 187.845 ;
        RECT -51.845 186.155 -51.515 186.485 ;
        RECT -51.845 184.795 -51.515 185.125 ;
        RECT -51.845 183.435 -51.515 183.765 ;
        RECT -51.845 182.075 -51.515 182.405 ;
        RECT -51.845 180.715 -51.515 181.045 ;
        RECT -51.845 179.355 -51.515 179.685 ;
        RECT -51.845 177.995 -51.515 178.325 ;
        RECT -51.845 176.635 -51.515 176.965 ;
        RECT -51.845 175.275 -51.515 175.605 ;
        RECT -51.845 173.915 -51.515 174.245 ;
        RECT -51.845 172.555 -51.515 172.885 ;
        RECT -51.845 171.195 -51.515 171.525 ;
        RECT -51.845 169.835 -51.515 170.165 ;
        RECT -51.845 168.475 -51.515 168.805 ;
        RECT -51.845 167.115 -51.515 167.445 ;
        RECT -51.845 165.755 -51.515 166.085 ;
        RECT -51.845 164.395 -51.515 164.725 ;
        RECT -51.845 163.035 -51.515 163.365 ;
        RECT -51.845 161.675 -51.515 162.005 ;
        RECT -51.845 160.315 -51.515 160.645 ;
        RECT -51.845 158.955 -51.515 159.285 ;
        RECT -51.845 157.595 -51.515 157.925 ;
        RECT -51.845 156.235 -51.515 156.565 ;
        RECT -51.845 154.875 -51.515 155.205 ;
        RECT -51.845 153.515 -51.515 153.845 ;
        RECT -51.845 152.155 -51.515 152.485 ;
        RECT -51.845 150.795 -51.515 151.125 ;
        RECT -51.845 149.435 -51.515 149.765 ;
        RECT -51.845 148.075 -51.515 148.405 ;
        RECT -51.845 146.715 -51.515 147.045 ;
        RECT -51.845 145.355 -51.515 145.685 ;
        RECT -51.845 143.995 -51.515 144.325 ;
        RECT -51.845 142.635 -51.515 142.965 ;
        RECT -51.845 141.275 -51.515 141.605 ;
        RECT -51.845 139.915 -51.515 140.245 ;
        RECT -51.845 138.555 -51.515 138.885 ;
        RECT -51.84 138.555 -51.52 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 97.755 -51.515 98.085 ;
        RECT -51.845 96.395 -51.515 96.725 ;
        RECT -51.845 95.035 -51.515 95.365 ;
        RECT -51.845 93.675 -51.515 94.005 ;
        RECT -51.845 92.315 -51.515 92.645 ;
        RECT -51.845 89.595 -51.515 89.925 ;
        RECT -51.845 88.235 -51.515 88.565 ;
        RECT -51.845 84.155 -51.515 84.485 ;
        RECT -51.845 82.795 -51.515 83.125 ;
        RECT -51.845 81.435 -51.515 81.765 ;
        RECT -51.845 80.075 -51.515 80.405 ;
        RECT -51.845 78.715 -51.515 79.045 ;
        RECT -51.845 77.355 -51.515 77.685 ;
        RECT -51.845 75.995 -51.515 76.325 ;
        RECT -51.845 74.635 -51.515 74.965 ;
        RECT -51.845 73.275 -51.515 73.605 ;
        RECT -51.845 71.915 -51.515 72.245 ;
        RECT -51.845 70.555 -51.515 70.885 ;
        RECT -51.845 69.195 -51.515 69.525 ;
        RECT -51.845 67.835 -51.515 68.165 ;
        RECT -51.845 66.475 -51.515 66.805 ;
        RECT -51.845 65.115 -51.515 65.445 ;
        RECT -51.845 63.755 -51.515 64.085 ;
        RECT -51.845 62.395 -51.515 62.725 ;
        RECT -51.845 61.035 -51.515 61.365 ;
        RECT -51.845 59.675 -51.515 60.005 ;
        RECT -51.845 58.315 -51.515 58.645 ;
        RECT -51.845 56.955 -51.515 57.285 ;
        RECT -51.845 55.595 -51.515 55.925 ;
        RECT -51.845 54.235 -51.515 54.565 ;
        RECT -51.845 52.875 -51.515 53.205 ;
        RECT -51.845 51.515 -51.515 51.845 ;
        RECT -51.845 50.155 -51.515 50.485 ;
        RECT -51.845 48.795 -51.515 49.125 ;
        RECT -51.845 47.435 -51.515 47.765 ;
        RECT -51.845 46.075 -51.515 46.405 ;
        RECT -51.845 44.715 -51.515 45.045 ;
        RECT -51.845 43.355 -51.515 43.685 ;
        RECT -51.845 41.995 -51.515 42.325 ;
        RECT -51.845 40.635 -51.515 40.965 ;
        RECT -51.845 39.275 -51.515 39.605 ;
        RECT -51.845 37.915 -51.515 38.245 ;
        RECT -51.845 36.555 -51.515 36.885 ;
        RECT -51.845 35.195 -51.515 35.525 ;
        RECT -51.845 33.835 -51.515 34.165 ;
        RECT -51.845 32.475 -51.515 32.805 ;
        RECT -51.845 31.115 -51.515 31.445 ;
        RECT -51.845 29.755 -51.515 30.085 ;
        RECT -51.845 28.395 -51.515 28.725 ;
        RECT -51.845 27.035 -51.515 27.365 ;
        RECT -51.845 25.675 -51.515 26.005 ;
        RECT -51.845 24.315 -51.515 24.645 ;
        RECT -51.845 22.955 -51.515 23.285 ;
        RECT -51.845 21.595 -51.515 21.925 ;
        RECT -51.845 20.235 -51.515 20.565 ;
        RECT -51.845 18.875 -51.515 19.205 ;
        RECT -51.845 17.515 -51.515 17.845 ;
        RECT -51.845 16.155 -51.515 16.485 ;
        RECT -51.845 14.795 -51.515 15.125 ;
        RECT -51.845 13.435 -51.515 13.765 ;
        RECT -51.845 12.075 -51.515 12.405 ;
        RECT -51.845 10.715 -51.515 11.045 ;
        RECT -51.845 9.355 -51.515 9.685 ;
        RECT -51.845 7.995 -51.515 8.325 ;
        RECT -51.845 6.635 -51.515 6.965 ;
        RECT -51.845 5.275 -51.515 5.605 ;
        RECT -51.845 3.915 -51.515 4.245 ;
        RECT -51.845 2.555 -51.515 2.885 ;
        RECT -51.845 1.195 -51.515 1.525 ;
        RECT -51.845 -0.165 -51.515 0.165 ;
        RECT -51.845 -1.525 -51.515 -1.195 ;
        RECT -51.845 -2.885 -51.515 -2.555 ;
        RECT -51.845 -4.245 -51.515 -3.915 ;
        RECT -51.845 -5.605 -51.515 -5.275 ;
        RECT -51.845 -6.965 -51.515 -6.635 ;
        RECT -51.845 -8.325 -51.515 -7.995 ;
        RECT -51.845 -9.685 -51.515 -9.355 ;
        RECT -51.845 -12.405 -51.515 -12.075 ;
        RECT -51.845 -13.765 -51.515 -13.435 ;
        RECT -51.845 -15.125 -51.515 -14.795 ;
        RECT -51.845 -16.485 -51.515 -16.155 ;
        RECT -51.845 -17.845 -51.515 -17.515 ;
        RECT -51.845 -19.205 -51.515 -18.875 ;
        RECT -51.845 -20.565 -51.515 -20.235 ;
        RECT -51.845 -21.925 -51.515 -21.595 ;
        RECT -51.845 -23.285 -51.515 -22.955 ;
        RECT -51.845 -24.645 -51.515 -24.315 ;
        RECT -51.845 -26.005 -51.515 -25.675 ;
        RECT -51.845 -27.365 -51.515 -27.035 ;
        RECT -51.845 -28.725 -51.515 -28.395 ;
        RECT -51.845 -30.085 -51.515 -29.755 ;
        RECT -51.845 -31.445 -51.515 -31.115 ;
        RECT -51.845 -32.805 -51.515 -32.475 ;
        RECT -51.845 -34.165 -51.515 -33.835 ;
        RECT -51.845 -35.525 -51.515 -35.195 ;
        RECT -51.845 -36.885 -51.515 -36.555 ;
        RECT -51.845 -38.245 -51.515 -37.915 ;
        RECT -51.845 -39.605 -51.515 -39.275 ;
        RECT -51.845 -40.965 -51.515 -40.635 ;
        RECT -51.845 -42.325 -51.515 -41.995 ;
        RECT -51.845 -43.685 -51.515 -43.355 ;
        RECT -51.845 -45.045 -51.515 -44.715 ;
        RECT -51.845 -46.405 -51.515 -46.075 ;
        RECT -51.845 -47.765 -51.515 -47.435 ;
        RECT -51.845 -49.125 -51.515 -48.795 ;
        RECT -51.845 -50.485 -51.515 -50.155 ;
        RECT -51.845 -51.845 -51.515 -51.515 ;
        RECT -51.845 -53.205 -51.515 -52.875 ;
        RECT -51.845 -54.565 -51.515 -54.235 ;
        RECT -51.845 -55.925 -51.515 -55.595 ;
        RECT -51.845 -57.285 -51.515 -56.955 ;
        RECT -51.845 -58.645 -51.515 -58.315 ;
        RECT -51.845 -60.005 -51.515 -59.675 ;
        RECT -51.845 -61.365 -51.515 -61.035 ;
        RECT -51.845 -62.725 -51.515 -62.395 ;
        RECT -51.845 -64.085 -51.515 -63.755 ;
        RECT -51.845 -65.445 -51.515 -65.115 ;
        RECT -51.845 -66.805 -51.515 -66.475 ;
        RECT -51.845 -68.165 -51.515 -67.835 ;
        RECT -51.845 -69.525 -51.515 -69.195 ;
        RECT -51.845 -70.885 -51.515 -70.555 ;
        RECT -51.845 -72.245 -51.515 -71.915 ;
        RECT -51.845 -73.605 -51.515 -73.275 ;
        RECT -51.845 -74.965 -51.515 -74.635 ;
        RECT -51.845 -76.325 -51.515 -75.995 ;
        RECT -51.845 -77.685 -51.515 -77.355 ;
        RECT -51.845 -79.045 -51.515 -78.715 ;
        RECT -51.845 -80.405 -51.515 -80.075 ;
        RECT -51.845 -81.765 -51.515 -81.435 ;
        RECT -51.845 -83.125 -51.515 -82.795 ;
        RECT -51.845 -84.485 -51.515 -84.155 ;
        RECT -51.845 -85.845 -51.515 -85.515 ;
        RECT -51.845 -87.205 -51.515 -86.875 ;
        RECT -51.845 -88.565 -51.515 -88.235 ;
        RECT -51.845 -89.925 -51.515 -89.595 ;
        RECT -51.845 -91.285 -51.515 -90.955 ;
        RECT -51.845 -92.645 -51.515 -92.315 ;
        RECT -51.845 -94.005 -51.515 -93.675 ;
        RECT -51.845 -95.365 -51.515 -95.035 ;
        RECT -51.845 -96.725 -51.515 -96.395 ;
        RECT -51.845 -98.085 -51.515 -97.755 ;
        RECT -51.845 -99.445 -51.515 -99.115 ;
        RECT -51.845 -100.805 -51.515 -100.475 ;
        RECT -51.845 -102.165 -51.515 -101.835 ;
        RECT -51.845 -103.525 -51.515 -103.195 ;
        RECT -51.845 -104.885 -51.515 -104.555 ;
        RECT -51.845 -106.245 -51.515 -105.915 ;
        RECT -51.845 -107.605 -51.515 -107.275 ;
        RECT -51.845 -108.965 -51.515 -108.635 ;
        RECT -51.845 -110.325 -51.515 -109.995 ;
        RECT -51.845 -111.685 -51.515 -111.355 ;
        RECT -51.845 -113.045 -51.515 -112.715 ;
        RECT -51.845 -114.405 -51.515 -114.075 ;
        RECT -51.845 -115.765 -51.515 -115.435 ;
        RECT -51.845 -117.125 -51.515 -116.795 ;
        RECT -51.845 -118.485 -51.515 -118.155 ;
        RECT -51.845 -119.845 -51.515 -119.515 ;
        RECT -51.845 -121.205 -51.515 -120.875 ;
        RECT -51.845 -122.565 -51.515 -122.235 ;
        RECT -51.845 -129.365 -51.515 -129.035 ;
        RECT -51.845 -130.725 -51.515 -130.395 ;
        RECT -51.845 -131.47 -51.515 -131.14 ;
        RECT -51.845 -133.445 -51.515 -133.115 ;
        RECT -51.845 -134.805 -51.515 -134.475 ;
        RECT -51.845 -136.165 -51.515 -135.835 ;
        RECT -51.845 -137.525 -51.515 -137.195 ;
        RECT -51.845 -140.245 -51.515 -139.915 ;
        RECT -51.845 -141.605 -51.515 -141.275 ;
        RECT -51.845 -142.965 -51.515 -142.635 ;
        RECT -51.845 -144.31 -51.515 -143.98 ;
        RECT -51.845 -145.685 -51.515 -145.355 ;
        RECT -51.845 -147.045 -51.515 -146.715 ;
        RECT -51.845 -149.765 -51.515 -149.435 ;
        RECT -51.845 -152.485 -51.515 -152.155 ;
        RECT -51.845 -153.845 -51.515 -153.515 ;
        RECT -51.845 -155.205 -51.515 -154.875 ;
        RECT -51.845 -156.565 -51.515 -156.235 ;
        RECT -51.845 -157.925 -51.515 -157.595 ;
        RECT -51.845 -159.285 -51.515 -158.955 ;
        RECT -51.845 -162.005 -51.515 -161.675 ;
        RECT -51.845 -163.365 -51.515 -163.035 ;
        RECT -51.845 -164.725 -51.515 -164.395 ;
        RECT -51.845 -166.085 -51.515 -165.755 ;
        RECT -51.845 -167.445 -51.515 -167.115 ;
        RECT -51.845 -168.805 -51.515 -168.475 ;
        RECT -51.845 -170.165 -51.515 -169.835 ;
        RECT -51.845 -171.525 -51.515 -171.195 ;
        RECT -51.845 -172.885 -51.515 -172.555 ;
        RECT -51.845 -174.245 -51.515 -173.915 ;
        RECT -51.845 -175.605 -51.515 -175.275 ;
        RECT -51.845 -176.965 -51.515 -176.635 ;
        RECT -51.845 -178.325 -51.515 -177.995 ;
        RECT -51.845 -179.685 -51.515 -179.355 ;
        RECT -51.845 -181.045 -51.515 -180.715 ;
        RECT -51.845 -182.405 -51.515 -182.075 ;
        RECT -51.845 -183.765 -51.515 -183.435 ;
        RECT -51.845 -185.125 -51.515 -184.795 ;
        RECT -51.845 -186.485 -51.515 -186.155 ;
        RECT -51.845 -187.845 -51.515 -187.515 ;
        RECT -51.845 -189.205 -51.515 -188.875 ;
        RECT -51.845 -190.565 -51.515 -190.235 ;
        RECT -51.845 -191.925 -51.515 -191.595 ;
        RECT -51.845 -193.285 -51.515 -192.955 ;
        RECT -51.845 -194.645 -51.515 -194.315 ;
        RECT -51.845 -196.005 -51.515 -195.675 ;
        RECT -51.845 -197.365 -51.515 -197.035 ;
        RECT -51.845 -198.725 -51.515 -198.395 ;
        RECT -51.845 -200.085 -51.515 -199.755 ;
        RECT -51.845 -201.445 -51.515 -201.115 ;
        RECT -51.845 -202.805 -51.515 -202.475 ;
        RECT -51.845 -204.165 -51.515 -203.835 ;
        RECT -51.845 -205.525 -51.515 -205.195 ;
        RECT -51.845 -206.885 -51.515 -206.555 ;
        RECT -51.845 -208.245 -51.515 -207.915 ;
        RECT -51.845 -209.605 -51.515 -209.275 ;
        RECT -51.845 -210.965 -51.515 -210.635 ;
        RECT -51.845 -212.325 -51.515 -211.995 ;
        RECT -51.845 -213.685 -51.515 -213.355 ;
        RECT -51.845 -215.045 -51.515 -214.715 ;
        RECT -51.845 -216.405 -51.515 -216.075 ;
        RECT -51.845 -217.765 -51.515 -217.435 ;
        RECT -51.845 -219.125 -51.515 -218.795 ;
        RECT -51.845 -220.485 -51.515 -220.155 ;
        RECT -51.845 -221.845 -51.515 -221.515 ;
        RECT -51.845 -223.205 -51.515 -222.875 ;
        RECT -51.845 -224.565 -51.515 -224.235 ;
        RECT -51.845 -226.155 -51.515 -225.825 ;
        RECT -51.845 -227.285 -51.515 -226.955 ;
        RECT -51.845 -228.645 -51.515 -228.315 ;
        RECT -51.845 -231.365 -51.515 -231.035 ;
        RECT -51.845 -234.085 -51.515 -233.755 ;
        RECT -51.845 -235.445 -51.515 -235.115 ;
        RECT -51.845 -236.805 -51.515 -236.475 ;
        RECT -51.845 -238.165 -51.515 -237.835 ;
        RECT -51.845 -243.81 -51.515 -242.68 ;
        RECT -51.84 -243.925 -51.52 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 246.76 -50.155 247.89 ;
        RECT -50.485 241.915 -50.155 242.245 ;
        RECT -50.485 240.555 -50.155 240.885 ;
        RECT -50.485 239.195 -50.155 239.525 ;
        RECT -50.485 237.835 -50.155 238.165 ;
        RECT -50.485 236.475 -50.155 236.805 ;
        RECT -50.485 235.115 -50.155 235.445 ;
        RECT -50.485 233.755 -50.155 234.085 ;
        RECT -50.485 232.395 -50.155 232.725 ;
        RECT -50.485 231.035 -50.155 231.365 ;
        RECT -50.485 229.675 -50.155 230.005 ;
        RECT -50.485 228.315 -50.155 228.645 ;
        RECT -50.485 226.955 -50.155 227.285 ;
        RECT -50.485 225.595 -50.155 225.925 ;
        RECT -50.485 224.235 -50.155 224.565 ;
        RECT -50.485 222.875 -50.155 223.205 ;
        RECT -50.485 221.515 -50.155 221.845 ;
        RECT -50.485 220.155 -50.155 220.485 ;
        RECT -50.485 218.795 -50.155 219.125 ;
        RECT -50.485 217.435 -50.155 217.765 ;
        RECT -50.485 216.075 -50.155 216.405 ;
        RECT -50.485 214.715 -50.155 215.045 ;
        RECT -50.485 213.355 -50.155 213.685 ;
        RECT -50.485 211.995 -50.155 212.325 ;
        RECT -50.485 210.635 -50.155 210.965 ;
        RECT -50.485 209.275 -50.155 209.605 ;
        RECT -50.485 207.915 -50.155 208.245 ;
        RECT -50.485 206.555 -50.155 206.885 ;
        RECT -50.485 205.195 -50.155 205.525 ;
        RECT -50.485 203.835 -50.155 204.165 ;
        RECT -50.485 202.475 -50.155 202.805 ;
        RECT -50.485 201.115 -50.155 201.445 ;
        RECT -50.485 199.755 -50.155 200.085 ;
        RECT -50.485 198.395 -50.155 198.725 ;
        RECT -50.485 197.035 -50.155 197.365 ;
        RECT -50.485 195.675 -50.155 196.005 ;
        RECT -50.485 194.315 -50.155 194.645 ;
        RECT -50.485 192.955 -50.155 193.285 ;
        RECT -50.485 191.595 -50.155 191.925 ;
        RECT -50.485 190.235 -50.155 190.565 ;
        RECT -50.485 188.875 -50.155 189.205 ;
        RECT -50.485 187.515 -50.155 187.845 ;
        RECT -50.485 186.155 -50.155 186.485 ;
        RECT -50.485 184.795 -50.155 185.125 ;
        RECT -50.485 183.435 -50.155 183.765 ;
        RECT -50.485 182.075 -50.155 182.405 ;
        RECT -50.485 180.715 -50.155 181.045 ;
        RECT -50.485 179.355 -50.155 179.685 ;
        RECT -50.485 177.995 -50.155 178.325 ;
        RECT -50.485 176.635 -50.155 176.965 ;
        RECT -50.485 175.275 -50.155 175.605 ;
        RECT -50.485 173.915 -50.155 174.245 ;
        RECT -50.485 172.555 -50.155 172.885 ;
        RECT -50.485 171.195 -50.155 171.525 ;
        RECT -50.485 169.835 -50.155 170.165 ;
        RECT -50.485 168.475 -50.155 168.805 ;
        RECT -50.485 167.115 -50.155 167.445 ;
        RECT -50.485 165.755 -50.155 166.085 ;
        RECT -50.485 164.395 -50.155 164.725 ;
        RECT -50.485 163.035 -50.155 163.365 ;
        RECT -50.485 161.675 -50.155 162.005 ;
        RECT -50.485 160.315 -50.155 160.645 ;
        RECT -50.485 158.955 -50.155 159.285 ;
        RECT -50.485 157.595 -50.155 157.925 ;
        RECT -50.485 156.235 -50.155 156.565 ;
        RECT -50.485 154.875 -50.155 155.205 ;
        RECT -50.485 153.515 -50.155 153.845 ;
        RECT -50.485 152.155 -50.155 152.485 ;
        RECT -50.485 150.795 -50.155 151.125 ;
        RECT -50.485 149.435 -50.155 149.765 ;
        RECT -50.485 148.075 -50.155 148.405 ;
        RECT -50.485 146.715 -50.155 147.045 ;
        RECT -50.485 145.355 -50.155 145.685 ;
        RECT -50.485 143.995 -50.155 144.325 ;
        RECT -50.485 142.635 -50.155 142.965 ;
        RECT -50.485 141.275 -50.155 141.605 ;
        RECT -50.485 139.915 -50.155 140.245 ;
        RECT -50.485 138.555 -50.155 138.885 ;
        RECT -50.48 138.555 -50.16 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 -15.125 -50.155 -14.795 ;
        RECT -50.485 -16.485 -50.155 -16.155 ;
        RECT -50.485 -17.845 -50.155 -17.515 ;
        RECT -50.485 -19.205 -50.155 -18.875 ;
        RECT -50.485 -20.565 -50.155 -20.235 ;
        RECT -50.485 -21.925 -50.155 -21.595 ;
        RECT -50.485 -23.285 -50.155 -22.955 ;
        RECT -50.485 -24.645 -50.155 -24.315 ;
        RECT -50.485 -26.005 -50.155 -25.675 ;
        RECT -50.485 -27.365 -50.155 -27.035 ;
        RECT -50.485 -28.725 -50.155 -28.395 ;
        RECT -50.485 -30.085 -50.155 -29.755 ;
        RECT -50.485 -31.445 -50.155 -31.115 ;
        RECT -50.485 -32.805 -50.155 -32.475 ;
        RECT -50.485 -34.165 -50.155 -33.835 ;
        RECT -50.485 -35.525 -50.155 -35.195 ;
        RECT -50.485 -36.885 -50.155 -36.555 ;
        RECT -50.485 -38.245 -50.155 -37.915 ;
        RECT -50.485 -39.605 -50.155 -39.275 ;
        RECT -50.485 -40.965 -50.155 -40.635 ;
        RECT -50.485 -42.325 -50.155 -41.995 ;
        RECT -50.485 -43.685 -50.155 -43.355 ;
        RECT -50.485 -45.045 -50.155 -44.715 ;
        RECT -50.485 -46.405 -50.155 -46.075 ;
        RECT -50.485 -47.765 -50.155 -47.435 ;
        RECT -50.485 -49.125 -50.155 -48.795 ;
        RECT -50.485 -50.485 -50.155 -50.155 ;
        RECT -50.485 -51.845 -50.155 -51.515 ;
        RECT -50.485 -53.205 -50.155 -52.875 ;
        RECT -50.485 -54.565 -50.155 -54.235 ;
        RECT -50.485 -55.925 -50.155 -55.595 ;
        RECT -50.485 -57.285 -50.155 -56.955 ;
        RECT -50.485 -58.645 -50.155 -58.315 ;
        RECT -50.485 -60.005 -50.155 -59.675 ;
        RECT -50.485 -61.365 -50.155 -61.035 ;
        RECT -50.485 -62.725 -50.155 -62.395 ;
        RECT -50.485 -64.085 -50.155 -63.755 ;
        RECT -50.485 -65.445 -50.155 -65.115 ;
        RECT -50.485 -66.805 -50.155 -66.475 ;
        RECT -50.485 -68.165 -50.155 -67.835 ;
        RECT -50.485 -69.525 -50.155 -69.195 ;
        RECT -50.485 -70.885 -50.155 -70.555 ;
        RECT -50.485 -72.245 -50.155 -71.915 ;
        RECT -50.485 -73.605 -50.155 -73.275 ;
        RECT -50.485 -74.965 -50.155 -74.635 ;
        RECT -50.485 -76.325 -50.155 -75.995 ;
        RECT -50.485 -77.685 -50.155 -77.355 ;
        RECT -50.485 -79.045 -50.155 -78.715 ;
        RECT -50.485 -80.405 -50.155 -80.075 ;
        RECT -50.485 -81.765 -50.155 -81.435 ;
        RECT -50.485 -83.125 -50.155 -82.795 ;
        RECT -50.485 -84.485 -50.155 -84.155 ;
        RECT -50.485 -85.845 -50.155 -85.515 ;
        RECT -50.485 -87.205 -50.155 -86.875 ;
        RECT -50.485 -88.565 -50.155 -88.235 ;
        RECT -50.485 -89.925 -50.155 -89.595 ;
        RECT -50.485 -91.285 -50.155 -90.955 ;
        RECT -50.485 -92.645 -50.155 -92.315 ;
        RECT -50.485 -94.005 -50.155 -93.675 ;
        RECT -50.485 -95.365 -50.155 -95.035 ;
        RECT -50.485 -96.725 -50.155 -96.395 ;
        RECT -50.485 -98.085 -50.155 -97.755 ;
        RECT -50.485 -99.445 -50.155 -99.115 ;
        RECT -50.485 -100.805 -50.155 -100.475 ;
        RECT -50.485 -102.165 -50.155 -101.835 ;
        RECT -50.485 -103.525 -50.155 -103.195 ;
        RECT -50.485 -104.885 -50.155 -104.555 ;
        RECT -50.485 -106.245 -50.155 -105.915 ;
        RECT -50.485 -107.605 -50.155 -107.275 ;
        RECT -50.485 -108.965 -50.155 -108.635 ;
        RECT -50.485 -110.325 -50.155 -109.995 ;
        RECT -50.485 -111.685 -50.155 -111.355 ;
        RECT -50.485 -113.045 -50.155 -112.715 ;
        RECT -50.485 -114.405 -50.155 -114.075 ;
        RECT -50.485 -115.765 -50.155 -115.435 ;
        RECT -50.485 -117.125 -50.155 -116.795 ;
        RECT -50.485 -118.485 -50.155 -118.155 ;
        RECT -50.485 -119.845 -50.155 -119.515 ;
        RECT -50.485 -121.205 -50.155 -120.875 ;
        RECT -50.485 -122.565 -50.155 -122.235 ;
        RECT -50.485 -129.365 -50.155 -129.035 ;
        RECT -50.485 -130.725 -50.155 -130.395 ;
        RECT -50.485 -131.47 -50.155 -131.14 ;
        RECT -50.485 -133.445 -50.155 -133.115 ;
        RECT -50.485 -134.805 -50.155 -134.475 ;
        RECT -50.485 -136.165 -50.155 -135.835 ;
        RECT -50.485 -137.525 -50.155 -137.195 ;
        RECT -50.485 -140.245 -50.155 -139.915 ;
        RECT -50.485 -141.605 -50.155 -141.275 ;
        RECT -50.485 -142.965 -50.155 -142.635 ;
        RECT -50.485 -144.31 -50.155 -143.98 ;
        RECT -50.485 -145.685 -50.155 -145.355 ;
        RECT -50.485 -147.045 -50.155 -146.715 ;
        RECT -50.485 -149.765 -50.155 -149.435 ;
        RECT -50.485 -152.485 -50.155 -152.155 ;
        RECT -50.485 -153.845 -50.155 -153.515 ;
        RECT -50.485 -155.205 -50.155 -154.875 ;
        RECT -50.485 -156.565 -50.155 -156.235 ;
        RECT -50.485 -157.925 -50.155 -157.595 ;
        RECT -50.485 -159.285 -50.155 -158.955 ;
        RECT -50.485 -162.005 -50.155 -161.675 ;
        RECT -50.485 -163.365 -50.155 -163.035 ;
        RECT -50.485 -164.725 -50.155 -164.395 ;
        RECT -50.485 -166.085 -50.155 -165.755 ;
        RECT -50.485 -167.445 -50.155 -167.115 ;
        RECT -50.485 -168.805 -50.155 -168.475 ;
        RECT -50.485 -170.165 -50.155 -169.835 ;
        RECT -50.485 -171.525 -50.155 -171.195 ;
        RECT -50.485 -172.885 -50.155 -172.555 ;
        RECT -50.485 -174.245 -50.155 -173.915 ;
        RECT -50.485 -175.605 -50.155 -175.275 ;
        RECT -50.485 -176.965 -50.155 -176.635 ;
        RECT -50.485 -178.325 -50.155 -177.995 ;
        RECT -50.485 -179.685 -50.155 -179.355 ;
        RECT -50.485 -181.045 -50.155 -180.715 ;
        RECT -50.485 -182.405 -50.155 -182.075 ;
        RECT -50.485 -183.765 -50.155 -183.435 ;
        RECT -50.485 -185.125 -50.155 -184.795 ;
        RECT -50.485 -186.485 -50.155 -186.155 ;
        RECT -50.485 -187.845 -50.155 -187.515 ;
        RECT -50.485 -189.205 -50.155 -188.875 ;
        RECT -50.485 -190.565 -50.155 -190.235 ;
        RECT -50.485 -191.925 -50.155 -191.595 ;
        RECT -50.485 -193.285 -50.155 -192.955 ;
        RECT -50.485 -194.645 -50.155 -194.315 ;
        RECT -50.485 -196.005 -50.155 -195.675 ;
        RECT -50.485 -197.365 -50.155 -197.035 ;
        RECT -50.485 -198.725 -50.155 -198.395 ;
        RECT -50.485 -200.085 -50.155 -199.755 ;
        RECT -50.485 -201.445 -50.155 -201.115 ;
        RECT -50.485 -202.805 -50.155 -202.475 ;
        RECT -50.485 -204.165 -50.155 -203.835 ;
        RECT -50.485 -205.525 -50.155 -205.195 ;
        RECT -50.485 -206.885 -50.155 -206.555 ;
        RECT -50.485 -208.245 -50.155 -207.915 ;
        RECT -50.485 -209.605 -50.155 -209.275 ;
        RECT -50.485 -210.965 -50.155 -210.635 ;
        RECT -50.485 -212.325 -50.155 -211.995 ;
        RECT -50.485 -213.685 -50.155 -213.355 ;
        RECT -50.485 -215.045 -50.155 -214.715 ;
        RECT -50.485 -216.405 -50.155 -216.075 ;
        RECT -50.485 -217.765 -50.155 -217.435 ;
        RECT -50.485 -219.125 -50.155 -218.795 ;
        RECT -50.485 -220.485 -50.155 -220.155 ;
        RECT -50.485 -221.845 -50.155 -221.515 ;
        RECT -50.485 -223.205 -50.155 -222.875 ;
        RECT -50.485 -224.565 -50.155 -224.235 ;
        RECT -50.485 -226.155 -50.155 -225.825 ;
        RECT -50.485 -227.285 -50.155 -226.955 ;
        RECT -50.485 -228.645 -50.155 -228.315 ;
        RECT -50.485 -230.005 -50.155 -229.675 ;
        RECT -50.485 -231.365 -50.155 -231.035 ;
        RECT -50.485 -234.085 -50.155 -233.755 ;
        RECT -50.485 -235.445 -50.155 -235.115 ;
        RECT -50.485 -236.805 -50.155 -236.475 ;
        RECT -50.485 -238.165 -50.155 -237.835 ;
        RECT -50.485 -243.81 -50.155 -242.68 ;
        RECT -50.48 -243.925 -50.16 98.085 ;
        RECT -50.485 97.755 -50.155 98.085 ;
        RECT -50.485 96.395 -50.155 96.725 ;
        RECT -50.485 95.035 -50.155 95.365 ;
        RECT -50.485 93.675 -50.155 94.005 ;
        RECT -50.485 92.315 -50.155 92.645 ;
        RECT -50.485 89.595 -50.155 89.925 ;
        RECT -50.485 88.235 -50.155 88.565 ;
        RECT -50.485 84.155 -50.155 84.485 ;
        RECT -50.485 82.795 -50.155 83.125 ;
        RECT -50.485 81.435 -50.155 81.765 ;
        RECT -50.485 80.075 -50.155 80.405 ;
        RECT -50.485 78.715 -50.155 79.045 ;
        RECT -50.485 77.355 -50.155 77.685 ;
        RECT -50.485 75.995 -50.155 76.325 ;
        RECT -50.485 74.635 -50.155 74.965 ;
        RECT -50.485 73.275 -50.155 73.605 ;
        RECT -50.485 71.915 -50.155 72.245 ;
        RECT -50.485 70.555 -50.155 70.885 ;
        RECT -50.485 69.195 -50.155 69.525 ;
        RECT -50.485 67.835 -50.155 68.165 ;
        RECT -50.485 66.475 -50.155 66.805 ;
        RECT -50.485 65.115 -50.155 65.445 ;
        RECT -50.485 63.755 -50.155 64.085 ;
        RECT -50.485 62.395 -50.155 62.725 ;
        RECT -50.485 61.035 -50.155 61.365 ;
        RECT -50.485 59.675 -50.155 60.005 ;
        RECT -50.485 58.315 -50.155 58.645 ;
        RECT -50.485 56.955 -50.155 57.285 ;
        RECT -50.485 55.595 -50.155 55.925 ;
        RECT -50.485 54.235 -50.155 54.565 ;
        RECT -50.485 52.875 -50.155 53.205 ;
        RECT -50.485 51.515 -50.155 51.845 ;
        RECT -50.485 50.155 -50.155 50.485 ;
        RECT -50.485 48.795 -50.155 49.125 ;
        RECT -50.485 47.435 -50.155 47.765 ;
        RECT -50.485 46.075 -50.155 46.405 ;
        RECT -50.485 44.715 -50.155 45.045 ;
        RECT -50.485 43.355 -50.155 43.685 ;
        RECT -50.485 41.995 -50.155 42.325 ;
        RECT -50.485 40.635 -50.155 40.965 ;
        RECT -50.485 39.275 -50.155 39.605 ;
        RECT -50.485 37.915 -50.155 38.245 ;
        RECT -50.485 36.555 -50.155 36.885 ;
        RECT -50.485 35.195 -50.155 35.525 ;
        RECT -50.485 33.835 -50.155 34.165 ;
        RECT -50.485 32.475 -50.155 32.805 ;
        RECT -50.485 31.115 -50.155 31.445 ;
        RECT -50.485 29.755 -50.155 30.085 ;
        RECT -50.485 28.395 -50.155 28.725 ;
        RECT -50.485 27.035 -50.155 27.365 ;
        RECT -50.485 25.675 -50.155 26.005 ;
        RECT -50.485 24.315 -50.155 24.645 ;
        RECT -50.485 22.955 -50.155 23.285 ;
        RECT -50.485 21.595 -50.155 21.925 ;
        RECT -50.485 20.235 -50.155 20.565 ;
        RECT -50.485 18.875 -50.155 19.205 ;
        RECT -50.485 17.515 -50.155 17.845 ;
        RECT -50.485 16.155 -50.155 16.485 ;
        RECT -50.485 14.795 -50.155 15.125 ;
        RECT -50.485 13.435 -50.155 13.765 ;
        RECT -50.485 12.075 -50.155 12.405 ;
        RECT -50.485 10.715 -50.155 11.045 ;
        RECT -50.485 9.355 -50.155 9.685 ;
        RECT -50.485 7.995 -50.155 8.325 ;
        RECT -50.485 6.635 -50.155 6.965 ;
        RECT -50.485 5.275 -50.155 5.605 ;
        RECT -50.485 3.915 -50.155 4.245 ;
        RECT -50.485 2.555 -50.155 2.885 ;
        RECT -50.485 1.195 -50.155 1.525 ;
        RECT -50.485 -0.165 -50.155 0.165 ;
        RECT -50.485 -1.525 -50.155 -1.195 ;
        RECT -50.485 -2.885 -50.155 -2.555 ;
        RECT -50.485 -4.245 -50.155 -3.915 ;
        RECT -50.485 -5.605 -50.155 -5.275 ;
        RECT -50.485 -6.965 -50.155 -6.635 ;
        RECT -50.485 -8.325 -50.155 -7.995 ;
        RECT -50.485 -9.685 -50.155 -9.355 ;
        RECT -50.485 -12.405 -50.155 -12.075 ;
        RECT -50.485 -13.765 -50.155 -13.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.285 246.76 -56.955 247.89 ;
        RECT -57.285 241.915 -56.955 242.245 ;
        RECT -57.285 240.555 -56.955 240.885 ;
        RECT -57.285 239.195 -56.955 239.525 ;
        RECT -57.285 237.835 -56.955 238.165 ;
        RECT -57.285 236.475 -56.955 236.805 ;
        RECT -57.285 235.115 -56.955 235.445 ;
        RECT -57.285 233.755 -56.955 234.085 ;
        RECT -57.285 232.395 -56.955 232.725 ;
        RECT -57.285 231.035 -56.955 231.365 ;
        RECT -57.285 229.675 -56.955 230.005 ;
        RECT -57.285 228.315 -56.955 228.645 ;
        RECT -57.285 226.955 -56.955 227.285 ;
        RECT -57.285 225.595 -56.955 225.925 ;
        RECT -57.285 224.235 -56.955 224.565 ;
        RECT -57.285 222.875 -56.955 223.205 ;
        RECT -57.285 221.515 -56.955 221.845 ;
        RECT -57.285 220.155 -56.955 220.485 ;
        RECT -57.285 218.795 -56.955 219.125 ;
        RECT -57.285 217.435 -56.955 217.765 ;
        RECT -57.285 216.075 -56.955 216.405 ;
        RECT -57.285 214.715 -56.955 215.045 ;
        RECT -57.285 213.355 -56.955 213.685 ;
        RECT -57.285 211.995 -56.955 212.325 ;
        RECT -57.285 210.635 -56.955 210.965 ;
        RECT -57.285 209.275 -56.955 209.605 ;
        RECT -57.285 207.915 -56.955 208.245 ;
        RECT -57.285 206.555 -56.955 206.885 ;
        RECT -57.285 205.195 -56.955 205.525 ;
        RECT -57.285 203.835 -56.955 204.165 ;
        RECT -57.285 202.475 -56.955 202.805 ;
        RECT -57.285 201.115 -56.955 201.445 ;
        RECT -57.285 199.755 -56.955 200.085 ;
        RECT -57.285 198.395 -56.955 198.725 ;
        RECT -57.285 197.035 -56.955 197.365 ;
        RECT -57.285 195.675 -56.955 196.005 ;
        RECT -57.285 194.315 -56.955 194.645 ;
        RECT -57.285 192.955 -56.955 193.285 ;
        RECT -57.285 191.595 -56.955 191.925 ;
        RECT -57.285 190.235 -56.955 190.565 ;
        RECT -57.285 188.875 -56.955 189.205 ;
        RECT -57.285 187.515 -56.955 187.845 ;
        RECT -57.285 186.155 -56.955 186.485 ;
        RECT -57.285 184.795 -56.955 185.125 ;
        RECT -57.285 183.435 -56.955 183.765 ;
        RECT -57.285 182.075 -56.955 182.405 ;
        RECT -57.285 180.715 -56.955 181.045 ;
        RECT -57.285 179.355 -56.955 179.685 ;
        RECT -57.285 177.995 -56.955 178.325 ;
        RECT -57.285 176.635 -56.955 176.965 ;
        RECT -57.285 175.275 -56.955 175.605 ;
        RECT -57.285 173.915 -56.955 174.245 ;
        RECT -57.285 172.555 -56.955 172.885 ;
        RECT -57.285 171.195 -56.955 171.525 ;
        RECT -57.285 169.835 -56.955 170.165 ;
        RECT -57.285 168.475 -56.955 168.805 ;
        RECT -57.285 167.115 -56.955 167.445 ;
        RECT -57.285 165.755 -56.955 166.085 ;
        RECT -57.285 164.395 -56.955 164.725 ;
        RECT -57.285 163.035 -56.955 163.365 ;
        RECT -57.285 161.675 -56.955 162.005 ;
        RECT -57.285 160.315 -56.955 160.645 ;
        RECT -57.285 158.955 -56.955 159.285 ;
        RECT -57.285 157.595 -56.955 157.925 ;
        RECT -57.285 156.235 -56.955 156.565 ;
        RECT -57.285 154.875 -56.955 155.205 ;
        RECT -57.285 153.515 -56.955 153.845 ;
        RECT -57.285 152.155 -56.955 152.485 ;
        RECT -57.285 150.795 -56.955 151.125 ;
        RECT -57.285 149.435 -56.955 149.765 ;
        RECT -57.285 148.075 -56.955 148.405 ;
        RECT -57.285 146.715 -56.955 147.045 ;
        RECT -57.285 145.355 -56.955 145.685 ;
        RECT -57.285 143.995 -56.955 144.325 ;
        RECT -57.285 142.635 -56.955 142.965 ;
        RECT -57.285 141.275 -56.955 141.605 ;
        RECT -57.285 139.915 -56.955 140.245 ;
        RECT -57.285 138.555 -56.955 138.885 ;
        RECT -57.285 136.42 -56.955 136.75 ;
        RECT -57.285 134.245 -56.955 134.575 ;
        RECT -57.285 133.395 -56.955 133.725 ;
        RECT -57.285 131.085 -56.955 131.415 ;
        RECT -57.285 130.235 -56.955 130.565 ;
        RECT -57.285 127.925 -56.955 128.255 ;
        RECT -57.285 127.075 -56.955 127.405 ;
        RECT -57.285 124.765 -56.955 125.095 ;
        RECT -57.285 123.915 -56.955 124.245 ;
        RECT -57.285 121.605 -56.955 121.935 ;
        RECT -57.285 120.755 -56.955 121.085 ;
        RECT -57.285 118.445 -56.955 118.775 ;
        RECT -57.285 117.595 -56.955 117.925 ;
        RECT -57.285 115.285 -56.955 115.615 ;
        RECT -57.285 114.435 -56.955 114.765 ;
        RECT -57.285 112.125 -56.955 112.455 ;
        RECT -57.285 111.275 -56.955 111.605 ;
        RECT -57.285 108.965 -56.955 109.295 ;
        RECT -57.285 108.115 -56.955 108.445 ;
        RECT -57.285 105.805 -56.955 106.135 ;
        RECT -57.285 104.955 -56.955 105.285 ;
        RECT -57.285 102.645 -56.955 102.975 ;
        RECT -57.285 101.795 -56.955 102.125 ;
        RECT -57.285 99.62 -56.955 99.95 ;
        RECT -57.285 97.755 -56.955 98.085 ;
        RECT -57.285 96.395 -56.955 96.725 ;
        RECT -57.285 95.035 -56.955 95.365 ;
        RECT -57.285 93.675 -56.955 94.005 ;
        RECT -57.285 92.315 -56.955 92.645 ;
        RECT -57.285 90.955 -56.955 91.285 ;
        RECT -57.285 89.595 -56.955 89.925 ;
        RECT -57.285 88.235 -56.955 88.565 ;
        RECT -57.285 86.875 -56.955 87.205 ;
        RECT -57.285 85.515 -56.955 85.845 ;
        RECT -57.285 84.155 -56.955 84.485 ;
        RECT -57.285 82.795 -56.955 83.125 ;
        RECT -57.285 81.435 -56.955 81.765 ;
        RECT -57.285 80.075 -56.955 80.405 ;
        RECT -57.285 78.715 -56.955 79.045 ;
        RECT -57.285 77.355 -56.955 77.685 ;
        RECT -57.285 75.995 -56.955 76.325 ;
        RECT -57.285 74.635 -56.955 74.965 ;
        RECT -57.285 73.275 -56.955 73.605 ;
        RECT -57.285 71.915 -56.955 72.245 ;
        RECT -57.285 70.555 -56.955 70.885 ;
        RECT -57.285 69.195 -56.955 69.525 ;
        RECT -57.285 67.835 -56.955 68.165 ;
        RECT -57.285 66.475 -56.955 66.805 ;
        RECT -57.285 65.115 -56.955 65.445 ;
        RECT -57.285 63.755 -56.955 64.085 ;
        RECT -57.285 62.395 -56.955 62.725 ;
        RECT -57.285 61.035 -56.955 61.365 ;
        RECT -57.285 59.675 -56.955 60.005 ;
        RECT -57.285 58.315 -56.955 58.645 ;
        RECT -57.285 56.955 -56.955 57.285 ;
        RECT -57.285 55.595 -56.955 55.925 ;
        RECT -57.285 54.235 -56.955 54.565 ;
        RECT -57.285 52.875 -56.955 53.205 ;
        RECT -57.285 51.515 -56.955 51.845 ;
        RECT -57.285 50.155 -56.955 50.485 ;
        RECT -57.285 48.795 -56.955 49.125 ;
        RECT -57.285 47.435 -56.955 47.765 ;
        RECT -57.285 46.075 -56.955 46.405 ;
        RECT -57.285 44.715 -56.955 45.045 ;
        RECT -57.285 43.355 -56.955 43.685 ;
        RECT -57.285 41.995 -56.955 42.325 ;
        RECT -57.285 40.635 -56.955 40.965 ;
        RECT -57.285 39.275 -56.955 39.605 ;
        RECT -57.285 37.915 -56.955 38.245 ;
        RECT -57.285 36.555 -56.955 36.885 ;
        RECT -57.285 35.195 -56.955 35.525 ;
        RECT -57.285 33.835 -56.955 34.165 ;
        RECT -57.285 32.475 -56.955 32.805 ;
        RECT -57.285 31.115 -56.955 31.445 ;
        RECT -57.285 29.755 -56.955 30.085 ;
        RECT -57.285 28.395 -56.955 28.725 ;
        RECT -57.285 27.035 -56.955 27.365 ;
        RECT -57.285 25.675 -56.955 26.005 ;
        RECT -57.285 24.315 -56.955 24.645 ;
        RECT -57.285 22.955 -56.955 23.285 ;
        RECT -57.285 21.595 -56.955 21.925 ;
        RECT -57.285 20.235 -56.955 20.565 ;
        RECT -57.285 18.875 -56.955 19.205 ;
        RECT -57.285 17.515 -56.955 17.845 ;
        RECT -57.285 16.155 -56.955 16.485 ;
        RECT -57.285 14.795 -56.955 15.125 ;
        RECT -57.285 13.435 -56.955 13.765 ;
        RECT -57.285 12.075 -56.955 12.405 ;
        RECT -57.285 10.715 -56.955 11.045 ;
        RECT -57.285 9.355 -56.955 9.685 ;
        RECT -57.285 7.995 -56.955 8.325 ;
        RECT -57.285 6.635 -56.955 6.965 ;
        RECT -57.285 5.275 -56.955 5.605 ;
        RECT -57.285 3.915 -56.955 4.245 ;
        RECT -57.285 2.555 -56.955 2.885 ;
        RECT -57.285 1.195 -56.955 1.525 ;
        RECT -57.285 -0.165 -56.955 0.165 ;
        RECT -57.285 -1.525 -56.955 -1.195 ;
        RECT -57.285 -2.885 -56.955 -2.555 ;
        RECT -57.285 -4.245 -56.955 -3.915 ;
        RECT -57.285 -5.605 -56.955 -5.275 ;
        RECT -57.285 -6.965 -56.955 -6.635 ;
        RECT -57.285 -8.325 -56.955 -7.995 ;
        RECT -57.285 -9.685 -56.955 -9.355 ;
        RECT -57.285 -11.045 -56.955 -10.715 ;
        RECT -57.285 -12.405 -56.955 -12.075 ;
        RECT -57.285 -13.765 -56.955 -13.435 ;
        RECT -57.285 -15.125 -56.955 -14.795 ;
        RECT -57.285 -16.485 -56.955 -16.155 ;
        RECT -57.285 -17.845 -56.955 -17.515 ;
        RECT -57.285 -19.205 -56.955 -18.875 ;
        RECT -57.285 -20.565 -56.955 -20.235 ;
        RECT -57.285 -21.925 -56.955 -21.595 ;
        RECT -57.285 -23.285 -56.955 -22.955 ;
        RECT -57.285 -24.645 -56.955 -24.315 ;
        RECT -57.285 -26.005 -56.955 -25.675 ;
        RECT -57.285 -27.365 -56.955 -27.035 ;
        RECT -57.285 -28.725 -56.955 -28.395 ;
        RECT -57.285 -30.085 -56.955 -29.755 ;
        RECT -57.285 -31.445 -56.955 -31.115 ;
        RECT -57.285 -32.805 -56.955 -32.475 ;
        RECT -57.285 -34.165 -56.955 -33.835 ;
        RECT -57.285 -35.525 -56.955 -35.195 ;
        RECT -57.285 -36.885 -56.955 -36.555 ;
        RECT -57.285 -38.245 -56.955 -37.915 ;
        RECT -57.285 -39.605 -56.955 -39.275 ;
        RECT -57.285 -40.965 -56.955 -40.635 ;
        RECT -57.285 -42.325 -56.955 -41.995 ;
        RECT -57.285 -43.685 -56.955 -43.355 ;
        RECT -57.285 -45.045 -56.955 -44.715 ;
        RECT -57.285 -46.405 -56.955 -46.075 ;
        RECT -57.285 -47.765 -56.955 -47.435 ;
        RECT -57.285 -49.125 -56.955 -48.795 ;
        RECT -57.285 -50.485 -56.955 -50.155 ;
        RECT -57.285 -51.845 -56.955 -51.515 ;
        RECT -57.285 -53.205 -56.955 -52.875 ;
        RECT -57.285 -54.565 -56.955 -54.235 ;
        RECT -57.285 -55.925 -56.955 -55.595 ;
        RECT -57.285 -57.285 -56.955 -56.955 ;
        RECT -57.285 -58.645 -56.955 -58.315 ;
        RECT -57.285 -60.005 -56.955 -59.675 ;
        RECT -57.285 -61.365 -56.955 -61.035 ;
        RECT -57.285 -62.725 -56.955 -62.395 ;
        RECT -57.285 -64.085 -56.955 -63.755 ;
        RECT -57.285 -65.445 -56.955 -65.115 ;
        RECT -57.285 -66.805 -56.955 -66.475 ;
        RECT -57.285 -68.165 -56.955 -67.835 ;
        RECT -57.285 -69.525 -56.955 -69.195 ;
        RECT -57.285 -70.885 -56.955 -70.555 ;
        RECT -57.285 -72.245 -56.955 -71.915 ;
        RECT -57.285 -73.605 -56.955 -73.275 ;
        RECT -57.285 -74.965 -56.955 -74.635 ;
        RECT -57.285 -76.325 -56.955 -75.995 ;
        RECT -57.285 -77.685 -56.955 -77.355 ;
        RECT -57.285 -79.045 -56.955 -78.715 ;
        RECT -57.285 -80.405 -56.955 -80.075 ;
        RECT -57.285 -81.765 -56.955 -81.435 ;
        RECT -57.285 -83.125 -56.955 -82.795 ;
        RECT -57.285 -84.485 -56.955 -84.155 ;
        RECT -57.285 -85.845 -56.955 -85.515 ;
        RECT -57.285 -87.205 -56.955 -86.875 ;
        RECT -57.285 -88.565 -56.955 -88.235 ;
        RECT -57.285 -89.925 -56.955 -89.595 ;
        RECT -57.285 -91.285 -56.955 -90.955 ;
        RECT -57.285 -92.645 -56.955 -92.315 ;
        RECT -57.285 -94.005 -56.955 -93.675 ;
        RECT -57.285 -95.365 -56.955 -95.035 ;
        RECT -57.285 -96.725 -56.955 -96.395 ;
        RECT -57.285 -98.085 -56.955 -97.755 ;
        RECT -57.285 -99.445 -56.955 -99.115 ;
        RECT -57.285 -100.805 -56.955 -100.475 ;
        RECT -57.285 -102.165 -56.955 -101.835 ;
        RECT -57.285 -103.525 -56.955 -103.195 ;
        RECT -57.285 -104.885 -56.955 -104.555 ;
        RECT -57.285 -106.245 -56.955 -105.915 ;
        RECT -57.285 -107.605 -56.955 -107.275 ;
        RECT -57.285 -108.965 -56.955 -108.635 ;
        RECT -57.285 -110.325 -56.955 -109.995 ;
        RECT -57.285 -111.685 -56.955 -111.355 ;
        RECT -57.285 -113.045 -56.955 -112.715 ;
        RECT -57.285 -114.405 -56.955 -114.075 ;
        RECT -57.285 -115.765 -56.955 -115.435 ;
        RECT -57.285 -117.125 -56.955 -116.795 ;
        RECT -57.285 -118.485 -56.955 -118.155 ;
        RECT -57.285 -119.845 -56.955 -119.515 ;
        RECT -57.285 -121.205 -56.955 -120.875 ;
        RECT -57.285 -122.565 -56.955 -122.235 ;
        RECT -57.285 -123.925 -56.955 -123.595 ;
        RECT -57.285 -129.365 -56.955 -129.035 ;
        RECT -57.285 -130.725 -56.955 -130.395 ;
        RECT -57.285 -131.47 -56.955 -131.14 ;
        RECT -57.285 -133.445 -56.955 -133.115 ;
        RECT -57.285 -134.805 -56.955 -134.475 ;
        RECT -57.285 -136.165 -56.955 -135.835 ;
        RECT -57.285 -137.525 -56.955 -137.195 ;
        RECT -57.285 -140.245 -56.955 -139.915 ;
        RECT -57.285 -141.605 -56.955 -141.275 ;
        RECT -57.285 -142.965 -56.955 -142.635 ;
        RECT -57.285 -144.31 -56.955 -143.98 ;
        RECT -57.285 -145.685 -56.955 -145.355 ;
        RECT -57.285 -147.045 -56.955 -146.715 ;
        RECT -57.285 -149.765 -56.955 -149.435 ;
        RECT -57.285 -152.485 -56.955 -152.155 ;
        RECT -57.285 -153.845 -56.955 -153.515 ;
        RECT -57.285 -155.205 -56.955 -154.875 ;
        RECT -57.285 -156.565 -56.955 -156.235 ;
        RECT -57.285 -157.925 -56.955 -157.595 ;
        RECT -57.285 -159.285 -56.955 -158.955 ;
        RECT -57.285 -162.005 -56.955 -161.675 ;
        RECT -57.285 -163.365 -56.955 -163.035 ;
        RECT -57.285 -164.725 -56.955 -164.395 ;
        RECT -57.285 -166.085 -56.955 -165.755 ;
        RECT -57.285 -167.445 -56.955 -167.115 ;
        RECT -57.285 -168.805 -56.955 -168.475 ;
        RECT -57.285 -170.165 -56.955 -169.835 ;
        RECT -57.285 -171.525 -56.955 -171.195 ;
        RECT -57.285 -172.885 -56.955 -172.555 ;
        RECT -57.285 -174.245 -56.955 -173.915 ;
        RECT -57.285 -175.605 -56.955 -175.275 ;
        RECT -57.285 -176.965 -56.955 -176.635 ;
        RECT -57.285 -178.325 -56.955 -177.995 ;
        RECT -57.285 -179.685 -56.955 -179.355 ;
        RECT -57.285 -181.045 -56.955 -180.715 ;
        RECT -57.285 -182.405 -56.955 -182.075 ;
        RECT -57.285 -183.765 -56.955 -183.435 ;
        RECT -57.285 -185.125 -56.955 -184.795 ;
        RECT -57.285 -186.485 -56.955 -186.155 ;
        RECT -57.285 -187.845 -56.955 -187.515 ;
        RECT -57.285 -189.205 -56.955 -188.875 ;
        RECT -57.285 -190.565 -56.955 -190.235 ;
        RECT -57.285 -191.925 -56.955 -191.595 ;
        RECT -57.285 -193.285 -56.955 -192.955 ;
        RECT -57.285 -194.645 -56.955 -194.315 ;
        RECT -57.285 -196.005 -56.955 -195.675 ;
        RECT -57.285 -197.365 -56.955 -197.035 ;
        RECT -57.285 -198.725 -56.955 -198.395 ;
        RECT -57.285 -200.085 -56.955 -199.755 ;
        RECT -57.285 -201.445 -56.955 -201.115 ;
        RECT -57.285 -202.805 -56.955 -202.475 ;
        RECT -57.285 -204.165 -56.955 -203.835 ;
        RECT -57.285 -205.525 -56.955 -205.195 ;
        RECT -57.285 -206.885 -56.955 -206.555 ;
        RECT -57.285 -208.245 -56.955 -207.915 ;
        RECT -57.285 -209.605 -56.955 -209.275 ;
        RECT -57.285 -210.965 -56.955 -210.635 ;
        RECT -57.285 -212.325 -56.955 -211.995 ;
        RECT -57.285 -213.685 -56.955 -213.355 ;
        RECT -57.285 -215.045 -56.955 -214.715 ;
        RECT -57.285 -216.405 -56.955 -216.075 ;
        RECT -57.285 -217.765 -56.955 -217.435 ;
        RECT -57.285 -219.125 -56.955 -218.795 ;
        RECT -57.285 -220.485 -56.955 -220.155 ;
        RECT -57.285 -221.845 -56.955 -221.515 ;
        RECT -57.285 -223.205 -56.955 -222.875 ;
        RECT -57.285 -224.565 -56.955 -224.235 ;
        RECT -57.285 -226.155 -56.955 -225.825 ;
        RECT -57.285 -227.285 -56.955 -226.955 ;
        RECT -57.285 -228.645 -56.955 -228.315 ;
        RECT -57.285 -231.365 -56.955 -231.035 ;
        RECT -57.285 -234.085 -56.955 -233.755 ;
        RECT -57.285 -235.445 -56.955 -235.115 ;
        RECT -57.285 -236.805 -56.955 -236.475 ;
        RECT -57.285 -238.165 -56.955 -237.835 ;
        RECT -57.285 -243.81 -56.955 -242.68 ;
        RECT -57.28 -243.925 -56.96 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 246.76 -55.595 247.89 ;
        RECT -55.925 241.915 -55.595 242.245 ;
        RECT -55.925 240.555 -55.595 240.885 ;
        RECT -55.925 239.195 -55.595 239.525 ;
        RECT -55.925 237.835 -55.595 238.165 ;
        RECT -55.925 236.475 -55.595 236.805 ;
        RECT -55.925 235.115 -55.595 235.445 ;
        RECT -55.925 233.755 -55.595 234.085 ;
        RECT -55.925 232.395 -55.595 232.725 ;
        RECT -55.925 231.035 -55.595 231.365 ;
        RECT -55.925 229.675 -55.595 230.005 ;
        RECT -55.925 228.315 -55.595 228.645 ;
        RECT -55.925 226.955 -55.595 227.285 ;
        RECT -55.925 225.595 -55.595 225.925 ;
        RECT -55.925 224.235 -55.595 224.565 ;
        RECT -55.925 222.875 -55.595 223.205 ;
        RECT -55.925 221.515 -55.595 221.845 ;
        RECT -55.925 220.155 -55.595 220.485 ;
        RECT -55.925 218.795 -55.595 219.125 ;
        RECT -55.925 217.435 -55.595 217.765 ;
        RECT -55.925 216.075 -55.595 216.405 ;
        RECT -55.925 214.715 -55.595 215.045 ;
        RECT -55.925 213.355 -55.595 213.685 ;
        RECT -55.925 211.995 -55.595 212.325 ;
        RECT -55.925 210.635 -55.595 210.965 ;
        RECT -55.925 209.275 -55.595 209.605 ;
        RECT -55.925 207.915 -55.595 208.245 ;
        RECT -55.925 206.555 -55.595 206.885 ;
        RECT -55.925 205.195 -55.595 205.525 ;
        RECT -55.925 203.835 -55.595 204.165 ;
        RECT -55.925 202.475 -55.595 202.805 ;
        RECT -55.925 201.115 -55.595 201.445 ;
        RECT -55.925 199.755 -55.595 200.085 ;
        RECT -55.925 198.395 -55.595 198.725 ;
        RECT -55.925 197.035 -55.595 197.365 ;
        RECT -55.925 195.675 -55.595 196.005 ;
        RECT -55.925 194.315 -55.595 194.645 ;
        RECT -55.925 192.955 -55.595 193.285 ;
        RECT -55.925 191.595 -55.595 191.925 ;
        RECT -55.925 190.235 -55.595 190.565 ;
        RECT -55.925 188.875 -55.595 189.205 ;
        RECT -55.925 187.515 -55.595 187.845 ;
        RECT -55.925 186.155 -55.595 186.485 ;
        RECT -55.925 184.795 -55.595 185.125 ;
        RECT -55.925 183.435 -55.595 183.765 ;
        RECT -55.925 182.075 -55.595 182.405 ;
        RECT -55.925 180.715 -55.595 181.045 ;
        RECT -55.925 179.355 -55.595 179.685 ;
        RECT -55.925 177.995 -55.595 178.325 ;
        RECT -55.925 176.635 -55.595 176.965 ;
        RECT -55.925 175.275 -55.595 175.605 ;
        RECT -55.925 173.915 -55.595 174.245 ;
        RECT -55.925 172.555 -55.595 172.885 ;
        RECT -55.925 171.195 -55.595 171.525 ;
        RECT -55.925 169.835 -55.595 170.165 ;
        RECT -55.925 168.475 -55.595 168.805 ;
        RECT -55.925 167.115 -55.595 167.445 ;
        RECT -55.925 165.755 -55.595 166.085 ;
        RECT -55.925 164.395 -55.595 164.725 ;
        RECT -55.925 163.035 -55.595 163.365 ;
        RECT -55.925 161.675 -55.595 162.005 ;
        RECT -55.925 160.315 -55.595 160.645 ;
        RECT -55.925 158.955 -55.595 159.285 ;
        RECT -55.925 157.595 -55.595 157.925 ;
        RECT -55.925 156.235 -55.595 156.565 ;
        RECT -55.925 154.875 -55.595 155.205 ;
        RECT -55.925 153.515 -55.595 153.845 ;
        RECT -55.925 152.155 -55.595 152.485 ;
        RECT -55.925 150.795 -55.595 151.125 ;
        RECT -55.925 149.435 -55.595 149.765 ;
        RECT -55.925 148.075 -55.595 148.405 ;
        RECT -55.925 146.715 -55.595 147.045 ;
        RECT -55.925 145.355 -55.595 145.685 ;
        RECT -55.925 143.995 -55.595 144.325 ;
        RECT -55.925 142.635 -55.595 142.965 ;
        RECT -55.925 141.275 -55.595 141.605 ;
        RECT -55.925 139.915 -55.595 140.245 ;
        RECT -55.925 138.555 -55.595 138.885 ;
        RECT -55.925 136.42 -55.595 136.75 ;
        RECT -55.925 134.245 -55.595 134.575 ;
        RECT -55.925 133.395 -55.595 133.725 ;
        RECT -55.925 131.085 -55.595 131.415 ;
        RECT -55.925 130.235 -55.595 130.565 ;
        RECT -55.925 127.925 -55.595 128.255 ;
        RECT -55.925 127.075 -55.595 127.405 ;
        RECT -55.925 124.765 -55.595 125.095 ;
        RECT -55.925 123.915 -55.595 124.245 ;
        RECT -55.925 121.605 -55.595 121.935 ;
        RECT -55.925 120.755 -55.595 121.085 ;
        RECT -55.925 118.445 -55.595 118.775 ;
        RECT -55.925 117.595 -55.595 117.925 ;
        RECT -55.925 115.285 -55.595 115.615 ;
        RECT -55.925 114.435 -55.595 114.765 ;
        RECT -55.925 112.125 -55.595 112.455 ;
        RECT -55.925 111.275 -55.595 111.605 ;
        RECT -55.925 108.965 -55.595 109.295 ;
        RECT -55.925 108.115 -55.595 108.445 ;
        RECT -55.925 105.805 -55.595 106.135 ;
        RECT -55.925 104.955 -55.595 105.285 ;
        RECT -55.925 102.645 -55.595 102.975 ;
        RECT -55.925 101.795 -55.595 102.125 ;
        RECT -55.925 99.62 -55.595 99.95 ;
        RECT -55.925 97.755 -55.595 98.085 ;
        RECT -55.925 96.395 -55.595 96.725 ;
        RECT -55.925 95.035 -55.595 95.365 ;
        RECT -55.925 93.675 -55.595 94.005 ;
        RECT -55.925 92.315 -55.595 92.645 ;
        RECT -55.925 90.955 -55.595 91.285 ;
        RECT -55.925 89.595 -55.595 89.925 ;
        RECT -55.925 88.235 -55.595 88.565 ;
        RECT -55.92 87.56 -55.6 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 -12.405 -55.595 -12.075 ;
        RECT -55.925 -13.765 -55.595 -13.435 ;
        RECT -55.925 -15.125 -55.595 -14.795 ;
        RECT -55.925 -16.485 -55.595 -16.155 ;
        RECT -55.925 -17.845 -55.595 -17.515 ;
        RECT -55.925 -19.205 -55.595 -18.875 ;
        RECT -55.925 -20.565 -55.595 -20.235 ;
        RECT -55.925 -21.925 -55.595 -21.595 ;
        RECT -55.925 -23.285 -55.595 -22.955 ;
        RECT -55.925 -24.645 -55.595 -24.315 ;
        RECT -55.925 -26.005 -55.595 -25.675 ;
        RECT -55.925 -27.365 -55.595 -27.035 ;
        RECT -55.925 -28.725 -55.595 -28.395 ;
        RECT -55.925 -30.085 -55.595 -29.755 ;
        RECT -55.925 -31.445 -55.595 -31.115 ;
        RECT -55.925 -32.805 -55.595 -32.475 ;
        RECT -55.925 -34.165 -55.595 -33.835 ;
        RECT -55.925 -35.525 -55.595 -35.195 ;
        RECT -55.925 -36.885 -55.595 -36.555 ;
        RECT -55.925 -38.245 -55.595 -37.915 ;
        RECT -55.925 -39.605 -55.595 -39.275 ;
        RECT -55.925 -40.965 -55.595 -40.635 ;
        RECT -55.925 -42.325 -55.595 -41.995 ;
        RECT -55.925 -43.685 -55.595 -43.355 ;
        RECT -55.925 -45.045 -55.595 -44.715 ;
        RECT -55.925 -46.405 -55.595 -46.075 ;
        RECT -55.925 -47.765 -55.595 -47.435 ;
        RECT -55.925 -49.125 -55.595 -48.795 ;
        RECT -55.925 -50.485 -55.595 -50.155 ;
        RECT -55.925 -51.845 -55.595 -51.515 ;
        RECT -55.925 -53.205 -55.595 -52.875 ;
        RECT -55.925 -54.565 -55.595 -54.235 ;
        RECT -55.925 -55.925 -55.595 -55.595 ;
        RECT -55.925 -57.285 -55.595 -56.955 ;
        RECT -55.925 -58.645 -55.595 -58.315 ;
        RECT -55.925 -60.005 -55.595 -59.675 ;
        RECT -55.925 -61.365 -55.595 -61.035 ;
        RECT -55.925 -62.725 -55.595 -62.395 ;
        RECT -55.925 -64.085 -55.595 -63.755 ;
        RECT -55.925 -65.445 -55.595 -65.115 ;
        RECT -55.925 -66.805 -55.595 -66.475 ;
        RECT -55.925 -68.165 -55.595 -67.835 ;
        RECT -55.925 -69.525 -55.595 -69.195 ;
        RECT -55.925 -70.885 -55.595 -70.555 ;
        RECT -55.925 -72.245 -55.595 -71.915 ;
        RECT -55.925 -73.605 -55.595 -73.275 ;
        RECT -55.925 -74.965 -55.595 -74.635 ;
        RECT -55.925 -76.325 -55.595 -75.995 ;
        RECT -55.925 -77.685 -55.595 -77.355 ;
        RECT -55.925 -79.045 -55.595 -78.715 ;
        RECT -55.925 -80.405 -55.595 -80.075 ;
        RECT -55.925 -81.765 -55.595 -81.435 ;
        RECT -55.925 -83.125 -55.595 -82.795 ;
        RECT -55.925 -84.485 -55.595 -84.155 ;
        RECT -55.925 -85.845 -55.595 -85.515 ;
        RECT -55.925 -87.205 -55.595 -86.875 ;
        RECT -55.925 -88.565 -55.595 -88.235 ;
        RECT -55.925 -89.925 -55.595 -89.595 ;
        RECT -55.925 -91.285 -55.595 -90.955 ;
        RECT -55.925 -92.645 -55.595 -92.315 ;
        RECT -55.925 -94.005 -55.595 -93.675 ;
        RECT -55.925 -95.365 -55.595 -95.035 ;
        RECT -55.925 -96.725 -55.595 -96.395 ;
        RECT -55.925 -98.085 -55.595 -97.755 ;
        RECT -55.925 -99.445 -55.595 -99.115 ;
        RECT -55.925 -100.805 -55.595 -100.475 ;
        RECT -55.925 -102.165 -55.595 -101.835 ;
        RECT -55.925 -103.525 -55.595 -103.195 ;
        RECT -55.925 -104.885 -55.595 -104.555 ;
        RECT -55.925 -106.245 -55.595 -105.915 ;
        RECT -55.925 -107.605 -55.595 -107.275 ;
        RECT -55.925 -108.965 -55.595 -108.635 ;
        RECT -55.925 -110.325 -55.595 -109.995 ;
        RECT -55.925 -111.685 -55.595 -111.355 ;
        RECT -55.925 -113.045 -55.595 -112.715 ;
        RECT -55.925 -114.405 -55.595 -114.075 ;
        RECT -55.925 -115.765 -55.595 -115.435 ;
        RECT -55.925 -117.125 -55.595 -116.795 ;
        RECT -55.925 -118.485 -55.595 -118.155 ;
        RECT -55.925 -119.845 -55.595 -119.515 ;
        RECT -55.925 -121.205 -55.595 -120.875 ;
        RECT -55.925 -122.565 -55.595 -122.235 ;
        RECT -55.925 -123.925 -55.595 -123.595 ;
        RECT -55.925 -129.365 -55.595 -129.035 ;
        RECT -55.925 -130.725 -55.595 -130.395 ;
        RECT -55.925 -131.47 -55.595 -131.14 ;
        RECT -55.925 -133.445 -55.595 -133.115 ;
        RECT -55.925 -134.805 -55.595 -134.475 ;
        RECT -55.925 -136.165 -55.595 -135.835 ;
        RECT -55.925 -137.525 -55.595 -137.195 ;
        RECT -55.925 -140.245 -55.595 -139.915 ;
        RECT -55.925 -141.605 -55.595 -141.275 ;
        RECT -55.925 -142.965 -55.595 -142.635 ;
        RECT -55.925 -144.31 -55.595 -143.98 ;
        RECT -55.925 -145.685 -55.595 -145.355 ;
        RECT -55.925 -147.045 -55.595 -146.715 ;
        RECT -55.925 -149.765 -55.595 -149.435 ;
        RECT -55.925 -152.485 -55.595 -152.155 ;
        RECT -55.925 -153.845 -55.595 -153.515 ;
        RECT -55.925 -155.205 -55.595 -154.875 ;
        RECT -55.925 -156.565 -55.595 -156.235 ;
        RECT -55.925 -157.925 -55.595 -157.595 ;
        RECT -55.925 -159.285 -55.595 -158.955 ;
        RECT -55.925 -162.005 -55.595 -161.675 ;
        RECT -55.925 -163.365 -55.595 -163.035 ;
        RECT -55.925 -164.725 -55.595 -164.395 ;
        RECT -55.925 -166.085 -55.595 -165.755 ;
        RECT -55.925 -167.445 -55.595 -167.115 ;
        RECT -55.925 -168.805 -55.595 -168.475 ;
        RECT -55.925 -170.165 -55.595 -169.835 ;
        RECT -55.925 -171.525 -55.595 -171.195 ;
        RECT -55.925 -172.885 -55.595 -172.555 ;
        RECT -55.925 -174.245 -55.595 -173.915 ;
        RECT -55.925 -175.605 -55.595 -175.275 ;
        RECT -55.925 -176.965 -55.595 -176.635 ;
        RECT -55.925 -178.325 -55.595 -177.995 ;
        RECT -55.925 -179.685 -55.595 -179.355 ;
        RECT -55.925 -181.045 -55.595 -180.715 ;
        RECT -55.925 -182.405 -55.595 -182.075 ;
        RECT -55.925 -183.765 -55.595 -183.435 ;
        RECT -55.925 -185.125 -55.595 -184.795 ;
        RECT -55.925 -186.485 -55.595 -186.155 ;
        RECT -55.925 -187.845 -55.595 -187.515 ;
        RECT -55.925 -189.205 -55.595 -188.875 ;
        RECT -55.925 -190.565 -55.595 -190.235 ;
        RECT -55.925 -191.925 -55.595 -191.595 ;
        RECT -55.925 -193.285 -55.595 -192.955 ;
        RECT -55.925 -194.645 -55.595 -194.315 ;
        RECT -55.925 -196.005 -55.595 -195.675 ;
        RECT -55.925 -197.365 -55.595 -197.035 ;
        RECT -55.925 -198.725 -55.595 -198.395 ;
        RECT -55.925 -200.085 -55.595 -199.755 ;
        RECT -55.925 -201.445 -55.595 -201.115 ;
        RECT -55.925 -202.805 -55.595 -202.475 ;
        RECT -55.925 -204.165 -55.595 -203.835 ;
        RECT -55.925 -205.525 -55.595 -205.195 ;
        RECT -55.925 -206.885 -55.595 -206.555 ;
        RECT -55.925 -208.245 -55.595 -207.915 ;
        RECT -55.925 -209.605 -55.595 -209.275 ;
        RECT -55.925 -210.965 -55.595 -210.635 ;
        RECT -55.925 -212.325 -55.595 -211.995 ;
        RECT -55.925 -213.685 -55.595 -213.355 ;
        RECT -55.925 -215.045 -55.595 -214.715 ;
        RECT -55.925 -216.405 -55.595 -216.075 ;
        RECT -55.925 -217.765 -55.595 -217.435 ;
        RECT -55.925 -219.125 -55.595 -218.795 ;
        RECT -55.925 -220.485 -55.595 -220.155 ;
        RECT -55.925 -221.845 -55.595 -221.515 ;
        RECT -55.925 -223.205 -55.595 -222.875 ;
        RECT -55.925 -224.565 -55.595 -224.235 ;
        RECT -55.925 -226.155 -55.595 -225.825 ;
        RECT -55.925 -227.285 -55.595 -226.955 ;
        RECT -55.925 -228.645 -55.595 -228.315 ;
        RECT -55.925 -230.005 -55.595 -229.675 ;
        RECT -55.925 -231.365 -55.595 -231.035 ;
        RECT -55.925 -234.085 -55.595 -233.755 ;
        RECT -55.925 -235.445 -55.595 -235.115 ;
        RECT -55.925 -236.805 -55.595 -236.475 ;
        RECT -55.925 -238.165 -55.595 -237.835 ;
        RECT -55.925 -243.81 -55.595 -242.68 ;
        RECT -55.92 -243.925 -55.6 -11.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 232.395 -54.235 232.725 ;
        RECT -54.565 231.035 -54.235 231.365 ;
        RECT -54.565 229.675 -54.235 230.005 ;
        RECT -54.565 228.315 -54.235 228.645 ;
        RECT -54.565 226.955 -54.235 227.285 ;
        RECT -54.565 225.595 -54.235 225.925 ;
        RECT -54.565 224.235 -54.235 224.565 ;
        RECT -54.565 222.875 -54.235 223.205 ;
        RECT -54.565 221.515 -54.235 221.845 ;
        RECT -54.565 220.155 -54.235 220.485 ;
        RECT -54.565 218.795 -54.235 219.125 ;
        RECT -54.565 217.435 -54.235 217.765 ;
        RECT -54.565 216.075 -54.235 216.405 ;
        RECT -54.565 214.715 -54.235 215.045 ;
        RECT -54.565 213.355 -54.235 213.685 ;
        RECT -54.565 211.995 -54.235 212.325 ;
        RECT -54.565 210.635 -54.235 210.965 ;
        RECT -54.565 209.275 -54.235 209.605 ;
        RECT -54.565 207.915 -54.235 208.245 ;
        RECT -54.565 206.555 -54.235 206.885 ;
        RECT -54.565 205.195 -54.235 205.525 ;
        RECT -54.565 203.835 -54.235 204.165 ;
        RECT -54.565 202.475 -54.235 202.805 ;
        RECT -54.565 201.115 -54.235 201.445 ;
        RECT -54.565 199.755 -54.235 200.085 ;
        RECT -54.565 198.395 -54.235 198.725 ;
        RECT -54.565 197.035 -54.235 197.365 ;
        RECT -54.565 195.675 -54.235 196.005 ;
        RECT -54.565 194.315 -54.235 194.645 ;
        RECT -54.565 192.955 -54.235 193.285 ;
        RECT -54.565 191.595 -54.235 191.925 ;
        RECT -54.565 190.235 -54.235 190.565 ;
        RECT -54.565 188.875 -54.235 189.205 ;
        RECT -54.565 187.515 -54.235 187.845 ;
        RECT -54.565 186.155 -54.235 186.485 ;
        RECT -54.565 184.795 -54.235 185.125 ;
        RECT -54.565 183.435 -54.235 183.765 ;
        RECT -54.565 182.075 -54.235 182.405 ;
        RECT -54.565 180.715 -54.235 181.045 ;
        RECT -54.565 179.355 -54.235 179.685 ;
        RECT -54.565 177.995 -54.235 178.325 ;
        RECT -54.565 176.635 -54.235 176.965 ;
        RECT -54.565 175.275 -54.235 175.605 ;
        RECT -54.565 173.915 -54.235 174.245 ;
        RECT -54.565 172.555 -54.235 172.885 ;
        RECT -54.565 171.195 -54.235 171.525 ;
        RECT -54.565 169.835 -54.235 170.165 ;
        RECT -54.565 168.475 -54.235 168.805 ;
        RECT -54.565 167.115 -54.235 167.445 ;
        RECT -54.565 165.755 -54.235 166.085 ;
        RECT -54.565 164.395 -54.235 164.725 ;
        RECT -54.565 163.035 -54.235 163.365 ;
        RECT -54.565 161.675 -54.235 162.005 ;
        RECT -54.565 160.315 -54.235 160.645 ;
        RECT -54.565 158.955 -54.235 159.285 ;
        RECT -54.565 157.595 -54.235 157.925 ;
        RECT -54.565 156.235 -54.235 156.565 ;
        RECT -54.565 154.875 -54.235 155.205 ;
        RECT -54.565 153.515 -54.235 153.845 ;
        RECT -54.565 152.155 -54.235 152.485 ;
        RECT -54.565 150.795 -54.235 151.125 ;
        RECT -54.565 149.435 -54.235 149.765 ;
        RECT -54.565 148.075 -54.235 148.405 ;
        RECT -54.565 146.715 -54.235 147.045 ;
        RECT -54.565 145.355 -54.235 145.685 ;
        RECT -54.565 143.995 -54.235 144.325 ;
        RECT -54.565 142.635 -54.235 142.965 ;
        RECT -54.565 141.275 -54.235 141.605 ;
        RECT -54.565 139.915 -54.235 140.245 ;
        RECT -54.565 138.555 -54.235 138.885 ;
        RECT -54.56 138.555 -54.24 248.005 ;
        RECT -54.565 246.76 -54.235 247.89 ;
        RECT -54.565 241.915 -54.235 242.245 ;
        RECT -54.565 240.555 -54.235 240.885 ;
        RECT -54.565 239.195 -54.235 239.525 ;
        RECT -54.565 237.835 -54.235 238.165 ;
        RECT -54.565 236.475 -54.235 236.805 ;
        RECT -54.565 235.115 -54.235 235.445 ;
        RECT -54.565 233.755 -54.235 234.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.365 246.76 -61.035 247.89 ;
        RECT -61.365 241.915 -61.035 242.245 ;
        RECT -61.365 240.555 -61.035 240.885 ;
        RECT -61.365 239.195 -61.035 239.525 ;
        RECT -61.365 237.835 -61.035 238.165 ;
        RECT -61.365 236.475 -61.035 236.805 ;
        RECT -61.365 235.115 -61.035 235.445 ;
        RECT -61.365 233.755 -61.035 234.085 ;
        RECT -61.365 232.395 -61.035 232.725 ;
        RECT -61.365 231.035 -61.035 231.365 ;
        RECT -61.365 229.675 -61.035 230.005 ;
        RECT -61.365 228.315 -61.035 228.645 ;
        RECT -61.365 226.955 -61.035 227.285 ;
        RECT -61.365 225.595 -61.035 225.925 ;
        RECT -61.365 224.235 -61.035 224.565 ;
        RECT -61.365 222.875 -61.035 223.205 ;
        RECT -61.365 221.515 -61.035 221.845 ;
        RECT -61.365 220.155 -61.035 220.485 ;
        RECT -61.365 218.795 -61.035 219.125 ;
        RECT -61.365 217.435 -61.035 217.765 ;
        RECT -61.365 216.075 -61.035 216.405 ;
        RECT -61.365 214.715 -61.035 215.045 ;
        RECT -61.365 213.355 -61.035 213.685 ;
        RECT -61.365 211.995 -61.035 212.325 ;
        RECT -61.365 210.635 -61.035 210.965 ;
        RECT -61.365 209.275 -61.035 209.605 ;
        RECT -61.365 207.915 -61.035 208.245 ;
        RECT -61.365 206.555 -61.035 206.885 ;
        RECT -61.365 205.195 -61.035 205.525 ;
        RECT -61.365 203.835 -61.035 204.165 ;
        RECT -61.365 202.475 -61.035 202.805 ;
        RECT -61.365 201.115 -61.035 201.445 ;
        RECT -61.365 199.755 -61.035 200.085 ;
        RECT -61.365 198.395 -61.035 198.725 ;
        RECT -61.365 197.035 -61.035 197.365 ;
        RECT -61.365 195.675 -61.035 196.005 ;
        RECT -61.365 194.315 -61.035 194.645 ;
        RECT -61.365 192.955 -61.035 193.285 ;
        RECT -61.365 191.595 -61.035 191.925 ;
        RECT -61.365 190.235 -61.035 190.565 ;
        RECT -61.365 188.875 -61.035 189.205 ;
        RECT -61.365 187.515 -61.035 187.845 ;
        RECT -61.365 186.155 -61.035 186.485 ;
        RECT -61.365 184.795 -61.035 185.125 ;
        RECT -61.365 183.435 -61.035 183.765 ;
        RECT -61.365 182.075 -61.035 182.405 ;
        RECT -61.365 180.715 -61.035 181.045 ;
        RECT -61.365 179.355 -61.035 179.685 ;
        RECT -61.365 177.995 -61.035 178.325 ;
        RECT -61.365 176.635 -61.035 176.965 ;
        RECT -61.365 175.275 -61.035 175.605 ;
        RECT -61.365 173.915 -61.035 174.245 ;
        RECT -61.365 172.555 -61.035 172.885 ;
        RECT -61.365 171.195 -61.035 171.525 ;
        RECT -61.365 169.835 -61.035 170.165 ;
        RECT -61.365 168.475 -61.035 168.805 ;
        RECT -61.365 167.115 -61.035 167.445 ;
        RECT -61.365 165.755 -61.035 166.085 ;
        RECT -61.365 164.395 -61.035 164.725 ;
        RECT -61.365 163.035 -61.035 163.365 ;
        RECT -61.365 161.675 -61.035 162.005 ;
        RECT -61.365 160.315 -61.035 160.645 ;
        RECT -61.365 158.955 -61.035 159.285 ;
        RECT -61.365 157.595 -61.035 157.925 ;
        RECT -61.365 156.235 -61.035 156.565 ;
        RECT -61.365 154.875 -61.035 155.205 ;
        RECT -61.365 153.515 -61.035 153.845 ;
        RECT -61.365 152.155 -61.035 152.485 ;
        RECT -61.365 150.795 -61.035 151.125 ;
        RECT -61.365 149.435 -61.035 149.765 ;
        RECT -61.365 148.075 -61.035 148.405 ;
        RECT -61.365 146.715 -61.035 147.045 ;
        RECT -61.365 145.355 -61.035 145.685 ;
        RECT -61.365 143.995 -61.035 144.325 ;
        RECT -61.365 142.635 -61.035 142.965 ;
        RECT -61.365 141.275 -61.035 141.605 ;
        RECT -61.365 139.915 -61.035 140.245 ;
        RECT -61.365 138.555 -61.035 138.885 ;
        RECT -61.365 97.755 -61.035 98.085 ;
        RECT -61.365 96.395 -61.035 96.725 ;
        RECT -61.365 95.035 -61.035 95.365 ;
        RECT -61.365 93.675 -61.035 94.005 ;
        RECT -61.365 92.315 -61.035 92.645 ;
        RECT -61.365 90.955 -61.035 91.285 ;
        RECT -61.365 89.595 -61.035 89.925 ;
        RECT -61.365 88.235 -61.035 88.565 ;
        RECT -61.365 86.875 -61.035 87.205 ;
        RECT -61.365 85.515 -61.035 85.845 ;
        RECT -61.365 84.155 -61.035 84.485 ;
        RECT -61.365 82.795 -61.035 83.125 ;
        RECT -61.365 81.435 -61.035 81.765 ;
        RECT -61.365 80.075 -61.035 80.405 ;
        RECT -61.365 78.715 -61.035 79.045 ;
        RECT -61.365 77.355 -61.035 77.685 ;
        RECT -61.365 75.995 -61.035 76.325 ;
        RECT -61.365 74.635 -61.035 74.965 ;
        RECT -61.365 73.275 -61.035 73.605 ;
        RECT -61.365 71.915 -61.035 72.245 ;
        RECT -61.365 70.555 -61.035 70.885 ;
        RECT -61.365 69.195 -61.035 69.525 ;
        RECT -61.365 67.835 -61.035 68.165 ;
        RECT -61.365 66.475 -61.035 66.805 ;
        RECT -61.365 65.115 -61.035 65.445 ;
        RECT -61.365 63.755 -61.035 64.085 ;
        RECT -61.365 62.395 -61.035 62.725 ;
        RECT -61.365 61.035 -61.035 61.365 ;
        RECT -61.365 59.675 -61.035 60.005 ;
        RECT -61.365 58.315 -61.035 58.645 ;
        RECT -61.365 56.955 -61.035 57.285 ;
        RECT -61.365 55.595 -61.035 55.925 ;
        RECT -61.365 54.235 -61.035 54.565 ;
        RECT -61.365 52.875 -61.035 53.205 ;
        RECT -61.365 51.515 -61.035 51.845 ;
        RECT -61.365 50.155 -61.035 50.485 ;
        RECT -61.365 48.795 -61.035 49.125 ;
        RECT -61.365 47.435 -61.035 47.765 ;
        RECT -61.365 46.075 -61.035 46.405 ;
        RECT -61.365 44.715 -61.035 45.045 ;
        RECT -61.365 43.355 -61.035 43.685 ;
        RECT -61.365 41.995 -61.035 42.325 ;
        RECT -61.365 40.635 -61.035 40.965 ;
        RECT -61.365 39.275 -61.035 39.605 ;
        RECT -61.365 37.915 -61.035 38.245 ;
        RECT -61.365 36.555 -61.035 36.885 ;
        RECT -61.365 35.195 -61.035 35.525 ;
        RECT -61.365 33.835 -61.035 34.165 ;
        RECT -61.365 32.475 -61.035 32.805 ;
        RECT -61.365 31.115 -61.035 31.445 ;
        RECT -61.365 29.755 -61.035 30.085 ;
        RECT -61.365 28.395 -61.035 28.725 ;
        RECT -61.365 27.035 -61.035 27.365 ;
        RECT -61.365 25.675 -61.035 26.005 ;
        RECT -61.365 24.315 -61.035 24.645 ;
        RECT -61.365 22.955 -61.035 23.285 ;
        RECT -61.365 21.595 -61.035 21.925 ;
        RECT -61.365 20.235 -61.035 20.565 ;
        RECT -61.365 18.875 -61.035 19.205 ;
        RECT -61.365 17.515 -61.035 17.845 ;
        RECT -61.365 16.155 -61.035 16.485 ;
        RECT -61.365 14.795 -61.035 15.125 ;
        RECT -61.365 13.435 -61.035 13.765 ;
        RECT -61.365 12.075 -61.035 12.405 ;
        RECT -61.365 10.715 -61.035 11.045 ;
        RECT -61.365 9.355 -61.035 9.685 ;
        RECT -61.365 7.995 -61.035 8.325 ;
        RECT -61.365 6.635 -61.035 6.965 ;
        RECT -61.365 5.275 -61.035 5.605 ;
        RECT -61.365 3.915 -61.035 4.245 ;
        RECT -61.365 2.555 -61.035 2.885 ;
        RECT -61.365 1.195 -61.035 1.525 ;
        RECT -61.365 -0.165 -61.035 0.165 ;
        RECT -61.365 -1.525 -61.035 -1.195 ;
        RECT -61.365 -2.885 -61.035 -2.555 ;
        RECT -61.365 -4.245 -61.035 -3.915 ;
        RECT -61.365 -5.605 -61.035 -5.275 ;
        RECT -61.365 -6.965 -61.035 -6.635 ;
        RECT -61.365 -8.325 -61.035 -7.995 ;
        RECT -61.365 -9.685 -61.035 -9.355 ;
        RECT -61.365 -11.045 -61.035 -10.715 ;
        RECT -61.365 -12.405 -61.035 -12.075 ;
        RECT -61.365 -13.765 -61.035 -13.435 ;
        RECT -61.365 -15.125 -61.035 -14.795 ;
        RECT -61.365 -16.485 -61.035 -16.155 ;
        RECT -61.365 -17.845 -61.035 -17.515 ;
        RECT -61.365 -19.205 -61.035 -18.875 ;
        RECT -61.365 -20.565 -61.035 -20.235 ;
        RECT -61.365 -21.925 -61.035 -21.595 ;
        RECT -61.365 -23.285 -61.035 -22.955 ;
        RECT -61.365 -24.645 -61.035 -24.315 ;
        RECT -61.365 -26.005 -61.035 -25.675 ;
        RECT -61.365 -27.365 -61.035 -27.035 ;
        RECT -61.365 -28.725 -61.035 -28.395 ;
        RECT -61.365 -30.085 -61.035 -29.755 ;
        RECT -61.365 -31.445 -61.035 -31.115 ;
        RECT -61.365 -32.805 -61.035 -32.475 ;
        RECT -61.365 -34.165 -61.035 -33.835 ;
        RECT -61.365 -35.525 -61.035 -35.195 ;
        RECT -61.365 -36.885 -61.035 -36.555 ;
        RECT -61.365 -38.245 -61.035 -37.915 ;
        RECT -61.365 -39.605 -61.035 -39.275 ;
        RECT -61.365 -40.965 -61.035 -40.635 ;
        RECT -61.365 -42.325 -61.035 -41.995 ;
        RECT -61.365 -43.685 -61.035 -43.355 ;
        RECT -61.365 -45.045 -61.035 -44.715 ;
        RECT -61.365 -46.405 -61.035 -46.075 ;
        RECT -61.365 -47.765 -61.035 -47.435 ;
        RECT -61.365 -49.125 -61.035 -48.795 ;
        RECT -61.365 -50.485 -61.035 -50.155 ;
        RECT -61.365 -51.845 -61.035 -51.515 ;
        RECT -61.365 -53.205 -61.035 -52.875 ;
        RECT -61.365 -54.565 -61.035 -54.235 ;
        RECT -61.365 -55.925 -61.035 -55.595 ;
        RECT -61.365 -57.285 -61.035 -56.955 ;
        RECT -61.365 -58.645 -61.035 -58.315 ;
        RECT -61.365 -60.005 -61.035 -59.675 ;
        RECT -61.365 -61.365 -61.035 -61.035 ;
        RECT -61.365 -62.725 -61.035 -62.395 ;
        RECT -61.365 -64.085 -61.035 -63.755 ;
        RECT -61.365 -65.445 -61.035 -65.115 ;
        RECT -61.365 -66.805 -61.035 -66.475 ;
        RECT -61.365 -68.165 -61.035 -67.835 ;
        RECT -61.365 -69.525 -61.035 -69.195 ;
        RECT -61.365 -70.885 -61.035 -70.555 ;
        RECT -61.365 -72.245 -61.035 -71.915 ;
        RECT -61.365 -73.605 -61.035 -73.275 ;
        RECT -61.365 -74.965 -61.035 -74.635 ;
        RECT -61.365 -76.325 -61.035 -75.995 ;
        RECT -61.365 -77.685 -61.035 -77.355 ;
        RECT -61.365 -79.045 -61.035 -78.715 ;
        RECT -61.365 -80.405 -61.035 -80.075 ;
        RECT -61.365 -81.765 -61.035 -81.435 ;
        RECT -61.365 -83.125 -61.035 -82.795 ;
        RECT -61.365 -84.485 -61.035 -84.155 ;
        RECT -61.365 -85.845 -61.035 -85.515 ;
        RECT -61.365 -87.205 -61.035 -86.875 ;
        RECT -61.365 -88.565 -61.035 -88.235 ;
        RECT -61.365 -89.925 -61.035 -89.595 ;
        RECT -61.365 -91.285 -61.035 -90.955 ;
        RECT -61.365 -92.645 -61.035 -92.315 ;
        RECT -61.365 -94.005 -61.035 -93.675 ;
        RECT -61.365 -95.365 -61.035 -95.035 ;
        RECT -61.365 -96.725 -61.035 -96.395 ;
        RECT -61.365 -98.085 -61.035 -97.755 ;
        RECT -61.365 -99.445 -61.035 -99.115 ;
        RECT -61.365 -100.805 -61.035 -100.475 ;
        RECT -61.365 -102.165 -61.035 -101.835 ;
        RECT -61.365 -103.525 -61.035 -103.195 ;
        RECT -61.365 -104.885 -61.035 -104.555 ;
        RECT -61.365 -106.245 -61.035 -105.915 ;
        RECT -61.365 -107.605 -61.035 -107.275 ;
        RECT -61.365 -108.965 -61.035 -108.635 ;
        RECT -61.365 -110.325 -61.035 -109.995 ;
        RECT -61.365 -111.685 -61.035 -111.355 ;
        RECT -61.365 -113.045 -61.035 -112.715 ;
        RECT -61.365 -114.405 -61.035 -114.075 ;
        RECT -61.365 -115.765 -61.035 -115.435 ;
        RECT -61.365 -117.125 -61.035 -116.795 ;
        RECT -61.365 -118.485 -61.035 -118.155 ;
        RECT -61.365 -119.845 -61.035 -119.515 ;
        RECT -61.365 -121.205 -61.035 -120.875 ;
        RECT -61.365 -122.565 -61.035 -122.235 ;
        RECT -61.365 -123.925 -61.035 -123.595 ;
        RECT -61.365 -125.285 -61.035 -124.955 ;
        RECT -61.365 -129.365 -61.035 -129.035 ;
        RECT -61.365 -130.725 -61.035 -130.395 ;
        RECT -61.365 -131.47 -61.035 -131.14 ;
        RECT -61.365 -133.445 -61.035 -133.115 ;
        RECT -61.365 -134.805 -61.035 -134.475 ;
        RECT -61.365 -136.165 -61.035 -135.835 ;
        RECT -61.365 -137.525 -61.035 -137.195 ;
        RECT -61.365 -140.245 -61.035 -139.915 ;
        RECT -61.365 -141.605 -61.035 -141.275 ;
        RECT -61.365 -142.965 -61.035 -142.635 ;
        RECT -61.365 -144.31 -61.035 -143.98 ;
        RECT -61.365 -145.685 -61.035 -145.355 ;
        RECT -61.365 -147.045 -61.035 -146.715 ;
        RECT -61.365 -149.765 -61.035 -149.435 ;
        RECT -61.365 -152.485 -61.035 -152.155 ;
        RECT -61.365 -153.845 -61.035 -153.515 ;
        RECT -61.365 -155.205 -61.035 -154.875 ;
        RECT -61.365 -156.565 -61.035 -156.235 ;
        RECT -61.365 -157.925 -61.035 -157.595 ;
        RECT -61.365 -159.285 -61.035 -158.955 ;
        RECT -61.365 -162.005 -61.035 -161.675 ;
        RECT -61.365 -163.365 -61.035 -163.035 ;
        RECT -61.365 -164.725 -61.035 -164.395 ;
        RECT -61.365 -166.085 -61.035 -165.755 ;
        RECT -61.365 -167.445 -61.035 -167.115 ;
        RECT -61.365 -168.805 -61.035 -168.475 ;
        RECT -61.365 -170.165 -61.035 -169.835 ;
        RECT -61.365 -171.525 -61.035 -171.195 ;
        RECT -61.365 -172.885 -61.035 -172.555 ;
        RECT -61.365 -174.245 -61.035 -173.915 ;
        RECT -61.365 -175.605 -61.035 -175.275 ;
        RECT -61.365 -176.965 -61.035 -176.635 ;
        RECT -61.365 -178.325 -61.035 -177.995 ;
        RECT -61.365 -179.685 -61.035 -179.355 ;
        RECT -61.365 -181.045 -61.035 -180.715 ;
        RECT -61.365 -182.405 -61.035 -182.075 ;
        RECT -61.365 -183.765 -61.035 -183.435 ;
        RECT -61.365 -185.125 -61.035 -184.795 ;
        RECT -61.365 -186.485 -61.035 -186.155 ;
        RECT -61.365 -187.845 -61.035 -187.515 ;
        RECT -61.365 -189.205 -61.035 -188.875 ;
        RECT -61.365 -190.565 -61.035 -190.235 ;
        RECT -61.365 -191.925 -61.035 -191.595 ;
        RECT -61.365 -193.285 -61.035 -192.955 ;
        RECT -61.365 -194.645 -61.035 -194.315 ;
        RECT -61.365 -196.005 -61.035 -195.675 ;
        RECT -61.365 -197.365 -61.035 -197.035 ;
        RECT -61.365 -198.725 -61.035 -198.395 ;
        RECT -61.365 -200.085 -61.035 -199.755 ;
        RECT -61.365 -201.445 -61.035 -201.115 ;
        RECT -61.365 -202.805 -61.035 -202.475 ;
        RECT -61.365 -204.165 -61.035 -203.835 ;
        RECT -61.365 -205.525 -61.035 -205.195 ;
        RECT -61.365 -206.885 -61.035 -206.555 ;
        RECT -61.365 -208.245 -61.035 -207.915 ;
        RECT -61.365 -209.605 -61.035 -209.275 ;
        RECT -61.365 -210.965 -61.035 -210.635 ;
        RECT -61.365 -212.325 -61.035 -211.995 ;
        RECT -61.365 -213.685 -61.035 -213.355 ;
        RECT -61.365 -215.045 -61.035 -214.715 ;
        RECT -61.365 -216.405 -61.035 -216.075 ;
        RECT -61.365 -217.765 -61.035 -217.435 ;
        RECT -61.365 -219.125 -61.035 -218.795 ;
        RECT -61.365 -220.485 -61.035 -220.155 ;
        RECT -61.365 -221.845 -61.035 -221.515 ;
        RECT -61.365 -223.205 -61.035 -222.875 ;
        RECT -61.365 -224.565 -61.035 -224.235 ;
        RECT -61.365 -226.155 -61.035 -225.825 ;
        RECT -61.365 -227.285 -61.035 -226.955 ;
        RECT -61.365 -228.645 -61.035 -228.315 ;
        RECT -61.365 -230.005 -61.035 -229.675 ;
        RECT -61.365 -234.085 -61.035 -233.755 ;
        RECT -61.365 -235.445 -61.035 -235.115 ;
        RECT -61.365 -236.805 -61.035 -236.475 ;
        RECT -61.365 -238.165 -61.035 -237.835 ;
        RECT -61.365 -243.81 -61.035 -242.68 ;
        RECT -61.36 -243.925 -61.04 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 246.76 -59.675 247.89 ;
        RECT -60.005 241.915 -59.675 242.245 ;
        RECT -60.005 240.555 -59.675 240.885 ;
        RECT -60.005 239.195 -59.675 239.525 ;
        RECT -60.005 237.835 -59.675 238.165 ;
        RECT -60.005 236.475 -59.675 236.805 ;
        RECT -60.005 235.115 -59.675 235.445 ;
        RECT -60.005 233.755 -59.675 234.085 ;
        RECT -60.005 232.395 -59.675 232.725 ;
        RECT -60.005 231.035 -59.675 231.365 ;
        RECT -60.005 229.675 -59.675 230.005 ;
        RECT -60.005 228.315 -59.675 228.645 ;
        RECT -60.005 226.955 -59.675 227.285 ;
        RECT -60.005 225.595 -59.675 225.925 ;
        RECT -60.005 224.235 -59.675 224.565 ;
        RECT -60.005 222.875 -59.675 223.205 ;
        RECT -60.005 221.515 -59.675 221.845 ;
        RECT -60.005 220.155 -59.675 220.485 ;
        RECT -60.005 218.795 -59.675 219.125 ;
        RECT -60.005 217.435 -59.675 217.765 ;
        RECT -60.005 216.075 -59.675 216.405 ;
        RECT -60.005 214.715 -59.675 215.045 ;
        RECT -60.005 213.355 -59.675 213.685 ;
        RECT -60.005 211.995 -59.675 212.325 ;
        RECT -60.005 210.635 -59.675 210.965 ;
        RECT -60.005 209.275 -59.675 209.605 ;
        RECT -60.005 207.915 -59.675 208.245 ;
        RECT -60.005 206.555 -59.675 206.885 ;
        RECT -60.005 205.195 -59.675 205.525 ;
        RECT -60.005 203.835 -59.675 204.165 ;
        RECT -60.005 202.475 -59.675 202.805 ;
        RECT -60.005 201.115 -59.675 201.445 ;
        RECT -60.005 199.755 -59.675 200.085 ;
        RECT -60.005 198.395 -59.675 198.725 ;
        RECT -60.005 197.035 -59.675 197.365 ;
        RECT -60.005 195.675 -59.675 196.005 ;
        RECT -60.005 194.315 -59.675 194.645 ;
        RECT -60.005 192.955 -59.675 193.285 ;
        RECT -60.005 191.595 -59.675 191.925 ;
        RECT -60.005 190.235 -59.675 190.565 ;
        RECT -60.005 188.875 -59.675 189.205 ;
        RECT -60.005 187.515 -59.675 187.845 ;
        RECT -60.005 186.155 -59.675 186.485 ;
        RECT -60.005 184.795 -59.675 185.125 ;
        RECT -60.005 183.435 -59.675 183.765 ;
        RECT -60.005 182.075 -59.675 182.405 ;
        RECT -60.005 180.715 -59.675 181.045 ;
        RECT -60.005 179.355 -59.675 179.685 ;
        RECT -60.005 177.995 -59.675 178.325 ;
        RECT -60.005 176.635 -59.675 176.965 ;
        RECT -60.005 175.275 -59.675 175.605 ;
        RECT -60.005 173.915 -59.675 174.245 ;
        RECT -60.005 172.555 -59.675 172.885 ;
        RECT -60.005 171.195 -59.675 171.525 ;
        RECT -60.005 169.835 -59.675 170.165 ;
        RECT -60.005 168.475 -59.675 168.805 ;
        RECT -60.005 167.115 -59.675 167.445 ;
        RECT -60.005 165.755 -59.675 166.085 ;
        RECT -60.005 164.395 -59.675 164.725 ;
        RECT -60.005 163.035 -59.675 163.365 ;
        RECT -60.005 161.675 -59.675 162.005 ;
        RECT -60.005 160.315 -59.675 160.645 ;
        RECT -60.005 158.955 -59.675 159.285 ;
        RECT -60.005 157.595 -59.675 157.925 ;
        RECT -60.005 156.235 -59.675 156.565 ;
        RECT -60.005 154.875 -59.675 155.205 ;
        RECT -60.005 153.515 -59.675 153.845 ;
        RECT -60.005 152.155 -59.675 152.485 ;
        RECT -60.005 150.795 -59.675 151.125 ;
        RECT -60.005 149.435 -59.675 149.765 ;
        RECT -60.005 148.075 -59.675 148.405 ;
        RECT -60.005 146.715 -59.675 147.045 ;
        RECT -60.005 145.355 -59.675 145.685 ;
        RECT -60.005 143.995 -59.675 144.325 ;
        RECT -60.005 142.635 -59.675 142.965 ;
        RECT -60.005 141.275 -59.675 141.605 ;
        RECT -60.005 139.915 -59.675 140.245 ;
        RECT -60.005 138.555 -59.675 138.885 ;
        RECT -60.005 136.42 -59.675 136.75 ;
        RECT -60.005 134.245 -59.675 134.575 ;
        RECT -60.005 133.395 -59.675 133.725 ;
        RECT -60.005 131.085 -59.675 131.415 ;
        RECT -60.005 130.235 -59.675 130.565 ;
        RECT -60.005 127.925 -59.675 128.255 ;
        RECT -60.005 127.075 -59.675 127.405 ;
        RECT -60.005 124.765 -59.675 125.095 ;
        RECT -60.005 123.915 -59.675 124.245 ;
        RECT -60.005 121.605 -59.675 121.935 ;
        RECT -60.005 120.755 -59.675 121.085 ;
        RECT -60.005 118.445 -59.675 118.775 ;
        RECT -60.005 117.595 -59.675 117.925 ;
        RECT -60.005 115.285 -59.675 115.615 ;
        RECT -60.005 114.435 -59.675 114.765 ;
        RECT -60.005 112.125 -59.675 112.455 ;
        RECT -60.005 111.275 -59.675 111.605 ;
        RECT -60.005 108.965 -59.675 109.295 ;
        RECT -60.005 108.115 -59.675 108.445 ;
        RECT -60.005 105.805 -59.675 106.135 ;
        RECT -60.005 104.955 -59.675 105.285 ;
        RECT -60.005 102.645 -59.675 102.975 ;
        RECT -60.005 101.795 -59.675 102.125 ;
        RECT -60.005 99.62 -59.675 99.95 ;
        RECT -60.005 97.755 -59.675 98.085 ;
        RECT -60.005 96.395 -59.675 96.725 ;
        RECT -60.005 95.035 -59.675 95.365 ;
        RECT -60.005 93.675 -59.675 94.005 ;
        RECT -60.005 92.315 -59.675 92.645 ;
        RECT -60.005 90.955 -59.675 91.285 ;
        RECT -60.005 89.595 -59.675 89.925 ;
        RECT -60.005 88.235 -59.675 88.565 ;
        RECT -60.005 86.875 -59.675 87.205 ;
        RECT -60.005 85.515 -59.675 85.845 ;
        RECT -60.005 84.155 -59.675 84.485 ;
        RECT -60.005 82.795 -59.675 83.125 ;
        RECT -60.005 81.435 -59.675 81.765 ;
        RECT -60.005 80.075 -59.675 80.405 ;
        RECT -60.005 78.715 -59.675 79.045 ;
        RECT -60.005 77.355 -59.675 77.685 ;
        RECT -60.005 75.995 -59.675 76.325 ;
        RECT -60.005 74.635 -59.675 74.965 ;
        RECT -60.005 73.275 -59.675 73.605 ;
        RECT -60.005 71.915 -59.675 72.245 ;
        RECT -60.005 70.555 -59.675 70.885 ;
        RECT -60.005 69.195 -59.675 69.525 ;
        RECT -60.005 67.835 -59.675 68.165 ;
        RECT -60.005 66.475 -59.675 66.805 ;
        RECT -60.005 65.115 -59.675 65.445 ;
        RECT -60.005 63.755 -59.675 64.085 ;
        RECT -60.005 62.395 -59.675 62.725 ;
        RECT -60.005 61.035 -59.675 61.365 ;
        RECT -60.005 59.675 -59.675 60.005 ;
        RECT -60.005 58.315 -59.675 58.645 ;
        RECT -60.005 56.955 -59.675 57.285 ;
        RECT -60.005 55.595 -59.675 55.925 ;
        RECT -60.005 54.235 -59.675 54.565 ;
        RECT -60.005 52.875 -59.675 53.205 ;
        RECT -60.005 51.515 -59.675 51.845 ;
        RECT -60.005 50.155 -59.675 50.485 ;
        RECT -60.005 48.795 -59.675 49.125 ;
        RECT -60.005 47.435 -59.675 47.765 ;
        RECT -60.005 46.075 -59.675 46.405 ;
        RECT -60.005 44.715 -59.675 45.045 ;
        RECT -60.005 43.355 -59.675 43.685 ;
        RECT -60.005 41.995 -59.675 42.325 ;
        RECT -60.005 40.635 -59.675 40.965 ;
        RECT -60.005 39.275 -59.675 39.605 ;
        RECT -60.005 37.915 -59.675 38.245 ;
        RECT -60.005 36.555 -59.675 36.885 ;
        RECT -60.005 35.195 -59.675 35.525 ;
        RECT -60.005 33.835 -59.675 34.165 ;
        RECT -60.005 32.475 -59.675 32.805 ;
        RECT -60.005 31.115 -59.675 31.445 ;
        RECT -60.005 29.755 -59.675 30.085 ;
        RECT -60.005 28.395 -59.675 28.725 ;
        RECT -60.005 27.035 -59.675 27.365 ;
        RECT -60.005 25.675 -59.675 26.005 ;
        RECT -60.005 24.315 -59.675 24.645 ;
        RECT -60.005 22.955 -59.675 23.285 ;
        RECT -60.005 21.595 -59.675 21.925 ;
        RECT -60.005 20.235 -59.675 20.565 ;
        RECT -60.005 18.875 -59.675 19.205 ;
        RECT -60.005 17.515 -59.675 17.845 ;
        RECT -60.005 16.155 -59.675 16.485 ;
        RECT -60.005 14.795 -59.675 15.125 ;
        RECT -60.005 13.435 -59.675 13.765 ;
        RECT -60.005 12.075 -59.675 12.405 ;
        RECT -60.005 10.715 -59.675 11.045 ;
        RECT -60.005 9.355 -59.675 9.685 ;
        RECT -60.005 7.995 -59.675 8.325 ;
        RECT -60.005 6.635 -59.675 6.965 ;
        RECT -60.005 5.275 -59.675 5.605 ;
        RECT -60.005 3.915 -59.675 4.245 ;
        RECT -60.005 2.555 -59.675 2.885 ;
        RECT -60.005 1.195 -59.675 1.525 ;
        RECT -60.005 -0.165 -59.675 0.165 ;
        RECT -60.005 -1.525 -59.675 -1.195 ;
        RECT -60.005 -2.885 -59.675 -2.555 ;
        RECT -60.005 -4.245 -59.675 -3.915 ;
        RECT -60.005 -5.605 -59.675 -5.275 ;
        RECT -60.005 -6.965 -59.675 -6.635 ;
        RECT -60.005 -8.325 -59.675 -7.995 ;
        RECT -60.005 -9.685 -59.675 -9.355 ;
        RECT -60.005 -11.045 -59.675 -10.715 ;
        RECT -60.005 -12.405 -59.675 -12.075 ;
        RECT -60.005 -13.765 -59.675 -13.435 ;
        RECT -60.005 -15.125 -59.675 -14.795 ;
        RECT -60.005 -16.485 -59.675 -16.155 ;
        RECT -60.005 -17.845 -59.675 -17.515 ;
        RECT -60.005 -19.205 -59.675 -18.875 ;
        RECT -60.005 -20.565 -59.675 -20.235 ;
        RECT -60.005 -21.925 -59.675 -21.595 ;
        RECT -60.005 -23.285 -59.675 -22.955 ;
        RECT -60.005 -24.645 -59.675 -24.315 ;
        RECT -60.005 -26.005 -59.675 -25.675 ;
        RECT -60.005 -27.365 -59.675 -27.035 ;
        RECT -60.005 -28.725 -59.675 -28.395 ;
        RECT -60.005 -30.085 -59.675 -29.755 ;
        RECT -60.005 -31.445 -59.675 -31.115 ;
        RECT -60.005 -32.805 -59.675 -32.475 ;
        RECT -60.005 -34.165 -59.675 -33.835 ;
        RECT -60.005 -35.525 -59.675 -35.195 ;
        RECT -60.005 -36.885 -59.675 -36.555 ;
        RECT -60.005 -38.245 -59.675 -37.915 ;
        RECT -60.005 -39.605 -59.675 -39.275 ;
        RECT -60.005 -40.965 -59.675 -40.635 ;
        RECT -60.005 -42.325 -59.675 -41.995 ;
        RECT -60.005 -43.685 -59.675 -43.355 ;
        RECT -60.005 -45.045 -59.675 -44.715 ;
        RECT -60.005 -46.405 -59.675 -46.075 ;
        RECT -60.005 -47.765 -59.675 -47.435 ;
        RECT -60.005 -49.125 -59.675 -48.795 ;
        RECT -60.005 -50.485 -59.675 -50.155 ;
        RECT -60.005 -51.845 -59.675 -51.515 ;
        RECT -60.005 -53.205 -59.675 -52.875 ;
        RECT -60.005 -54.565 -59.675 -54.235 ;
        RECT -60.005 -55.925 -59.675 -55.595 ;
        RECT -60.005 -57.285 -59.675 -56.955 ;
        RECT -60.005 -58.645 -59.675 -58.315 ;
        RECT -60.005 -60.005 -59.675 -59.675 ;
        RECT -60.005 -61.365 -59.675 -61.035 ;
        RECT -60.005 -62.725 -59.675 -62.395 ;
        RECT -60.005 -64.085 -59.675 -63.755 ;
        RECT -60.005 -65.445 -59.675 -65.115 ;
        RECT -60.005 -66.805 -59.675 -66.475 ;
        RECT -60.005 -68.165 -59.675 -67.835 ;
        RECT -60.005 -69.525 -59.675 -69.195 ;
        RECT -60.005 -70.885 -59.675 -70.555 ;
        RECT -60.005 -72.245 -59.675 -71.915 ;
        RECT -60.005 -73.605 -59.675 -73.275 ;
        RECT -60.005 -74.965 -59.675 -74.635 ;
        RECT -60.005 -76.325 -59.675 -75.995 ;
        RECT -60.005 -77.685 -59.675 -77.355 ;
        RECT -60.005 -79.045 -59.675 -78.715 ;
        RECT -60.005 -80.405 -59.675 -80.075 ;
        RECT -60.005 -81.765 -59.675 -81.435 ;
        RECT -60.005 -83.125 -59.675 -82.795 ;
        RECT -60.005 -84.485 -59.675 -84.155 ;
        RECT -60.005 -85.845 -59.675 -85.515 ;
        RECT -60.005 -87.205 -59.675 -86.875 ;
        RECT -60.005 -88.565 -59.675 -88.235 ;
        RECT -60.005 -89.925 -59.675 -89.595 ;
        RECT -60.005 -91.285 -59.675 -90.955 ;
        RECT -60.005 -92.645 -59.675 -92.315 ;
        RECT -60.005 -94.005 -59.675 -93.675 ;
        RECT -60.005 -95.365 -59.675 -95.035 ;
        RECT -60.005 -96.725 -59.675 -96.395 ;
        RECT -60.005 -98.085 -59.675 -97.755 ;
        RECT -60.005 -99.445 -59.675 -99.115 ;
        RECT -60.005 -100.805 -59.675 -100.475 ;
        RECT -60.005 -102.165 -59.675 -101.835 ;
        RECT -60.005 -103.525 -59.675 -103.195 ;
        RECT -60.005 -104.885 -59.675 -104.555 ;
        RECT -60.005 -106.245 -59.675 -105.915 ;
        RECT -60.005 -107.605 -59.675 -107.275 ;
        RECT -60.005 -108.965 -59.675 -108.635 ;
        RECT -60.005 -110.325 -59.675 -109.995 ;
        RECT -60.005 -111.685 -59.675 -111.355 ;
        RECT -60.005 -113.045 -59.675 -112.715 ;
        RECT -60.005 -114.405 -59.675 -114.075 ;
        RECT -60.005 -115.765 -59.675 -115.435 ;
        RECT -60.005 -117.125 -59.675 -116.795 ;
        RECT -60.005 -118.485 -59.675 -118.155 ;
        RECT -60.005 -119.845 -59.675 -119.515 ;
        RECT -60.005 -121.205 -59.675 -120.875 ;
        RECT -60.005 -122.565 -59.675 -122.235 ;
        RECT -60.005 -123.925 -59.675 -123.595 ;
        RECT -60.005 -125.285 -59.675 -124.955 ;
        RECT -60.005 -129.365 -59.675 -129.035 ;
        RECT -60.005 -130.725 -59.675 -130.395 ;
        RECT -60.005 -131.47 -59.675 -131.14 ;
        RECT -60.005 -133.445 -59.675 -133.115 ;
        RECT -60.005 -134.805 -59.675 -134.475 ;
        RECT -60.005 -136.165 -59.675 -135.835 ;
        RECT -60.005 -137.525 -59.675 -137.195 ;
        RECT -60.005 -140.245 -59.675 -139.915 ;
        RECT -60.005 -141.605 -59.675 -141.275 ;
        RECT -60.005 -142.965 -59.675 -142.635 ;
        RECT -60.005 -144.31 -59.675 -143.98 ;
        RECT -60.005 -145.685 -59.675 -145.355 ;
        RECT -60.005 -147.045 -59.675 -146.715 ;
        RECT -60.005 -149.765 -59.675 -149.435 ;
        RECT -60.005 -153.845 -59.675 -153.515 ;
        RECT -60.005 -155.205 -59.675 -154.875 ;
        RECT -60.005 -156.565 -59.675 -156.235 ;
        RECT -60.005 -157.925 -59.675 -157.595 ;
        RECT -60.005 -159.285 -59.675 -158.955 ;
        RECT -60.005 -162.005 -59.675 -161.675 ;
        RECT -60.005 -163.365 -59.675 -163.035 ;
        RECT -60.005 -164.725 -59.675 -164.395 ;
        RECT -60.005 -166.085 -59.675 -165.755 ;
        RECT -60.005 -167.445 -59.675 -167.115 ;
        RECT -60.005 -168.805 -59.675 -168.475 ;
        RECT -60.005 -170.165 -59.675 -169.835 ;
        RECT -60.005 -171.525 -59.675 -171.195 ;
        RECT -60.005 -172.885 -59.675 -172.555 ;
        RECT -60.005 -174.245 -59.675 -173.915 ;
        RECT -60.005 -175.605 -59.675 -175.275 ;
        RECT -60.005 -176.965 -59.675 -176.635 ;
        RECT -60.005 -178.325 -59.675 -177.995 ;
        RECT -60.005 -179.685 -59.675 -179.355 ;
        RECT -60.005 -181.045 -59.675 -180.715 ;
        RECT -60.005 -182.405 -59.675 -182.075 ;
        RECT -60.005 -183.765 -59.675 -183.435 ;
        RECT -60.005 -185.125 -59.675 -184.795 ;
        RECT -60.005 -186.485 -59.675 -186.155 ;
        RECT -60.005 -187.845 -59.675 -187.515 ;
        RECT -60.005 -189.205 -59.675 -188.875 ;
        RECT -60.005 -190.565 -59.675 -190.235 ;
        RECT -60.005 -191.925 -59.675 -191.595 ;
        RECT -60.005 -193.285 -59.675 -192.955 ;
        RECT -60.005 -194.645 -59.675 -194.315 ;
        RECT -60.005 -196.005 -59.675 -195.675 ;
        RECT -60.005 -197.365 -59.675 -197.035 ;
        RECT -60.005 -198.725 -59.675 -198.395 ;
        RECT -60.005 -200.085 -59.675 -199.755 ;
        RECT -60.005 -201.445 -59.675 -201.115 ;
        RECT -60.005 -202.805 -59.675 -202.475 ;
        RECT -60.005 -204.165 -59.675 -203.835 ;
        RECT -60.005 -205.525 -59.675 -205.195 ;
        RECT -60.005 -206.885 -59.675 -206.555 ;
        RECT -60.005 -208.245 -59.675 -207.915 ;
        RECT -60.005 -209.605 -59.675 -209.275 ;
        RECT -60.005 -210.965 -59.675 -210.635 ;
        RECT -60.005 -212.325 -59.675 -211.995 ;
        RECT -60.005 -213.685 -59.675 -213.355 ;
        RECT -60.005 -215.045 -59.675 -214.715 ;
        RECT -60.005 -216.405 -59.675 -216.075 ;
        RECT -60.005 -217.765 -59.675 -217.435 ;
        RECT -60.005 -219.125 -59.675 -218.795 ;
        RECT -60.005 -220.485 -59.675 -220.155 ;
        RECT -60.005 -221.845 -59.675 -221.515 ;
        RECT -60.005 -223.205 -59.675 -222.875 ;
        RECT -60.005 -224.565 -59.675 -224.235 ;
        RECT -60.005 -227.285 -59.675 -226.955 ;
        RECT -60.005 -228.645 -59.675 -228.315 ;
        RECT -60.005 -234.085 -59.675 -233.755 ;
        RECT -60.005 -235.445 -59.675 -235.115 ;
        RECT -60.005 -236.805 -59.675 -236.475 ;
        RECT -60.005 -238.165 -59.675 -237.835 ;
        RECT -60.005 -243.81 -59.675 -242.68 ;
        RECT -60 -243.925 -59.68 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.645 -201.445 -58.315 -201.115 ;
        RECT -58.645 -202.805 -58.315 -202.475 ;
        RECT -58.645 -204.165 -58.315 -203.835 ;
        RECT -58.645 -205.525 -58.315 -205.195 ;
        RECT -58.645 -206.885 -58.315 -206.555 ;
        RECT -58.645 -208.245 -58.315 -207.915 ;
        RECT -58.645 -209.605 -58.315 -209.275 ;
        RECT -58.645 -210.965 -58.315 -210.635 ;
        RECT -58.645 -212.325 -58.315 -211.995 ;
        RECT -58.645 -213.685 -58.315 -213.355 ;
        RECT -58.645 -215.045 -58.315 -214.715 ;
        RECT -58.645 -216.405 -58.315 -216.075 ;
        RECT -58.645 -217.765 -58.315 -217.435 ;
        RECT -58.645 -219.125 -58.315 -218.795 ;
        RECT -58.645 -220.485 -58.315 -220.155 ;
        RECT -58.645 -221.845 -58.315 -221.515 ;
        RECT -58.645 -223.205 -58.315 -222.875 ;
        RECT -58.645 -224.565 -58.315 -224.235 ;
        RECT -58.645 -226.155 -58.315 -225.825 ;
        RECT -58.645 -227.285 -58.315 -226.955 ;
        RECT -58.645 -228.645 -58.315 -228.315 ;
        RECT -58.64 -229.32 -58.32 248.005 ;
        RECT -58.645 246.76 -58.315 247.89 ;
        RECT -58.645 241.915 -58.315 242.245 ;
        RECT -58.645 240.555 -58.315 240.885 ;
        RECT -58.645 239.195 -58.315 239.525 ;
        RECT -58.645 237.835 -58.315 238.165 ;
        RECT -58.645 236.475 -58.315 236.805 ;
        RECT -58.645 235.115 -58.315 235.445 ;
        RECT -58.645 233.755 -58.315 234.085 ;
        RECT -58.645 232.395 -58.315 232.725 ;
        RECT -58.645 231.035 -58.315 231.365 ;
        RECT -58.645 229.675 -58.315 230.005 ;
        RECT -58.645 228.315 -58.315 228.645 ;
        RECT -58.645 226.955 -58.315 227.285 ;
        RECT -58.645 225.595 -58.315 225.925 ;
        RECT -58.645 224.235 -58.315 224.565 ;
        RECT -58.645 222.875 -58.315 223.205 ;
        RECT -58.645 221.515 -58.315 221.845 ;
        RECT -58.645 220.155 -58.315 220.485 ;
        RECT -58.645 218.795 -58.315 219.125 ;
        RECT -58.645 217.435 -58.315 217.765 ;
        RECT -58.645 216.075 -58.315 216.405 ;
        RECT -58.645 214.715 -58.315 215.045 ;
        RECT -58.645 213.355 -58.315 213.685 ;
        RECT -58.645 211.995 -58.315 212.325 ;
        RECT -58.645 210.635 -58.315 210.965 ;
        RECT -58.645 209.275 -58.315 209.605 ;
        RECT -58.645 207.915 -58.315 208.245 ;
        RECT -58.645 206.555 -58.315 206.885 ;
        RECT -58.645 205.195 -58.315 205.525 ;
        RECT -58.645 203.835 -58.315 204.165 ;
        RECT -58.645 202.475 -58.315 202.805 ;
        RECT -58.645 201.115 -58.315 201.445 ;
        RECT -58.645 199.755 -58.315 200.085 ;
        RECT -58.645 198.395 -58.315 198.725 ;
        RECT -58.645 197.035 -58.315 197.365 ;
        RECT -58.645 195.675 -58.315 196.005 ;
        RECT -58.645 194.315 -58.315 194.645 ;
        RECT -58.645 192.955 -58.315 193.285 ;
        RECT -58.645 191.595 -58.315 191.925 ;
        RECT -58.645 190.235 -58.315 190.565 ;
        RECT -58.645 188.875 -58.315 189.205 ;
        RECT -58.645 187.515 -58.315 187.845 ;
        RECT -58.645 186.155 -58.315 186.485 ;
        RECT -58.645 184.795 -58.315 185.125 ;
        RECT -58.645 183.435 -58.315 183.765 ;
        RECT -58.645 182.075 -58.315 182.405 ;
        RECT -58.645 180.715 -58.315 181.045 ;
        RECT -58.645 179.355 -58.315 179.685 ;
        RECT -58.645 177.995 -58.315 178.325 ;
        RECT -58.645 176.635 -58.315 176.965 ;
        RECT -58.645 175.275 -58.315 175.605 ;
        RECT -58.645 173.915 -58.315 174.245 ;
        RECT -58.645 172.555 -58.315 172.885 ;
        RECT -58.645 171.195 -58.315 171.525 ;
        RECT -58.645 169.835 -58.315 170.165 ;
        RECT -58.645 168.475 -58.315 168.805 ;
        RECT -58.645 167.115 -58.315 167.445 ;
        RECT -58.645 165.755 -58.315 166.085 ;
        RECT -58.645 164.395 -58.315 164.725 ;
        RECT -58.645 163.035 -58.315 163.365 ;
        RECT -58.645 161.675 -58.315 162.005 ;
        RECT -58.645 160.315 -58.315 160.645 ;
        RECT -58.645 158.955 -58.315 159.285 ;
        RECT -58.645 157.595 -58.315 157.925 ;
        RECT -58.645 156.235 -58.315 156.565 ;
        RECT -58.645 154.875 -58.315 155.205 ;
        RECT -58.645 153.515 -58.315 153.845 ;
        RECT -58.645 152.155 -58.315 152.485 ;
        RECT -58.645 150.795 -58.315 151.125 ;
        RECT -58.645 149.435 -58.315 149.765 ;
        RECT -58.645 148.075 -58.315 148.405 ;
        RECT -58.645 146.715 -58.315 147.045 ;
        RECT -58.645 145.355 -58.315 145.685 ;
        RECT -58.645 143.995 -58.315 144.325 ;
        RECT -58.645 142.635 -58.315 142.965 ;
        RECT -58.645 141.275 -58.315 141.605 ;
        RECT -58.645 139.915 -58.315 140.245 ;
        RECT -58.645 138.555 -58.315 138.885 ;
        RECT -58.645 136.42 -58.315 136.75 ;
        RECT -58.645 134.245 -58.315 134.575 ;
        RECT -58.645 133.395 -58.315 133.725 ;
        RECT -58.645 131.085 -58.315 131.415 ;
        RECT -58.645 130.235 -58.315 130.565 ;
        RECT -58.645 127.925 -58.315 128.255 ;
        RECT -58.645 127.075 -58.315 127.405 ;
        RECT -58.645 124.765 -58.315 125.095 ;
        RECT -58.645 123.915 -58.315 124.245 ;
        RECT -58.645 121.605 -58.315 121.935 ;
        RECT -58.645 120.755 -58.315 121.085 ;
        RECT -58.645 118.445 -58.315 118.775 ;
        RECT -58.645 117.595 -58.315 117.925 ;
        RECT -58.645 115.285 -58.315 115.615 ;
        RECT -58.645 114.435 -58.315 114.765 ;
        RECT -58.645 112.125 -58.315 112.455 ;
        RECT -58.645 111.275 -58.315 111.605 ;
        RECT -58.645 108.965 -58.315 109.295 ;
        RECT -58.645 108.115 -58.315 108.445 ;
        RECT -58.645 105.805 -58.315 106.135 ;
        RECT -58.645 104.955 -58.315 105.285 ;
        RECT -58.645 102.645 -58.315 102.975 ;
        RECT -58.645 101.795 -58.315 102.125 ;
        RECT -58.645 99.62 -58.315 99.95 ;
        RECT -58.645 97.755 -58.315 98.085 ;
        RECT -58.645 96.395 -58.315 96.725 ;
        RECT -58.645 95.035 -58.315 95.365 ;
        RECT -58.645 93.675 -58.315 94.005 ;
        RECT -58.645 92.315 -58.315 92.645 ;
        RECT -58.645 90.955 -58.315 91.285 ;
        RECT -58.645 89.595 -58.315 89.925 ;
        RECT -58.645 88.235 -58.315 88.565 ;
        RECT -58.645 86.875 -58.315 87.205 ;
        RECT -58.645 85.515 -58.315 85.845 ;
        RECT -58.645 84.155 -58.315 84.485 ;
        RECT -58.645 82.795 -58.315 83.125 ;
        RECT -58.645 81.435 -58.315 81.765 ;
        RECT -58.645 80.075 -58.315 80.405 ;
        RECT -58.645 78.715 -58.315 79.045 ;
        RECT -58.645 77.355 -58.315 77.685 ;
        RECT -58.645 75.995 -58.315 76.325 ;
        RECT -58.645 74.635 -58.315 74.965 ;
        RECT -58.645 73.275 -58.315 73.605 ;
        RECT -58.645 71.915 -58.315 72.245 ;
        RECT -58.645 70.555 -58.315 70.885 ;
        RECT -58.645 69.195 -58.315 69.525 ;
        RECT -58.645 67.835 -58.315 68.165 ;
        RECT -58.645 66.475 -58.315 66.805 ;
        RECT -58.645 65.115 -58.315 65.445 ;
        RECT -58.645 63.755 -58.315 64.085 ;
        RECT -58.645 62.395 -58.315 62.725 ;
        RECT -58.645 61.035 -58.315 61.365 ;
        RECT -58.645 59.675 -58.315 60.005 ;
        RECT -58.645 58.315 -58.315 58.645 ;
        RECT -58.645 56.955 -58.315 57.285 ;
        RECT -58.645 55.595 -58.315 55.925 ;
        RECT -58.645 54.235 -58.315 54.565 ;
        RECT -58.645 52.875 -58.315 53.205 ;
        RECT -58.645 51.515 -58.315 51.845 ;
        RECT -58.645 50.155 -58.315 50.485 ;
        RECT -58.645 48.795 -58.315 49.125 ;
        RECT -58.645 47.435 -58.315 47.765 ;
        RECT -58.645 46.075 -58.315 46.405 ;
        RECT -58.645 44.715 -58.315 45.045 ;
        RECT -58.645 43.355 -58.315 43.685 ;
        RECT -58.645 41.995 -58.315 42.325 ;
        RECT -58.645 40.635 -58.315 40.965 ;
        RECT -58.645 39.275 -58.315 39.605 ;
        RECT -58.645 37.915 -58.315 38.245 ;
        RECT -58.645 36.555 -58.315 36.885 ;
        RECT -58.645 35.195 -58.315 35.525 ;
        RECT -58.645 33.835 -58.315 34.165 ;
        RECT -58.645 32.475 -58.315 32.805 ;
        RECT -58.645 31.115 -58.315 31.445 ;
        RECT -58.645 29.755 -58.315 30.085 ;
        RECT -58.645 28.395 -58.315 28.725 ;
        RECT -58.645 27.035 -58.315 27.365 ;
        RECT -58.645 25.675 -58.315 26.005 ;
        RECT -58.645 24.315 -58.315 24.645 ;
        RECT -58.645 22.955 -58.315 23.285 ;
        RECT -58.645 21.595 -58.315 21.925 ;
        RECT -58.645 20.235 -58.315 20.565 ;
        RECT -58.645 18.875 -58.315 19.205 ;
        RECT -58.645 17.515 -58.315 17.845 ;
        RECT -58.645 16.155 -58.315 16.485 ;
        RECT -58.645 14.795 -58.315 15.125 ;
        RECT -58.645 13.435 -58.315 13.765 ;
        RECT -58.645 12.075 -58.315 12.405 ;
        RECT -58.645 10.715 -58.315 11.045 ;
        RECT -58.645 9.355 -58.315 9.685 ;
        RECT -58.645 7.995 -58.315 8.325 ;
        RECT -58.645 6.635 -58.315 6.965 ;
        RECT -58.645 5.275 -58.315 5.605 ;
        RECT -58.645 3.915 -58.315 4.245 ;
        RECT -58.645 2.555 -58.315 2.885 ;
        RECT -58.645 1.195 -58.315 1.525 ;
        RECT -58.645 -0.165 -58.315 0.165 ;
        RECT -58.645 -1.525 -58.315 -1.195 ;
        RECT -58.645 -2.885 -58.315 -2.555 ;
        RECT -58.645 -4.245 -58.315 -3.915 ;
        RECT -58.645 -5.605 -58.315 -5.275 ;
        RECT -58.645 -6.965 -58.315 -6.635 ;
        RECT -58.645 -8.325 -58.315 -7.995 ;
        RECT -58.645 -9.685 -58.315 -9.355 ;
        RECT -58.645 -11.045 -58.315 -10.715 ;
        RECT -58.645 -12.405 -58.315 -12.075 ;
        RECT -58.645 -13.765 -58.315 -13.435 ;
        RECT -58.645 -15.125 -58.315 -14.795 ;
        RECT -58.645 -16.485 -58.315 -16.155 ;
        RECT -58.645 -17.845 -58.315 -17.515 ;
        RECT -58.645 -19.205 -58.315 -18.875 ;
        RECT -58.645 -20.565 -58.315 -20.235 ;
        RECT -58.645 -21.925 -58.315 -21.595 ;
        RECT -58.645 -23.285 -58.315 -22.955 ;
        RECT -58.645 -24.645 -58.315 -24.315 ;
        RECT -58.645 -26.005 -58.315 -25.675 ;
        RECT -58.645 -27.365 -58.315 -27.035 ;
        RECT -58.645 -28.725 -58.315 -28.395 ;
        RECT -58.645 -30.085 -58.315 -29.755 ;
        RECT -58.645 -31.445 -58.315 -31.115 ;
        RECT -58.645 -32.805 -58.315 -32.475 ;
        RECT -58.645 -34.165 -58.315 -33.835 ;
        RECT -58.645 -35.525 -58.315 -35.195 ;
        RECT -58.645 -36.885 -58.315 -36.555 ;
        RECT -58.645 -38.245 -58.315 -37.915 ;
        RECT -58.645 -39.605 -58.315 -39.275 ;
        RECT -58.645 -40.965 -58.315 -40.635 ;
        RECT -58.645 -42.325 -58.315 -41.995 ;
        RECT -58.645 -43.685 -58.315 -43.355 ;
        RECT -58.645 -45.045 -58.315 -44.715 ;
        RECT -58.645 -46.405 -58.315 -46.075 ;
        RECT -58.645 -47.765 -58.315 -47.435 ;
        RECT -58.645 -49.125 -58.315 -48.795 ;
        RECT -58.645 -50.485 -58.315 -50.155 ;
        RECT -58.645 -51.845 -58.315 -51.515 ;
        RECT -58.645 -53.205 -58.315 -52.875 ;
        RECT -58.645 -54.565 -58.315 -54.235 ;
        RECT -58.645 -55.925 -58.315 -55.595 ;
        RECT -58.645 -57.285 -58.315 -56.955 ;
        RECT -58.645 -58.645 -58.315 -58.315 ;
        RECT -58.645 -60.005 -58.315 -59.675 ;
        RECT -58.645 -61.365 -58.315 -61.035 ;
        RECT -58.645 -62.725 -58.315 -62.395 ;
        RECT -58.645 -64.085 -58.315 -63.755 ;
        RECT -58.645 -65.445 -58.315 -65.115 ;
        RECT -58.645 -66.805 -58.315 -66.475 ;
        RECT -58.645 -68.165 -58.315 -67.835 ;
        RECT -58.645 -69.525 -58.315 -69.195 ;
        RECT -58.645 -70.885 -58.315 -70.555 ;
        RECT -58.645 -72.245 -58.315 -71.915 ;
        RECT -58.645 -73.605 -58.315 -73.275 ;
        RECT -58.645 -74.965 -58.315 -74.635 ;
        RECT -58.645 -76.325 -58.315 -75.995 ;
        RECT -58.645 -77.685 -58.315 -77.355 ;
        RECT -58.645 -79.045 -58.315 -78.715 ;
        RECT -58.645 -80.405 -58.315 -80.075 ;
        RECT -58.645 -81.765 -58.315 -81.435 ;
        RECT -58.645 -83.125 -58.315 -82.795 ;
        RECT -58.645 -84.485 -58.315 -84.155 ;
        RECT -58.645 -85.845 -58.315 -85.515 ;
        RECT -58.645 -87.205 -58.315 -86.875 ;
        RECT -58.645 -88.565 -58.315 -88.235 ;
        RECT -58.645 -89.925 -58.315 -89.595 ;
        RECT -58.645 -91.285 -58.315 -90.955 ;
        RECT -58.645 -92.645 -58.315 -92.315 ;
        RECT -58.645 -94.005 -58.315 -93.675 ;
        RECT -58.645 -95.365 -58.315 -95.035 ;
        RECT -58.645 -96.725 -58.315 -96.395 ;
        RECT -58.645 -98.085 -58.315 -97.755 ;
        RECT -58.645 -99.445 -58.315 -99.115 ;
        RECT -58.645 -100.805 -58.315 -100.475 ;
        RECT -58.645 -102.165 -58.315 -101.835 ;
        RECT -58.645 -103.525 -58.315 -103.195 ;
        RECT -58.645 -104.885 -58.315 -104.555 ;
        RECT -58.645 -106.245 -58.315 -105.915 ;
        RECT -58.645 -107.605 -58.315 -107.275 ;
        RECT -58.645 -108.965 -58.315 -108.635 ;
        RECT -58.645 -110.325 -58.315 -109.995 ;
        RECT -58.645 -111.685 -58.315 -111.355 ;
        RECT -58.645 -113.045 -58.315 -112.715 ;
        RECT -58.645 -114.405 -58.315 -114.075 ;
        RECT -58.645 -115.765 -58.315 -115.435 ;
        RECT -58.645 -117.125 -58.315 -116.795 ;
        RECT -58.645 -118.485 -58.315 -118.155 ;
        RECT -58.645 -119.845 -58.315 -119.515 ;
        RECT -58.645 -121.205 -58.315 -120.875 ;
        RECT -58.645 -122.565 -58.315 -122.235 ;
        RECT -58.645 -123.925 -58.315 -123.595 ;
        RECT -58.645 -129.365 -58.315 -129.035 ;
        RECT -58.645 -130.725 -58.315 -130.395 ;
        RECT -58.645 -131.47 -58.315 -131.14 ;
        RECT -58.645 -133.445 -58.315 -133.115 ;
        RECT -58.645 -134.805 -58.315 -134.475 ;
        RECT -58.645 -136.165 -58.315 -135.835 ;
        RECT -58.645 -137.525 -58.315 -137.195 ;
        RECT -58.645 -140.245 -58.315 -139.915 ;
        RECT -58.645 -141.605 -58.315 -141.275 ;
        RECT -58.645 -142.965 -58.315 -142.635 ;
        RECT -58.645 -144.31 -58.315 -143.98 ;
        RECT -58.645 -145.685 -58.315 -145.355 ;
        RECT -58.645 -147.045 -58.315 -146.715 ;
        RECT -58.645 -149.765 -58.315 -149.435 ;
        RECT -58.645 -153.845 -58.315 -153.515 ;
        RECT -58.645 -155.205 -58.315 -154.875 ;
        RECT -58.645 -156.565 -58.315 -156.235 ;
        RECT -58.645 -157.925 -58.315 -157.595 ;
        RECT -58.645 -159.285 -58.315 -158.955 ;
        RECT -58.645 -162.005 -58.315 -161.675 ;
        RECT -58.645 -163.365 -58.315 -163.035 ;
        RECT -58.645 -164.725 -58.315 -164.395 ;
        RECT -58.645 -166.085 -58.315 -165.755 ;
        RECT -58.645 -167.445 -58.315 -167.115 ;
        RECT -58.645 -168.805 -58.315 -168.475 ;
        RECT -58.645 -170.165 -58.315 -169.835 ;
        RECT -58.645 -171.525 -58.315 -171.195 ;
        RECT -58.645 -172.885 -58.315 -172.555 ;
        RECT -58.645 -174.245 -58.315 -173.915 ;
        RECT -58.645 -175.605 -58.315 -175.275 ;
        RECT -58.645 -176.965 -58.315 -176.635 ;
        RECT -58.645 -178.325 -58.315 -177.995 ;
        RECT -58.645 -179.685 -58.315 -179.355 ;
        RECT -58.645 -181.045 -58.315 -180.715 ;
        RECT -58.645 -182.405 -58.315 -182.075 ;
        RECT -58.645 -183.765 -58.315 -183.435 ;
        RECT -58.645 -185.125 -58.315 -184.795 ;
        RECT -58.645 -186.485 -58.315 -186.155 ;
        RECT -58.645 -187.845 -58.315 -187.515 ;
        RECT -58.645 -189.205 -58.315 -188.875 ;
        RECT -58.645 -190.565 -58.315 -190.235 ;
        RECT -58.645 -191.925 -58.315 -191.595 ;
        RECT -58.645 -193.285 -58.315 -192.955 ;
        RECT -58.645 -194.645 -58.315 -194.315 ;
        RECT -58.645 -196.005 -58.315 -195.675 ;
        RECT -58.645 -197.365 -58.315 -197.035 ;
        RECT -58.645 -198.725 -58.315 -198.395 ;
        RECT -58.645 -200.085 -58.315 -199.755 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.805 -234.085 -66.475 -233.755 ;
        RECT -66.805 -235.445 -66.475 -235.115 ;
        RECT -66.805 -236.805 -66.475 -236.475 ;
        RECT -66.805 -238.165 -66.475 -237.835 ;
        RECT -66.805 -243.81 -66.475 -242.68 ;
        RECT -66.8 -243.925 -66.48 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.445 246.76 -65.115 247.89 ;
        RECT -65.445 241.915 -65.115 242.245 ;
        RECT -65.445 240.555 -65.115 240.885 ;
        RECT -65.445 239.195 -65.115 239.525 ;
        RECT -65.445 237.835 -65.115 238.165 ;
        RECT -65.445 236.475 -65.115 236.805 ;
        RECT -65.445 235.115 -65.115 235.445 ;
        RECT -65.445 233.755 -65.115 234.085 ;
        RECT -65.445 232.395 -65.115 232.725 ;
        RECT -65.445 231.035 -65.115 231.365 ;
        RECT -65.445 229.675 -65.115 230.005 ;
        RECT -65.445 228.315 -65.115 228.645 ;
        RECT -65.445 226.955 -65.115 227.285 ;
        RECT -65.445 225.595 -65.115 225.925 ;
        RECT -65.445 224.235 -65.115 224.565 ;
        RECT -65.445 222.875 -65.115 223.205 ;
        RECT -65.445 221.515 -65.115 221.845 ;
        RECT -65.445 220.155 -65.115 220.485 ;
        RECT -65.445 218.795 -65.115 219.125 ;
        RECT -65.445 217.435 -65.115 217.765 ;
        RECT -65.445 216.075 -65.115 216.405 ;
        RECT -65.445 214.715 -65.115 215.045 ;
        RECT -65.445 213.355 -65.115 213.685 ;
        RECT -65.445 211.995 -65.115 212.325 ;
        RECT -65.445 210.635 -65.115 210.965 ;
        RECT -65.445 209.275 -65.115 209.605 ;
        RECT -65.445 207.915 -65.115 208.245 ;
        RECT -65.445 206.555 -65.115 206.885 ;
        RECT -65.445 205.195 -65.115 205.525 ;
        RECT -65.445 203.835 -65.115 204.165 ;
        RECT -65.445 202.475 -65.115 202.805 ;
        RECT -65.445 201.115 -65.115 201.445 ;
        RECT -65.445 199.755 -65.115 200.085 ;
        RECT -65.445 198.395 -65.115 198.725 ;
        RECT -65.445 197.035 -65.115 197.365 ;
        RECT -65.445 195.675 -65.115 196.005 ;
        RECT -65.445 194.315 -65.115 194.645 ;
        RECT -65.445 192.955 -65.115 193.285 ;
        RECT -65.445 191.595 -65.115 191.925 ;
        RECT -65.445 190.235 -65.115 190.565 ;
        RECT -65.445 188.875 -65.115 189.205 ;
        RECT -65.445 187.515 -65.115 187.845 ;
        RECT -65.445 186.155 -65.115 186.485 ;
        RECT -65.445 184.795 -65.115 185.125 ;
        RECT -65.445 183.435 -65.115 183.765 ;
        RECT -65.445 182.075 -65.115 182.405 ;
        RECT -65.445 180.715 -65.115 181.045 ;
        RECT -65.445 179.355 -65.115 179.685 ;
        RECT -65.445 177.995 -65.115 178.325 ;
        RECT -65.445 176.635 -65.115 176.965 ;
        RECT -65.445 175.275 -65.115 175.605 ;
        RECT -65.445 173.915 -65.115 174.245 ;
        RECT -65.445 172.555 -65.115 172.885 ;
        RECT -65.445 171.195 -65.115 171.525 ;
        RECT -65.445 169.835 -65.115 170.165 ;
        RECT -65.445 168.475 -65.115 168.805 ;
        RECT -65.445 167.115 -65.115 167.445 ;
        RECT -65.445 165.755 -65.115 166.085 ;
        RECT -65.445 164.395 -65.115 164.725 ;
        RECT -65.445 163.035 -65.115 163.365 ;
        RECT -65.445 161.675 -65.115 162.005 ;
        RECT -65.445 160.315 -65.115 160.645 ;
        RECT -65.445 158.955 -65.115 159.285 ;
        RECT -65.445 157.595 -65.115 157.925 ;
        RECT -65.445 156.235 -65.115 156.565 ;
        RECT -65.445 154.875 -65.115 155.205 ;
        RECT -65.445 153.515 -65.115 153.845 ;
        RECT -65.445 152.155 -65.115 152.485 ;
        RECT -65.445 150.795 -65.115 151.125 ;
        RECT -65.445 149.435 -65.115 149.765 ;
        RECT -65.445 148.075 -65.115 148.405 ;
        RECT -65.445 146.715 -65.115 147.045 ;
        RECT -65.445 145.355 -65.115 145.685 ;
        RECT -65.445 143.995 -65.115 144.325 ;
        RECT -65.445 142.635 -65.115 142.965 ;
        RECT -65.445 141.275 -65.115 141.605 ;
        RECT -65.445 139.915 -65.115 140.245 ;
        RECT -65.445 138.555 -65.115 138.885 ;
        RECT -65.445 137.195 -65.115 137.525 ;
        RECT -65.445 135.835 -65.115 136.165 ;
        RECT -65.445 134.475 -65.115 134.805 ;
        RECT -65.445 133.115 -65.115 133.445 ;
        RECT -65.445 131.755 -65.115 132.085 ;
        RECT -65.445 130.395 -65.115 130.725 ;
        RECT -65.445 129.035 -65.115 129.365 ;
        RECT -65.445 127.675 -65.115 128.005 ;
        RECT -65.445 126.315 -65.115 126.645 ;
        RECT -65.445 124.955 -65.115 125.285 ;
        RECT -65.445 123.595 -65.115 123.925 ;
        RECT -65.445 122.235 -65.115 122.565 ;
        RECT -65.445 120.875 -65.115 121.205 ;
        RECT -65.445 119.515 -65.115 119.845 ;
        RECT -65.445 118.155 -65.115 118.485 ;
        RECT -65.445 116.795 -65.115 117.125 ;
        RECT -65.445 115.435 -65.115 115.765 ;
        RECT -65.445 114.075 -65.115 114.405 ;
        RECT -65.445 112.715 -65.115 113.045 ;
        RECT -65.445 111.355 -65.115 111.685 ;
        RECT -65.445 109.995 -65.115 110.325 ;
        RECT -65.445 108.635 -65.115 108.965 ;
        RECT -65.445 107.275 -65.115 107.605 ;
        RECT -65.445 105.915 -65.115 106.245 ;
        RECT -65.445 104.555 -65.115 104.885 ;
        RECT -65.445 103.195 -65.115 103.525 ;
        RECT -65.445 101.835 -65.115 102.165 ;
        RECT -65.445 100.475 -65.115 100.805 ;
        RECT -65.445 99.115 -65.115 99.445 ;
        RECT -65.445 97.755 -65.115 98.085 ;
        RECT -65.445 96.395 -65.115 96.725 ;
        RECT -65.445 95.035 -65.115 95.365 ;
        RECT -65.445 93.675 -65.115 94.005 ;
        RECT -65.445 92.315 -65.115 92.645 ;
        RECT -65.445 90.955 -65.115 91.285 ;
        RECT -65.445 89.595 -65.115 89.925 ;
        RECT -65.445 88.235 -65.115 88.565 ;
        RECT -65.445 86.875 -65.115 87.205 ;
        RECT -65.445 85.515 -65.115 85.845 ;
        RECT -65.445 84.155 -65.115 84.485 ;
        RECT -65.445 82.795 -65.115 83.125 ;
        RECT -65.445 81.435 -65.115 81.765 ;
        RECT -65.445 80.075 -65.115 80.405 ;
        RECT -65.445 78.715 -65.115 79.045 ;
        RECT -65.445 77.355 -65.115 77.685 ;
        RECT -65.445 75.995 -65.115 76.325 ;
        RECT -65.445 74.635 -65.115 74.965 ;
        RECT -65.445 73.275 -65.115 73.605 ;
        RECT -65.445 71.915 -65.115 72.245 ;
        RECT -65.445 70.555 -65.115 70.885 ;
        RECT -65.445 69.195 -65.115 69.525 ;
        RECT -65.445 67.835 -65.115 68.165 ;
        RECT -65.445 66.475 -65.115 66.805 ;
        RECT -65.445 65.115 -65.115 65.445 ;
        RECT -65.445 63.755 -65.115 64.085 ;
        RECT -65.445 62.395 -65.115 62.725 ;
        RECT -65.445 61.035 -65.115 61.365 ;
        RECT -65.445 59.675 -65.115 60.005 ;
        RECT -65.445 58.315 -65.115 58.645 ;
        RECT -65.445 56.955 -65.115 57.285 ;
        RECT -65.445 55.595 -65.115 55.925 ;
        RECT -65.445 54.235 -65.115 54.565 ;
        RECT -65.445 52.875 -65.115 53.205 ;
        RECT -65.445 51.515 -65.115 51.845 ;
        RECT -65.445 50.155 -65.115 50.485 ;
        RECT -65.445 48.795 -65.115 49.125 ;
        RECT -65.445 47.435 -65.115 47.765 ;
        RECT -65.445 46.075 -65.115 46.405 ;
        RECT -65.445 44.715 -65.115 45.045 ;
        RECT -65.445 43.355 -65.115 43.685 ;
        RECT -65.445 41.995 -65.115 42.325 ;
        RECT -65.445 40.635 -65.115 40.965 ;
        RECT -65.445 39.275 -65.115 39.605 ;
        RECT -65.445 37.915 -65.115 38.245 ;
        RECT -65.445 36.555 -65.115 36.885 ;
        RECT -65.445 35.195 -65.115 35.525 ;
        RECT -65.445 33.835 -65.115 34.165 ;
        RECT -65.445 32.475 -65.115 32.805 ;
        RECT -65.445 31.115 -65.115 31.445 ;
        RECT -65.445 29.755 -65.115 30.085 ;
        RECT -65.445 28.395 -65.115 28.725 ;
        RECT -65.445 27.035 -65.115 27.365 ;
        RECT -65.445 25.675 -65.115 26.005 ;
        RECT -65.445 24.315 -65.115 24.645 ;
        RECT -65.445 22.955 -65.115 23.285 ;
        RECT -65.445 21.595 -65.115 21.925 ;
        RECT -65.445 20.235 -65.115 20.565 ;
        RECT -65.445 18.875 -65.115 19.205 ;
        RECT -65.445 17.515 -65.115 17.845 ;
        RECT -65.445 16.155 -65.115 16.485 ;
        RECT -65.445 14.795 -65.115 15.125 ;
        RECT -65.445 13.435 -65.115 13.765 ;
        RECT -65.445 12.075 -65.115 12.405 ;
        RECT -65.445 10.715 -65.115 11.045 ;
        RECT -65.445 9.355 -65.115 9.685 ;
        RECT -65.445 7.995 -65.115 8.325 ;
        RECT -65.445 6.635 -65.115 6.965 ;
        RECT -65.445 5.275 -65.115 5.605 ;
        RECT -65.445 3.915 -65.115 4.245 ;
        RECT -65.445 2.555 -65.115 2.885 ;
        RECT -65.445 1.195 -65.115 1.525 ;
        RECT -65.445 -0.165 -65.115 0.165 ;
        RECT -65.445 -1.525 -65.115 -1.195 ;
        RECT -65.445 -2.885 -65.115 -2.555 ;
        RECT -65.445 -4.245 -65.115 -3.915 ;
        RECT -65.445 -5.605 -65.115 -5.275 ;
        RECT -65.445 -6.965 -65.115 -6.635 ;
        RECT -65.445 -8.325 -65.115 -7.995 ;
        RECT -65.445 -9.685 -65.115 -9.355 ;
        RECT -65.445 -11.045 -65.115 -10.715 ;
        RECT -65.445 -12.405 -65.115 -12.075 ;
        RECT -65.445 -13.765 -65.115 -13.435 ;
        RECT -65.445 -15.125 -65.115 -14.795 ;
        RECT -65.445 -16.485 -65.115 -16.155 ;
        RECT -65.445 -17.845 -65.115 -17.515 ;
        RECT -65.445 -19.205 -65.115 -18.875 ;
        RECT -65.445 -20.565 -65.115 -20.235 ;
        RECT -65.445 -21.925 -65.115 -21.595 ;
        RECT -65.445 -23.285 -65.115 -22.955 ;
        RECT -65.445 -24.645 -65.115 -24.315 ;
        RECT -65.445 -26.005 -65.115 -25.675 ;
        RECT -65.445 -27.365 -65.115 -27.035 ;
        RECT -65.445 -28.725 -65.115 -28.395 ;
        RECT -65.445 -30.085 -65.115 -29.755 ;
        RECT -65.445 -31.445 -65.115 -31.115 ;
        RECT -65.445 -32.805 -65.115 -32.475 ;
        RECT -65.445 -34.165 -65.115 -33.835 ;
        RECT -65.445 -35.525 -65.115 -35.195 ;
        RECT -65.445 -36.885 -65.115 -36.555 ;
        RECT -65.445 -38.245 -65.115 -37.915 ;
        RECT -65.445 -39.605 -65.115 -39.275 ;
        RECT -65.445 -40.965 -65.115 -40.635 ;
        RECT -65.445 -42.325 -65.115 -41.995 ;
        RECT -65.445 -43.685 -65.115 -43.355 ;
        RECT -65.445 -45.045 -65.115 -44.715 ;
        RECT -65.445 -46.405 -65.115 -46.075 ;
        RECT -65.445 -47.765 -65.115 -47.435 ;
        RECT -65.445 -49.125 -65.115 -48.795 ;
        RECT -65.445 -50.485 -65.115 -50.155 ;
        RECT -65.445 -51.845 -65.115 -51.515 ;
        RECT -65.445 -53.205 -65.115 -52.875 ;
        RECT -65.445 -54.565 -65.115 -54.235 ;
        RECT -65.445 -55.925 -65.115 -55.595 ;
        RECT -65.445 -57.285 -65.115 -56.955 ;
        RECT -65.445 -58.645 -65.115 -58.315 ;
        RECT -65.445 -60.005 -65.115 -59.675 ;
        RECT -65.445 -61.365 -65.115 -61.035 ;
        RECT -65.445 -62.725 -65.115 -62.395 ;
        RECT -65.445 -64.085 -65.115 -63.755 ;
        RECT -65.445 -65.445 -65.115 -65.115 ;
        RECT -65.445 -66.805 -65.115 -66.475 ;
        RECT -65.445 -68.165 -65.115 -67.835 ;
        RECT -65.445 -69.525 -65.115 -69.195 ;
        RECT -65.445 -70.885 -65.115 -70.555 ;
        RECT -65.445 -72.245 -65.115 -71.915 ;
        RECT -65.445 -73.605 -65.115 -73.275 ;
        RECT -65.445 -74.965 -65.115 -74.635 ;
        RECT -65.445 -76.325 -65.115 -75.995 ;
        RECT -65.445 -77.685 -65.115 -77.355 ;
        RECT -65.445 -79.045 -65.115 -78.715 ;
        RECT -65.445 -80.405 -65.115 -80.075 ;
        RECT -65.445 -81.765 -65.115 -81.435 ;
        RECT -65.445 -83.125 -65.115 -82.795 ;
        RECT -65.445 -84.485 -65.115 -84.155 ;
        RECT -65.445 -85.845 -65.115 -85.515 ;
        RECT -65.445 -87.205 -65.115 -86.875 ;
        RECT -65.445 -88.565 -65.115 -88.235 ;
        RECT -65.445 -89.925 -65.115 -89.595 ;
        RECT -65.445 -91.285 -65.115 -90.955 ;
        RECT -65.445 -92.645 -65.115 -92.315 ;
        RECT -65.445 -94.005 -65.115 -93.675 ;
        RECT -65.445 -95.365 -65.115 -95.035 ;
        RECT -65.445 -96.725 -65.115 -96.395 ;
        RECT -65.445 -98.085 -65.115 -97.755 ;
        RECT -65.445 -99.445 -65.115 -99.115 ;
        RECT -65.445 -100.805 -65.115 -100.475 ;
        RECT -65.445 -102.165 -65.115 -101.835 ;
        RECT -65.445 -103.525 -65.115 -103.195 ;
        RECT -65.445 -104.885 -65.115 -104.555 ;
        RECT -65.445 -106.245 -65.115 -105.915 ;
        RECT -65.445 -107.605 -65.115 -107.275 ;
        RECT -65.445 -108.965 -65.115 -108.635 ;
        RECT -65.445 -110.325 -65.115 -109.995 ;
        RECT -65.445 -111.685 -65.115 -111.355 ;
        RECT -65.445 -113.045 -65.115 -112.715 ;
        RECT -65.445 -114.405 -65.115 -114.075 ;
        RECT -65.445 -115.765 -65.115 -115.435 ;
        RECT -65.445 -117.125 -65.115 -116.795 ;
        RECT -65.445 -118.485 -65.115 -118.155 ;
        RECT -65.445 -119.845 -65.115 -119.515 ;
        RECT -65.445 -121.205 -65.115 -120.875 ;
        RECT -65.445 -122.565 -65.115 -122.235 ;
        RECT -65.445 -123.925 -65.115 -123.595 ;
        RECT -65.445 -125.285 -65.115 -124.955 ;
        RECT -65.445 -126.645 -65.115 -126.315 ;
        RECT -65.445 -129.365 -65.115 -129.035 ;
        RECT -65.445 -130.725 -65.115 -130.395 ;
        RECT -65.445 -131.47 -65.115 -131.14 ;
        RECT -65.445 -133.445 -65.115 -133.115 ;
        RECT -65.445 -134.805 -65.115 -134.475 ;
        RECT -65.445 -136.165 -65.115 -135.835 ;
        RECT -65.445 -137.525 -65.115 -137.195 ;
        RECT -65.445 -140.245 -65.115 -139.915 ;
        RECT -65.445 -141.605 -65.115 -141.275 ;
        RECT -65.445 -142.965 -65.115 -142.635 ;
        RECT -65.445 -144.31 -65.115 -143.98 ;
        RECT -65.445 -145.685 -65.115 -145.355 ;
        RECT -65.445 -147.045 -65.115 -146.715 ;
        RECT -65.445 -149.765 -65.115 -149.435 ;
        RECT -65.445 -152.485 -65.115 -152.155 ;
        RECT -65.445 -153.845 -65.115 -153.515 ;
        RECT -65.445 -155.205 -65.115 -154.875 ;
        RECT -65.445 -156.565 -65.115 -156.235 ;
        RECT -65.445 -157.925 -65.115 -157.595 ;
        RECT -65.445 -159.285 -65.115 -158.955 ;
        RECT -65.445 -162.005 -65.115 -161.675 ;
        RECT -65.445 -163.365 -65.115 -163.035 ;
        RECT -65.445 -164.725 -65.115 -164.395 ;
        RECT -65.445 -166.085 -65.115 -165.755 ;
        RECT -65.445 -167.445 -65.115 -167.115 ;
        RECT -65.445 -168.805 -65.115 -168.475 ;
        RECT -65.445 -170.165 -65.115 -169.835 ;
        RECT -65.445 -171.525 -65.115 -171.195 ;
        RECT -65.445 -172.885 -65.115 -172.555 ;
        RECT -65.445 -174.245 -65.115 -173.915 ;
        RECT -65.445 -175.605 -65.115 -175.275 ;
        RECT -65.445 -176.965 -65.115 -176.635 ;
        RECT -65.445 -178.325 -65.115 -177.995 ;
        RECT -65.445 -179.685 -65.115 -179.355 ;
        RECT -65.445 -181.045 -65.115 -180.715 ;
        RECT -65.445 -182.405 -65.115 -182.075 ;
        RECT -65.445 -183.765 -65.115 -183.435 ;
        RECT -65.445 -185.125 -65.115 -184.795 ;
        RECT -65.445 -186.485 -65.115 -186.155 ;
        RECT -65.445 -187.845 -65.115 -187.515 ;
        RECT -65.445 -189.205 -65.115 -188.875 ;
        RECT -65.445 -190.565 -65.115 -190.235 ;
        RECT -65.445 -191.925 -65.115 -191.595 ;
        RECT -65.445 -193.285 -65.115 -192.955 ;
        RECT -65.445 -194.645 -65.115 -194.315 ;
        RECT -65.445 -196.005 -65.115 -195.675 ;
        RECT -65.445 -197.365 -65.115 -197.035 ;
        RECT -65.445 -198.725 -65.115 -198.395 ;
        RECT -65.445 -200.085 -65.115 -199.755 ;
        RECT -65.445 -201.445 -65.115 -201.115 ;
        RECT -65.445 -202.805 -65.115 -202.475 ;
        RECT -65.445 -204.165 -65.115 -203.835 ;
        RECT -65.445 -205.525 -65.115 -205.195 ;
        RECT -65.445 -206.885 -65.115 -206.555 ;
        RECT -65.445 -208.245 -65.115 -207.915 ;
        RECT -65.445 -209.605 -65.115 -209.275 ;
        RECT -65.445 -210.965 -65.115 -210.635 ;
        RECT -65.445 -212.325 -65.115 -211.995 ;
        RECT -65.445 -213.685 -65.115 -213.355 ;
        RECT -65.445 -215.045 -65.115 -214.715 ;
        RECT -65.445 -216.405 -65.115 -216.075 ;
        RECT -65.445 -217.765 -65.115 -217.435 ;
        RECT -65.445 -219.125 -65.115 -218.795 ;
        RECT -65.445 -220.485 -65.115 -220.155 ;
        RECT -65.445 -221.845 -65.115 -221.515 ;
        RECT -65.445 -223.205 -65.115 -222.875 ;
        RECT -65.445 -224.565 -65.115 -224.235 ;
        RECT -65.445 -226.155 -65.115 -225.825 ;
        RECT -65.445 -227.285 -65.115 -226.955 ;
        RECT -65.445 -228.645 -65.115 -228.315 ;
        RECT -65.44 -229.32 -65.12 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.085 246.76 -63.755 247.89 ;
        RECT -64.085 241.915 -63.755 242.245 ;
        RECT -64.085 240.555 -63.755 240.885 ;
        RECT -64.085 239.195 -63.755 239.525 ;
        RECT -64.085 237.835 -63.755 238.165 ;
        RECT -64.085 236.475 -63.755 236.805 ;
        RECT -64.085 235.115 -63.755 235.445 ;
        RECT -64.085 233.755 -63.755 234.085 ;
        RECT -64.085 232.395 -63.755 232.725 ;
        RECT -64.085 231.035 -63.755 231.365 ;
        RECT -64.085 229.675 -63.755 230.005 ;
        RECT -64.085 228.315 -63.755 228.645 ;
        RECT -64.085 226.955 -63.755 227.285 ;
        RECT -64.085 225.595 -63.755 225.925 ;
        RECT -64.085 224.235 -63.755 224.565 ;
        RECT -64.085 222.875 -63.755 223.205 ;
        RECT -64.085 221.515 -63.755 221.845 ;
        RECT -64.085 220.155 -63.755 220.485 ;
        RECT -64.085 218.795 -63.755 219.125 ;
        RECT -64.085 217.435 -63.755 217.765 ;
        RECT -64.085 216.075 -63.755 216.405 ;
        RECT -64.085 214.715 -63.755 215.045 ;
        RECT -64.085 213.355 -63.755 213.685 ;
        RECT -64.085 211.995 -63.755 212.325 ;
        RECT -64.085 210.635 -63.755 210.965 ;
        RECT -64.085 209.275 -63.755 209.605 ;
        RECT -64.085 207.915 -63.755 208.245 ;
        RECT -64.085 206.555 -63.755 206.885 ;
        RECT -64.085 205.195 -63.755 205.525 ;
        RECT -64.085 203.835 -63.755 204.165 ;
        RECT -64.085 202.475 -63.755 202.805 ;
        RECT -64.085 201.115 -63.755 201.445 ;
        RECT -64.085 199.755 -63.755 200.085 ;
        RECT -64.085 198.395 -63.755 198.725 ;
        RECT -64.085 197.035 -63.755 197.365 ;
        RECT -64.085 195.675 -63.755 196.005 ;
        RECT -64.085 194.315 -63.755 194.645 ;
        RECT -64.085 192.955 -63.755 193.285 ;
        RECT -64.085 191.595 -63.755 191.925 ;
        RECT -64.085 190.235 -63.755 190.565 ;
        RECT -64.085 188.875 -63.755 189.205 ;
        RECT -64.085 187.515 -63.755 187.845 ;
        RECT -64.085 186.155 -63.755 186.485 ;
        RECT -64.085 184.795 -63.755 185.125 ;
        RECT -64.085 183.435 -63.755 183.765 ;
        RECT -64.085 182.075 -63.755 182.405 ;
        RECT -64.085 180.715 -63.755 181.045 ;
        RECT -64.085 179.355 -63.755 179.685 ;
        RECT -64.085 177.995 -63.755 178.325 ;
        RECT -64.085 176.635 -63.755 176.965 ;
        RECT -64.085 175.275 -63.755 175.605 ;
        RECT -64.085 173.915 -63.755 174.245 ;
        RECT -64.085 172.555 -63.755 172.885 ;
        RECT -64.085 171.195 -63.755 171.525 ;
        RECT -64.085 169.835 -63.755 170.165 ;
        RECT -64.085 168.475 -63.755 168.805 ;
        RECT -64.085 167.115 -63.755 167.445 ;
        RECT -64.085 165.755 -63.755 166.085 ;
        RECT -64.085 164.395 -63.755 164.725 ;
        RECT -64.085 163.035 -63.755 163.365 ;
        RECT -64.085 161.675 -63.755 162.005 ;
        RECT -64.085 160.315 -63.755 160.645 ;
        RECT -64.085 158.955 -63.755 159.285 ;
        RECT -64.085 157.595 -63.755 157.925 ;
        RECT -64.085 156.235 -63.755 156.565 ;
        RECT -64.085 154.875 -63.755 155.205 ;
        RECT -64.085 153.515 -63.755 153.845 ;
        RECT -64.085 152.155 -63.755 152.485 ;
        RECT -64.085 150.795 -63.755 151.125 ;
        RECT -64.085 149.435 -63.755 149.765 ;
        RECT -64.085 148.075 -63.755 148.405 ;
        RECT -64.085 146.715 -63.755 147.045 ;
        RECT -64.085 145.355 -63.755 145.685 ;
        RECT -64.085 143.995 -63.755 144.325 ;
        RECT -64.085 142.635 -63.755 142.965 ;
        RECT -64.085 141.275 -63.755 141.605 ;
        RECT -64.085 139.915 -63.755 140.245 ;
        RECT -64.085 138.555 -63.755 138.885 ;
        RECT -64.085 137.195 -63.755 137.525 ;
        RECT -64.085 135.835 -63.755 136.165 ;
        RECT -64.085 134.475 -63.755 134.805 ;
        RECT -64.085 133.115 -63.755 133.445 ;
        RECT -64.085 131.755 -63.755 132.085 ;
        RECT -64.085 130.395 -63.755 130.725 ;
        RECT -64.085 129.035 -63.755 129.365 ;
        RECT -64.085 127.675 -63.755 128.005 ;
        RECT -64.085 126.315 -63.755 126.645 ;
        RECT -64.085 124.955 -63.755 125.285 ;
        RECT -64.085 123.595 -63.755 123.925 ;
        RECT -64.085 122.235 -63.755 122.565 ;
        RECT -64.085 120.875 -63.755 121.205 ;
        RECT -64.085 119.515 -63.755 119.845 ;
        RECT -64.085 118.155 -63.755 118.485 ;
        RECT -64.085 116.795 -63.755 117.125 ;
        RECT -64.085 115.435 -63.755 115.765 ;
        RECT -64.085 114.075 -63.755 114.405 ;
        RECT -64.085 112.715 -63.755 113.045 ;
        RECT -64.085 111.355 -63.755 111.685 ;
        RECT -64.085 109.995 -63.755 110.325 ;
        RECT -64.085 108.635 -63.755 108.965 ;
        RECT -64.085 107.275 -63.755 107.605 ;
        RECT -64.085 105.915 -63.755 106.245 ;
        RECT -64.085 104.555 -63.755 104.885 ;
        RECT -64.085 103.195 -63.755 103.525 ;
        RECT -64.085 101.835 -63.755 102.165 ;
        RECT -64.085 100.475 -63.755 100.805 ;
        RECT -64.085 99.115 -63.755 99.445 ;
        RECT -64.085 97.755 -63.755 98.085 ;
        RECT -64.085 96.395 -63.755 96.725 ;
        RECT -64.085 95.035 -63.755 95.365 ;
        RECT -64.085 93.675 -63.755 94.005 ;
        RECT -64.085 92.315 -63.755 92.645 ;
        RECT -64.085 90.955 -63.755 91.285 ;
        RECT -64.085 89.595 -63.755 89.925 ;
        RECT -64.085 88.235 -63.755 88.565 ;
        RECT -64.085 86.875 -63.755 87.205 ;
        RECT -64.085 85.515 -63.755 85.845 ;
        RECT -64.085 84.155 -63.755 84.485 ;
        RECT -64.085 82.795 -63.755 83.125 ;
        RECT -64.085 81.435 -63.755 81.765 ;
        RECT -64.085 80.075 -63.755 80.405 ;
        RECT -64.085 78.715 -63.755 79.045 ;
        RECT -64.085 77.355 -63.755 77.685 ;
        RECT -64.085 75.995 -63.755 76.325 ;
        RECT -64.085 74.635 -63.755 74.965 ;
        RECT -64.085 73.275 -63.755 73.605 ;
        RECT -64.085 71.915 -63.755 72.245 ;
        RECT -64.085 70.555 -63.755 70.885 ;
        RECT -64.085 69.195 -63.755 69.525 ;
        RECT -64.085 67.835 -63.755 68.165 ;
        RECT -64.085 66.475 -63.755 66.805 ;
        RECT -64.085 65.115 -63.755 65.445 ;
        RECT -64.085 63.755 -63.755 64.085 ;
        RECT -64.085 62.395 -63.755 62.725 ;
        RECT -64.085 61.035 -63.755 61.365 ;
        RECT -64.085 59.675 -63.755 60.005 ;
        RECT -64.085 58.315 -63.755 58.645 ;
        RECT -64.085 56.955 -63.755 57.285 ;
        RECT -64.085 55.595 -63.755 55.925 ;
        RECT -64.085 54.235 -63.755 54.565 ;
        RECT -64.085 52.875 -63.755 53.205 ;
        RECT -64.085 51.515 -63.755 51.845 ;
        RECT -64.085 50.155 -63.755 50.485 ;
        RECT -64.085 48.795 -63.755 49.125 ;
        RECT -64.085 47.435 -63.755 47.765 ;
        RECT -64.085 46.075 -63.755 46.405 ;
        RECT -64.085 44.715 -63.755 45.045 ;
        RECT -64.085 43.355 -63.755 43.685 ;
        RECT -64.085 41.995 -63.755 42.325 ;
        RECT -64.085 40.635 -63.755 40.965 ;
        RECT -64.085 39.275 -63.755 39.605 ;
        RECT -64.085 37.915 -63.755 38.245 ;
        RECT -64.085 36.555 -63.755 36.885 ;
        RECT -64.085 35.195 -63.755 35.525 ;
        RECT -64.085 33.835 -63.755 34.165 ;
        RECT -64.085 32.475 -63.755 32.805 ;
        RECT -64.085 31.115 -63.755 31.445 ;
        RECT -64.085 29.755 -63.755 30.085 ;
        RECT -64.085 28.395 -63.755 28.725 ;
        RECT -64.085 27.035 -63.755 27.365 ;
        RECT -64.085 25.675 -63.755 26.005 ;
        RECT -64.085 24.315 -63.755 24.645 ;
        RECT -64.085 22.955 -63.755 23.285 ;
        RECT -64.085 21.595 -63.755 21.925 ;
        RECT -64.085 20.235 -63.755 20.565 ;
        RECT -64.085 18.875 -63.755 19.205 ;
        RECT -64.085 17.515 -63.755 17.845 ;
        RECT -64.085 16.155 -63.755 16.485 ;
        RECT -64.085 14.795 -63.755 15.125 ;
        RECT -64.085 13.435 -63.755 13.765 ;
        RECT -64.085 12.075 -63.755 12.405 ;
        RECT -64.085 10.715 -63.755 11.045 ;
        RECT -64.085 9.355 -63.755 9.685 ;
        RECT -64.085 7.995 -63.755 8.325 ;
        RECT -64.085 6.635 -63.755 6.965 ;
        RECT -64.085 5.275 -63.755 5.605 ;
        RECT -64.085 3.915 -63.755 4.245 ;
        RECT -64.085 2.555 -63.755 2.885 ;
        RECT -64.085 1.195 -63.755 1.525 ;
        RECT -64.085 -0.165 -63.755 0.165 ;
        RECT -64.085 -1.525 -63.755 -1.195 ;
        RECT -64.085 -2.885 -63.755 -2.555 ;
        RECT -64.085 -4.245 -63.755 -3.915 ;
        RECT -64.085 -5.605 -63.755 -5.275 ;
        RECT -64.085 -6.965 -63.755 -6.635 ;
        RECT -64.085 -8.325 -63.755 -7.995 ;
        RECT -64.085 -9.685 -63.755 -9.355 ;
        RECT -64.085 -11.045 -63.755 -10.715 ;
        RECT -64.085 -12.405 -63.755 -12.075 ;
        RECT -64.085 -13.765 -63.755 -13.435 ;
        RECT -64.085 -15.125 -63.755 -14.795 ;
        RECT -64.085 -16.485 -63.755 -16.155 ;
        RECT -64.085 -17.845 -63.755 -17.515 ;
        RECT -64.085 -19.205 -63.755 -18.875 ;
        RECT -64.085 -20.565 -63.755 -20.235 ;
        RECT -64.085 -21.925 -63.755 -21.595 ;
        RECT -64.085 -23.285 -63.755 -22.955 ;
        RECT -64.085 -24.645 -63.755 -24.315 ;
        RECT -64.085 -26.005 -63.755 -25.675 ;
        RECT -64.085 -27.365 -63.755 -27.035 ;
        RECT -64.085 -28.725 -63.755 -28.395 ;
        RECT -64.085 -30.085 -63.755 -29.755 ;
        RECT -64.085 -31.445 -63.755 -31.115 ;
        RECT -64.085 -32.805 -63.755 -32.475 ;
        RECT -64.085 -34.165 -63.755 -33.835 ;
        RECT -64.085 -35.525 -63.755 -35.195 ;
        RECT -64.085 -36.885 -63.755 -36.555 ;
        RECT -64.085 -38.245 -63.755 -37.915 ;
        RECT -64.085 -39.605 -63.755 -39.275 ;
        RECT -64.085 -40.965 -63.755 -40.635 ;
        RECT -64.085 -42.325 -63.755 -41.995 ;
        RECT -64.085 -43.685 -63.755 -43.355 ;
        RECT -64.085 -45.045 -63.755 -44.715 ;
        RECT -64.085 -46.405 -63.755 -46.075 ;
        RECT -64.085 -47.765 -63.755 -47.435 ;
        RECT -64.085 -49.125 -63.755 -48.795 ;
        RECT -64.085 -50.485 -63.755 -50.155 ;
        RECT -64.085 -51.845 -63.755 -51.515 ;
        RECT -64.085 -53.205 -63.755 -52.875 ;
        RECT -64.085 -54.565 -63.755 -54.235 ;
        RECT -64.085 -55.925 -63.755 -55.595 ;
        RECT -64.085 -57.285 -63.755 -56.955 ;
        RECT -64.085 -58.645 -63.755 -58.315 ;
        RECT -64.085 -60.005 -63.755 -59.675 ;
        RECT -64.085 -61.365 -63.755 -61.035 ;
        RECT -64.085 -62.725 -63.755 -62.395 ;
        RECT -64.085 -64.085 -63.755 -63.755 ;
        RECT -64.085 -65.445 -63.755 -65.115 ;
        RECT -64.085 -66.805 -63.755 -66.475 ;
        RECT -64.085 -68.165 -63.755 -67.835 ;
        RECT -64.085 -69.525 -63.755 -69.195 ;
        RECT -64.085 -70.885 -63.755 -70.555 ;
        RECT -64.085 -72.245 -63.755 -71.915 ;
        RECT -64.085 -73.605 -63.755 -73.275 ;
        RECT -64.085 -74.965 -63.755 -74.635 ;
        RECT -64.085 -76.325 -63.755 -75.995 ;
        RECT -64.085 -77.685 -63.755 -77.355 ;
        RECT -64.085 -79.045 -63.755 -78.715 ;
        RECT -64.085 -80.405 -63.755 -80.075 ;
        RECT -64.085 -81.765 -63.755 -81.435 ;
        RECT -64.085 -83.125 -63.755 -82.795 ;
        RECT -64.085 -84.485 -63.755 -84.155 ;
        RECT -64.085 -85.845 -63.755 -85.515 ;
        RECT -64.085 -87.205 -63.755 -86.875 ;
        RECT -64.085 -88.565 -63.755 -88.235 ;
        RECT -64.085 -89.925 -63.755 -89.595 ;
        RECT -64.085 -91.285 -63.755 -90.955 ;
        RECT -64.085 -92.645 -63.755 -92.315 ;
        RECT -64.085 -94.005 -63.755 -93.675 ;
        RECT -64.085 -95.365 -63.755 -95.035 ;
        RECT -64.085 -96.725 -63.755 -96.395 ;
        RECT -64.085 -98.085 -63.755 -97.755 ;
        RECT -64.085 -99.445 -63.755 -99.115 ;
        RECT -64.085 -100.805 -63.755 -100.475 ;
        RECT -64.085 -102.165 -63.755 -101.835 ;
        RECT -64.085 -103.525 -63.755 -103.195 ;
        RECT -64.085 -104.885 -63.755 -104.555 ;
        RECT -64.085 -106.245 -63.755 -105.915 ;
        RECT -64.085 -107.605 -63.755 -107.275 ;
        RECT -64.085 -108.965 -63.755 -108.635 ;
        RECT -64.085 -110.325 -63.755 -109.995 ;
        RECT -64.085 -111.685 -63.755 -111.355 ;
        RECT -64.085 -113.045 -63.755 -112.715 ;
        RECT -64.085 -114.405 -63.755 -114.075 ;
        RECT -64.085 -115.765 -63.755 -115.435 ;
        RECT -64.085 -117.125 -63.755 -116.795 ;
        RECT -64.085 -118.485 -63.755 -118.155 ;
        RECT -64.085 -119.845 -63.755 -119.515 ;
        RECT -64.085 -121.205 -63.755 -120.875 ;
        RECT -64.085 -122.565 -63.755 -122.235 ;
        RECT -64.085 -123.925 -63.755 -123.595 ;
        RECT -64.085 -125.285 -63.755 -124.955 ;
        RECT -64.085 -129.365 -63.755 -129.035 ;
        RECT -64.085 -130.725 -63.755 -130.395 ;
        RECT -64.085 -131.47 -63.755 -131.14 ;
        RECT -64.085 -133.445 -63.755 -133.115 ;
        RECT -64.085 -134.805 -63.755 -134.475 ;
        RECT -64.085 -136.165 -63.755 -135.835 ;
        RECT -64.085 -137.525 -63.755 -137.195 ;
        RECT -64.085 -140.245 -63.755 -139.915 ;
        RECT -64.085 -141.605 -63.755 -141.275 ;
        RECT -64.085 -142.965 -63.755 -142.635 ;
        RECT -64.085 -144.31 -63.755 -143.98 ;
        RECT -64.085 -145.685 -63.755 -145.355 ;
        RECT -64.085 -147.045 -63.755 -146.715 ;
        RECT -64.085 -149.765 -63.755 -149.435 ;
        RECT -64.085 -152.485 -63.755 -152.155 ;
        RECT -64.085 -153.845 -63.755 -153.515 ;
        RECT -64.085 -155.205 -63.755 -154.875 ;
        RECT -64.085 -156.565 -63.755 -156.235 ;
        RECT -64.085 -157.925 -63.755 -157.595 ;
        RECT -64.085 -159.285 -63.755 -158.955 ;
        RECT -64.085 -162.005 -63.755 -161.675 ;
        RECT -64.085 -163.365 -63.755 -163.035 ;
        RECT -64.085 -164.725 -63.755 -164.395 ;
        RECT -64.085 -166.085 -63.755 -165.755 ;
        RECT -64.085 -167.445 -63.755 -167.115 ;
        RECT -64.085 -168.805 -63.755 -168.475 ;
        RECT -64.085 -170.165 -63.755 -169.835 ;
        RECT -64.085 -171.525 -63.755 -171.195 ;
        RECT -64.085 -172.885 -63.755 -172.555 ;
        RECT -64.085 -174.245 -63.755 -173.915 ;
        RECT -64.085 -175.605 -63.755 -175.275 ;
        RECT -64.085 -176.965 -63.755 -176.635 ;
        RECT -64.085 -178.325 -63.755 -177.995 ;
        RECT -64.085 -179.685 -63.755 -179.355 ;
        RECT -64.085 -181.045 -63.755 -180.715 ;
        RECT -64.085 -182.405 -63.755 -182.075 ;
        RECT -64.085 -183.765 -63.755 -183.435 ;
        RECT -64.085 -185.125 -63.755 -184.795 ;
        RECT -64.085 -186.485 -63.755 -186.155 ;
        RECT -64.085 -187.845 -63.755 -187.515 ;
        RECT -64.085 -189.205 -63.755 -188.875 ;
        RECT -64.085 -190.565 -63.755 -190.235 ;
        RECT -64.085 -191.925 -63.755 -191.595 ;
        RECT -64.085 -193.285 -63.755 -192.955 ;
        RECT -64.085 -194.645 -63.755 -194.315 ;
        RECT -64.085 -196.005 -63.755 -195.675 ;
        RECT -64.085 -197.365 -63.755 -197.035 ;
        RECT -64.085 -198.725 -63.755 -198.395 ;
        RECT -64.085 -200.085 -63.755 -199.755 ;
        RECT -64.085 -201.445 -63.755 -201.115 ;
        RECT -64.085 -202.805 -63.755 -202.475 ;
        RECT -64.085 -204.165 -63.755 -203.835 ;
        RECT -64.085 -205.525 -63.755 -205.195 ;
        RECT -64.085 -206.885 -63.755 -206.555 ;
        RECT -64.085 -208.245 -63.755 -207.915 ;
        RECT -64.085 -209.605 -63.755 -209.275 ;
        RECT -64.085 -210.965 -63.755 -210.635 ;
        RECT -64.085 -212.325 -63.755 -211.995 ;
        RECT -64.085 -213.685 -63.755 -213.355 ;
        RECT -64.085 -215.045 -63.755 -214.715 ;
        RECT -64.085 -216.405 -63.755 -216.075 ;
        RECT -64.085 -217.765 -63.755 -217.435 ;
        RECT -64.085 -219.125 -63.755 -218.795 ;
        RECT -64.085 -220.485 -63.755 -220.155 ;
        RECT -64.085 -221.845 -63.755 -221.515 ;
        RECT -64.085 -223.205 -63.755 -222.875 ;
        RECT -64.085 -224.565 -63.755 -224.235 ;
        RECT -64.085 -226.155 -63.755 -225.825 ;
        RECT -64.085 -227.285 -63.755 -226.955 ;
        RECT -64.085 -228.645 -63.755 -228.315 ;
        RECT -64.085 -234.085 -63.755 -233.755 ;
        RECT -64.085 -235.445 -63.755 -235.115 ;
        RECT -64.085 -236.805 -63.755 -236.475 ;
        RECT -64.085 -238.165 -63.755 -237.835 ;
        RECT -64.085 -243.81 -63.755 -242.68 ;
        RECT -64.08 -243.925 -63.76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.725 -196.005 -62.395 -195.675 ;
        RECT -62.725 -197.365 -62.395 -197.035 ;
        RECT -62.725 -198.725 -62.395 -198.395 ;
        RECT -62.725 -200.085 -62.395 -199.755 ;
        RECT -62.725 -201.445 -62.395 -201.115 ;
        RECT -62.725 -202.805 -62.395 -202.475 ;
        RECT -62.725 -204.165 -62.395 -203.835 ;
        RECT -62.725 -205.525 -62.395 -205.195 ;
        RECT -62.725 -206.885 -62.395 -206.555 ;
        RECT -62.725 -208.245 -62.395 -207.915 ;
        RECT -62.725 -209.605 -62.395 -209.275 ;
        RECT -62.725 -210.965 -62.395 -210.635 ;
        RECT -62.725 -212.325 -62.395 -211.995 ;
        RECT -62.725 -213.685 -62.395 -213.355 ;
        RECT -62.725 -215.045 -62.395 -214.715 ;
        RECT -62.725 -216.405 -62.395 -216.075 ;
        RECT -62.725 -217.765 -62.395 -217.435 ;
        RECT -62.725 -219.125 -62.395 -218.795 ;
        RECT -62.725 -220.485 -62.395 -220.155 ;
        RECT -62.725 -221.845 -62.395 -221.515 ;
        RECT -62.725 -223.205 -62.395 -222.875 ;
        RECT -62.725 -224.565 -62.395 -224.235 ;
        RECT -62.725 -226.155 -62.395 -225.825 ;
        RECT -62.725 -227.285 -62.395 -226.955 ;
        RECT -62.725 -228.645 -62.395 -228.315 ;
        RECT -62.725 -230.005 -62.395 -229.675 ;
        RECT -62.725 -231.365 -62.395 -231.035 ;
        RECT -62.725 -234.085 -62.395 -233.755 ;
        RECT -62.725 -235.445 -62.395 -235.115 ;
        RECT -62.725 -236.805 -62.395 -236.475 ;
        RECT -62.725 -238.165 -62.395 -237.835 ;
        RECT -62.725 -243.81 -62.395 -242.68 ;
        RECT -62.72 -243.925 -62.4 248.005 ;
        RECT -62.725 246.76 -62.395 247.89 ;
        RECT -62.725 241.915 -62.395 242.245 ;
        RECT -62.725 240.555 -62.395 240.885 ;
        RECT -62.725 239.195 -62.395 239.525 ;
        RECT -62.725 237.835 -62.395 238.165 ;
        RECT -62.725 236.475 -62.395 236.805 ;
        RECT -62.725 235.115 -62.395 235.445 ;
        RECT -62.725 233.755 -62.395 234.085 ;
        RECT -62.725 232.395 -62.395 232.725 ;
        RECT -62.725 231.035 -62.395 231.365 ;
        RECT -62.725 229.675 -62.395 230.005 ;
        RECT -62.725 228.315 -62.395 228.645 ;
        RECT -62.725 226.955 -62.395 227.285 ;
        RECT -62.725 225.595 -62.395 225.925 ;
        RECT -62.725 224.235 -62.395 224.565 ;
        RECT -62.725 222.875 -62.395 223.205 ;
        RECT -62.725 221.515 -62.395 221.845 ;
        RECT -62.725 220.155 -62.395 220.485 ;
        RECT -62.725 218.795 -62.395 219.125 ;
        RECT -62.725 217.435 -62.395 217.765 ;
        RECT -62.725 216.075 -62.395 216.405 ;
        RECT -62.725 214.715 -62.395 215.045 ;
        RECT -62.725 213.355 -62.395 213.685 ;
        RECT -62.725 211.995 -62.395 212.325 ;
        RECT -62.725 210.635 -62.395 210.965 ;
        RECT -62.725 209.275 -62.395 209.605 ;
        RECT -62.725 207.915 -62.395 208.245 ;
        RECT -62.725 206.555 -62.395 206.885 ;
        RECT -62.725 205.195 -62.395 205.525 ;
        RECT -62.725 203.835 -62.395 204.165 ;
        RECT -62.725 202.475 -62.395 202.805 ;
        RECT -62.725 201.115 -62.395 201.445 ;
        RECT -62.725 199.755 -62.395 200.085 ;
        RECT -62.725 198.395 -62.395 198.725 ;
        RECT -62.725 197.035 -62.395 197.365 ;
        RECT -62.725 195.675 -62.395 196.005 ;
        RECT -62.725 194.315 -62.395 194.645 ;
        RECT -62.725 192.955 -62.395 193.285 ;
        RECT -62.725 191.595 -62.395 191.925 ;
        RECT -62.725 190.235 -62.395 190.565 ;
        RECT -62.725 188.875 -62.395 189.205 ;
        RECT -62.725 187.515 -62.395 187.845 ;
        RECT -62.725 186.155 -62.395 186.485 ;
        RECT -62.725 184.795 -62.395 185.125 ;
        RECT -62.725 183.435 -62.395 183.765 ;
        RECT -62.725 182.075 -62.395 182.405 ;
        RECT -62.725 180.715 -62.395 181.045 ;
        RECT -62.725 179.355 -62.395 179.685 ;
        RECT -62.725 177.995 -62.395 178.325 ;
        RECT -62.725 176.635 -62.395 176.965 ;
        RECT -62.725 175.275 -62.395 175.605 ;
        RECT -62.725 173.915 -62.395 174.245 ;
        RECT -62.725 172.555 -62.395 172.885 ;
        RECT -62.725 171.195 -62.395 171.525 ;
        RECT -62.725 169.835 -62.395 170.165 ;
        RECT -62.725 168.475 -62.395 168.805 ;
        RECT -62.725 167.115 -62.395 167.445 ;
        RECT -62.725 165.755 -62.395 166.085 ;
        RECT -62.725 164.395 -62.395 164.725 ;
        RECT -62.725 163.035 -62.395 163.365 ;
        RECT -62.725 161.675 -62.395 162.005 ;
        RECT -62.725 160.315 -62.395 160.645 ;
        RECT -62.725 158.955 -62.395 159.285 ;
        RECT -62.725 157.595 -62.395 157.925 ;
        RECT -62.725 156.235 -62.395 156.565 ;
        RECT -62.725 154.875 -62.395 155.205 ;
        RECT -62.725 153.515 -62.395 153.845 ;
        RECT -62.725 152.155 -62.395 152.485 ;
        RECT -62.725 150.795 -62.395 151.125 ;
        RECT -62.725 149.435 -62.395 149.765 ;
        RECT -62.725 148.075 -62.395 148.405 ;
        RECT -62.725 146.715 -62.395 147.045 ;
        RECT -62.725 145.355 -62.395 145.685 ;
        RECT -62.725 143.995 -62.395 144.325 ;
        RECT -62.725 142.635 -62.395 142.965 ;
        RECT -62.725 141.275 -62.395 141.605 ;
        RECT -62.725 139.915 -62.395 140.245 ;
        RECT -62.725 138.555 -62.395 138.885 ;
        RECT -62.725 137.195 -62.395 137.525 ;
        RECT -62.725 135.835 -62.395 136.165 ;
        RECT -62.725 134.475 -62.395 134.805 ;
        RECT -62.725 133.115 -62.395 133.445 ;
        RECT -62.725 131.755 -62.395 132.085 ;
        RECT -62.725 130.395 -62.395 130.725 ;
        RECT -62.725 129.035 -62.395 129.365 ;
        RECT -62.725 127.675 -62.395 128.005 ;
        RECT -62.725 126.315 -62.395 126.645 ;
        RECT -62.725 124.955 -62.395 125.285 ;
        RECT -62.725 123.595 -62.395 123.925 ;
        RECT -62.725 122.235 -62.395 122.565 ;
        RECT -62.725 120.875 -62.395 121.205 ;
        RECT -62.725 119.515 -62.395 119.845 ;
        RECT -62.725 118.155 -62.395 118.485 ;
        RECT -62.725 116.795 -62.395 117.125 ;
        RECT -62.725 115.435 -62.395 115.765 ;
        RECT -62.725 114.075 -62.395 114.405 ;
        RECT -62.725 112.715 -62.395 113.045 ;
        RECT -62.725 111.355 -62.395 111.685 ;
        RECT -62.725 109.995 -62.395 110.325 ;
        RECT -62.725 108.635 -62.395 108.965 ;
        RECT -62.725 107.275 -62.395 107.605 ;
        RECT -62.725 105.915 -62.395 106.245 ;
        RECT -62.725 104.555 -62.395 104.885 ;
        RECT -62.725 103.195 -62.395 103.525 ;
        RECT -62.725 101.835 -62.395 102.165 ;
        RECT -62.725 100.475 -62.395 100.805 ;
        RECT -62.725 99.115 -62.395 99.445 ;
        RECT -62.725 97.755 -62.395 98.085 ;
        RECT -62.725 96.395 -62.395 96.725 ;
        RECT -62.725 95.035 -62.395 95.365 ;
        RECT -62.725 93.675 -62.395 94.005 ;
        RECT -62.725 92.315 -62.395 92.645 ;
        RECT -62.725 90.955 -62.395 91.285 ;
        RECT -62.725 89.595 -62.395 89.925 ;
        RECT -62.725 88.235 -62.395 88.565 ;
        RECT -62.725 86.875 -62.395 87.205 ;
        RECT -62.725 85.515 -62.395 85.845 ;
        RECT -62.725 84.155 -62.395 84.485 ;
        RECT -62.725 82.795 -62.395 83.125 ;
        RECT -62.725 81.435 -62.395 81.765 ;
        RECT -62.725 80.075 -62.395 80.405 ;
        RECT -62.725 78.715 -62.395 79.045 ;
        RECT -62.725 77.355 -62.395 77.685 ;
        RECT -62.725 75.995 -62.395 76.325 ;
        RECT -62.725 74.635 -62.395 74.965 ;
        RECT -62.725 73.275 -62.395 73.605 ;
        RECT -62.725 71.915 -62.395 72.245 ;
        RECT -62.725 70.555 -62.395 70.885 ;
        RECT -62.725 69.195 -62.395 69.525 ;
        RECT -62.725 67.835 -62.395 68.165 ;
        RECT -62.725 66.475 -62.395 66.805 ;
        RECT -62.725 65.115 -62.395 65.445 ;
        RECT -62.725 63.755 -62.395 64.085 ;
        RECT -62.725 62.395 -62.395 62.725 ;
        RECT -62.725 61.035 -62.395 61.365 ;
        RECT -62.725 59.675 -62.395 60.005 ;
        RECT -62.725 58.315 -62.395 58.645 ;
        RECT -62.725 56.955 -62.395 57.285 ;
        RECT -62.725 55.595 -62.395 55.925 ;
        RECT -62.725 54.235 -62.395 54.565 ;
        RECT -62.725 52.875 -62.395 53.205 ;
        RECT -62.725 51.515 -62.395 51.845 ;
        RECT -62.725 50.155 -62.395 50.485 ;
        RECT -62.725 48.795 -62.395 49.125 ;
        RECT -62.725 47.435 -62.395 47.765 ;
        RECT -62.725 46.075 -62.395 46.405 ;
        RECT -62.725 44.715 -62.395 45.045 ;
        RECT -62.725 43.355 -62.395 43.685 ;
        RECT -62.725 41.995 -62.395 42.325 ;
        RECT -62.725 40.635 -62.395 40.965 ;
        RECT -62.725 39.275 -62.395 39.605 ;
        RECT -62.725 37.915 -62.395 38.245 ;
        RECT -62.725 36.555 -62.395 36.885 ;
        RECT -62.725 35.195 -62.395 35.525 ;
        RECT -62.725 33.835 -62.395 34.165 ;
        RECT -62.725 32.475 -62.395 32.805 ;
        RECT -62.725 31.115 -62.395 31.445 ;
        RECT -62.725 29.755 -62.395 30.085 ;
        RECT -62.725 28.395 -62.395 28.725 ;
        RECT -62.725 27.035 -62.395 27.365 ;
        RECT -62.725 25.675 -62.395 26.005 ;
        RECT -62.725 24.315 -62.395 24.645 ;
        RECT -62.725 22.955 -62.395 23.285 ;
        RECT -62.725 21.595 -62.395 21.925 ;
        RECT -62.725 20.235 -62.395 20.565 ;
        RECT -62.725 18.875 -62.395 19.205 ;
        RECT -62.725 17.515 -62.395 17.845 ;
        RECT -62.725 16.155 -62.395 16.485 ;
        RECT -62.725 14.795 -62.395 15.125 ;
        RECT -62.725 13.435 -62.395 13.765 ;
        RECT -62.725 12.075 -62.395 12.405 ;
        RECT -62.725 10.715 -62.395 11.045 ;
        RECT -62.725 9.355 -62.395 9.685 ;
        RECT -62.725 7.995 -62.395 8.325 ;
        RECT -62.725 6.635 -62.395 6.965 ;
        RECT -62.725 5.275 -62.395 5.605 ;
        RECT -62.725 3.915 -62.395 4.245 ;
        RECT -62.725 2.555 -62.395 2.885 ;
        RECT -62.725 1.195 -62.395 1.525 ;
        RECT -62.725 -0.165 -62.395 0.165 ;
        RECT -62.725 -1.525 -62.395 -1.195 ;
        RECT -62.725 -2.885 -62.395 -2.555 ;
        RECT -62.725 -4.245 -62.395 -3.915 ;
        RECT -62.725 -5.605 -62.395 -5.275 ;
        RECT -62.725 -6.965 -62.395 -6.635 ;
        RECT -62.725 -8.325 -62.395 -7.995 ;
        RECT -62.725 -9.685 -62.395 -9.355 ;
        RECT -62.725 -11.045 -62.395 -10.715 ;
        RECT -62.725 -12.405 -62.395 -12.075 ;
        RECT -62.725 -13.765 -62.395 -13.435 ;
        RECT -62.725 -15.125 -62.395 -14.795 ;
        RECT -62.725 -16.485 -62.395 -16.155 ;
        RECT -62.725 -17.845 -62.395 -17.515 ;
        RECT -62.725 -19.205 -62.395 -18.875 ;
        RECT -62.725 -20.565 -62.395 -20.235 ;
        RECT -62.725 -21.925 -62.395 -21.595 ;
        RECT -62.725 -23.285 -62.395 -22.955 ;
        RECT -62.725 -24.645 -62.395 -24.315 ;
        RECT -62.725 -26.005 -62.395 -25.675 ;
        RECT -62.725 -27.365 -62.395 -27.035 ;
        RECT -62.725 -28.725 -62.395 -28.395 ;
        RECT -62.725 -30.085 -62.395 -29.755 ;
        RECT -62.725 -31.445 -62.395 -31.115 ;
        RECT -62.725 -32.805 -62.395 -32.475 ;
        RECT -62.725 -34.165 -62.395 -33.835 ;
        RECT -62.725 -35.525 -62.395 -35.195 ;
        RECT -62.725 -36.885 -62.395 -36.555 ;
        RECT -62.725 -38.245 -62.395 -37.915 ;
        RECT -62.725 -39.605 -62.395 -39.275 ;
        RECT -62.725 -40.965 -62.395 -40.635 ;
        RECT -62.725 -42.325 -62.395 -41.995 ;
        RECT -62.725 -43.685 -62.395 -43.355 ;
        RECT -62.725 -45.045 -62.395 -44.715 ;
        RECT -62.725 -46.405 -62.395 -46.075 ;
        RECT -62.725 -47.765 -62.395 -47.435 ;
        RECT -62.725 -49.125 -62.395 -48.795 ;
        RECT -62.725 -50.485 -62.395 -50.155 ;
        RECT -62.725 -51.845 -62.395 -51.515 ;
        RECT -62.725 -53.205 -62.395 -52.875 ;
        RECT -62.725 -54.565 -62.395 -54.235 ;
        RECT -62.725 -55.925 -62.395 -55.595 ;
        RECT -62.725 -57.285 -62.395 -56.955 ;
        RECT -62.725 -58.645 -62.395 -58.315 ;
        RECT -62.725 -60.005 -62.395 -59.675 ;
        RECT -62.725 -61.365 -62.395 -61.035 ;
        RECT -62.725 -62.725 -62.395 -62.395 ;
        RECT -62.725 -64.085 -62.395 -63.755 ;
        RECT -62.725 -65.445 -62.395 -65.115 ;
        RECT -62.725 -66.805 -62.395 -66.475 ;
        RECT -62.725 -68.165 -62.395 -67.835 ;
        RECT -62.725 -69.525 -62.395 -69.195 ;
        RECT -62.725 -70.885 -62.395 -70.555 ;
        RECT -62.725 -72.245 -62.395 -71.915 ;
        RECT -62.725 -73.605 -62.395 -73.275 ;
        RECT -62.725 -74.965 -62.395 -74.635 ;
        RECT -62.725 -76.325 -62.395 -75.995 ;
        RECT -62.725 -77.685 -62.395 -77.355 ;
        RECT -62.725 -79.045 -62.395 -78.715 ;
        RECT -62.725 -80.405 -62.395 -80.075 ;
        RECT -62.725 -81.765 -62.395 -81.435 ;
        RECT -62.725 -83.125 -62.395 -82.795 ;
        RECT -62.725 -84.485 -62.395 -84.155 ;
        RECT -62.725 -85.845 -62.395 -85.515 ;
        RECT -62.725 -87.205 -62.395 -86.875 ;
        RECT -62.725 -88.565 -62.395 -88.235 ;
        RECT -62.725 -89.925 -62.395 -89.595 ;
        RECT -62.725 -91.285 -62.395 -90.955 ;
        RECT -62.725 -92.645 -62.395 -92.315 ;
        RECT -62.725 -94.005 -62.395 -93.675 ;
        RECT -62.725 -95.365 -62.395 -95.035 ;
        RECT -62.725 -96.725 -62.395 -96.395 ;
        RECT -62.725 -98.085 -62.395 -97.755 ;
        RECT -62.725 -99.445 -62.395 -99.115 ;
        RECT -62.725 -100.805 -62.395 -100.475 ;
        RECT -62.725 -102.165 -62.395 -101.835 ;
        RECT -62.725 -103.525 -62.395 -103.195 ;
        RECT -62.725 -104.885 -62.395 -104.555 ;
        RECT -62.725 -106.245 -62.395 -105.915 ;
        RECT -62.725 -107.605 -62.395 -107.275 ;
        RECT -62.725 -108.965 -62.395 -108.635 ;
        RECT -62.725 -110.325 -62.395 -109.995 ;
        RECT -62.725 -111.685 -62.395 -111.355 ;
        RECT -62.725 -113.045 -62.395 -112.715 ;
        RECT -62.725 -114.405 -62.395 -114.075 ;
        RECT -62.725 -115.765 -62.395 -115.435 ;
        RECT -62.725 -117.125 -62.395 -116.795 ;
        RECT -62.725 -118.485 -62.395 -118.155 ;
        RECT -62.725 -119.845 -62.395 -119.515 ;
        RECT -62.725 -121.205 -62.395 -120.875 ;
        RECT -62.725 -122.565 -62.395 -122.235 ;
        RECT -62.725 -123.925 -62.395 -123.595 ;
        RECT -62.725 -125.285 -62.395 -124.955 ;
        RECT -62.725 -129.365 -62.395 -129.035 ;
        RECT -62.725 -130.725 -62.395 -130.395 ;
        RECT -62.725 -131.47 -62.395 -131.14 ;
        RECT -62.725 -133.445 -62.395 -133.115 ;
        RECT -62.725 -134.805 -62.395 -134.475 ;
        RECT -62.725 -136.165 -62.395 -135.835 ;
        RECT -62.725 -137.525 -62.395 -137.195 ;
        RECT -62.725 -140.245 -62.395 -139.915 ;
        RECT -62.725 -141.605 -62.395 -141.275 ;
        RECT -62.725 -142.965 -62.395 -142.635 ;
        RECT -62.725 -144.31 -62.395 -143.98 ;
        RECT -62.725 -145.685 -62.395 -145.355 ;
        RECT -62.725 -147.045 -62.395 -146.715 ;
        RECT -62.725 -149.765 -62.395 -149.435 ;
        RECT -62.725 -152.485 -62.395 -152.155 ;
        RECT -62.725 -153.845 -62.395 -153.515 ;
        RECT -62.725 -155.205 -62.395 -154.875 ;
        RECT -62.725 -156.565 -62.395 -156.235 ;
        RECT -62.725 -157.925 -62.395 -157.595 ;
        RECT -62.725 -159.285 -62.395 -158.955 ;
        RECT -62.725 -162.005 -62.395 -161.675 ;
        RECT -62.725 -163.365 -62.395 -163.035 ;
        RECT -62.725 -164.725 -62.395 -164.395 ;
        RECT -62.725 -166.085 -62.395 -165.755 ;
        RECT -62.725 -167.445 -62.395 -167.115 ;
        RECT -62.725 -168.805 -62.395 -168.475 ;
        RECT -62.725 -170.165 -62.395 -169.835 ;
        RECT -62.725 -171.525 -62.395 -171.195 ;
        RECT -62.725 -172.885 -62.395 -172.555 ;
        RECT -62.725 -174.245 -62.395 -173.915 ;
        RECT -62.725 -175.605 -62.395 -175.275 ;
        RECT -62.725 -176.965 -62.395 -176.635 ;
        RECT -62.725 -178.325 -62.395 -177.995 ;
        RECT -62.725 -179.685 -62.395 -179.355 ;
        RECT -62.725 -181.045 -62.395 -180.715 ;
        RECT -62.725 -182.405 -62.395 -182.075 ;
        RECT -62.725 -183.765 -62.395 -183.435 ;
        RECT -62.725 -185.125 -62.395 -184.795 ;
        RECT -62.725 -186.485 -62.395 -186.155 ;
        RECT -62.725 -187.845 -62.395 -187.515 ;
        RECT -62.725 -189.205 -62.395 -188.875 ;
        RECT -62.725 -190.565 -62.395 -190.235 ;
        RECT -62.725 -191.925 -62.395 -191.595 ;
        RECT -62.725 -193.285 -62.395 -192.955 ;
        RECT -62.725 -194.645 -62.395 -194.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.525 246.76 -69.195 247.89 ;
        RECT -69.525 241.915 -69.195 242.245 ;
        RECT -69.525 240.555 -69.195 240.885 ;
        RECT -69.525 239.195 -69.195 239.525 ;
        RECT -69.525 237.835 -69.195 238.165 ;
        RECT -69.525 236.475 -69.195 236.805 ;
        RECT -69.525 235.115 -69.195 235.445 ;
        RECT -69.525 233.755 -69.195 234.085 ;
        RECT -69.525 232.395 -69.195 232.725 ;
        RECT -69.525 231.035 -69.195 231.365 ;
        RECT -69.525 229.675 -69.195 230.005 ;
        RECT -69.525 228.315 -69.195 228.645 ;
        RECT -69.525 226.955 -69.195 227.285 ;
        RECT -69.525 225.595 -69.195 225.925 ;
        RECT -69.525 224.235 -69.195 224.565 ;
        RECT -69.525 222.875 -69.195 223.205 ;
        RECT -69.525 221.515 -69.195 221.845 ;
        RECT -69.525 220.155 -69.195 220.485 ;
        RECT -69.525 218.795 -69.195 219.125 ;
        RECT -69.525 217.435 -69.195 217.765 ;
        RECT -69.525 216.075 -69.195 216.405 ;
        RECT -69.525 214.715 -69.195 215.045 ;
        RECT -69.525 213.355 -69.195 213.685 ;
        RECT -69.525 211.995 -69.195 212.325 ;
        RECT -69.525 210.635 -69.195 210.965 ;
        RECT -69.525 209.275 -69.195 209.605 ;
        RECT -69.525 207.915 -69.195 208.245 ;
        RECT -69.525 206.555 -69.195 206.885 ;
        RECT -69.525 205.195 -69.195 205.525 ;
        RECT -69.525 203.835 -69.195 204.165 ;
        RECT -69.525 202.475 -69.195 202.805 ;
        RECT -69.525 201.115 -69.195 201.445 ;
        RECT -69.525 199.755 -69.195 200.085 ;
        RECT -69.525 198.395 -69.195 198.725 ;
        RECT -69.525 197.035 -69.195 197.365 ;
        RECT -69.525 195.675 -69.195 196.005 ;
        RECT -69.525 194.315 -69.195 194.645 ;
        RECT -69.525 192.955 -69.195 193.285 ;
        RECT -69.525 191.595 -69.195 191.925 ;
        RECT -69.525 190.235 -69.195 190.565 ;
        RECT -69.525 188.875 -69.195 189.205 ;
        RECT -69.525 187.515 -69.195 187.845 ;
        RECT -69.525 186.155 -69.195 186.485 ;
        RECT -69.525 184.795 -69.195 185.125 ;
        RECT -69.525 183.435 -69.195 183.765 ;
        RECT -69.525 182.075 -69.195 182.405 ;
        RECT -69.525 180.715 -69.195 181.045 ;
        RECT -69.525 179.355 -69.195 179.685 ;
        RECT -69.525 177.995 -69.195 178.325 ;
        RECT -69.525 176.635 -69.195 176.965 ;
        RECT -69.525 175.275 -69.195 175.605 ;
        RECT -69.525 173.915 -69.195 174.245 ;
        RECT -69.525 172.555 -69.195 172.885 ;
        RECT -69.525 171.195 -69.195 171.525 ;
        RECT -69.525 169.835 -69.195 170.165 ;
        RECT -69.525 168.475 -69.195 168.805 ;
        RECT -69.525 167.115 -69.195 167.445 ;
        RECT -69.525 165.755 -69.195 166.085 ;
        RECT -69.525 164.395 -69.195 164.725 ;
        RECT -69.525 163.035 -69.195 163.365 ;
        RECT -69.525 161.675 -69.195 162.005 ;
        RECT -69.525 160.315 -69.195 160.645 ;
        RECT -69.525 158.955 -69.195 159.285 ;
        RECT -69.525 157.595 -69.195 157.925 ;
        RECT -69.525 156.235 -69.195 156.565 ;
        RECT -69.525 154.875 -69.195 155.205 ;
        RECT -69.525 153.515 -69.195 153.845 ;
        RECT -69.525 152.155 -69.195 152.485 ;
        RECT -69.525 150.795 -69.195 151.125 ;
        RECT -69.525 149.435 -69.195 149.765 ;
        RECT -69.525 148.075 -69.195 148.405 ;
        RECT -69.525 146.715 -69.195 147.045 ;
        RECT -69.525 145.355 -69.195 145.685 ;
        RECT -69.525 143.995 -69.195 144.325 ;
        RECT -69.525 142.635 -69.195 142.965 ;
        RECT -69.525 141.275 -69.195 141.605 ;
        RECT -69.525 139.915 -69.195 140.245 ;
        RECT -69.525 138.555 -69.195 138.885 ;
        RECT -69.525 137.195 -69.195 137.525 ;
        RECT -69.525 135.835 -69.195 136.165 ;
        RECT -69.525 134.475 -69.195 134.805 ;
        RECT -69.525 133.115 -69.195 133.445 ;
        RECT -69.525 131.755 -69.195 132.085 ;
        RECT -69.525 130.395 -69.195 130.725 ;
        RECT -69.525 129.035 -69.195 129.365 ;
        RECT -69.525 127.675 -69.195 128.005 ;
        RECT -69.525 126.315 -69.195 126.645 ;
        RECT -69.525 124.955 -69.195 125.285 ;
        RECT -69.525 123.595 -69.195 123.925 ;
        RECT -69.525 122.235 -69.195 122.565 ;
        RECT -69.525 120.875 -69.195 121.205 ;
        RECT -69.525 119.515 -69.195 119.845 ;
        RECT -69.525 118.155 -69.195 118.485 ;
        RECT -69.525 116.795 -69.195 117.125 ;
        RECT -69.525 115.435 -69.195 115.765 ;
        RECT -69.525 114.075 -69.195 114.405 ;
        RECT -69.525 112.715 -69.195 113.045 ;
        RECT -69.525 111.355 -69.195 111.685 ;
        RECT -69.525 109.995 -69.195 110.325 ;
        RECT -69.525 108.635 -69.195 108.965 ;
        RECT -69.525 107.275 -69.195 107.605 ;
        RECT -69.525 105.915 -69.195 106.245 ;
        RECT -69.525 104.555 -69.195 104.885 ;
        RECT -69.525 103.195 -69.195 103.525 ;
        RECT -69.525 101.835 -69.195 102.165 ;
        RECT -69.525 100.475 -69.195 100.805 ;
        RECT -69.525 99.115 -69.195 99.445 ;
        RECT -69.525 97.755 -69.195 98.085 ;
        RECT -69.525 96.395 -69.195 96.725 ;
        RECT -69.525 95.035 -69.195 95.365 ;
        RECT -69.525 93.675 -69.195 94.005 ;
        RECT -69.525 92.315 -69.195 92.645 ;
        RECT -69.525 90.955 -69.195 91.285 ;
        RECT -69.525 89.595 -69.195 89.925 ;
        RECT -69.525 88.235 -69.195 88.565 ;
        RECT -69.525 86.875 -69.195 87.205 ;
        RECT -69.525 85.515 -69.195 85.845 ;
        RECT -69.525 84.155 -69.195 84.485 ;
        RECT -69.525 82.795 -69.195 83.125 ;
        RECT -69.525 81.435 -69.195 81.765 ;
        RECT -69.525 80.075 -69.195 80.405 ;
        RECT -69.525 78.715 -69.195 79.045 ;
        RECT -69.525 77.355 -69.195 77.685 ;
        RECT -69.525 75.995 -69.195 76.325 ;
        RECT -69.525 74.635 -69.195 74.965 ;
        RECT -69.525 73.275 -69.195 73.605 ;
        RECT -69.525 71.915 -69.195 72.245 ;
        RECT -69.525 70.555 -69.195 70.885 ;
        RECT -69.525 69.195 -69.195 69.525 ;
        RECT -69.525 67.835 -69.195 68.165 ;
        RECT -69.525 66.475 -69.195 66.805 ;
        RECT -69.525 65.115 -69.195 65.445 ;
        RECT -69.525 63.755 -69.195 64.085 ;
        RECT -69.525 62.395 -69.195 62.725 ;
        RECT -69.525 61.035 -69.195 61.365 ;
        RECT -69.525 59.675 -69.195 60.005 ;
        RECT -69.525 58.315 -69.195 58.645 ;
        RECT -69.525 56.955 -69.195 57.285 ;
        RECT -69.525 55.595 -69.195 55.925 ;
        RECT -69.525 54.235 -69.195 54.565 ;
        RECT -69.525 52.875 -69.195 53.205 ;
        RECT -69.525 51.515 -69.195 51.845 ;
        RECT -69.525 50.155 -69.195 50.485 ;
        RECT -69.525 48.795 -69.195 49.125 ;
        RECT -69.525 47.435 -69.195 47.765 ;
        RECT -69.525 46.075 -69.195 46.405 ;
        RECT -69.525 44.715 -69.195 45.045 ;
        RECT -69.525 43.355 -69.195 43.685 ;
        RECT -69.525 41.995 -69.195 42.325 ;
        RECT -69.525 40.635 -69.195 40.965 ;
        RECT -69.525 39.275 -69.195 39.605 ;
        RECT -69.525 37.915 -69.195 38.245 ;
        RECT -69.525 36.555 -69.195 36.885 ;
        RECT -69.525 35.195 -69.195 35.525 ;
        RECT -69.525 33.835 -69.195 34.165 ;
        RECT -69.525 32.475 -69.195 32.805 ;
        RECT -69.525 31.115 -69.195 31.445 ;
        RECT -69.525 29.755 -69.195 30.085 ;
        RECT -69.525 28.395 -69.195 28.725 ;
        RECT -69.525 27.035 -69.195 27.365 ;
        RECT -69.525 25.675 -69.195 26.005 ;
        RECT -69.525 24.315 -69.195 24.645 ;
        RECT -69.525 22.955 -69.195 23.285 ;
        RECT -69.525 21.595 -69.195 21.925 ;
        RECT -69.525 20.235 -69.195 20.565 ;
        RECT -69.525 18.875 -69.195 19.205 ;
        RECT -69.525 17.515 -69.195 17.845 ;
        RECT -69.525 16.155 -69.195 16.485 ;
        RECT -69.525 14.795 -69.195 15.125 ;
        RECT -69.525 13.435 -69.195 13.765 ;
        RECT -69.525 12.075 -69.195 12.405 ;
        RECT -69.525 10.715 -69.195 11.045 ;
        RECT -69.525 9.355 -69.195 9.685 ;
        RECT -69.525 7.995 -69.195 8.325 ;
        RECT -69.525 6.635 -69.195 6.965 ;
        RECT -69.525 5.275 -69.195 5.605 ;
        RECT -69.525 3.915 -69.195 4.245 ;
        RECT -69.525 2.555 -69.195 2.885 ;
        RECT -69.525 1.195 -69.195 1.525 ;
        RECT -69.525 -0.165 -69.195 0.165 ;
        RECT -69.525 -1.525 -69.195 -1.195 ;
        RECT -69.525 -2.885 -69.195 -2.555 ;
        RECT -69.525 -4.245 -69.195 -3.915 ;
        RECT -69.525 -5.605 -69.195 -5.275 ;
        RECT -69.525 -6.965 -69.195 -6.635 ;
        RECT -69.525 -8.325 -69.195 -7.995 ;
        RECT -69.525 -9.685 -69.195 -9.355 ;
        RECT -69.525 -11.045 -69.195 -10.715 ;
        RECT -69.525 -12.405 -69.195 -12.075 ;
        RECT -69.525 -13.765 -69.195 -13.435 ;
        RECT -69.525 -15.125 -69.195 -14.795 ;
        RECT -69.525 -16.485 -69.195 -16.155 ;
        RECT -69.525 -17.845 -69.195 -17.515 ;
        RECT -69.525 -19.205 -69.195 -18.875 ;
        RECT -69.525 -20.565 -69.195 -20.235 ;
        RECT -69.525 -21.925 -69.195 -21.595 ;
        RECT -69.525 -23.285 -69.195 -22.955 ;
        RECT -69.525 -24.645 -69.195 -24.315 ;
        RECT -69.525 -26.005 -69.195 -25.675 ;
        RECT -69.525 -27.365 -69.195 -27.035 ;
        RECT -69.525 -28.725 -69.195 -28.395 ;
        RECT -69.525 -30.085 -69.195 -29.755 ;
        RECT -69.525 -31.445 -69.195 -31.115 ;
        RECT -69.525 -32.805 -69.195 -32.475 ;
        RECT -69.525 -34.165 -69.195 -33.835 ;
        RECT -69.525 -35.525 -69.195 -35.195 ;
        RECT -69.525 -36.885 -69.195 -36.555 ;
        RECT -69.525 -38.245 -69.195 -37.915 ;
        RECT -69.525 -39.605 -69.195 -39.275 ;
        RECT -69.525 -40.965 -69.195 -40.635 ;
        RECT -69.525 -42.325 -69.195 -41.995 ;
        RECT -69.525 -43.685 -69.195 -43.355 ;
        RECT -69.525 -45.045 -69.195 -44.715 ;
        RECT -69.525 -46.405 -69.195 -46.075 ;
        RECT -69.525 -47.765 -69.195 -47.435 ;
        RECT -69.525 -49.125 -69.195 -48.795 ;
        RECT -69.525 -50.485 -69.195 -50.155 ;
        RECT -69.525 -51.845 -69.195 -51.515 ;
        RECT -69.525 -53.205 -69.195 -52.875 ;
        RECT -69.525 -54.565 -69.195 -54.235 ;
        RECT -69.525 -55.925 -69.195 -55.595 ;
        RECT -69.525 -57.285 -69.195 -56.955 ;
        RECT -69.525 -58.645 -69.195 -58.315 ;
        RECT -69.525 -60.005 -69.195 -59.675 ;
        RECT -69.525 -61.365 -69.195 -61.035 ;
        RECT -69.525 -62.725 -69.195 -62.395 ;
        RECT -69.525 -64.085 -69.195 -63.755 ;
        RECT -69.525 -65.445 -69.195 -65.115 ;
        RECT -69.525 -66.805 -69.195 -66.475 ;
        RECT -69.525 -68.165 -69.195 -67.835 ;
        RECT -69.525 -69.525 -69.195 -69.195 ;
        RECT -69.525 -70.885 -69.195 -70.555 ;
        RECT -69.525 -72.245 -69.195 -71.915 ;
        RECT -69.525 -73.605 -69.195 -73.275 ;
        RECT -69.525 -74.965 -69.195 -74.635 ;
        RECT -69.525 -76.325 -69.195 -75.995 ;
        RECT -69.525 -77.685 -69.195 -77.355 ;
        RECT -69.525 -79.045 -69.195 -78.715 ;
        RECT -69.525 -80.405 -69.195 -80.075 ;
        RECT -69.525 -81.765 -69.195 -81.435 ;
        RECT -69.525 -83.125 -69.195 -82.795 ;
        RECT -69.525 -84.485 -69.195 -84.155 ;
        RECT -69.525 -85.845 -69.195 -85.515 ;
        RECT -69.525 -87.205 -69.195 -86.875 ;
        RECT -69.525 -88.565 -69.195 -88.235 ;
        RECT -69.525 -89.925 -69.195 -89.595 ;
        RECT -69.525 -91.285 -69.195 -90.955 ;
        RECT -69.525 -92.645 -69.195 -92.315 ;
        RECT -69.525 -94.005 -69.195 -93.675 ;
        RECT -69.525 -95.365 -69.195 -95.035 ;
        RECT -69.525 -96.725 -69.195 -96.395 ;
        RECT -69.525 -98.085 -69.195 -97.755 ;
        RECT -69.525 -99.445 -69.195 -99.115 ;
        RECT -69.525 -100.805 -69.195 -100.475 ;
        RECT -69.525 -102.165 -69.195 -101.835 ;
        RECT -69.525 -103.525 -69.195 -103.195 ;
        RECT -69.525 -104.885 -69.195 -104.555 ;
        RECT -69.525 -106.245 -69.195 -105.915 ;
        RECT -69.525 -107.605 -69.195 -107.275 ;
        RECT -69.525 -108.965 -69.195 -108.635 ;
        RECT -69.525 -110.325 -69.195 -109.995 ;
        RECT -69.525 -111.685 -69.195 -111.355 ;
        RECT -69.525 -113.045 -69.195 -112.715 ;
        RECT -69.525 -114.405 -69.195 -114.075 ;
        RECT -69.525 -115.765 -69.195 -115.435 ;
        RECT -69.525 -117.125 -69.195 -116.795 ;
        RECT -69.525 -118.485 -69.195 -118.155 ;
        RECT -69.525 -119.845 -69.195 -119.515 ;
        RECT -69.525 -121.205 -69.195 -120.875 ;
        RECT -69.525 -122.565 -69.195 -122.235 ;
        RECT -69.525 -123.925 -69.195 -123.595 ;
        RECT -69.525 -125.285 -69.195 -124.955 ;
        RECT -69.525 -126.645 -69.195 -126.315 ;
        RECT -69.525 -128.005 -69.195 -127.675 ;
        RECT -69.525 -129.365 -69.195 -129.035 ;
        RECT -69.525 -130.725 -69.195 -130.395 ;
        RECT -69.525 -131.47 -69.195 -131.14 ;
        RECT -69.525 -133.445 -69.195 -133.115 ;
        RECT -69.525 -134.805 -69.195 -134.475 ;
        RECT -69.525 -136.165 -69.195 -135.835 ;
        RECT -69.525 -137.525 -69.195 -137.195 ;
        RECT -69.525 -140.245 -69.195 -139.915 ;
        RECT -69.525 -141.605 -69.195 -141.275 ;
        RECT -69.525 -142.965 -69.195 -142.635 ;
        RECT -69.525 -144.31 -69.195 -143.98 ;
        RECT -69.525 -145.685 -69.195 -145.355 ;
        RECT -69.525 -147.045 -69.195 -146.715 ;
        RECT -69.525 -149.765 -69.195 -149.435 ;
        RECT -69.525 -152.485 -69.195 -152.155 ;
        RECT -69.525 -153.845 -69.195 -153.515 ;
        RECT -69.525 -155.205 -69.195 -154.875 ;
        RECT -69.525 -156.565 -69.195 -156.235 ;
        RECT -69.525 -157.925 -69.195 -157.595 ;
        RECT -69.525 -159.285 -69.195 -158.955 ;
        RECT -69.525 -162.005 -69.195 -161.675 ;
        RECT -69.525 -163.365 -69.195 -163.035 ;
        RECT -69.525 -164.725 -69.195 -164.395 ;
        RECT -69.525 -166.085 -69.195 -165.755 ;
        RECT -69.525 -167.445 -69.195 -167.115 ;
        RECT -69.525 -168.805 -69.195 -168.475 ;
        RECT -69.525 -170.165 -69.195 -169.835 ;
        RECT -69.525 -171.525 -69.195 -171.195 ;
        RECT -69.525 -172.885 -69.195 -172.555 ;
        RECT -69.525 -174.245 -69.195 -173.915 ;
        RECT -69.525 -175.605 -69.195 -175.275 ;
        RECT -69.525 -176.965 -69.195 -176.635 ;
        RECT -69.525 -178.325 -69.195 -177.995 ;
        RECT -69.525 -179.685 -69.195 -179.355 ;
        RECT -69.525 -181.045 -69.195 -180.715 ;
        RECT -69.525 -182.405 -69.195 -182.075 ;
        RECT -69.525 -183.765 -69.195 -183.435 ;
        RECT -69.525 -185.125 -69.195 -184.795 ;
        RECT -69.525 -186.485 -69.195 -186.155 ;
        RECT -69.525 -187.845 -69.195 -187.515 ;
        RECT -69.525 -189.205 -69.195 -188.875 ;
        RECT -69.525 -190.565 -69.195 -190.235 ;
        RECT -69.525 -191.925 -69.195 -191.595 ;
        RECT -69.525 -193.285 -69.195 -192.955 ;
        RECT -69.525 -194.645 -69.195 -194.315 ;
        RECT -69.525 -196.005 -69.195 -195.675 ;
        RECT -69.525 -197.365 -69.195 -197.035 ;
        RECT -69.525 -198.725 -69.195 -198.395 ;
        RECT -69.525 -200.085 -69.195 -199.755 ;
        RECT -69.525 -201.445 -69.195 -201.115 ;
        RECT -69.525 -202.805 -69.195 -202.475 ;
        RECT -69.525 -204.165 -69.195 -203.835 ;
        RECT -69.525 -205.525 -69.195 -205.195 ;
        RECT -69.525 -206.885 -69.195 -206.555 ;
        RECT -69.525 -208.245 -69.195 -207.915 ;
        RECT -69.525 -209.605 -69.195 -209.275 ;
        RECT -69.525 -210.965 -69.195 -210.635 ;
        RECT -69.525 -212.325 -69.195 -211.995 ;
        RECT -69.525 -213.685 -69.195 -213.355 ;
        RECT -69.525 -215.045 -69.195 -214.715 ;
        RECT -69.525 -216.405 -69.195 -216.075 ;
        RECT -69.525 -217.765 -69.195 -217.435 ;
        RECT -69.525 -219.125 -69.195 -218.795 ;
        RECT -69.525 -220.485 -69.195 -220.155 ;
        RECT -69.525 -221.845 -69.195 -221.515 ;
        RECT -69.525 -223.205 -69.195 -222.875 ;
        RECT -69.525 -224.565 -69.195 -224.235 ;
        RECT -69.525 -226.155 -69.195 -225.825 ;
        RECT -69.525 -227.285 -69.195 -226.955 ;
        RECT -69.525 -228.645 -69.195 -228.315 ;
        RECT -69.525 -230.005 -69.195 -229.675 ;
        RECT -69.525 -234.085 -69.195 -233.755 ;
        RECT -69.525 -235.445 -69.195 -235.115 ;
        RECT -69.525 -236.805 -69.195 -236.475 ;
        RECT -69.525 -238.165 -69.195 -237.835 ;
        RECT -69.525 -243.81 -69.195 -242.68 ;
        RECT -69.52 -243.925 -69.2 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.165 246.76 -67.835 247.89 ;
        RECT -68.165 241.915 -67.835 242.245 ;
        RECT -68.165 240.555 -67.835 240.885 ;
        RECT -68.165 239.195 -67.835 239.525 ;
        RECT -68.165 237.835 -67.835 238.165 ;
        RECT -68.165 236.475 -67.835 236.805 ;
        RECT -68.165 235.115 -67.835 235.445 ;
        RECT -68.165 233.755 -67.835 234.085 ;
        RECT -68.165 232.395 -67.835 232.725 ;
        RECT -68.165 231.035 -67.835 231.365 ;
        RECT -68.165 229.675 -67.835 230.005 ;
        RECT -68.165 228.315 -67.835 228.645 ;
        RECT -68.165 226.955 -67.835 227.285 ;
        RECT -68.165 225.595 -67.835 225.925 ;
        RECT -68.165 224.235 -67.835 224.565 ;
        RECT -68.165 222.875 -67.835 223.205 ;
        RECT -68.165 221.515 -67.835 221.845 ;
        RECT -68.165 220.155 -67.835 220.485 ;
        RECT -68.165 218.795 -67.835 219.125 ;
        RECT -68.165 217.435 -67.835 217.765 ;
        RECT -68.165 216.075 -67.835 216.405 ;
        RECT -68.165 214.715 -67.835 215.045 ;
        RECT -68.165 213.355 -67.835 213.685 ;
        RECT -68.165 211.995 -67.835 212.325 ;
        RECT -68.165 210.635 -67.835 210.965 ;
        RECT -68.165 209.275 -67.835 209.605 ;
        RECT -68.165 207.915 -67.835 208.245 ;
        RECT -68.165 206.555 -67.835 206.885 ;
        RECT -68.165 205.195 -67.835 205.525 ;
        RECT -68.165 203.835 -67.835 204.165 ;
        RECT -68.165 202.475 -67.835 202.805 ;
        RECT -68.165 201.115 -67.835 201.445 ;
        RECT -68.165 199.755 -67.835 200.085 ;
        RECT -68.165 198.395 -67.835 198.725 ;
        RECT -68.165 197.035 -67.835 197.365 ;
        RECT -68.165 195.675 -67.835 196.005 ;
        RECT -68.165 194.315 -67.835 194.645 ;
        RECT -68.165 192.955 -67.835 193.285 ;
        RECT -68.165 191.595 -67.835 191.925 ;
        RECT -68.165 190.235 -67.835 190.565 ;
        RECT -68.165 188.875 -67.835 189.205 ;
        RECT -68.165 187.515 -67.835 187.845 ;
        RECT -68.165 186.155 -67.835 186.485 ;
        RECT -68.165 184.795 -67.835 185.125 ;
        RECT -68.165 183.435 -67.835 183.765 ;
        RECT -68.165 182.075 -67.835 182.405 ;
        RECT -68.165 180.715 -67.835 181.045 ;
        RECT -68.165 179.355 -67.835 179.685 ;
        RECT -68.165 177.995 -67.835 178.325 ;
        RECT -68.165 176.635 -67.835 176.965 ;
        RECT -68.165 175.275 -67.835 175.605 ;
        RECT -68.165 173.915 -67.835 174.245 ;
        RECT -68.165 172.555 -67.835 172.885 ;
        RECT -68.165 171.195 -67.835 171.525 ;
        RECT -68.165 169.835 -67.835 170.165 ;
        RECT -68.165 168.475 -67.835 168.805 ;
        RECT -68.165 167.115 -67.835 167.445 ;
        RECT -68.165 165.755 -67.835 166.085 ;
        RECT -68.165 164.395 -67.835 164.725 ;
        RECT -68.165 163.035 -67.835 163.365 ;
        RECT -68.165 161.675 -67.835 162.005 ;
        RECT -68.165 160.315 -67.835 160.645 ;
        RECT -68.165 158.955 -67.835 159.285 ;
        RECT -68.165 157.595 -67.835 157.925 ;
        RECT -68.165 156.235 -67.835 156.565 ;
        RECT -68.165 154.875 -67.835 155.205 ;
        RECT -68.165 153.515 -67.835 153.845 ;
        RECT -68.165 152.155 -67.835 152.485 ;
        RECT -68.165 150.795 -67.835 151.125 ;
        RECT -68.165 149.435 -67.835 149.765 ;
        RECT -68.165 148.075 -67.835 148.405 ;
        RECT -68.165 146.715 -67.835 147.045 ;
        RECT -68.165 145.355 -67.835 145.685 ;
        RECT -68.165 143.995 -67.835 144.325 ;
        RECT -68.165 142.635 -67.835 142.965 ;
        RECT -68.165 141.275 -67.835 141.605 ;
        RECT -68.165 139.915 -67.835 140.245 ;
        RECT -68.165 138.555 -67.835 138.885 ;
        RECT -68.165 137.195 -67.835 137.525 ;
        RECT -68.165 135.835 -67.835 136.165 ;
        RECT -68.165 134.475 -67.835 134.805 ;
        RECT -68.165 133.115 -67.835 133.445 ;
        RECT -68.165 131.755 -67.835 132.085 ;
        RECT -68.165 130.395 -67.835 130.725 ;
        RECT -68.165 129.035 -67.835 129.365 ;
        RECT -68.165 127.675 -67.835 128.005 ;
        RECT -68.165 126.315 -67.835 126.645 ;
        RECT -68.165 124.955 -67.835 125.285 ;
        RECT -68.165 123.595 -67.835 123.925 ;
        RECT -68.165 122.235 -67.835 122.565 ;
        RECT -68.165 120.875 -67.835 121.205 ;
        RECT -68.165 119.515 -67.835 119.845 ;
        RECT -68.165 118.155 -67.835 118.485 ;
        RECT -68.165 116.795 -67.835 117.125 ;
        RECT -68.165 115.435 -67.835 115.765 ;
        RECT -68.165 114.075 -67.835 114.405 ;
        RECT -68.165 112.715 -67.835 113.045 ;
        RECT -68.165 111.355 -67.835 111.685 ;
        RECT -68.165 109.995 -67.835 110.325 ;
        RECT -68.165 108.635 -67.835 108.965 ;
        RECT -68.165 107.275 -67.835 107.605 ;
        RECT -68.165 105.915 -67.835 106.245 ;
        RECT -68.165 104.555 -67.835 104.885 ;
        RECT -68.165 103.195 -67.835 103.525 ;
        RECT -68.165 101.835 -67.835 102.165 ;
        RECT -68.165 100.475 -67.835 100.805 ;
        RECT -68.165 99.115 -67.835 99.445 ;
        RECT -68.165 97.755 -67.835 98.085 ;
        RECT -68.165 96.395 -67.835 96.725 ;
        RECT -68.165 95.035 -67.835 95.365 ;
        RECT -68.165 93.675 -67.835 94.005 ;
        RECT -68.165 92.315 -67.835 92.645 ;
        RECT -68.165 90.955 -67.835 91.285 ;
        RECT -68.165 89.595 -67.835 89.925 ;
        RECT -68.165 88.235 -67.835 88.565 ;
        RECT -68.165 86.875 -67.835 87.205 ;
        RECT -68.165 85.515 -67.835 85.845 ;
        RECT -68.165 84.155 -67.835 84.485 ;
        RECT -68.165 82.795 -67.835 83.125 ;
        RECT -68.165 81.435 -67.835 81.765 ;
        RECT -68.165 80.075 -67.835 80.405 ;
        RECT -68.165 78.715 -67.835 79.045 ;
        RECT -68.165 77.355 -67.835 77.685 ;
        RECT -68.165 75.995 -67.835 76.325 ;
        RECT -68.165 74.635 -67.835 74.965 ;
        RECT -68.165 73.275 -67.835 73.605 ;
        RECT -68.165 71.915 -67.835 72.245 ;
        RECT -68.165 70.555 -67.835 70.885 ;
        RECT -68.165 69.195 -67.835 69.525 ;
        RECT -68.165 67.835 -67.835 68.165 ;
        RECT -68.165 66.475 -67.835 66.805 ;
        RECT -68.165 65.115 -67.835 65.445 ;
        RECT -68.165 63.755 -67.835 64.085 ;
        RECT -68.165 62.395 -67.835 62.725 ;
        RECT -68.165 61.035 -67.835 61.365 ;
        RECT -68.165 59.675 -67.835 60.005 ;
        RECT -68.165 58.315 -67.835 58.645 ;
        RECT -68.165 56.955 -67.835 57.285 ;
        RECT -68.165 55.595 -67.835 55.925 ;
        RECT -68.165 54.235 -67.835 54.565 ;
        RECT -68.165 52.875 -67.835 53.205 ;
        RECT -68.165 51.515 -67.835 51.845 ;
        RECT -68.165 50.155 -67.835 50.485 ;
        RECT -68.165 48.795 -67.835 49.125 ;
        RECT -68.165 47.435 -67.835 47.765 ;
        RECT -68.165 46.075 -67.835 46.405 ;
        RECT -68.165 44.715 -67.835 45.045 ;
        RECT -68.165 43.355 -67.835 43.685 ;
        RECT -68.165 41.995 -67.835 42.325 ;
        RECT -68.165 40.635 -67.835 40.965 ;
        RECT -68.165 39.275 -67.835 39.605 ;
        RECT -68.165 37.915 -67.835 38.245 ;
        RECT -68.165 36.555 -67.835 36.885 ;
        RECT -68.165 35.195 -67.835 35.525 ;
        RECT -68.165 33.835 -67.835 34.165 ;
        RECT -68.165 32.475 -67.835 32.805 ;
        RECT -68.165 31.115 -67.835 31.445 ;
        RECT -68.165 29.755 -67.835 30.085 ;
        RECT -68.165 28.395 -67.835 28.725 ;
        RECT -68.165 27.035 -67.835 27.365 ;
        RECT -68.165 25.675 -67.835 26.005 ;
        RECT -68.165 24.315 -67.835 24.645 ;
        RECT -68.165 22.955 -67.835 23.285 ;
        RECT -68.165 21.595 -67.835 21.925 ;
        RECT -68.165 20.235 -67.835 20.565 ;
        RECT -68.165 18.875 -67.835 19.205 ;
        RECT -68.165 17.515 -67.835 17.845 ;
        RECT -68.165 16.155 -67.835 16.485 ;
        RECT -68.165 14.795 -67.835 15.125 ;
        RECT -68.165 13.435 -67.835 13.765 ;
        RECT -68.165 12.075 -67.835 12.405 ;
        RECT -68.165 10.715 -67.835 11.045 ;
        RECT -68.165 9.355 -67.835 9.685 ;
        RECT -68.165 7.995 -67.835 8.325 ;
        RECT -68.165 6.635 -67.835 6.965 ;
        RECT -68.165 5.275 -67.835 5.605 ;
        RECT -68.165 3.915 -67.835 4.245 ;
        RECT -68.165 2.555 -67.835 2.885 ;
        RECT -68.165 1.195 -67.835 1.525 ;
        RECT -68.165 -0.165 -67.835 0.165 ;
        RECT -68.165 -1.525 -67.835 -1.195 ;
        RECT -68.165 -2.885 -67.835 -2.555 ;
        RECT -68.165 -4.245 -67.835 -3.915 ;
        RECT -68.165 -5.605 -67.835 -5.275 ;
        RECT -68.165 -6.965 -67.835 -6.635 ;
        RECT -68.165 -8.325 -67.835 -7.995 ;
        RECT -68.165 -9.685 -67.835 -9.355 ;
        RECT -68.165 -11.045 -67.835 -10.715 ;
        RECT -68.165 -12.405 -67.835 -12.075 ;
        RECT -68.165 -13.765 -67.835 -13.435 ;
        RECT -68.165 -15.125 -67.835 -14.795 ;
        RECT -68.165 -16.485 -67.835 -16.155 ;
        RECT -68.165 -17.845 -67.835 -17.515 ;
        RECT -68.165 -19.205 -67.835 -18.875 ;
        RECT -68.165 -20.565 -67.835 -20.235 ;
        RECT -68.165 -21.925 -67.835 -21.595 ;
        RECT -68.165 -23.285 -67.835 -22.955 ;
        RECT -68.165 -24.645 -67.835 -24.315 ;
        RECT -68.165 -26.005 -67.835 -25.675 ;
        RECT -68.165 -27.365 -67.835 -27.035 ;
        RECT -68.165 -28.725 -67.835 -28.395 ;
        RECT -68.165 -30.085 -67.835 -29.755 ;
        RECT -68.165 -31.445 -67.835 -31.115 ;
        RECT -68.165 -32.805 -67.835 -32.475 ;
        RECT -68.165 -34.165 -67.835 -33.835 ;
        RECT -68.165 -35.525 -67.835 -35.195 ;
        RECT -68.165 -36.885 -67.835 -36.555 ;
        RECT -68.165 -38.245 -67.835 -37.915 ;
        RECT -68.165 -39.605 -67.835 -39.275 ;
        RECT -68.165 -40.965 -67.835 -40.635 ;
        RECT -68.165 -42.325 -67.835 -41.995 ;
        RECT -68.165 -43.685 -67.835 -43.355 ;
        RECT -68.165 -45.045 -67.835 -44.715 ;
        RECT -68.165 -46.405 -67.835 -46.075 ;
        RECT -68.165 -47.765 -67.835 -47.435 ;
        RECT -68.165 -49.125 -67.835 -48.795 ;
        RECT -68.165 -50.485 -67.835 -50.155 ;
        RECT -68.165 -51.845 -67.835 -51.515 ;
        RECT -68.165 -53.205 -67.835 -52.875 ;
        RECT -68.165 -54.565 -67.835 -54.235 ;
        RECT -68.165 -55.925 -67.835 -55.595 ;
        RECT -68.165 -57.285 -67.835 -56.955 ;
        RECT -68.165 -58.645 -67.835 -58.315 ;
        RECT -68.165 -60.005 -67.835 -59.675 ;
        RECT -68.165 -61.365 -67.835 -61.035 ;
        RECT -68.165 -62.725 -67.835 -62.395 ;
        RECT -68.165 -64.085 -67.835 -63.755 ;
        RECT -68.165 -65.445 -67.835 -65.115 ;
        RECT -68.165 -66.805 -67.835 -66.475 ;
        RECT -68.165 -68.165 -67.835 -67.835 ;
        RECT -68.165 -69.525 -67.835 -69.195 ;
        RECT -68.165 -70.885 -67.835 -70.555 ;
        RECT -68.165 -72.245 -67.835 -71.915 ;
        RECT -68.165 -73.605 -67.835 -73.275 ;
        RECT -68.165 -74.965 -67.835 -74.635 ;
        RECT -68.165 -76.325 -67.835 -75.995 ;
        RECT -68.165 -77.685 -67.835 -77.355 ;
        RECT -68.165 -79.045 -67.835 -78.715 ;
        RECT -68.165 -80.405 -67.835 -80.075 ;
        RECT -68.165 -81.765 -67.835 -81.435 ;
        RECT -68.165 -83.125 -67.835 -82.795 ;
        RECT -68.165 -84.485 -67.835 -84.155 ;
        RECT -68.165 -85.845 -67.835 -85.515 ;
        RECT -68.165 -87.205 -67.835 -86.875 ;
        RECT -68.165 -88.565 -67.835 -88.235 ;
        RECT -68.165 -89.925 -67.835 -89.595 ;
        RECT -68.165 -91.285 -67.835 -90.955 ;
        RECT -68.165 -92.645 -67.835 -92.315 ;
        RECT -68.165 -94.005 -67.835 -93.675 ;
        RECT -68.165 -95.365 -67.835 -95.035 ;
        RECT -68.165 -96.725 -67.835 -96.395 ;
        RECT -68.165 -98.085 -67.835 -97.755 ;
        RECT -68.165 -99.445 -67.835 -99.115 ;
        RECT -68.165 -100.805 -67.835 -100.475 ;
        RECT -68.165 -102.165 -67.835 -101.835 ;
        RECT -68.165 -103.525 -67.835 -103.195 ;
        RECT -68.165 -104.885 -67.835 -104.555 ;
        RECT -68.165 -106.245 -67.835 -105.915 ;
        RECT -68.165 -107.605 -67.835 -107.275 ;
        RECT -68.165 -108.965 -67.835 -108.635 ;
        RECT -68.165 -110.325 -67.835 -109.995 ;
        RECT -68.165 -111.685 -67.835 -111.355 ;
        RECT -68.165 -113.045 -67.835 -112.715 ;
        RECT -68.165 -114.405 -67.835 -114.075 ;
        RECT -68.165 -115.765 -67.835 -115.435 ;
        RECT -68.165 -117.125 -67.835 -116.795 ;
        RECT -68.165 -118.485 -67.835 -118.155 ;
        RECT -68.165 -119.845 -67.835 -119.515 ;
        RECT -68.165 -121.205 -67.835 -120.875 ;
        RECT -68.165 -122.565 -67.835 -122.235 ;
        RECT -68.165 -123.925 -67.835 -123.595 ;
        RECT -68.165 -125.285 -67.835 -124.955 ;
        RECT -68.165 -126.645 -67.835 -126.315 ;
        RECT -68.165 -129.365 -67.835 -129.035 ;
        RECT -68.165 -130.725 -67.835 -130.395 ;
        RECT -68.165 -131.47 -67.835 -131.14 ;
        RECT -68.165 -133.445 -67.835 -133.115 ;
        RECT -68.165 -134.805 -67.835 -134.475 ;
        RECT -68.165 -136.165 -67.835 -135.835 ;
        RECT -68.165 -137.525 -67.835 -137.195 ;
        RECT -68.165 -140.245 -67.835 -139.915 ;
        RECT -68.165 -141.605 -67.835 -141.275 ;
        RECT -68.165 -142.965 -67.835 -142.635 ;
        RECT -68.165 -144.31 -67.835 -143.98 ;
        RECT -68.165 -145.685 -67.835 -145.355 ;
        RECT -68.165 -147.045 -67.835 -146.715 ;
        RECT -68.165 -149.765 -67.835 -149.435 ;
        RECT -68.16 -151.8 -67.84 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.165 -234.085 -67.835 -233.755 ;
        RECT -68.165 -235.445 -67.835 -235.115 ;
        RECT -68.165 -236.805 -67.835 -236.475 ;
        RECT -68.165 -238.165 -67.835 -237.835 ;
        RECT -68.165 -243.81 -67.835 -242.68 ;
        RECT -68.16 -243.925 -67.84 -231.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.805 -122.565 -66.475 -122.235 ;
        RECT -66.805 -123.925 -66.475 -123.595 ;
        RECT -66.805 -125.285 -66.475 -124.955 ;
        RECT -66.805 -126.645 -66.475 -126.315 ;
        RECT -66.805 -129.365 -66.475 -129.035 ;
        RECT -66.805 -130.725 -66.475 -130.395 ;
        RECT -66.805 -131.47 -66.475 -131.14 ;
        RECT -66.805 -133.445 -66.475 -133.115 ;
        RECT -66.805 -134.805 -66.475 -134.475 ;
        RECT -66.805 -136.165 -66.475 -135.835 ;
        RECT -66.805 -137.525 -66.475 -137.195 ;
        RECT -66.805 -140.245 -66.475 -139.915 ;
        RECT -66.805 -141.605 -66.475 -141.275 ;
        RECT -66.805 -142.965 -66.475 -142.635 ;
        RECT -66.805 -144.31 -66.475 -143.98 ;
        RECT -66.805 -145.685 -66.475 -145.355 ;
        RECT -66.805 -147.045 -66.475 -146.715 ;
        RECT -66.805 -149.765 -66.475 -149.435 ;
        RECT -66.8 -149.765 -66.48 248.005 ;
        RECT -66.805 246.76 -66.475 247.89 ;
        RECT -66.805 241.915 -66.475 242.245 ;
        RECT -66.805 240.555 -66.475 240.885 ;
        RECT -66.805 239.195 -66.475 239.525 ;
        RECT -66.805 237.835 -66.475 238.165 ;
        RECT -66.805 236.475 -66.475 236.805 ;
        RECT -66.805 235.115 -66.475 235.445 ;
        RECT -66.805 233.755 -66.475 234.085 ;
        RECT -66.805 232.395 -66.475 232.725 ;
        RECT -66.805 231.035 -66.475 231.365 ;
        RECT -66.805 229.675 -66.475 230.005 ;
        RECT -66.805 228.315 -66.475 228.645 ;
        RECT -66.805 226.955 -66.475 227.285 ;
        RECT -66.805 225.595 -66.475 225.925 ;
        RECT -66.805 224.235 -66.475 224.565 ;
        RECT -66.805 222.875 -66.475 223.205 ;
        RECT -66.805 221.515 -66.475 221.845 ;
        RECT -66.805 220.155 -66.475 220.485 ;
        RECT -66.805 218.795 -66.475 219.125 ;
        RECT -66.805 217.435 -66.475 217.765 ;
        RECT -66.805 216.075 -66.475 216.405 ;
        RECT -66.805 214.715 -66.475 215.045 ;
        RECT -66.805 213.355 -66.475 213.685 ;
        RECT -66.805 211.995 -66.475 212.325 ;
        RECT -66.805 210.635 -66.475 210.965 ;
        RECT -66.805 209.275 -66.475 209.605 ;
        RECT -66.805 207.915 -66.475 208.245 ;
        RECT -66.805 206.555 -66.475 206.885 ;
        RECT -66.805 205.195 -66.475 205.525 ;
        RECT -66.805 203.835 -66.475 204.165 ;
        RECT -66.805 202.475 -66.475 202.805 ;
        RECT -66.805 201.115 -66.475 201.445 ;
        RECT -66.805 199.755 -66.475 200.085 ;
        RECT -66.805 198.395 -66.475 198.725 ;
        RECT -66.805 197.035 -66.475 197.365 ;
        RECT -66.805 195.675 -66.475 196.005 ;
        RECT -66.805 194.315 -66.475 194.645 ;
        RECT -66.805 192.955 -66.475 193.285 ;
        RECT -66.805 191.595 -66.475 191.925 ;
        RECT -66.805 190.235 -66.475 190.565 ;
        RECT -66.805 188.875 -66.475 189.205 ;
        RECT -66.805 187.515 -66.475 187.845 ;
        RECT -66.805 186.155 -66.475 186.485 ;
        RECT -66.805 184.795 -66.475 185.125 ;
        RECT -66.805 183.435 -66.475 183.765 ;
        RECT -66.805 182.075 -66.475 182.405 ;
        RECT -66.805 180.715 -66.475 181.045 ;
        RECT -66.805 179.355 -66.475 179.685 ;
        RECT -66.805 177.995 -66.475 178.325 ;
        RECT -66.805 176.635 -66.475 176.965 ;
        RECT -66.805 175.275 -66.475 175.605 ;
        RECT -66.805 173.915 -66.475 174.245 ;
        RECT -66.805 172.555 -66.475 172.885 ;
        RECT -66.805 171.195 -66.475 171.525 ;
        RECT -66.805 169.835 -66.475 170.165 ;
        RECT -66.805 168.475 -66.475 168.805 ;
        RECT -66.805 167.115 -66.475 167.445 ;
        RECT -66.805 165.755 -66.475 166.085 ;
        RECT -66.805 164.395 -66.475 164.725 ;
        RECT -66.805 163.035 -66.475 163.365 ;
        RECT -66.805 161.675 -66.475 162.005 ;
        RECT -66.805 160.315 -66.475 160.645 ;
        RECT -66.805 158.955 -66.475 159.285 ;
        RECT -66.805 157.595 -66.475 157.925 ;
        RECT -66.805 156.235 -66.475 156.565 ;
        RECT -66.805 154.875 -66.475 155.205 ;
        RECT -66.805 153.515 -66.475 153.845 ;
        RECT -66.805 152.155 -66.475 152.485 ;
        RECT -66.805 150.795 -66.475 151.125 ;
        RECT -66.805 149.435 -66.475 149.765 ;
        RECT -66.805 148.075 -66.475 148.405 ;
        RECT -66.805 146.715 -66.475 147.045 ;
        RECT -66.805 145.355 -66.475 145.685 ;
        RECT -66.805 143.995 -66.475 144.325 ;
        RECT -66.805 142.635 -66.475 142.965 ;
        RECT -66.805 141.275 -66.475 141.605 ;
        RECT -66.805 139.915 -66.475 140.245 ;
        RECT -66.805 138.555 -66.475 138.885 ;
        RECT -66.805 137.195 -66.475 137.525 ;
        RECT -66.805 135.835 -66.475 136.165 ;
        RECT -66.805 134.475 -66.475 134.805 ;
        RECT -66.805 133.115 -66.475 133.445 ;
        RECT -66.805 131.755 -66.475 132.085 ;
        RECT -66.805 130.395 -66.475 130.725 ;
        RECT -66.805 129.035 -66.475 129.365 ;
        RECT -66.805 127.675 -66.475 128.005 ;
        RECT -66.805 126.315 -66.475 126.645 ;
        RECT -66.805 124.955 -66.475 125.285 ;
        RECT -66.805 123.595 -66.475 123.925 ;
        RECT -66.805 122.235 -66.475 122.565 ;
        RECT -66.805 120.875 -66.475 121.205 ;
        RECT -66.805 119.515 -66.475 119.845 ;
        RECT -66.805 118.155 -66.475 118.485 ;
        RECT -66.805 116.795 -66.475 117.125 ;
        RECT -66.805 115.435 -66.475 115.765 ;
        RECT -66.805 114.075 -66.475 114.405 ;
        RECT -66.805 112.715 -66.475 113.045 ;
        RECT -66.805 111.355 -66.475 111.685 ;
        RECT -66.805 109.995 -66.475 110.325 ;
        RECT -66.805 108.635 -66.475 108.965 ;
        RECT -66.805 107.275 -66.475 107.605 ;
        RECT -66.805 105.915 -66.475 106.245 ;
        RECT -66.805 104.555 -66.475 104.885 ;
        RECT -66.805 103.195 -66.475 103.525 ;
        RECT -66.805 101.835 -66.475 102.165 ;
        RECT -66.805 100.475 -66.475 100.805 ;
        RECT -66.805 99.115 -66.475 99.445 ;
        RECT -66.805 97.755 -66.475 98.085 ;
        RECT -66.805 96.395 -66.475 96.725 ;
        RECT -66.805 95.035 -66.475 95.365 ;
        RECT -66.805 93.675 -66.475 94.005 ;
        RECT -66.805 92.315 -66.475 92.645 ;
        RECT -66.805 90.955 -66.475 91.285 ;
        RECT -66.805 89.595 -66.475 89.925 ;
        RECT -66.805 88.235 -66.475 88.565 ;
        RECT -66.805 86.875 -66.475 87.205 ;
        RECT -66.805 85.515 -66.475 85.845 ;
        RECT -66.805 84.155 -66.475 84.485 ;
        RECT -66.805 82.795 -66.475 83.125 ;
        RECT -66.805 81.435 -66.475 81.765 ;
        RECT -66.805 80.075 -66.475 80.405 ;
        RECT -66.805 78.715 -66.475 79.045 ;
        RECT -66.805 77.355 -66.475 77.685 ;
        RECT -66.805 75.995 -66.475 76.325 ;
        RECT -66.805 74.635 -66.475 74.965 ;
        RECT -66.805 73.275 -66.475 73.605 ;
        RECT -66.805 71.915 -66.475 72.245 ;
        RECT -66.805 70.555 -66.475 70.885 ;
        RECT -66.805 69.195 -66.475 69.525 ;
        RECT -66.805 67.835 -66.475 68.165 ;
        RECT -66.805 66.475 -66.475 66.805 ;
        RECT -66.805 65.115 -66.475 65.445 ;
        RECT -66.805 63.755 -66.475 64.085 ;
        RECT -66.805 62.395 -66.475 62.725 ;
        RECT -66.805 61.035 -66.475 61.365 ;
        RECT -66.805 59.675 -66.475 60.005 ;
        RECT -66.805 58.315 -66.475 58.645 ;
        RECT -66.805 56.955 -66.475 57.285 ;
        RECT -66.805 55.595 -66.475 55.925 ;
        RECT -66.805 54.235 -66.475 54.565 ;
        RECT -66.805 52.875 -66.475 53.205 ;
        RECT -66.805 51.515 -66.475 51.845 ;
        RECT -66.805 50.155 -66.475 50.485 ;
        RECT -66.805 48.795 -66.475 49.125 ;
        RECT -66.805 47.435 -66.475 47.765 ;
        RECT -66.805 46.075 -66.475 46.405 ;
        RECT -66.805 44.715 -66.475 45.045 ;
        RECT -66.805 43.355 -66.475 43.685 ;
        RECT -66.805 41.995 -66.475 42.325 ;
        RECT -66.805 40.635 -66.475 40.965 ;
        RECT -66.805 39.275 -66.475 39.605 ;
        RECT -66.805 37.915 -66.475 38.245 ;
        RECT -66.805 36.555 -66.475 36.885 ;
        RECT -66.805 35.195 -66.475 35.525 ;
        RECT -66.805 33.835 -66.475 34.165 ;
        RECT -66.805 32.475 -66.475 32.805 ;
        RECT -66.805 31.115 -66.475 31.445 ;
        RECT -66.805 29.755 -66.475 30.085 ;
        RECT -66.805 28.395 -66.475 28.725 ;
        RECT -66.805 27.035 -66.475 27.365 ;
        RECT -66.805 25.675 -66.475 26.005 ;
        RECT -66.805 24.315 -66.475 24.645 ;
        RECT -66.805 22.955 -66.475 23.285 ;
        RECT -66.805 21.595 -66.475 21.925 ;
        RECT -66.805 20.235 -66.475 20.565 ;
        RECT -66.805 18.875 -66.475 19.205 ;
        RECT -66.805 17.515 -66.475 17.845 ;
        RECT -66.805 16.155 -66.475 16.485 ;
        RECT -66.805 14.795 -66.475 15.125 ;
        RECT -66.805 13.435 -66.475 13.765 ;
        RECT -66.805 12.075 -66.475 12.405 ;
        RECT -66.805 10.715 -66.475 11.045 ;
        RECT -66.805 9.355 -66.475 9.685 ;
        RECT -66.805 7.995 -66.475 8.325 ;
        RECT -66.805 6.635 -66.475 6.965 ;
        RECT -66.805 5.275 -66.475 5.605 ;
        RECT -66.805 3.915 -66.475 4.245 ;
        RECT -66.805 2.555 -66.475 2.885 ;
        RECT -66.805 1.195 -66.475 1.525 ;
        RECT -66.805 -0.165 -66.475 0.165 ;
        RECT -66.805 -1.525 -66.475 -1.195 ;
        RECT -66.805 -2.885 -66.475 -2.555 ;
        RECT -66.805 -4.245 -66.475 -3.915 ;
        RECT -66.805 -5.605 -66.475 -5.275 ;
        RECT -66.805 -6.965 -66.475 -6.635 ;
        RECT -66.805 -8.325 -66.475 -7.995 ;
        RECT -66.805 -9.685 -66.475 -9.355 ;
        RECT -66.805 -11.045 -66.475 -10.715 ;
        RECT -66.805 -12.405 -66.475 -12.075 ;
        RECT -66.805 -13.765 -66.475 -13.435 ;
        RECT -66.805 -15.125 -66.475 -14.795 ;
        RECT -66.805 -16.485 -66.475 -16.155 ;
        RECT -66.805 -17.845 -66.475 -17.515 ;
        RECT -66.805 -19.205 -66.475 -18.875 ;
        RECT -66.805 -20.565 -66.475 -20.235 ;
        RECT -66.805 -21.925 -66.475 -21.595 ;
        RECT -66.805 -23.285 -66.475 -22.955 ;
        RECT -66.805 -24.645 -66.475 -24.315 ;
        RECT -66.805 -26.005 -66.475 -25.675 ;
        RECT -66.805 -27.365 -66.475 -27.035 ;
        RECT -66.805 -28.725 -66.475 -28.395 ;
        RECT -66.805 -30.085 -66.475 -29.755 ;
        RECT -66.805 -31.445 -66.475 -31.115 ;
        RECT -66.805 -32.805 -66.475 -32.475 ;
        RECT -66.805 -34.165 -66.475 -33.835 ;
        RECT -66.805 -35.525 -66.475 -35.195 ;
        RECT -66.805 -36.885 -66.475 -36.555 ;
        RECT -66.805 -38.245 -66.475 -37.915 ;
        RECT -66.805 -39.605 -66.475 -39.275 ;
        RECT -66.805 -40.965 -66.475 -40.635 ;
        RECT -66.805 -42.325 -66.475 -41.995 ;
        RECT -66.805 -43.685 -66.475 -43.355 ;
        RECT -66.805 -45.045 -66.475 -44.715 ;
        RECT -66.805 -46.405 -66.475 -46.075 ;
        RECT -66.805 -47.765 -66.475 -47.435 ;
        RECT -66.805 -49.125 -66.475 -48.795 ;
        RECT -66.805 -50.485 -66.475 -50.155 ;
        RECT -66.805 -51.845 -66.475 -51.515 ;
        RECT -66.805 -53.205 -66.475 -52.875 ;
        RECT -66.805 -54.565 -66.475 -54.235 ;
        RECT -66.805 -55.925 -66.475 -55.595 ;
        RECT -66.805 -57.285 -66.475 -56.955 ;
        RECT -66.805 -58.645 -66.475 -58.315 ;
        RECT -66.805 -60.005 -66.475 -59.675 ;
        RECT -66.805 -61.365 -66.475 -61.035 ;
        RECT -66.805 -62.725 -66.475 -62.395 ;
        RECT -66.805 -64.085 -66.475 -63.755 ;
        RECT -66.805 -65.445 -66.475 -65.115 ;
        RECT -66.805 -66.805 -66.475 -66.475 ;
        RECT -66.805 -68.165 -66.475 -67.835 ;
        RECT -66.805 -69.525 -66.475 -69.195 ;
        RECT -66.805 -70.885 -66.475 -70.555 ;
        RECT -66.805 -72.245 -66.475 -71.915 ;
        RECT -66.805 -73.605 -66.475 -73.275 ;
        RECT -66.805 -74.965 -66.475 -74.635 ;
        RECT -66.805 -76.325 -66.475 -75.995 ;
        RECT -66.805 -77.685 -66.475 -77.355 ;
        RECT -66.805 -79.045 -66.475 -78.715 ;
        RECT -66.805 -80.405 -66.475 -80.075 ;
        RECT -66.805 -81.765 -66.475 -81.435 ;
        RECT -66.805 -83.125 -66.475 -82.795 ;
        RECT -66.805 -84.485 -66.475 -84.155 ;
        RECT -66.805 -85.845 -66.475 -85.515 ;
        RECT -66.805 -87.205 -66.475 -86.875 ;
        RECT -66.805 -88.565 -66.475 -88.235 ;
        RECT -66.805 -89.925 -66.475 -89.595 ;
        RECT -66.805 -91.285 -66.475 -90.955 ;
        RECT -66.805 -92.645 -66.475 -92.315 ;
        RECT -66.805 -94.005 -66.475 -93.675 ;
        RECT -66.805 -95.365 -66.475 -95.035 ;
        RECT -66.805 -96.725 -66.475 -96.395 ;
        RECT -66.805 -98.085 -66.475 -97.755 ;
        RECT -66.805 -99.445 -66.475 -99.115 ;
        RECT -66.805 -100.805 -66.475 -100.475 ;
        RECT -66.805 -102.165 -66.475 -101.835 ;
        RECT -66.805 -103.525 -66.475 -103.195 ;
        RECT -66.805 -104.885 -66.475 -104.555 ;
        RECT -66.805 -106.245 -66.475 -105.915 ;
        RECT -66.805 -107.605 -66.475 -107.275 ;
        RECT -66.805 -108.965 -66.475 -108.635 ;
        RECT -66.805 -110.325 -66.475 -109.995 ;
        RECT -66.805 -111.685 -66.475 -111.355 ;
        RECT -66.805 -113.045 -66.475 -112.715 ;
        RECT -66.805 -114.405 -66.475 -114.075 ;
        RECT -66.805 -115.765 -66.475 -115.435 ;
        RECT -66.805 -117.125 -66.475 -116.795 ;
        RECT -66.805 -118.485 -66.475 -118.155 ;
        RECT -66.805 -119.845 -66.475 -119.515 ;
        RECT -66.805 -121.205 -66.475 -120.875 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.605 246.76 -73.275 247.89 ;
        RECT -73.605 241.915 -73.275 242.245 ;
        RECT -73.605 240.555 -73.275 240.885 ;
        RECT -73.605 239.195 -73.275 239.525 ;
        RECT -73.605 237.835 -73.275 238.165 ;
        RECT -73.605 236.475 -73.275 236.805 ;
        RECT -73.605 235.115 -73.275 235.445 ;
        RECT -73.605 233.755 -73.275 234.085 ;
        RECT -73.605 232.395 -73.275 232.725 ;
        RECT -73.605 231.035 -73.275 231.365 ;
        RECT -73.605 229.675 -73.275 230.005 ;
        RECT -73.605 228.315 -73.275 228.645 ;
        RECT -73.605 226.955 -73.275 227.285 ;
        RECT -73.605 225.595 -73.275 225.925 ;
        RECT -73.605 224.235 -73.275 224.565 ;
        RECT -73.605 222.875 -73.275 223.205 ;
        RECT -73.605 221.515 -73.275 221.845 ;
        RECT -73.605 220.155 -73.275 220.485 ;
        RECT -73.605 218.795 -73.275 219.125 ;
        RECT -73.605 217.435 -73.275 217.765 ;
        RECT -73.605 216.075 -73.275 216.405 ;
        RECT -73.605 214.715 -73.275 215.045 ;
        RECT -73.605 213.355 -73.275 213.685 ;
        RECT -73.605 211.995 -73.275 212.325 ;
        RECT -73.605 210.635 -73.275 210.965 ;
        RECT -73.605 209.275 -73.275 209.605 ;
        RECT -73.605 207.915 -73.275 208.245 ;
        RECT -73.605 206.555 -73.275 206.885 ;
        RECT -73.605 205.195 -73.275 205.525 ;
        RECT -73.605 203.835 -73.275 204.165 ;
        RECT -73.605 202.475 -73.275 202.805 ;
        RECT -73.605 201.115 -73.275 201.445 ;
        RECT -73.605 199.755 -73.275 200.085 ;
        RECT -73.605 198.395 -73.275 198.725 ;
        RECT -73.605 197.035 -73.275 197.365 ;
        RECT -73.605 195.675 -73.275 196.005 ;
        RECT -73.605 194.315 -73.275 194.645 ;
        RECT -73.605 192.955 -73.275 193.285 ;
        RECT -73.605 191.595 -73.275 191.925 ;
        RECT -73.605 190.235 -73.275 190.565 ;
        RECT -73.605 188.875 -73.275 189.205 ;
        RECT -73.605 187.515 -73.275 187.845 ;
        RECT -73.605 186.155 -73.275 186.485 ;
        RECT -73.605 184.795 -73.275 185.125 ;
        RECT -73.605 183.435 -73.275 183.765 ;
        RECT -73.605 182.075 -73.275 182.405 ;
        RECT -73.605 180.715 -73.275 181.045 ;
        RECT -73.605 179.355 -73.275 179.685 ;
        RECT -73.605 177.995 -73.275 178.325 ;
        RECT -73.605 176.635 -73.275 176.965 ;
        RECT -73.605 175.275 -73.275 175.605 ;
        RECT -73.605 173.915 -73.275 174.245 ;
        RECT -73.605 172.555 -73.275 172.885 ;
        RECT -73.605 171.195 -73.275 171.525 ;
        RECT -73.605 169.835 -73.275 170.165 ;
        RECT -73.605 168.475 -73.275 168.805 ;
        RECT -73.605 167.115 -73.275 167.445 ;
        RECT -73.605 165.755 -73.275 166.085 ;
        RECT -73.605 164.395 -73.275 164.725 ;
        RECT -73.605 163.035 -73.275 163.365 ;
        RECT -73.605 161.675 -73.275 162.005 ;
        RECT -73.605 160.315 -73.275 160.645 ;
        RECT -73.605 158.955 -73.275 159.285 ;
        RECT -73.605 157.595 -73.275 157.925 ;
        RECT -73.605 156.235 -73.275 156.565 ;
        RECT -73.605 154.875 -73.275 155.205 ;
        RECT -73.605 153.515 -73.275 153.845 ;
        RECT -73.605 152.155 -73.275 152.485 ;
        RECT -73.605 150.795 -73.275 151.125 ;
        RECT -73.605 149.435 -73.275 149.765 ;
        RECT -73.605 148.075 -73.275 148.405 ;
        RECT -73.605 146.715 -73.275 147.045 ;
        RECT -73.605 145.355 -73.275 145.685 ;
        RECT -73.605 143.995 -73.275 144.325 ;
        RECT -73.605 142.635 -73.275 142.965 ;
        RECT -73.605 141.275 -73.275 141.605 ;
        RECT -73.605 139.915 -73.275 140.245 ;
        RECT -73.605 138.555 -73.275 138.885 ;
        RECT -73.605 137.195 -73.275 137.525 ;
        RECT -73.605 135.835 -73.275 136.165 ;
        RECT -73.605 134.475 -73.275 134.805 ;
        RECT -73.605 133.115 -73.275 133.445 ;
        RECT -73.605 131.755 -73.275 132.085 ;
        RECT -73.605 130.395 -73.275 130.725 ;
        RECT -73.605 129.035 -73.275 129.365 ;
        RECT -73.605 127.675 -73.275 128.005 ;
        RECT -73.605 126.315 -73.275 126.645 ;
        RECT -73.605 124.955 -73.275 125.285 ;
        RECT -73.605 123.595 -73.275 123.925 ;
        RECT -73.605 122.235 -73.275 122.565 ;
        RECT -73.605 120.875 -73.275 121.205 ;
        RECT -73.605 119.515 -73.275 119.845 ;
        RECT -73.605 118.155 -73.275 118.485 ;
        RECT -73.605 116.795 -73.275 117.125 ;
        RECT -73.605 115.435 -73.275 115.765 ;
        RECT -73.605 114.075 -73.275 114.405 ;
        RECT -73.605 112.715 -73.275 113.045 ;
        RECT -73.605 111.355 -73.275 111.685 ;
        RECT -73.605 109.995 -73.275 110.325 ;
        RECT -73.605 108.635 -73.275 108.965 ;
        RECT -73.605 107.275 -73.275 107.605 ;
        RECT -73.605 105.915 -73.275 106.245 ;
        RECT -73.605 104.555 -73.275 104.885 ;
        RECT -73.605 103.195 -73.275 103.525 ;
        RECT -73.605 101.835 -73.275 102.165 ;
        RECT -73.605 100.475 -73.275 100.805 ;
        RECT -73.605 99.115 -73.275 99.445 ;
        RECT -73.605 97.755 -73.275 98.085 ;
        RECT -73.605 96.395 -73.275 96.725 ;
        RECT -73.605 95.035 -73.275 95.365 ;
        RECT -73.605 93.675 -73.275 94.005 ;
        RECT -73.605 92.315 -73.275 92.645 ;
        RECT -73.605 90.955 -73.275 91.285 ;
        RECT -73.605 89.595 -73.275 89.925 ;
        RECT -73.605 88.235 -73.275 88.565 ;
        RECT -73.605 86.875 -73.275 87.205 ;
        RECT -73.605 85.515 -73.275 85.845 ;
        RECT -73.605 84.155 -73.275 84.485 ;
        RECT -73.605 82.795 -73.275 83.125 ;
        RECT -73.605 81.435 -73.275 81.765 ;
        RECT -73.605 80.075 -73.275 80.405 ;
        RECT -73.605 78.715 -73.275 79.045 ;
        RECT -73.605 77.355 -73.275 77.685 ;
        RECT -73.605 75.995 -73.275 76.325 ;
        RECT -73.605 74.635 -73.275 74.965 ;
        RECT -73.605 73.275 -73.275 73.605 ;
        RECT -73.605 71.915 -73.275 72.245 ;
        RECT -73.605 70.555 -73.275 70.885 ;
        RECT -73.605 69.195 -73.275 69.525 ;
        RECT -73.605 67.835 -73.275 68.165 ;
        RECT -73.605 66.475 -73.275 66.805 ;
        RECT -73.605 65.115 -73.275 65.445 ;
        RECT -73.605 63.755 -73.275 64.085 ;
        RECT -73.605 62.395 -73.275 62.725 ;
        RECT -73.605 61.035 -73.275 61.365 ;
        RECT -73.605 59.675 -73.275 60.005 ;
        RECT -73.605 58.315 -73.275 58.645 ;
        RECT -73.605 56.955 -73.275 57.285 ;
        RECT -73.605 55.595 -73.275 55.925 ;
        RECT -73.605 54.235 -73.275 54.565 ;
        RECT -73.605 52.875 -73.275 53.205 ;
        RECT -73.605 51.515 -73.275 51.845 ;
        RECT -73.605 50.155 -73.275 50.485 ;
        RECT -73.605 48.795 -73.275 49.125 ;
        RECT -73.605 47.435 -73.275 47.765 ;
        RECT -73.605 46.075 -73.275 46.405 ;
        RECT -73.605 44.715 -73.275 45.045 ;
        RECT -73.605 43.355 -73.275 43.685 ;
        RECT -73.605 41.995 -73.275 42.325 ;
        RECT -73.605 40.635 -73.275 40.965 ;
        RECT -73.605 39.275 -73.275 39.605 ;
        RECT -73.605 37.915 -73.275 38.245 ;
        RECT -73.605 36.555 -73.275 36.885 ;
        RECT -73.605 35.195 -73.275 35.525 ;
        RECT -73.605 33.835 -73.275 34.165 ;
        RECT -73.605 32.475 -73.275 32.805 ;
        RECT -73.605 31.115 -73.275 31.445 ;
        RECT -73.605 29.755 -73.275 30.085 ;
        RECT -73.605 28.395 -73.275 28.725 ;
        RECT -73.605 27.035 -73.275 27.365 ;
        RECT -73.605 25.675 -73.275 26.005 ;
        RECT -73.605 24.315 -73.275 24.645 ;
        RECT -73.605 22.955 -73.275 23.285 ;
        RECT -73.605 21.595 -73.275 21.925 ;
        RECT -73.605 20.235 -73.275 20.565 ;
        RECT -73.605 18.875 -73.275 19.205 ;
        RECT -73.605 17.515 -73.275 17.845 ;
        RECT -73.605 16.155 -73.275 16.485 ;
        RECT -73.605 14.795 -73.275 15.125 ;
        RECT -73.605 13.435 -73.275 13.765 ;
        RECT -73.605 12.075 -73.275 12.405 ;
        RECT -73.605 10.715 -73.275 11.045 ;
        RECT -73.605 9.355 -73.275 9.685 ;
        RECT -73.605 7.995 -73.275 8.325 ;
        RECT -73.605 6.635 -73.275 6.965 ;
        RECT -73.605 5.275 -73.275 5.605 ;
        RECT -73.605 3.915 -73.275 4.245 ;
        RECT -73.605 2.555 -73.275 2.885 ;
        RECT -73.605 1.195 -73.275 1.525 ;
        RECT -73.605 -0.165 -73.275 0.165 ;
        RECT -73.605 -1.525 -73.275 -1.195 ;
        RECT -73.605 -2.885 -73.275 -2.555 ;
        RECT -73.605 -4.245 -73.275 -3.915 ;
        RECT -73.605 -5.605 -73.275 -5.275 ;
        RECT -73.605 -6.965 -73.275 -6.635 ;
        RECT -73.605 -8.325 -73.275 -7.995 ;
        RECT -73.605 -9.685 -73.275 -9.355 ;
        RECT -73.605 -11.045 -73.275 -10.715 ;
        RECT -73.605 -12.405 -73.275 -12.075 ;
        RECT -73.605 -13.765 -73.275 -13.435 ;
        RECT -73.605 -15.125 -73.275 -14.795 ;
        RECT -73.605 -16.485 -73.275 -16.155 ;
        RECT -73.605 -17.845 -73.275 -17.515 ;
        RECT -73.605 -19.205 -73.275 -18.875 ;
        RECT -73.605 -20.565 -73.275 -20.235 ;
        RECT -73.605 -21.925 -73.275 -21.595 ;
        RECT -73.605 -23.285 -73.275 -22.955 ;
        RECT -73.605 -24.645 -73.275 -24.315 ;
        RECT -73.605 -26.005 -73.275 -25.675 ;
        RECT -73.605 -27.365 -73.275 -27.035 ;
        RECT -73.605 -28.725 -73.275 -28.395 ;
        RECT -73.605 -30.085 -73.275 -29.755 ;
        RECT -73.605 -31.445 -73.275 -31.115 ;
        RECT -73.605 -32.805 -73.275 -32.475 ;
        RECT -73.605 -34.165 -73.275 -33.835 ;
        RECT -73.605 -35.525 -73.275 -35.195 ;
        RECT -73.605 -36.885 -73.275 -36.555 ;
        RECT -73.605 -38.245 -73.275 -37.915 ;
        RECT -73.605 -39.605 -73.275 -39.275 ;
        RECT -73.605 -40.965 -73.275 -40.635 ;
        RECT -73.605 -42.325 -73.275 -41.995 ;
        RECT -73.605 -43.685 -73.275 -43.355 ;
        RECT -73.605 -45.045 -73.275 -44.715 ;
        RECT -73.605 -46.405 -73.275 -46.075 ;
        RECT -73.605 -47.765 -73.275 -47.435 ;
        RECT -73.605 -49.125 -73.275 -48.795 ;
        RECT -73.605 -50.485 -73.275 -50.155 ;
        RECT -73.605 -51.845 -73.275 -51.515 ;
        RECT -73.605 -53.205 -73.275 -52.875 ;
        RECT -73.605 -54.565 -73.275 -54.235 ;
        RECT -73.605 -55.925 -73.275 -55.595 ;
        RECT -73.605 -57.285 -73.275 -56.955 ;
        RECT -73.605 -58.645 -73.275 -58.315 ;
        RECT -73.605 -60.005 -73.275 -59.675 ;
        RECT -73.605 -61.365 -73.275 -61.035 ;
        RECT -73.605 -62.725 -73.275 -62.395 ;
        RECT -73.605 -64.085 -73.275 -63.755 ;
        RECT -73.605 -65.445 -73.275 -65.115 ;
        RECT -73.605 -66.805 -73.275 -66.475 ;
        RECT -73.605 -68.165 -73.275 -67.835 ;
        RECT -73.605 -69.525 -73.275 -69.195 ;
        RECT -73.605 -70.885 -73.275 -70.555 ;
        RECT -73.605 -72.245 -73.275 -71.915 ;
        RECT -73.605 -73.605 -73.275 -73.275 ;
        RECT -73.605 -74.965 -73.275 -74.635 ;
        RECT -73.605 -76.325 -73.275 -75.995 ;
        RECT -73.605 -77.685 -73.275 -77.355 ;
        RECT -73.605 -79.045 -73.275 -78.715 ;
        RECT -73.605 -80.405 -73.275 -80.075 ;
        RECT -73.605 -81.765 -73.275 -81.435 ;
        RECT -73.605 -83.125 -73.275 -82.795 ;
        RECT -73.605 -84.485 -73.275 -84.155 ;
        RECT -73.605 -85.845 -73.275 -85.515 ;
        RECT -73.605 -87.205 -73.275 -86.875 ;
        RECT -73.605 -88.565 -73.275 -88.235 ;
        RECT -73.605 -89.925 -73.275 -89.595 ;
        RECT -73.605 -91.285 -73.275 -90.955 ;
        RECT -73.605 -92.645 -73.275 -92.315 ;
        RECT -73.605 -94.005 -73.275 -93.675 ;
        RECT -73.605 -95.365 -73.275 -95.035 ;
        RECT -73.605 -96.725 -73.275 -96.395 ;
        RECT -73.605 -98.085 -73.275 -97.755 ;
        RECT -73.605 -99.445 -73.275 -99.115 ;
        RECT -73.605 -100.805 -73.275 -100.475 ;
        RECT -73.605 -102.165 -73.275 -101.835 ;
        RECT -73.605 -103.525 -73.275 -103.195 ;
        RECT -73.605 -104.885 -73.275 -104.555 ;
        RECT -73.605 -106.245 -73.275 -105.915 ;
        RECT -73.605 -107.605 -73.275 -107.275 ;
        RECT -73.605 -108.965 -73.275 -108.635 ;
        RECT -73.605 -110.325 -73.275 -109.995 ;
        RECT -73.605 -111.685 -73.275 -111.355 ;
        RECT -73.605 -113.045 -73.275 -112.715 ;
        RECT -73.605 -114.405 -73.275 -114.075 ;
        RECT -73.605 -115.765 -73.275 -115.435 ;
        RECT -73.605 -117.125 -73.275 -116.795 ;
        RECT -73.605 -118.485 -73.275 -118.155 ;
        RECT -73.605 -119.845 -73.275 -119.515 ;
        RECT -73.605 -121.205 -73.275 -120.875 ;
        RECT -73.605 -122.565 -73.275 -122.235 ;
        RECT -73.605 -123.925 -73.275 -123.595 ;
        RECT -73.605 -125.285 -73.275 -124.955 ;
        RECT -73.605 -126.645 -73.275 -126.315 ;
        RECT -73.605 -128.005 -73.275 -127.675 ;
        RECT -73.605 -129.365 -73.275 -129.035 ;
        RECT -73.605 -130.725 -73.275 -130.395 ;
        RECT -73.605 -132.085 -73.275 -131.755 ;
        RECT -73.605 -133.445 -73.275 -133.115 ;
        RECT -73.605 -134.805 -73.275 -134.475 ;
        RECT -73.605 -136.165 -73.275 -135.835 ;
        RECT -73.605 -137.525 -73.275 -137.195 ;
        RECT -73.605 -138.885 -73.275 -138.555 ;
        RECT -73.605 -140.245 -73.275 -139.915 ;
        RECT -73.605 -141.605 -73.275 -141.275 ;
        RECT -73.605 -142.965 -73.275 -142.635 ;
        RECT -73.605 -144.325 -73.275 -143.995 ;
        RECT -73.605 -145.685 -73.275 -145.355 ;
        RECT -73.605 -147.045 -73.275 -146.715 ;
        RECT -73.605 -148.405 -73.275 -148.075 ;
        RECT -73.605 -149.765 -73.275 -149.435 ;
        RECT -73.605 -151.125 -73.275 -150.795 ;
        RECT -73.605 -152.485 -73.275 -152.155 ;
        RECT -73.605 -153.845 -73.275 -153.515 ;
        RECT -73.605 -155.205 -73.275 -154.875 ;
        RECT -73.605 -156.565 -73.275 -156.235 ;
        RECT -73.605 -157.925 -73.275 -157.595 ;
        RECT -73.605 -159.285 -73.275 -158.955 ;
        RECT -73.605 -160.645 -73.275 -160.315 ;
        RECT -73.605 -162.005 -73.275 -161.675 ;
        RECT -73.605 -163.365 -73.275 -163.035 ;
        RECT -73.605 -164.725 -73.275 -164.395 ;
        RECT -73.605 -166.085 -73.275 -165.755 ;
        RECT -73.605 -167.445 -73.275 -167.115 ;
        RECT -73.605 -168.805 -73.275 -168.475 ;
        RECT -73.605 -170.165 -73.275 -169.835 ;
        RECT -73.605 -171.525 -73.275 -171.195 ;
        RECT -73.605 -172.885 -73.275 -172.555 ;
        RECT -73.605 -174.245 -73.275 -173.915 ;
        RECT -73.605 -175.605 -73.275 -175.275 ;
        RECT -73.605 -176.965 -73.275 -176.635 ;
        RECT -73.605 -178.325 -73.275 -177.995 ;
        RECT -73.605 -179.685 -73.275 -179.355 ;
        RECT -73.605 -181.045 -73.275 -180.715 ;
        RECT -73.605 -182.405 -73.275 -182.075 ;
        RECT -73.605 -183.765 -73.275 -183.435 ;
        RECT -73.605 -185.125 -73.275 -184.795 ;
        RECT -73.605 -186.485 -73.275 -186.155 ;
        RECT -73.605 -187.845 -73.275 -187.515 ;
        RECT -73.605 -189.205 -73.275 -188.875 ;
        RECT -73.605 -190.565 -73.275 -190.235 ;
        RECT -73.605 -191.925 -73.275 -191.595 ;
        RECT -73.605 -193.285 -73.275 -192.955 ;
        RECT -73.605 -194.645 -73.275 -194.315 ;
        RECT -73.605 -196.005 -73.275 -195.675 ;
        RECT -73.605 -197.365 -73.275 -197.035 ;
        RECT -73.605 -198.725 -73.275 -198.395 ;
        RECT -73.605 -200.085 -73.275 -199.755 ;
        RECT -73.605 -201.445 -73.275 -201.115 ;
        RECT -73.605 -202.805 -73.275 -202.475 ;
        RECT -73.605 -204.165 -73.275 -203.835 ;
        RECT -73.605 -205.525 -73.275 -205.195 ;
        RECT -73.605 -206.885 -73.275 -206.555 ;
        RECT -73.605 -208.245 -73.275 -207.915 ;
        RECT -73.605 -209.605 -73.275 -209.275 ;
        RECT -73.605 -210.965 -73.275 -210.635 ;
        RECT -73.605 -212.325 -73.275 -211.995 ;
        RECT -73.605 -213.685 -73.275 -213.355 ;
        RECT -73.605 -215.045 -73.275 -214.715 ;
        RECT -73.605 -216.405 -73.275 -216.075 ;
        RECT -73.605 -217.765 -73.275 -217.435 ;
        RECT -73.605 -219.125 -73.275 -218.795 ;
        RECT -73.605 -220.485 -73.275 -220.155 ;
        RECT -73.605 -221.845 -73.275 -221.515 ;
        RECT -73.605 -223.205 -73.275 -222.875 ;
        RECT -73.605 -224.565 -73.275 -224.235 ;
        RECT -73.605 -226.155 -73.275 -225.825 ;
        RECT -73.605 -227.285 -73.275 -226.955 ;
        RECT -73.605 -228.645 -73.275 -228.315 ;
        RECT -73.605 -230.005 -73.275 -229.675 ;
        RECT -73.605 -234.085 -73.275 -233.755 ;
        RECT -73.605 -235.445 -73.275 -235.115 ;
        RECT -73.605 -236.805 -73.275 -236.475 ;
        RECT -73.605 -238.165 -73.275 -237.835 ;
        RECT -73.605 -243.81 -73.275 -242.68 ;
        RECT -73.6 -243.925 -73.28 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.245 246.76 -71.915 247.89 ;
        RECT -72.245 241.915 -71.915 242.245 ;
        RECT -72.245 240.555 -71.915 240.885 ;
        RECT -72.245 239.195 -71.915 239.525 ;
        RECT -72.245 237.835 -71.915 238.165 ;
        RECT -72.245 236.475 -71.915 236.805 ;
        RECT -72.245 235.115 -71.915 235.445 ;
        RECT -72.245 233.755 -71.915 234.085 ;
        RECT -72.245 232.395 -71.915 232.725 ;
        RECT -72.245 231.035 -71.915 231.365 ;
        RECT -72.245 229.675 -71.915 230.005 ;
        RECT -72.245 228.315 -71.915 228.645 ;
        RECT -72.245 226.955 -71.915 227.285 ;
        RECT -72.245 225.595 -71.915 225.925 ;
        RECT -72.245 224.235 -71.915 224.565 ;
        RECT -72.245 222.875 -71.915 223.205 ;
        RECT -72.245 221.515 -71.915 221.845 ;
        RECT -72.245 220.155 -71.915 220.485 ;
        RECT -72.245 218.795 -71.915 219.125 ;
        RECT -72.245 217.435 -71.915 217.765 ;
        RECT -72.245 216.075 -71.915 216.405 ;
        RECT -72.245 214.715 -71.915 215.045 ;
        RECT -72.245 213.355 -71.915 213.685 ;
        RECT -72.245 211.995 -71.915 212.325 ;
        RECT -72.245 210.635 -71.915 210.965 ;
        RECT -72.245 209.275 -71.915 209.605 ;
        RECT -72.245 207.915 -71.915 208.245 ;
        RECT -72.245 206.555 -71.915 206.885 ;
        RECT -72.245 205.195 -71.915 205.525 ;
        RECT -72.245 203.835 -71.915 204.165 ;
        RECT -72.245 202.475 -71.915 202.805 ;
        RECT -72.245 201.115 -71.915 201.445 ;
        RECT -72.245 199.755 -71.915 200.085 ;
        RECT -72.245 198.395 -71.915 198.725 ;
        RECT -72.245 197.035 -71.915 197.365 ;
        RECT -72.245 195.675 -71.915 196.005 ;
        RECT -72.245 194.315 -71.915 194.645 ;
        RECT -72.245 192.955 -71.915 193.285 ;
        RECT -72.245 191.595 -71.915 191.925 ;
        RECT -72.245 190.235 -71.915 190.565 ;
        RECT -72.245 188.875 -71.915 189.205 ;
        RECT -72.245 187.515 -71.915 187.845 ;
        RECT -72.245 186.155 -71.915 186.485 ;
        RECT -72.245 184.795 -71.915 185.125 ;
        RECT -72.245 183.435 -71.915 183.765 ;
        RECT -72.245 182.075 -71.915 182.405 ;
        RECT -72.245 180.715 -71.915 181.045 ;
        RECT -72.245 179.355 -71.915 179.685 ;
        RECT -72.245 177.995 -71.915 178.325 ;
        RECT -72.245 176.635 -71.915 176.965 ;
        RECT -72.245 175.275 -71.915 175.605 ;
        RECT -72.245 173.915 -71.915 174.245 ;
        RECT -72.245 172.555 -71.915 172.885 ;
        RECT -72.245 171.195 -71.915 171.525 ;
        RECT -72.245 169.835 -71.915 170.165 ;
        RECT -72.245 168.475 -71.915 168.805 ;
        RECT -72.245 167.115 -71.915 167.445 ;
        RECT -72.245 165.755 -71.915 166.085 ;
        RECT -72.245 164.395 -71.915 164.725 ;
        RECT -72.245 163.035 -71.915 163.365 ;
        RECT -72.245 161.675 -71.915 162.005 ;
        RECT -72.245 160.315 -71.915 160.645 ;
        RECT -72.245 158.955 -71.915 159.285 ;
        RECT -72.245 157.595 -71.915 157.925 ;
        RECT -72.245 156.235 -71.915 156.565 ;
        RECT -72.245 154.875 -71.915 155.205 ;
        RECT -72.245 153.515 -71.915 153.845 ;
        RECT -72.245 152.155 -71.915 152.485 ;
        RECT -72.245 150.795 -71.915 151.125 ;
        RECT -72.245 149.435 -71.915 149.765 ;
        RECT -72.245 148.075 -71.915 148.405 ;
        RECT -72.245 146.715 -71.915 147.045 ;
        RECT -72.245 145.355 -71.915 145.685 ;
        RECT -72.245 143.995 -71.915 144.325 ;
        RECT -72.245 142.635 -71.915 142.965 ;
        RECT -72.245 141.275 -71.915 141.605 ;
        RECT -72.245 139.915 -71.915 140.245 ;
        RECT -72.245 138.555 -71.915 138.885 ;
        RECT -72.245 137.195 -71.915 137.525 ;
        RECT -72.245 135.835 -71.915 136.165 ;
        RECT -72.245 134.475 -71.915 134.805 ;
        RECT -72.245 133.115 -71.915 133.445 ;
        RECT -72.245 131.755 -71.915 132.085 ;
        RECT -72.245 130.395 -71.915 130.725 ;
        RECT -72.245 129.035 -71.915 129.365 ;
        RECT -72.245 127.675 -71.915 128.005 ;
        RECT -72.245 126.315 -71.915 126.645 ;
        RECT -72.245 124.955 -71.915 125.285 ;
        RECT -72.245 123.595 -71.915 123.925 ;
        RECT -72.245 122.235 -71.915 122.565 ;
        RECT -72.245 120.875 -71.915 121.205 ;
        RECT -72.245 119.515 -71.915 119.845 ;
        RECT -72.245 118.155 -71.915 118.485 ;
        RECT -72.245 116.795 -71.915 117.125 ;
        RECT -72.245 115.435 -71.915 115.765 ;
        RECT -72.245 114.075 -71.915 114.405 ;
        RECT -72.245 112.715 -71.915 113.045 ;
        RECT -72.245 111.355 -71.915 111.685 ;
        RECT -72.245 109.995 -71.915 110.325 ;
        RECT -72.245 108.635 -71.915 108.965 ;
        RECT -72.245 107.275 -71.915 107.605 ;
        RECT -72.245 105.915 -71.915 106.245 ;
        RECT -72.245 104.555 -71.915 104.885 ;
        RECT -72.245 103.195 -71.915 103.525 ;
        RECT -72.245 101.835 -71.915 102.165 ;
        RECT -72.245 100.475 -71.915 100.805 ;
        RECT -72.245 99.115 -71.915 99.445 ;
        RECT -72.245 97.755 -71.915 98.085 ;
        RECT -72.245 96.395 -71.915 96.725 ;
        RECT -72.245 95.035 -71.915 95.365 ;
        RECT -72.245 93.675 -71.915 94.005 ;
        RECT -72.245 92.315 -71.915 92.645 ;
        RECT -72.245 90.955 -71.915 91.285 ;
        RECT -72.245 89.595 -71.915 89.925 ;
        RECT -72.245 88.235 -71.915 88.565 ;
        RECT -72.245 86.875 -71.915 87.205 ;
        RECT -72.245 85.515 -71.915 85.845 ;
        RECT -72.245 84.155 -71.915 84.485 ;
        RECT -72.245 82.795 -71.915 83.125 ;
        RECT -72.245 81.435 -71.915 81.765 ;
        RECT -72.245 80.075 -71.915 80.405 ;
        RECT -72.245 78.715 -71.915 79.045 ;
        RECT -72.245 77.355 -71.915 77.685 ;
        RECT -72.245 75.995 -71.915 76.325 ;
        RECT -72.245 74.635 -71.915 74.965 ;
        RECT -72.245 73.275 -71.915 73.605 ;
        RECT -72.245 71.915 -71.915 72.245 ;
        RECT -72.245 70.555 -71.915 70.885 ;
        RECT -72.245 69.195 -71.915 69.525 ;
        RECT -72.245 67.835 -71.915 68.165 ;
        RECT -72.245 66.475 -71.915 66.805 ;
        RECT -72.245 65.115 -71.915 65.445 ;
        RECT -72.245 63.755 -71.915 64.085 ;
        RECT -72.245 62.395 -71.915 62.725 ;
        RECT -72.245 61.035 -71.915 61.365 ;
        RECT -72.245 59.675 -71.915 60.005 ;
        RECT -72.245 58.315 -71.915 58.645 ;
        RECT -72.245 56.955 -71.915 57.285 ;
        RECT -72.245 55.595 -71.915 55.925 ;
        RECT -72.245 54.235 -71.915 54.565 ;
        RECT -72.245 52.875 -71.915 53.205 ;
        RECT -72.245 51.515 -71.915 51.845 ;
        RECT -72.245 50.155 -71.915 50.485 ;
        RECT -72.245 48.795 -71.915 49.125 ;
        RECT -72.245 47.435 -71.915 47.765 ;
        RECT -72.245 46.075 -71.915 46.405 ;
        RECT -72.245 44.715 -71.915 45.045 ;
        RECT -72.245 43.355 -71.915 43.685 ;
        RECT -72.245 41.995 -71.915 42.325 ;
        RECT -72.245 40.635 -71.915 40.965 ;
        RECT -72.245 39.275 -71.915 39.605 ;
        RECT -72.245 37.915 -71.915 38.245 ;
        RECT -72.245 36.555 -71.915 36.885 ;
        RECT -72.245 35.195 -71.915 35.525 ;
        RECT -72.245 33.835 -71.915 34.165 ;
        RECT -72.245 32.475 -71.915 32.805 ;
        RECT -72.245 31.115 -71.915 31.445 ;
        RECT -72.245 29.755 -71.915 30.085 ;
        RECT -72.245 28.395 -71.915 28.725 ;
        RECT -72.245 27.035 -71.915 27.365 ;
        RECT -72.245 25.675 -71.915 26.005 ;
        RECT -72.245 24.315 -71.915 24.645 ;
        RECT -72.245 22.955 -71.915 23.285 ;
        RECT -72.245 21.595 -71.915 21.925 ;
        RECT -72.245 20.235 -71.915 20.565 ;
        RECT -72.245 18.875 -71.915 19.205 ;
        RECT -72.245 17.515 -71.915 17.845 ;
        RECT -72.245 16.155 -71.915 16.485 ;
        RECT -72.245 14.795 -71.915 15.125 ;
        RECT -72.245 13.435 -71.915 13.765 ;
        RECT -72.245 12.075 -71.915 12.405 ;
        RECT -72.245 10.715 -71.915 11.045 ;
        RECT -72.245 9.355 -71.915 9.685 ;
        RECT -72.245 7.995 -71.915 8.325 ;
        RECT -72.245 6.635 -71.915 6.965 ;
        RECT -72.245 5.275 -71.915 5.605 ;
        RECT -72.245 3.915 -71.915 4.245 ;
        RECT -72.245 2.555 -71.915 2.885 ;
        RECT -72.245 1.195 -71.915 1.525 ;
        RECT -72.245 -0.165 -71.915 0.165 ;
        RECT -72.245 -1.525 -71.915 -1.195 ;
        RECT -72.245 -2.885 -71.915 -2.555 ;
        RECT -72.245 -4.245 -71.915 -3.915 ;
        RECT -72.245 -5.605 -71.915 -5.275 ;
        RECT -72.245 -6.965 -71.915 -6.635 ;
        RECT -72.245 -8.325 -71.915 -7.995 ;
        RECT -72.245 -9.685 -71.915 -9.355 ;
        RECT -72.245 -11.045 -71.915 -10.715 ;
        RECT -72.245 -12.405 -71.915 -12.075 ;
        RECT -72.245 -13.765 -71.915 -13.435 ;
        RECT -72.245 -15.125 -71.915 -14.795 ;
        RECT -72.245 -16.485 -71.915 -16.155 ;
        RECT -72.245 -17.845 -71.915 -17.515 ;
        RECT -72.245 -19.205 -71.915 -18.875 ;
        RECT -72.245 -20.565 -71.915 -20.235 ;
        RECT -72.245 -21.925 -71.915 -21.595 ;
        RECT -72.245 -23.285 -71.915 -22.955 ;
        RECT -72.245 -24.645 -71.915 -24.315 ;
        RECT -72.245 -26.005 -71.915 -25.675 ;
        RECT -72.245 -27.365 -71.915 -27.035 ;
        RECT -72.245 -28.725 -71.915 -28.395 ;
        RECT -72.245 -30.085 -71.915 -29.755 ;
        RECT -72.245 -31.445 -71.915 -31.115 ;
        RECT -72.245 -32.805 -71.915 -32.475 ;
        RECT -72.245 -34.165 -71.915 -33.835 ;
        RECT -72.245 -35.525 -71.915 -35.195 ;
        RECT -72.245 -36.885 -71.915 -36.555 ;
        RECT -72.245 -38.245 -71.915 -37.915 ;
        RECT -72.245 -39.605 -71.915 -39.275 ;
        RECT -72.245 -40.965 -71.915 -40.635 ;
        RECT -72.245 -42.325 -71.915 -41.995 ;
        RECT -72.245 -43.685 -71.915 -43.355 ;
        RECT -72.245 -45.045 -71.915 -44.715 ;
        RECT -72.245 -46.405 -71.915 -46.075 ;
        RECT -72.245 -47.765 -71.915 -47.435 ;
        RECT -72.245 -49.125 -71.915 -48.795 ;
        RECT -72.245 -50.485 -71.915 -50.155 ;
        RECT -72.245 -51.845 -71.915 -51.515 ;
        RECT -72.245 -53.205 -71.915 -52.875 ;
        RECT -72.245 -54.565 -71.915 -54.235 ;
        RECT -72.245 -55.925 -71.915 -55.595 ;
        RECT -72.245 -57.285 -71.915 -56.955 ;
        RECT -72.245 -58.645 -71.915 -58.315 ;
        RECT -72.245 -60.005 -71.915 -59.675 ;
        RECT -72.245 -61.365 -71.915 -61.035 ;
        RECT -72.245 -62.725 -71.915 -62.395 ;
        RECT -72.245 -64.085 -71.915 -63.755 ;
        RECT -72.245 -65.445 -71.915 -65.115 ;
        RECT -72.245 -66.805 -71.915 -66.475 ;
        RECT -72.245 -68.165 -71.915 -67.835 ;
        RECT -72.245 -69.525 -71.915 -69.195 ;
        RECT -72.245 -70.885 -71.915 -70.555 ;
        RECT -72.245 -72.245 -71.915 -71.915 ;
        RECT -72.245 -73.605 -71.915 -73.275 ;
        RECT -72.245 -74.965 -71.915 -74.635 ;
        RECT -72.245 -76.325 -71.915 -75.995 ;
        RECT -72.245 -77.685 -71.915 -77.355 ;
        RECT -72.245 -79.045 -71.915 -78.715 ;
        RECT -72.245 -80.405 -71.915 -80.075 ;
        RECT -72.245 -81.765 -71.915 -81.435 ;
        RECT -72.245 -83.125 -71.915 -82.795 ;
        RECT -72.245 -84.485 -71.915 -84.155 ;
        RECT -72.245 -85.845 -71.915 -85.515 ;
        RECT -72.245 -87.205 -71.915 -86.875 ;
        RECT -72.245 -88.565 -71.915 -88.235 ;
        RECT -72.245 -89.925 -71.915 -89.595 ;
        RECT -72.245 -91.285 -71.915 -90.955 ;
        RECT -72.245 -92.645 -71.915 -92.315 ;
        RECT -72.245 -94.005 -71.915 -93.675 ;
        RECT -72.245 -95.365 -71.915 -95.035 ;
        RECT -72.245 -96.725 -71.915 -96.395 ;
        RECT -72.245 -98.085 -71.915 -97.755 ;
        RECT -72.245 -99.445 -71.915 -99.115 ;
        RECT -72.245 -100.805 -71.915 -100.475 ;
        RECT -72.245 -102.165 -71.915 -101.835 ;
        RECT -72.245 -103.525 -71.915 -103.195 ;
        RECT -72.245 -104.885 -71.915 -104.555 ;
        RECT -72.245 -106.245 -71.915 -105.915 ;
        RECT -72.245 -107.605 -71.915 -107.275 ;
        RECT -72.245 -108.965 -71.915 -108.635 ;
        RECT -72.245 -110.325 -71.915 -109.995 ;
        RECT -72.245 -111.685 -71.915 -111.355 ;
        RECT -72.245 -113.045 -71.915 -112.715 ;
        RECT -72.245 -114.405 -71.915 -114.075 ;
        RECT -72.245 -115.765 -71.915 -115.435 ;
        RECT -72.245 -117.125 -71.915 -116.795 ;
        RECT -72.245 -118.485 -71.915 -118.155 ;
        RECT -72.245 -119.845 -71.915 -119.515 ;
        RECT -72.245 -121.205 -71.915 -120.875 ;
        RECT -72.245 -122.565 -71.915 -122.235 ;
        RECT -72.245 -123.925 -71.915 -123.595 ;
        RECT -72.245 -125.285 -71.915 -124.955 ;
        RECT -72.245 -126.645 -71.915 -126.315 ;
        RECT -72.245 -128.005 -71.915 -127.675 ;
        RECT -72.245 -129.365 -71.915 -129.035 ;
        RECT -72.245 -130.725 -71.915 -130.395 ;
        RECT -72.245 -132.085 -71.915 -131.755 ;
        RECT -72.245 -133.445 -71.915 -133.115 ;
        RECT -72.245 -134.805 -71.915 -134.475 ;
        RECT -72.245 -136.165 -71.915 -135.835 ;
        RECT -72.245 -137.525 -71.915 -137.195 ;
        RECT -72.245 -138.885 -71.915 -138.555 ;
        RECT -72.245 -140.245 -71.915 -139.915 ;
        RECT -72.245 -141.605 -71.915 -141.275 ;
        RECT -72.245 -142.965 -71.915 -142.635 ;
        RECT -72.245 -144.325 -71.915 -143.995 ;
        RECT -72.245 -145.685 -71.915 -145.355 ;
        RECT -72.245 -147.045 -71.915 -146.715 ;
        RECT -72.245 -148.405 -71.915 -148.075 ;
        RECT -72.245 -149.765 -71.915 -149.435 ;
        RECT -72.245 -151.125 -71.915 -150.795 ;
        RECT -72.245 -152.485 -71.915 -152.155 ;
        RECT -72.245 -153.845 -71.915 -153.515 ;
        RECT -72.245 -155.205 -71.915 -154.875 ;
        RECT -72.245 -156.565 -71.915 -156.235 ;
        RECT -72.245 -157.925 -71.915 -157.595 ;
        RECT -72.245 -159.285 -71.915 -158.955 ;
        RECT -72.245 -160.645 -71.915 -160.315 ;
        RECT -72.245 -162.005 -71.915 -161.675 ;
        RECT -72.245 -163.365 -71.915 -163.035 ;
        RECT -72.245 -164.725 -71.915 -164.395 ;
        RECT -72.245 -166.085 -71.915 -165.755 ;
        RECT -72.245 -167.445 -71.915 -167.115 ;
        RECT -72.245 -168.805 -71.915 -168.475 ;
        RECT -72.245 -170.165 -71.915 -169.835 ;
        RECT -72.245 -171.525 -71.915 -171.195 ;
        RECT -72.245 -172.885 -71.915 -172.555 ;
        RECT -72.245 -174.245 -71.915 -173.915 ;
        RECT -72.245 -175.605 -71.915 -175.275 ;
        RECT -72.245 -176.965 -71.915 -176.635 ;
        RECT -72.245 -178.325 -71.915 -177.995 ;
        RECT -72.245 -179.685 -71.915 -179.355 ;
        RECT -72.245 -181.045 -71.915 -180.715 ;
        RECT -72.245 -182.405 -71.915 -182.075 ;
        RECT -72.245 -183.765 -71.915 -183.435 ;
        RECT -72.245 -185.125 -71.915 -184.795 ;
        RECT -72.245 -186.485 -71.915 -186.155 ;
        RECT -72.245 -187.845 -71.915 -187.515 ;
        RECT -72.245 -189.205 -71.915 -188.875 ;
        RECT -72.245 -190.565 -71.915 -190.235 ;
        RECT -72.245 -191.925 -71.915 -191.595 ;
        RECT -72.245 -193.285 -71.915 -192.955 ;
        RECT -72.245 -194.645 -71.915 -194.315 ;
        RECT -72.245 -196.005 -71.915 -195.675 ;
        RECT -72.245 -197.365 -71.915 -197.035 ;
        RECT -72.245 -198.725 -71.915 -198.395 ;
        RECT -72.245 -200.085 -71.915 -199.755 ;
        RECT -72.245 -201.445 -71.915 -201.115 ;
        RECT -72.245 -202.805 -71.915 -202.475 ;
        RECT -72.245 -204.165 -71.915 -203.835 ;
        RECT -72.245 -205.525 -71.915 -205.195 ;
        RECT -72.245 -206.885 -71.915 -206.555 ;
        RECT -72.245 -208.245 -71.915 -207.915 ;
        RECT -72.245 -209.605 -71.915 -209.275 ;
        RECT -72.245 -210.965 -71.915 -210.635 ;
        RECT -72.245 -212.325 -71.915 -211.995 ;
        RECT -72.245 -213.685 -71.915 -213.355 ;
        RECT -72.245 -215.045 -71.915 -214.715 ;
        RECT -72.245 -216.405 -71.915 -216.075 ;
        RECT -72.245 -217.765 -71.915 -217.435 ;
        RECT -72.245 -219.125 -71.915 -218.795 ;
        RECT -72.245 -220.485 -71.915 -220.155 ;
        RECT -72.245 -221.845 -71.915 -221.515 ;
        RECT -72.245 -223.205 -71.915 -222.875 ;
        RECT -72.245 -224.565 -71.915 -224.235 ;
        RECT -72.245 -227.285 -71.915 -226.955 ;
        RECT -72.245 -228.645 -71.915 -228.315 ;
        RECT -72.245 -234.085 -71.915 -233.755 ;
        RECT -72.245 -235.445 -71.915 -235.115 ;
        RECT -72.245 -236.805 -71.915 -236.475 ;
        RECT -72.245 -238.165 -71.915 -237.835 ;
        RECT -72.245 -243.81 -71.915 -242.68 ;
        RECT -72.24 -243.925 -71.92 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.885 -221.845 -70.555 -221.515 ;
        RECT -70.885 -223.205 -70.555 -222.875 ;
        RECT -70.885 -224.565 -70.555 -224.235 ;
        RECT -70.885 -226.155 -70.555 -225.825 ;
        RECT -70.885 -227.285 -70.555 -226.955 ;
        RECT -70.885 -228.645 -70.555 -228.315 ;
        RECT -70.885 -234.085 -70.555 -233.755 ;
        RECT -70.885 -235.445 -70.555 -235.115 ;
        RECT -70.885 -236.805 -70.555 -236.475 ;
        RECT -70.885 -238.165 -70.555 -237.835 ;
        RECT -70.885 -243.81 -70.555 -242.68 ;
        RECT -70.88 -243.925 -70.56 248.005 ;
        RECT -70.885 246.76 -70.555 247.89 ;
        RECT -70.885 241.915 -70.555 242.245 ;
        RECT -70.885 240.555 -70.555 240.885 ;
        RECT -70.885 239.195 -70.555 239.525 ;
        RECT -70.885 237.835 -70.555 238.165 ;
        RECT -70.885 236.475 -70.555 236.805 ;
        RECT -70.885 235.115 -70.555 235.445 ;
        RECT -70.885 233.755 -70.555 234.085 ;
        RECT -70.885 232.395 -70.555 232.725 ;
        RECT -70.885 231.035 -70.555 231.365 ;
        RECT -70.885 229.675 -70.555 230.005 ;
        RECT -70.885 228.315 -70.555 228.645 ;
        RECT -70.885 226.955 -70.555 227.285 ;
        RECT -70.885 225.595 -70.555 225.925 ;
        RECT -70.885 224.235 -70.555 224.565 ;
        RECT -70.885 222.875 -70.555 223.205 ;
        RECT -70.885 221.515 -70.555 221.845 ;
        RECT -70.885 220.155 -70.555 220.485 ;
        RECT -70.885 218.795 -70.555 219.125 ;
        RECT -70.885 217.435 -70.555 217.765 ;
        RECT -70.885 216.075 -70.555 216.405 ;
        RECT -70.885 214.715 -70.555 215.045 ;
        RECT -70.885 213.355 -70.555 213.685 ;
        RECT -70.885 211.995 -70.555 212.325 ;
        RECT -70.885 210.635 -70.555 210.965 ;
        RECT -70.885 209.275 -70.555 209.605 ;
        RECT -70.885 207.915 -70.555 208.245 ;
        RECT -70.885 206.555 -70.555 206.885 ;
        RECT -70.885 205.195 -70.555 205.525 ;
        RECT -70.885 203.835 -70.555 204.165 ;
        RECT -70.885 202.475 -70.555 202.805 ;
        RECT -70.885 201.115 -70.555 201.445 ;
        RECT -70.885 199.755 -70.555 200.085 ;
        RECT -70.885 198.395 -70.555 198.725 ;
        RECT -70.885 197.035 -70.555 197.365 ;
        RECT -70.885 195.675 -70.555 196.005 ;
        RECT -70.885 194.315 -70.555 194.645 ;
        RECT -70.885 192.955 -70.555 193.285 ;
        RECT -70.885 191.595 -70.555 191.925 ;
        RECT -70.885 190.235 -70.555 190.565 ;
        RECT -70.885 188.875 -70.555 189.205 ;
        RECT -70.885 187.515 -70.555 187.845 ;
        RECT -70.885 186.155 -70.555 186.485 ;
        RECT -70.885 184.795 -70.555 185.125 ;
        RECT -70.885 183.435 -70.555 183.765 ;
        RECT -70.885 182.075 -70.555 182.405 ;
        RECT -70.885 180.715 -70.555 181.045 ;
        RECT -70.885 179.355 -70.555 179.685 ;
        RECT -70.885 177.995 -70.555 178.325 ;
        RECT -70.885 176.635 -70.555 176.965 ;
        RECT -70.885 175.275 -70.555 175.605 ;
        RECT -70.885 173.915 -70.555 174.245 ;
        RECT -70.885 172.555 -70.555 172.885 ;
        RECT -70.885 171.195 -70.555 171.525 ;
        RECT -70.885 169.835 -70.555 170.165 ;
        RECT -70.885 168.475 -70.555 168.805 ;
        RECT -70.885 167.115 -70.555 167.445 ;
        RECT -70.885 165.755 -70.555 166.085 ;
        RECT -70.885 164.395 -70.555 164.725 ;
        RECT -70.885 163.035 -70.555 163.365 ;
        RECT -70.885 161.675 -70.555 162.005 ;
        RECT -70.885 160.315 -70.555 160.645 ;
        RECT -70.885 158.955 -70.555 159.285 ;
        RECT -70.885 157.595 -70.555 157.925 ;
        RECT -70.885 156.235 -70.555 156.565 ;
        RECT -70.885 154.875 -70.555 155.205 ;
        RECT -70.885 153.515 -70.555 153.845 ;
        RECT -70.885 152.155 -70.555 152.485 ;
        RECT -70.885 150.795 -70.555 151.125 ;
        RECT -70.885 149.435 -70.555 149.765 ;
        RECT -70.885 148.075 -70.555 148.405 ;
        RECT -70.885 146.715 -70.555 147.045 ;
        RECT -70.885 145.355 -70.555 145.685 ;
        RECT -70.885 143.995 -70.555 144.325 ;
        RECT -70.885 142.635 -70.555 142.965 ;
        RECT -70.885 141.275 -70.555 141.605 ;
        RECT -70.885 139.915 -70.555 140.245 ;
        RECT -70.885 138.555 -70.555 138.885 ;
        RECT -70.885 137.195 -70.555 137.525 ;
        RECT -70.885 135.835 -70.555 136.165 ;
        RECT -70.885 134.475 -70.555 134.805 ;
        RECT -70.885 133.115 -70.555 133.445 ;
        RECT -70.885 131.755 -70.555 132.085 ;
        RECT -70.885 130.395 -70.555 130.725 ;
        RECT -70.885 129.035 -70.555 129.365 ;
        RECT -70.885 127.675 -70.555 128.005 ;
        RECT -70.885 126.315 -70.555 126.645 ;
        RECT -70.885 124.955 -70.555 125.285 ;
        RECT -70.885 123.595 -70.555 123.925 ;
        RECT -70.885 122.235 -70.555 122.565 ;
        RECT -70.885 120.875 -70.555 121.205 ;
        RECT -70.885 119.515 -70.555 119.845 ;
        RECT -70.885 118.155 -70.555 118.485 ;
        RECT -70.885 116.795 -70.555 117.125 ;
        RECT -70.885 115.435 -70.555 115.765 ;
        RECT -70.885 114.075 -70.555 114.405 ;
        RECT -70.885 112.715 -70.555 113.045 ;
        RECT -70.885 111.355 -70.555 111.685 ;
        RECT -70.885 109.995 -70.555 110.325 ;
        RECT -70.885 108.635 -70.555 108.965 ;
        RECT -70.885 107.275 -70.555 107.605 ;
        RECT -70.885 105.915 -70.555 106.245 ;
        RECT -70.885 104.555 -70.555 104.885 ;
        RECT -70.885 103.195 -70.555 103.525 ;
        RECT -70.885 101.835 -70.555 102.165 ;
        RECT -70.885 100.475 -70.555 100.805 ;
        RECT -70.885 99.115 -70.555 99.445 ;
        RECT -70.885 97.755 -70.555 98.085 ;
        RECT -70.885 96.395 -70.555 96.725 ;
        RECT -70.885 95.035 -70.555 95.365 ;
        RECT -70.885 93.675 -70.555 94.005 ;
        RECT -70.885 92.315 -70.555 92.645 ;
        RECT -70.885 90.955 -70.555 91.285 ;
        RECT -70.885 89.595 -70.555 89.925 ;
        RECT -70.885 88.235 -70.555 88.565 ;
        RECT -70.885 86.875 -70.555 87.205 ;
        RECT -70.885 85.515 -70.555 85.845 ;
        RECT -70.885 84.155 -70.555 84.485 ;
        RECT -70.885 82.795 -70.555 83.125 ;
        RECT -70.885 81.435 -70.555 81.765 ;
        RECT -70.885 80.075 -70.555 80.405 ;
        RECT -70.885 78.715 -70.555 79.045 ;
        RECT -70.885 77.355 -70.555 77.685 ;
        RECT -70.885 75.995 -70.555 76.325 ;
        RECT -70.885 74.635 -70.555 74.965 ;
        RECT -70.885 73.275 -70.555 73.605 ;
        RECT -70.885 71.915 -70.555 72.245 ;
        RECT -70.885 70.555 -70.555 70.885 ;
        RECT -70.885 69.195 -70.555 69.525 ;
        RECT -70.885 67.835 -70.555 68.165 ;
        RECT -70.885 66.475 -70.555 66.805 ;
        RECT -70.885 65.115 -70.555 65.445 ;
        RECT -70.885 63.755 -70.555 64.085 ;
        RECT -70.885 62.395 -70.555 62.725 ;
        RECT -70.885 61.035 -70.555 61.365 ;
        RECT -70.885 59.675 -70.555 60.005 ;
        RECT -70.885 58.315 -70.555 58.645 ;
        RECT -70.885 56.955 -70.555 57.285 ;
        RECT -70.885 55.595 -70.555 55.925 ;
        RECT -70.885 54.235 -70.555 54.565 ;
        RECT -70.885 52.875 -70.555 53.205 ;
        RECT -70.885 51.515 -70.555 51.845 ;
        RECT -70.885 50.155 -70.555 50.485 ;
        RECT -70.885 48.795 -70.555 49.125 ;
        RECT -70.885 47.435 -70.555 47.765 ;
        RECT -70.885 46.075 -70.555 46.405 ;
        RECT -70.885 44.715 -70.555 45.045 ;
        RECT -70.885 43.355 -70.555 43.685 ;
        RECT -70.885 41.995 -70.555 42.325 ;
        RECT -70.885 40.635 -70.555 40.965 ;
        RECT -70.885 39.275 -70.555 39.605 ;
        RECT -70.885 37.915 -70.555 38.245 ;
        RECT -70.885 36.555 -70.555 36.885 ;
        RECT -70.885 35.195 -70.555 35.525 ;
        RECT -70.885 33.835 -70.555 34.165 ;
        RECT -70.885 32.475 -70.555 32.805 ;
        RECT -70.885 31.115 -70.555 31.445 ;
        RECT -70.885 29.755 -70.555 30.085 ;
        RECT -70.885 28.395 -70.555 28.725 ;
        RECT -70.885 27.035 -70.555 27.365 ;
        RECT -70.885 25.675 -70.555 26.005 ;
        RECT -70.885 24.315 -70.555 24.645 ;
        RECT -70.885 22.955 -70.555 23.285 ;
        RECT -70.885 21.595 -70.555 21.925 ;
        RECT -70.885 20.235 -70.555 20.565 ;
        RECT -70.885 18.875 -70.555 19.205 ;
        RECT -70.885 17.515 -70.555 17.845 ;
        RECT -70.885 16.155 -70.555 16.485 ;
        RECT -70.885 14.795 -70.555 15.125 ;
        RECT -70.885 13.435 -70.555 13.765 ;
        RECT -70.885 12.075 -70.555 12.405 ;
        RECT -70.885 10.715 -70.555 11.045 ;
        RECT -70.885 9.355 -70.555 9.685 ;
        RECT -70.885 7.995 -70.555 8.325 ;
        RECT -70.885 6.635 -70.555 6.965 ;
        RECT -70.885 5.275 -70.555 5.605 ;
        RECT -70.885 3.915 -70.555 4.245 ;
        RECT -70.885 2.555 -70.555 2.885 ;
        RECT -70.885 1.195 -70.555 1.525 ;
        RECT -70.885 -0.165 -70.555 0.165 ;
        RECT -70.885 -1.525 -70.555 -1.195 ;
        RECT -70.885 -2.885 -70.555 -2.555 ;
        RECT -70.885 -4.245 -70.555 -3.915 ;
        RECT -70.885 -5.605 -70.555 -5.275 ;
        RECT -70.885 -6.965 -70.555 -6.635 ;
        RECT -70.885 -8.325 -70.555 -7.995 ;
        RECT -70.885 -9.685 -70.555 -9.355 ;
        RECT -70.885 -11.045 -70.555 -10.715 ;
        RECT -70.885 -12.405 -70.555 -12.075 ;
        RECT -70.885 -13.765 -70.555 -13.435 ;
        RECT -70.885 -15.125 -70.555 -14.795 ;
        RECT -70.885 -16.485 -70.555 -16.155 ;
        RECT -70.885 -17.845 -70.555 -17.515 ;
        RECT -70.885 -19.205 -70.555 -18.875 ;
        RECT -70.885 -20.565 -70.555 -20.235 ;
        RECT -70.885 -21.925 -70.555 -21.595 ;
        RECT -70.885 -23.285 -70.555 -22.955 ;
        RECT -70.885 -24.645 -70.555 -24.315 ;
        RECT -70.885 -26.005 -70.555 -25.675 ;
        RECT -70.885 -27.365 -70.555 -27.035 ;
        RECT -70.885 -28.725 -70.555 -28.395 ;
        RECT -70.885 -30.085 -70.555 -29.755 ;
        RECT -70.885 -31.445 -70.555 -31.115 ;
        RECT -70.885 -32.805 -70.555 -32.475 ;
        RECT -70.885 -34.165 -70.555 -33.835 ;
        RECT -70.885 -35.525 -70.555 -35.195 ;
        RECT -70.885 -36.885 -70.555 -36.555 ;
        RECT -70.885 -38.245 -70.555 -37.915 ;
        RECT -70.885 -39.605 -70.555 -39.275 ;
        RECT -70.885 -40.965 -70.555 -40.635 ;
        RECT -70.885 -42.325 -70.555 -41.995 ;
        RECT -70.885 -43.685 -70.555 -43.355 ;
        RECT -70.885 -45.045 -70.555 -44.715 ;
        RECT -70.885 -46.405 -70.555 -46.075 ;
        RECT -70.885 -47.765 -70.555 -47.435 ;
        RECT -70.885 -49.125 -70.555 -48.795 ;
        RECT -70.885 -50.485 -70.555 -50.155 ;
        RECT -70.885 -51.845 -70.555 -51.515 ;
        RECT -70.885 -53.205 -70.555 -52.875 ;
        RECT -70.885 -54.565 -70.555 -54.235 ;
        RECT -70.885 -55.925 -70.555 -55.595 ;
        RECT -70.885 -57.285 -70.555 -56.955 ;
        RECT -70.885 -58.645 -70.555 -58.315 ;
        RECT -70.885 -60.005 -70.555 -59.675 ;
        RECT -70.885 -61.365 -70.555 -61.035 ;
        RECT -70.885 -62.725 -70.555 -62.395 ;
        RECT -70.885 -64.085 -70.555 -63.755 ;
        RECT -70.885 -65.445 -70.555 -65.115 ;
        RECT -70.885 -66.805 -70.555 -66.475 ;
        RECT -70.885 -68.165 -70.555 -67.835 ;
        RECT -70.885 -69.525 -70.555 -69.195 ;
        RECT -70.885 -70.885 -70.555 -70.555 ;
        RECT -70.885 -72.245 -70.555 -71.915 ;
        RECT -70.885 -73.605 -70.555 -73.275 ;
        RECT -70.885 -74.965 -70.555 -74.635 ;
        RECT -70.885 -76.325 -70.555 -75.995 ;
        RECT -70.885 -77.685 -70.555 -77.355 ;
        RECT -70.885 -79.045 -70.555 -78.715 ;
        RECT -70.885 -80.405 -70.555 -80.075 ;
        RECT -70.885 -81.765 -70.555 -81.435 ;
        RECT -70.885 -83.125 -70.555 -82.795 ;
        RECT -70.885 -84.485 -70.555 -84.155 ;
        RECT -70.885 -85.845 -70.555 -85.515 ;
        RECT -70.885 -87.205 -70.555 -86.875 ;
        RECT -70.885 -88.565 -70.555 -88.235 ;
        RECT -70.885 -89.925 -70.555 -89.595 ;
        RECT -70.885 -91.285 -70.555 -90.955 ;
        RECT -70.885 -92.645 -70.555 -92.315 ;
        RECT -70.885 -94.005 -70.555 -93.675 ;
        RECT -70.885 -95.365 -70.555 -95.035 ;
        RECT -70.885 -96.725 -70.555 -96.395 ;
        RECT -70.885 -98.085 -70.555 -97.755 ;
        RECT -70.885 -99.445 -70.555 -99.115 ;
        RECT -70.885 -100.805 -70.555 -100.475 ;
        RECT -70.885 -102.165 -70.555 -101.835 ;
        RECT -70.885 -103.525 -70.555 -103.195 ;
        RECT -70.885 -104.885 -70.555 -104.555 ;
        RECT -70.885 -106.245 -70.555 -105.915 ;
        RECT -70.885 -107.605 -70.555 -107.275 ;
        RECT -70.885 -108.965 -70.555 -108.635 ;
        RECT -70.885 -110.325 -70.555 -109.995 ;
        RECT -70.885 -111.685 -70.555 -111.355 ;
        RECT -70.885 -113.045 -70.555 -112.715 ;
        RECT -70.885 -114.405 -70.555 -114.075 ;
        RECT -70.885 -115.765 -70.555 -115.435 ;
        RECT -70.885 -117.125 -70.555 -116.795 ;
        RECT -70.885 -118.485 -70.555 -118.155 ;
        RECT -70.885 -119.845 -70.555 -119.515 ;
        RECT -70.885 -121.205 -70.555 -120.875 ;
        RECT -70.885 -122.565 -70.555 -122.235 ;
        RECT -70.885 -123.925 -70.555 -123.595 ;
        RECT -70.885 -125.285 -70.555 -124.955 ;
        RECT -70.885 -126.645 -70.555 -126.315 ;
        RECT -70.885 -128.005 -70.555 -127.675 ;
        RECT -70.885 -129.365 -70.555 -129.035 ;
        RECT -70.885 -130.725 -70.555 -130.395 ;
        RECT -70.885 -133.445 -70.555 -133.115 ;
        RECT -70.885 -134.805 -70.555 -134.475 ;
        RECT -70.885 -136.165 -70.555 -135.835 ;
        RECT -70.885 -137.525 -70.555 -137.195 ;
        RECT -70.885 -140.245 -70.555 -139.915 ;
        RECT -70.885 -141.605 -70.555 -141.275 ;
        RECT -70.885 -142.965 -70.555 -142.635 ;
        RECT -70.885 -145.685 -70.555 -145.355 ;
        RECT -70.885 -147.045 -70.555 -146.715 ;
        RECT -70.885 -149.765 -70.555 -149.435 ;
        RECT -70.885 -152.485 -70.555 -152.155 ;
        RECT -70.885 -153.845 -70.555 -153.515 ;
        RECT -70.885 -155.205 -70.555 -154.875 ;
        RECT -70.885 -156.565 -70.555 -156.235 ;
        RECT -70.885 -157.925 -70.555 -157.595 ;
        RECT -70.885 -159.285 -70.555 -158.955 ;
        RECT -70.885 -162.005 -70.555 -161.675 ;
        RECT -70.885 -163.365 -70.555 -163.035 ;
        RECT -70.885 -164.725 -70.555 -164.395 ;
        RECT -70.885 -166.085 -70.555 -165.755 ;
        RECT -70.885 -167.445 -70.555 -167.115 ;
        RECT -70.885 -168.805 -70.555 -168.475 ;
        RECT -70.885 -170.165 -70.555 -169.835 ;
        RECT -70.885 -171.525 -70.555 -171.195 ;
        RECT -70.885 -172.885 -70.555 -172.555 ;
        RECT -70.885 -174.245 -70.555 -173.915 ;
        RECT -70.885 -175.605 -70.555 -175.275 ;
        RECT -70.885 -176.965 -70.555 -176.635 ;
        RECT -70.885 -178.325 -70.555 -177.995 ;
        RECT -70.885 -179.685 -70.555 -179.355 ;
        RECT -70.885 -181.045 -70.555 -180.715 ;
        RECT -70.885 -182.405 -70.555 -182.075 ;
        RECT -70.885 -183.765 -70.555 -183.435 ;
        RECT -70.885 -185.125 -70.555 -184.795 ;
        RECT -70.885 -186.485 -70.555 -186.155 ;
        RECT -70.885 -187.845 -70.555 -187.515 ;
        RECT -70.885 -189.205 -70.555 -188.875 ;
        RECT -70.885 -190.565 -70.555 -190.235 ;
        RECT -70.885 -191.925 -70.555 -191.595 ;
        RECT -70.885 -193.285 -70.555 -192.955 ;
        RECT -70.885 -194.645 -70.555 -194.315 ;
        RECT -70.885 -196.005 -70.555 -195.675 ;
        RECT -70.885 -197.365 -70.555 -197.035 ;
        RECT -70.885 -198.725 -70.555 -198.395 ;
        RECT -70.885 -200.085 -70.555 -199.755 ;
        RECT -70.885 -201.445 -70.555 -201.115 ;
        RECT -70.885 -202.805 -70.555 -202.475 ;
        RECT -70.885 -204.165 -70.555 -203.835 ;
        RECT -70.885 -205.525 -70.555 -205.195 ;
        RECT -70.885 -206.885 -70.555 -206.555 ;
        RECT -70.885 -208.245 -70.555 -207.915 ;
        RECT -70.885 -209.605 -70.555 -209.275 ;
        RECT -70.885 -210.965 -70.555 -210.635 ;
        RECT -70.885 -212.325 -70.555 -211.995 ;
        RECT -70.885 -213.685 -70.555 -213.355 ;
        RECT -70.885 -215.045 -70.555 -214.715 ;
        RECT -70.885 -216.405 -70.555 -216.075 ;
        RECT -70.885 -217.765 -70.555 -217.435 ;
        RECT -70.885 -219.125 -70.555 -218.795 ;
        RECT -70.885 -220.485 -70.555 -220.155 ;
    END
    PORT
      LAYER met3 ;
        RECT -77.685 246.76 -77.355 247.89 ;
        RECT -77.685 241.915 -77.355 242.245 ;
        RECT -77.685 240.555 -77.355 240.885 ;
        RECT -77.685 239.195 -77.355 239.525 ;
        RECT -77.685 237.835 -77.355 238.165 ;
        RECT -77.685 236.475 -77.355 236.805 ;
        RECT -77.685 235.115 -77.355 235.445 ;
        RECT -77.685 233.755 -77.355 234.085 ;
        RECT -77.685 232.395 -77.355 232.725 ;
        RECT -77.685 231.035 -77.355 231.365 ;
        RECT -77.685 229.675 -77.355 230.005 ;
        RECT -77.685 228.315 -77.355 228.645 ;
        RECT -77.685 226.955 -77.355 227.285 ;
        RECT -77.685 225.595 -77.355 225.925 ;
        RECT -77.685 224.235 -77.355 224.565 ;
        RECT -77.685 222.875 -77.355 223.205 ;
        RECT -77.685 221.515 -77.355 221.845 ;
        RECT -77.685 220.155 -77.355 220.485 ;
        RECT -77.685 218.795 -77.355 219.125 ;
        RECT -77.685 217.435 -77.355 217.765 ;
        RECT -77.685 216.075 -77.355 216.405 ;
        RECT -77.685 214.715 -77.355 215.045 ;
        RECT -77.685 213.355 -77.355 213.685 ;
        RECT -77.685 211.995 -77.355 212.325 ;
        RECT -77.685 210.635 -77.355 210.965 ;
        RECT -77.685 209.275 -77.355 209.605 ;
        RECT -77.685 207.915 -77.355 208.245 ;
        RECT -77.685 206.555 -77.355 206.885 ;
        RECT -77.685 205.195 -77.355 205.525 ;
        RECT -77.685 203.835 -77.355 204.165 ;
        RECT -77.685 202.475 -77.355 202.805 ;
        RECT -77.685 201.115 -77.355 201.445 ;
        RECT -77.685 199.755 -77.355 200.085 ;
        RECT -77.685 198.395 -77.355 198.725 ;
        RECT -77.685 197.035 -77.355 197.365 ;
        RECT -77.685 195.675 -77.355 196.005 ;
        RECT -77.685 194.315 -77.355 194.645 ;
        RECT -77.685 192.955 -77.355 193.285 ;
        RECT -77.685 191.595 -77.355 191.925 ;
        RECT -77.685 190.235 -77.355 190.565 ;
        RECT -77.685 188.875 -77.355 189.205 ;
        RECT -77.685 187.515 -77.355 187.845 ;
        RECT -77.685 186.155 -77.355 186.485 ;
        RECT -77.685 184.795 -77.355 185.125 ;
        RECT -77.685 183.435 -77.355 183.765 ;
        RECT -77.685 182.075 -77.355 182.405 ;
        RECT -77.685 180.715 -77.355 181.045 ;
        RECT -77.685 179.355 -77.355 179.685 ;
        RECT -77.685 177.995 -77.355 178.325 ;
        RECT -77.685 176.635 -77.355 176.965 ;
        RECT -77.685 175.275 -77.355 175.605 ;
        RECT -77.685 173.915 -77.355 174.245 ;
        RECT -77.685 172.555 -77.355 172.885 ;
        RECT -77.685 171.195 -77.355 171.525 ;
        RECT -77.685 169.835 -77.355 170.165 ;
        RECT -77.685 168.475 -77.355 168.805 ;
        RECT -77.685 167.115 -77.355 167.445 ;
        RECT -77.685 165.755 -77.355 166.085 ;
        RECT -77.685 164.395 -77.355 164.725 ;
        RECT -77.685 163.035 -77.355 163.365 ;
        RECT -77.685 161.675 -77.355 162.005 ;
        RECT -77.685 160.315 -77.355 160.645 ;
        RECT -77.685 158.955 -77.355 159.285 ;
        RECT -77.685 157.595 -77.355 157.925 ;
        RECT -77.685 156.235 -77.355 156.565 ;
        RECT -77.685 154.875 -77.355 155.205 ;
        RECT -77.685 153.515 -77.355 153.845 ;
        RECT -77.685 152.155 -77.355 152.485 ;
        RECT -77.685 150.795 -77.355 151.125 ;
        RECT -77.685 149.435 -77.355 149.765 ;
        RECT -77.685 148.075 -77.355 148.405 ;
        RECT -77.685 146.715 -77.355 147.045 ;
        RECT -77.685 145.355 -77.355 145.685 ;
        RECT -77.685 143.995 -77.355 144.325 ;
        RECT -77.685 142.635 -77.355 142.965 ;
        RECT -77.685 141.275 -77.355 141.605 ;
        RECT -77.685 139.915 -77.355 140.245 ;
        RECT -77.685 138.555 -77.355 138.885 ;
        RECT -77.685 137.195 -77.355 137.525 ;
        RECT -77.685 135.835 -77.355 136.165 ;
        RECT -77.685 134.475 -77.355 134.805 ;
        RECT -77.685 133.115 -77.355 133.445 ;
        RECT -77.685 131.755 -77.355 132.085 ;
        RECT -77.685 130.395 -77.355 130.725 ;
        RECT -77.685 129.035 -77.355 129.365 ;
        RECT -77.685 127.675 -77.355 128.005 ;
        RECT -77.685 126.315 -77.355 126.645 ;
        RECT -77.685 124.955 -77.355 125.285 ;
        RECT -77.685 123.595 -77.355 123.925 ;
        RECT -77.685 122.235 -77.355 122.565 ;
        RECT -77.685 120.875 -77.355 121.205 ;
        RECT -77.685 119.515 -77.355 119.845 ;
        RECT -77.685 118.155 -77.355 118.485 ;
        RECT -77.685 116.795 -77.355 117.125 ;
        RECT -77.685 115.435 -77.355 115.765 ;
        RECT -77.685 114.075 -77.355 114.405 ;
        RECT -77.685 112.715 -77.355 113.045 ;
        RECT -77.685 111.355 -77.355 111.685 ;
        RECT -77.685 109.995 -77.355 110.325 ;
        RECT -77.685 108.635 -77.355 108.965 ;
        RECT -77.685 107.275 -77.355 107.605 ;
        RECT -77.685 105.915 -77.355 106.245 ;
        RECT -77.685 104.555 -77.355 104.885 ;
        RECT -77.685 103.195 -77.355 103.525 ;
        RECT -77.685 101.835 -77.355 102.165 ;
        RECT -77.685 100.475 -77.355 100.805 ;
        RECT -77.685 99.115 -77.355 99.445 ;
        RECT -77.685 97.755 -77.355 98.085 ;
        RECT -77.685 96.395 -77.355 96.725 ;
        RECT -77.685 95.035 -77.355 95.365 ;
        RECT -77.685 93.675 -77.355 94.005 ;
        RECT -77.685 92.315 -77.355 92.645 ;
        RECT -77.685 90.955 -77.355 91.285 ;
        RECT -77.685 89.595 -77.355 89.925 ;
        RECT -77.685 88.235 -77.355 88.565 ;
        RECT -77.685 86.875 -77.355 87.205 ;
        RECT -77.685 85.515 -77.355 85.845 ;
        RECT -77.685 84.155 -77.355 84.485 ;
        RECT -77.685 82.795 -77.355 83.125 ;
        RECT -77.685 81.435 -77.355 81.765 ;
        RECT -77.685 80.075 -77.355 80.405 ;
        RECT -77.685 78.715 -77.355 79.045 ;
        RECT -77.685 77.355 -77.355 77.685 ;
        RECT -77.685 75.995 -77.355 76.325 ;
        RECT -77.685 74.635 -77.355 74.965 ;
        RECT -77.685 73.275 -77.355 73.605 ;
        RECT -77.685 71.915 -77.355 72.245 ;
        RECT -77.685 70.555 -77.355 70.885 ;
        RECT -77.685 69.195 -77.355 69.525 ;
        RECT -77.685 67.835 -77.355 68.165 ;
        RECT -77.685 66.475 -77.355 66.805 ;
        RECT -77.685 65.115 -77.355 65.445 ;
        RECT -77.685 63.755 -77.355 64.085 ;
        RECT -77.685 62.395 -77.355 62.725 ;
        RECT -77.685 61.035 -77.355 61.365 ;
        RECT -77.685 59.675 -77.355 60.005 ;
        RECT -77.685 58.315 -77.355 58.645 ;
        RECT -77.685 56.955 -77.355 57.285 ;
        RECT -77.685 55.595 -77.355 55.925 ;
        RECT -77.685 54.235 -77.355 54.565 ;
        RECT -77.685 52.875 -77.355 53.205 ;
        RECT -77.685 51.515 -77.355 51.845 ;
        RECT -77.685 50.155 -77.355 50.485 ;
        RECT -77.685 48.795 -77.355 49.125 ;
        RECT -77.685 47.435 -77.355 47.765 ;
        RECT -77.685 46.075 -77.355 46.405 ;
        RECT -77.685 44.715 -77.355 45.045 ;
        RECT -77.685 43.355 -77.355 43.685 ;
        RECT -77.685 41.995 -77.355 42.325 ;
        RECT -77.685 40.635 -77.355 40.965 ;
        RECT -77.685 39.275 -77.355 39.605 ;
        RECT -77.685 37.915 -77.355 38.245 ;
        RECT -77.685 36.555 -77.355 36.885 ;
        RECT -77.685 35.195 -77.355 35.525 ;
        RECT -77.685 33.835 -77.355 34.165 ;
        RECT -77.685 32.475 -77.355 32.805 ;
        RECT -77.685 31.115 -77.355 31.445 ;
        RECT -77.685 29.755 -77.355 30.085 ;
        RECT -77.685 28.395 -77.355 28.725 ;
        RECT -77.685 27.035 -77.355 27.365 ;
        RECT -77.685 25.675 -77.355 26.005 ;
        RECT -77.685 24.315 -77.355 24.645 ;
        RECT -77.685 22.955 -77.355 23.285 ;
        RECT -77.685 21.595 -77.355 21.925 ;
        RECT -77.685 20.235 -77.355 20.565 ;
        RECT -77.685 18.875 -77.355 19.205 ;
        RECT -77.685 17.515 -77.355 17.845 ;
        RECT -77.685 16.155 -77.355 16.485 ;
        RECT -77.685 14.795 -77.355 15.125 ;
        RECT -77.685 13.435 -77.355 13.765 ;
        RECT -77.685 12.075 -77.355 12.405 ;
        RECT -77.685 10.715 -77.355 11.045 ;
        RECT -77.685 9.355 -77.355 9.685 ;
        RECT -77.685 7.995 -77.355 8.325 ;
        RECT -77.685 6.635 -77.355 6.965 ;
        RECT -77.685 5.275 -77.355 5.605 ;
        RECT -77.685 3.915 -77.355 4.245 ;
        RECT -77.685 2.555 -77.355 2.885 ;
        RECT -77.685 1.195 -77.355 1.525 ;
        RECT -77.685 -0.165 -77.355 0.165 ;
        RECT -77.685 -1.525 -77.355 -1.195 ;
        RECT -77.685 -2.885 -77.355 -2.555 ;
        RECT -77.685 -4.245 -77.355 -3.915 ;
        RECT -77.685 -5.605 -77.355 -5.275 ;
        RECT -77.685 -6.965 -77.355 -6.635 ;
        RECT -77.685 -8.325 -77.355 -7.995 ;
        RECT -77.685 -9.685 -77.355 -9.355 ;
        RECT -77.685 -11.045 -77.355 -10.715 ;
        RECT -77.685 -12.405 -77.355 -12.075 ;
        RECT -77.685 -13.765 -77.355 -13.435 ;
        RECT -77.685 -15.125 -77.355 -14.795 ;
        RECT -77.685 -16.485 -77.355 -16.155 ;
        RECT -77.685 -17.845 -77.355 -17.515 ;
        RECT -77.685 -19.205 -77.355 -18.875 ;
        RECT -77.685 -20.565 -77.355 -20.235 ;
        RECT -77.685 -21.925 -77.355 -21.595 ;
        RECT -77.685 -23.285 -77.355 -22.955 ;
        RECT -77.685 -24.645 -77.355 -24.315 ;
        RECT -77.685 -26.005 -77.355 -25.675 ;
        RECT -77.685 -27.365 -77.355 -27.035 ;
        RECT -77.685 -28.725 -77.355 -28.395 ;
        RECT -77.685 -30.085 -77.355 -29.755 ;
        RECT -77.685 -31.445 -77.355 -31.115 ;
        RECT -77.685 -32.805 -77.355 -32.475 ;
        RECT -77.685 -34.165 -77.355 -33.835 ;
        RECT -77.685 -35.525 -77.355 -35.195 ;
        RECT -77.685 -36.885 -77.355 -36.555 ;
        RECT -77.685 -38.245 -77.355 -37.915 ;
        RECT -77.685 -39.605 -77.355 -39.275 ;
        RECT -77.685 -40.965 -77.355 -40.635 ;
        RECT -77.685 -42.325 -77.355 -41.995 ;
        RECT -77.685 -43.685 -77.355 -43.355 ;
        RECT -77.685 -45.045 -77.355 -44.715 ;
        RECT -77.685 -46.405 -77.355 -46.075 ;
        RECT -77.685 -47.765 -77.355 -47.435 ;
        RECT -77.685 -49.125 -77.355 -48.795 ;
        RECT -77.685 -50.485 -77.355 -50.155 ;
        RECT -77.685 -51.845 -77.355 -51.515 ;
        RECT -77.685 -53.205 -77.355 -52.875 ;
        RECT -77.685 -54.565 -77.355 -54.235 ;
        RECT -77.685 -55.925 -77.355 -55.595 ;
        RECT -77.685 -57.285 -77.355 -56.955 ;
        RECT -77.685 -58.645 -77.355 -58.315 ;
        RECT -77.685 -60.005 -77.355 -59.675 ;
        RECT -77.685 -61.365 -77.355 -61.035 ;
        RECT -77.685 -62.725 -77.355 -62.395 ;
        RECT -77.685 -64.085 -77.355 -63.755 ;
        RECT -77.685 -65.445 -77.355 -65.115 ;
        RECT -77.685 -66.805 -77.355 -66.475 ;
        RECT -77.685 -68.165 -77.355 -67.835 ;
        RECT -77.685 -69.525 -77.355 -69.195 ;
        RECT -77.685 -70.885 -77.355 -70.555 ;
        RECT -77.685 -72.245 -77.355 -71.915 ;
        RECT -77.685 -73.605 -77.355 -73.275 ;
        RECT -77.685 -74.965 -77.355 -74.635 ;
        RECT -77.685 -76.325 -77.355 -75.995 ;
        RECT -77.685 -77.685 -77.355 -77.355 ;
        RECT -77.685 -79.045 -77.355 -78.715 ;
        RECT -77.685 -80.405 -77.355 -80.075 ;
        RECT -77.685 -81.765 -77.355 -81.435 ;
        RECT -77.685 -83.125 -77.355 -82.795 ;
        RECT -77.685 -84.485 -77.355 -84.155 ;
        RECT -77.685 -85.845 -77.355 -85.515 ;
        RECT -77.685 -87.205 -77.355 -86.875 ;
        RECT -77.685 -88.565 -77.355 -88.235 ;
        RECT -77.685 -89.925 -77.355 -89.595 ;
        RECT -77.685 -91.285 -77.355 -90.955 ;
        RECT -77.685 -92.645 -77.355 -92.315 ;
        RECT -77.685 -94.005 -77.355 -93.675 ;
        RECT -77.685 -95.365 -77.355 -95.035 ;
        RECT -77.685 -96.725 -77.355 -96.395 ;
        RECT -77.685 -98.085 -77.355 -97.755 ;
        RECT -77.685 -99.445 -77.355 -99.115 ;
        RECT -77.685 -100.805 -77.355 -100.475 ;
        RECT -77.685 -102.165 -77.355 -101.835 ;
        RECT -77.685 -103.525 -77.355 -103.195 ;
        RECT -77.685 -104.885 -77.355 -104.555 ;
        RECT -77.685 -106.245 -77.355 -105.915 ;
        RECT -77.685 -107.605 -77.355 -107.275 ;
        RECT -77.685 -108.965 -77.355 -108.635 ;
        RECT -77.685 -110.325 -77.355 -109.995 ;
        RECT -77.685 -111.685 -77.355 -111.355 ;
        RECT -77.685 -113.045 -77.355 -112.715 ;
        RECT -77.685 -114.405 -77.355 -114.075 ;
        RECT -77.685 -115.765 -77.355 -115.435 ;
        RECT -77.685 -117.125 -77.355 -116.795 ;
        RECT -77.685 -118.485 -77.355 -118.155 ;
        RECT -77.685 -119.845 -77.355 -119.515 ;
        RECT -77.685 -121.205 -77.355 -120.875 ;
        RECT -77.685 -122.565 -77.355 -122.235 ;
        RECT -77.685 -123.925 -77.355 -123.595 ;
        RECT -77.685 -125.285 -77.355 -124.955 ;
        RECT -77.685 -126.645 -77.355 -126.315 ;
        RECT -77.685 -128.005 -77.355 -127.675 ;
        RECT -77.685 -129.365 -77.355 -129.035 ;
        RECT -77.685 -130.725 -77.355 -130.395 ;
        RECT -77.685 -132.085 -77.355 -131.755 ;
        RECT -77.685 -133.445 -77.355 -133.115 ;
        RECT -77.685 -134.805 -77.355 -134.475 ;
        RECT -77.685 -136.165 -77.355 -135.835 ;
        RECT -77.685 -137.525 -77.355 -137.195 ;
        RECT -77.685 -138.885 -77.355 -138.555 ;
        RECT -77.685 -140.245 -77.355 -139.915 ;
        RECT -77.685 -141.605 -77.355 -141.275 ;
        RECT -77.685 -142.965 -77.355 -142.635 ;
        RECT -77.685 -144.325 -77.355 -143.995 ;
        RECT -77.685 -145.685 -77.355 -145.355 ;
        RECT -77.685 -147.045 -77.355 -146.715 ;
        RECT -77.685 -148.405 -77.355 -148.075 ;
        RECT -77.685 -149.765 -77.355 -149.435 ;
        RECT -77.685 -151.125 -77.355 -150.795 ;
        RECT -77.685 -152.485 -77.355 -152.155 ;
        RECT -77.685 -153.845 -77.355 -153.515 ;
        RECT -77.685 -155.205 -77.355 -154.875 ;
        RECT -77.685 -156.565 -77.355 -156.235 ;
        RECT -77.685 -157.925 -77.355 -157.595 ;
        RECT -77.685 -159.285 -77.355 -158.955 ;
        RECT -77.685 -160.645 -77.355 -160.315 ;
        RECT -77.685 -162.005 -77.355 -161.675 ;
        RECT -77.685 -163.365 -77.355 -163.035 ;
        RECT -77.685 -164.725 -77.355 -164.395 ;
        RECT -77.685 -166.085 -77.355 -165.755 ;
        RECT -77.685 -167.445 -77.355 -167.115 ;
        RECT -77.685 -168.805 -77.355 -168.475 ;
        RECT -77.685 -170.165 -77.355 -169.835 ;
        RECT -77.685 -171.525 -77.355 -171.195 ;
        RECT -77.685 -172.885 -77.355 -172.555 ;
        RECT -77.685 -174.245 -77.355 -173.915 ;
        RECT -77.685 -175.605 -77.355 -175.275 ;
        RECT -77.685 -176.965 -77.355 -176.635 ;
        RECT -77.685 -178.325 -77.355 -177.995 ;
        RECT -77.685 -179.685 -77.355 -179.355 ;
        RECT -77.685 -181.045 -77.355 -180.715 ;
        RECT -77.685 -182.405 -77.355 -182.075 ;
        RECT -77.685 -183.765 -77.355 -183.435 ;
        RECT -77.685 -185.125 -77.355 -184.795 ;
        RECT -77.685 -186.485 -77.355 -186.155 ;
        RECT -77.685 -187.845 -77.355 -187.515 ;
        RECT -77.685 -189.205 -77.355 -188.875 ;
        RECT -77.685 -190.565 -77.355 -190.235 ;
        RECT -77.685 -191.925 -77.355 -191.595 ;
        RECT -77.685 -193.285 -77.355 -192.955 ;
        RECT -77.685 -194.645 -77.355 -194.315 ;
        RECT -77.685 -196.005 -77.355 -195.675 ;
        RECT -77.685 -197.365 -77.355 -197.035 ;
        RECT -77.685 -198.725 -77.355 -198.395 ;
        RECT -77.685 -200.085 -77.355 -199.755 ;
        RECT -77.685 -201.445 -77.355 -201.115 ;
        RECT -77.685 -202.805 -77.355 -202.475 ;
        RECT -77.685 -204.165 -77.355 -203.835 ;
        RECT -77.685 -205.525 -77.355 -205.195 ;
        RECT -77.685 -206.885 -77.355 -206.555 ;
        RECT -77.685 -208.245 -77.355 -207.915 ;
        RECT -77.685 -209.605 -77.355 -209.275 ;
        RECT -77.685 -210.965 -77.355 -210.635 ;
        RECT -77.685 -212.325 -77.355 -211.995 ;
        RECT -77.685 -213.685 -77.355 -213.355 ;
        RECT -77.685 -215.045 -77.355 -214.715 ;
        RECT -77.685 -216.405 -77.355 -216.075 ;
        RECT -77.685 -217.765 -77.355 -217.435 ;
        RECT -77.685 -219.125 -77.355 -218.795 ;
        RECT -77.685 -220.485 -77.355 -220.155 ;
        RECT -77.685 -221.845 -77.355 -221.515 ;
        RECT -77.685 -223.205 -77.355 -222.875 ;
        RECT -77.685 -224.565 -77.355 -224.235 ;
        RECT -77.685 -226.155 -77.355 -225.825 ;
        RECT -77.685 -227.285 -77.355 -226.955 ;
        RECT -77.685 -228.645 -77.355 -228.315 ;
        RECT -77.68 -229.32 -77.36 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -76.325 246.76 -75.995 247.89 ;
        RECT -76.325 241.915 -75.995 242.245 ;
        RECT -76.325 240.555 -75.995 240.885 ;
        RECT -76.325 239.195 -75.995 239.525 ;
        RECT -76.325 237.835 -75.995 238.165 ;
        RECT -76.325 236.475 -75.995 236.805 ;
        RECT -76.325 235.115 -75.995 235.445 ;
        RECT -76.325 233.755 -75.995 234.085 ;
        RECT -76.325 232.395 -75.995 232.725 ;
        RECT -76.325 231.035 -75.995 231.365 ;
        RECT -76.325 229.675 -75.995 230.005 ;
        RECT -76.325 228.315 -75.995 228.645 ;
        RECT -76.325 226.955 -75.995 227.285 ;
        RECT -76.325 225.595 -75.995 225.925 ;
        RECT -76.325 224.235 -75.995 224.565 ;
        RECT -76.325 222.875 -75.995 223.205 ;
        RECT -76.325 221.515 -75.995 221.845 ;
        RECT -76.325 220.155 -75.995 220.485 ;
        RECT -76.325 218.795 -75.995 219.125 ;
        RECT -76.325 217.435 -75.995 217.765 ;
        RECT -76.325 216.075 -75.995 216.405 ;
        RECT -76.325 214.715 -75.995 215.045 ;
        RECT -76.325 213.355 -75.995 213.685 ;
        RECT -76.325 211.995 -75.995 212.325 ;
        RECT -76.325 210.635 -75.995 210.965 ;
        RECT -76.325 209.275 -75.995 209.605 ;
        RECT -76.325 207.915 -75.995 208.245 ;
        RECT -76.325 206.555 -75.995 206.885 ;
        RECT -76.325 205.195 -75.995 205.525 ;
        RECT -76.325 203.835 -75.995 204.165 ;
        RECT -76.325 202.475 -75.995 202.805 ;
        RECT -76.325 201.115 -75.995 201.445 ;
        RECT -76.325 199.755 -75.995 200.085 ;
        RECT -76.325 198.395 -75.995 198.725 ;
        RECT -76.325 197.035 -75.995 197.365 ;
        RECT -76.325 195.675 -75.995 196.005 ;
        RECT -76.325 194.315 -75.995 194.645 ;
        RECT -76.325 192.955 -75.995 193.285 ;
        RECT -76.325 191.595 -75.995 191.925 ;
        RECT -76.325 190.235 -75.995 190.565 ;
        RECT -76.325 188.875 -75.995 189.205 ;
        RECT -76.325 187.515 -75.995 187.845 ;
        RECT -76.325 186.155 -75.995 186.485 ;
        RECT -76.325 184.795 -75.995 185.125 ;
        RECT -76.325 183.435 -75.995 183.765 ;
        RECT -76.325 182.075 -75.995 182.405 ;
        RECT -76.325 180.715 -75.995 181.045 ;
        RECT -76.325 179.355 -75.995 179.685 ;
        RECT -76.325 177.995 -75.995 178.325 ;
        RECT -76.325 176.635 -75.995 176.965 ;
        RECT -76.325 175.275 -75.995 175.605 ;
        RECT -76.325 173.915 -75.995 174.245 ;
        RECT -76.325 172.555 -75.995 172.885 ;
        RECT -76.325 171.195 -75.995 171.525 ;
        RECT -76.325 169.835 -75.995 170.165 ;
        RECT -76.325 168.475 -75.995 168.805 ;
        RECT -76.325 167.115 -75.995 167.445 ;
        RECT -76.325 165.755 -75.995 166.085 ;
        RECT -76.325 164.395 -75.995 164.725 ;
        RECT -76.325 163.035 -75.995 163.365 ;
        RECT -76.325 161.675 -75.995 162.005 ;
        RECT -76.325 160.315 -75.995 160.645 ;
        RECT -76.325 158.955 -75.995 159.285 ;
        RECT -76.325 157.595 -75.995 157.925 ;
        RECT -76.325 156.235 -75.995 156.565 ;
        RECT -76.325 154.875 -75.995 155.205 ;
        RECT -76.325 153.515 -75.995 153.845 ;
        RECT -76.325 152.155 -75.995 152.485 ;
        RECT -76.325 150.795 -75.995 151.125 ;
        RECT -76.325 149.435 -75.995 149.765 ;
        RECT -76.325 148.075 -75.995 148.405 ;
        RECT -76.325 146.715 -75.995 147.045 ;
        RECT -76.325 145.355 -75.995 145.685 ;
        RECT -76.325 143.995 -75.995 144.325 ;
        RECT -76.325 142.635 -75.995 142.965 ;
        RECT -76.325 141.275 -75.995 141.605 ;
        RECT -76.325 139.915 -75.995 140.245 ;
        RECT -76.325 138.555 -75.995 138.885 ;
        RECT -76.325 137.195 -75.995 137.525 ;
        RECT -76.325 135.835 -75.995 136.165 ;
        RECT -76.325 134.475 -75.995 134.805 ;
        RECT -76.325 133.115 -75.995 133.445 ;
        RECT -76.325 131.755 -75.995 132.085 ;
        RECT -76.325 130.395 -75.995 130.725 ;
        RECT -76.325 129.035 -75.995 129.365 ;
        RECT -76.325 127.675 -75.995 128.005 ;
        RECT -76.325 126.315 -75.995 126.645 ;
        RECT -76.325 124.955 -75.995 125.285 ;
        RECT -76.325 123.595 -75.995 123.925 ;
        RECT -76.325 122.235 -75.995 122.565 ;
        RECT -76.325 120.875 -75.995 121.205 ;
        RECT -76.325 119.515 -75.995 119.845 ;
        RECT -76.325 118.155 -75.995 118.485 ;
        RECT -76.325 116.795 -75.995 117.125 ;
        RECT -76.325 115.435 -75.995 115.765 ;
        RECT -76.325 114.075 -75.995 114.405 ;
        RECT -76.325 112.715 -75.995 113.045 ;
        RECT -76.325 111.355 -75.995 111.685 ;
        RECT -76.325 109.995 -75.995 110.325 ;
        RECT -76.325 108.635 -75.995 108.965 ;
        RECT -76.325 107.275 -75.995 107.605 ;
        RECT -76.325 105.915 -75.995 106.245 ;
        RECT -76.325 104.555 -75.995 104.885 ;
        RECT -76.325 103.195 -75.995 103.525 ;
        RECT -76.325 101.835 -75.995 102.165 ;
        RECT -76.325 100.475 -75.995 100.805 ;
        RECT -76.325 99.115 -75.995 99.445 ;
        RECT -76.325 97.755 -75.995 98.085 ;
        RECT -76.325 96.395 -75.995 96.725 ;
        RECT -76.325 95.035 -75.995 95.365 ;
        RECT -76.325 93.675 -75.995 94.005 ;
        RECT -76.325 92.315 -75.995 92.645 ;
        RECT -76.325 90.955 -75.995 91.285 ;
        RECT -76.325 89.595 -75.995 89.925 ;
        RECT -76.325 88.235 -75.995 88.565 ;
        RECT -76.325 86.875 -75.995 87.205 ;
        RECT -76.325 85.515 -75.995 85.845 ;
        RECT -76.325 84.155 -75.995 84.485 ;
        RECT -76.325 82.795 -75.995 83.125 ;
        RECT -76.325 81.435 -75.995 81.765 ;
        RECT -76.325 80.075 -75.995 80.405 ;
        RECT -76.325 78.715 -75.995 79.045 ;
        RECT -76.325 77.355 -75.995 77.685 ;
        RECT -76.325 75.995 -75.995 76.325 ;
        RECT -76.325 74.635 -75.995 74.965 ;
        RECT -76.325 73.275 -75.995 73.605 ;
        RECT -76.325 71.915 -75.995 72.245 ;
        RECT -76.325 70.555 -75.995 70.885 ;
        RECT -76.325 69.195 -75.995 69.525 ;
        RECT -76.325 67.835 -75.995 68.165 ;
        RECT -76.325 66.475 -75.995 66.805 ;
        RECT -76.325 65.115 -75.995 65.445 ;
        RECT -76.325 63.755 -75.995 64.085 ;
        RECT -76.325 62.395 -75.995 62.725 ;
        RECT -76.325 61.035 -75.995 61.365 ;
        RECT -76.325 59.675 -75.995 60.005 ;
        RECT -76.325 58.315 -75.995 58.645 ;
        RECT -76.325 56.955 -75.995 57.285 ;
        RECT -76.325 55.595 -75.995 55.925 ;
        RECT -76.325 54.235 -75.995 54.565 ;
        RECT -76.325 52.875 -75.995 53.205 ;
        RECT -76.325 51.515 -75.995 51.845 ;
        RECT -76.325 50.155 -75.995 50.485 ;
        RECT -76.325 48.795 -75.995 49.125 ;
        RECT -76.325 47.435 -75.995 47.765 ;
        RECT -76.325 46.075 -75.995 46.405 ;
        RECT -76.325 44.715 -75.995 45.045 ;
        RECT -76.325 43.355 -75.995 43.685 ;
        RECT -76.325 41.995 -75.995 42.325 ;
        RECT -76.325 40.635 -75.995 40.965 ;
        RECT -76.325 39.275 -75.995 39.605 ;
        RECT -76.325 37.915 -75.995 38.245 ;
        RECT -76.325 36.555 -75.995 36.885 ;
        RECT -76.325 35.195 -75.995 35.525 ;
        RECT -76.325 33.835 -75.995 34.165 ;
        RECT -76.325 32.475 -75.995 32.805 ;
        RECT -76.325 31.115 -75.995 31.445 ;
        RECT -76.325 29.755 -75.995 30.085 ;
        RECT -76.325 28.395 -75.995 28.725 ;
        RECT -76.325 27.035 -75.995 27.365 ;
        RECT -76.325 25.675 -75.995 26.005 ;
        RECT -76.325 24.315 -75.995 24.645 ;
        RECT -76.325 22.955 -75.995 23.285 ;
        RECT -76.325 21.595 -75.995 21.925 ;
        RECT -76.325 20.235 -75.995 20.565 ;
        RECT -76.325 18.875 -75.995 19.205 ;
        RECT -76.325 17.515 -75.995 17.845 ;
        RECT -76.325 16.155 -75.995 16.485 ;
        RECT -76.325 14.795 -75.995 15.125 ;
        RECT -76.325 13.435 -75.995 13.765 ;
        RECT -76.325 12.075 -75.995 12.405 ;
        RECT -76.325 10.715 -75.995 11.045 ;
        RECT -76.325 9.355 -75.995 9.685 ;
        RECT -76.325 7.995 -75.995 8.325 ;
        RECT -76.325 6.635 -75.995 6.965 ;
        RECT -76.325 5.275 -75.995 5.605 ;
        RECT -76.325 3.915 -75.995 4.245 ;
        RECT -76.325 2.555 -75.995 2.885 ;
        RECT -76.325 1.195 -75.995 1.525 ;
        RECT -76.325 -0.165 -75.995 0.165 ;
        RECT -76.325 -1.525 -75.995 -1.195 ;
        RECT -76.325 -2.885 -75.995 -2.555 ;
        RECT -76.325 -4.245 -75.995 -3.915 ;
        RECT -76.325 -5.605 -75.995 -5.275 ;
        RECT -76.325 -6.965 -75.995 -6.635 ;
        RECT -76.325 -8.325 -75.995 -7.995 ;
        RECT -76.325 -9.685 -75.995 -9.355 ;
        RECT -76.325 -11.045 -75.995 -10.715 ;
        RECT -76.325 -12.405 -75.995 -12.075 ;
        RECT -76.325 -13.765 -75.995 -13.435 ;
        RECT -76.325 -15.125 -75.995 -14.795 ;
        RECT -76.325 -16.485 -75.995 -16.155 ;
        RECT -76.325 -17.845 -75.995 -17.515 ;
        RECT -76.325 -19.205 -75.995 -18.875 ;
        RECT -76.325 -20.565 -75.995 -20.235 ;
        RECT -76.325 -21.925 -75.995 -21.595 ;
        RECT -76.325 -23.285 -75.995 -22.955 ;
        RECT -76.325 -24.645 -75.995 -24.315 ;
        RECT -76.325 -26.005 -75.995 -25.675 ;
        RECT -76.325 -27.365 -75.995 -27.035 ;
        RECT -76.325 -28.725 -75.995 -28.395 ;
        RECT -76.325 -30.085 -75.995 -29.755 ;
        RECT -76.325 -31.445 -75.995 -31.115 ;
        RECT -76.325 -32.805 -75.995 -32.475 ;
        RECT -76.325 -34.165 -75.995 -33.835 ;
        RECT -76.325 -35.525 -75.995 -35.195 ;
        RECT -76.325 -36.885 -75.995 -36.555 ;
        RECT -76.325 -38.245 -75.995 -37.915 ;
        RECT -76.325 -39.605 -75.995 -39.275 ;
        RECT -76.325 -40.965 -75.995 -40.635 ;
        RECT -76.325 -42.325 -75.995 -41.995 ;
        RECT -76.325 -43.685 -75.995 -43.355 ;
        RECT -76.325 -45.045 -75.995 -44.715 ;
        RECT -76.325 -46.405 -75.995 -46.075 ;
        RECT -76.325 -47.765 -75.995 -47.435 ;
        RECT -76.325 -49.125 -75.995 -48.795 ;
        RECT -76.325 -50.485 -75.995 -50.155 ;
        RECT -76.325 -51.845 -75.995 -51.515 ;
        RECT -76.325 -53.205 -75.995 -52.875 ;
        RECT -76.325 -54.565 -75.995 -54.235 ;
        RECT -76.325 -55.925 -75.995 -55.595 ;
        RECT -76.325 -57.285 -75.995 -56.955 ;
        RECT -76.325 -58.645 -75.995 -58.315 ;
        RECT -76.325 -60.005 -75.995 -59.675 ;
        RECT -76.325 -61.365 -75.995 -61.035 ;
        RECT -76.325 -62.725 -75.995 -62.395 ;
        RECT -76.325 -64.085 -75.995 -63.755 ;
        RECT -76.325 -65.445 -75.995 -65.115 ;
        RECT -76.325 -66.805 -75.995 -66.475 ;
        RECT -76.325 -68.165 -75.995 -67.835 ;
        RECT -76.325 -69.525 -75.995 -69.195 ;
        RECT -76.325 -70.885 -75.995 -70.555 ;
        RECT -76.325 -72.245 -75.995 -71.915 ;
        RECT -76.325 -73.605 -75.995 -73.275 ;
        RECT -76.325 -74.965 -75.995 -74.635 ;
        RECT -76.325 -76.325 -75.995 -75.995 ;
        RECT -76.325 -77.685 -75.995 -77.355 ;
        RECT -76.325 -79.045 -75.995 -78.715 ;
        RECT -76.325 -80.405 -75.995 -80.075 ;
        RECT -76.325 -81.765 -75.995 -81.435 ;
        RECT -76.325 -83.125 -75.995 -82.795 ;
        RECT -76.325 -84.485 -75.995 -84.155 ;
        RECT -76.325 -85.845 -75.995 -85.515 ;
        RECT -76.325 -87.205 -75.995 -86.875 ;
        RECT -76.325 -88.565 -75.995 -88.235 ;
        RECT -76.325 -89.925 -75.995 -89.595 ;
        RECT -76.325 -91.285 -75.995 -90.955 ;
        RECT -76.325 -92.645 -75.995 -92.315 ;
        RECT -76.325 -94.005 -75.995 -93.675 ;
        RECT -76.325 -95.365 -75.995 -95.035 ;
        RECT -76.325 -96.725 -75.995 -96.395 ;
        RECT -76.325 -98.085 -75.995 -97.755 ;
        RECT -76.325 -99.445 -75.995 -99.115 ;
        RECT -76.325 -100.805 -75.995 -100.475 ;
        RECT -76.325 -102.165 -75.995 -101.835 ;
        RECT -76.325 -103.525 -75.995 -103.195 ;
        RECT -76.325 -104.885 -75.995 -104.555 ;
        RECT -76.325 -106.245 -75.995 -105.915 ;
        RECT -76.325 -107.605 -75.995 -107.275 ;
        RECT -76.325 -108.965 -75.995 -108.635 ;
        RECT -76.325 -110.325 -75.995 -109.995 ;
        RECT -76.325 -111.685 -75.995 -111.355 ;
        RECT -76.325 -113.045 -75.995 -112.715 ;
        RECT -76.325 -114.405 -75.995 -114.075 ;
        RECT -76.325 -115.765 -75.995 -115.435 ;
        RECT -76.325 -117.125 -75.995 -116.795 ;
        RECT -76.325 -118.485 -75.995 -118.155 ;
        RECT -76.325 -119.845 -75.995 -119.515 ;
        RECT -76.325 -121.205 -75.995 -120.875 ;
        RECT -76.325 -122.565 -75.995 -122.235 ;
        RECT -76.325 -123.925 -75.995 -123.595 ;
        RECT -76.325 -125.285 -75.995 -124.955 ;
        RECT -76.325 -126.645 -75.995 -126.315 ;
        RECT -76.325 -128.005 -75.995 -127.675 ;
        RECT -76.325 -129.365 -75.995 -129.035 ;
        RECT -76.325 -130.725 -75.995 -130.395 ;
        RECT -76.325 -132.085 -75.995 -131.755 ;
        RECT -76.325 -133.445 -75.995 -133.115 ;
        RECT -76.325 -134.805 -75.995 -134.475 ;
        RECT -76.325 -136.165 -75.995 -135.835 ;
        RECT -76.325 -137.525 -75.995 -137.195 ;
        RECT -76.325 -138.885 -75.995 -138.555 ;
        RECT -76.325 -140.245 -75.995 -139.915 ;
        RECT -76.325 -141.605 -75.995 -141.275 ;
        RECT -76.325 -142.965 -75.995 -142.635 ;
        RECT -76.325 -144.325 -75.995 -143.995 ;
        RECT -76.325 -145.685 -75.995 -145.355 ;
        RECT -76.325 -147.045 -75.995 -146.715 ;
        RECT -76.325 -148.405 -75.995 -148.075 ;
        RECT -76.325 -149.765 -75.995 -149.435 ;
        RECT -76.325 -151.125 -75.995 -150.795 ;
        RECT -76.325 -152.485 -75.995 -152.155 ;
        RECT -76.325 -153.845 -75.995 -153.515 ;
        RECT -76.325 -155.205 -75.995 -154.875 ;
        RECT -76.325 -156.565 -75.995 -156.235 ;
        RECT -76.325 -157.925 -75.995 -157.595 ;
        RECT -76.325 -159.285 -75.995 -158.955 ;
        RECT -76.325 -160.645 -75.995 -160.315 ;
        RECT -76.325 -162.005 -75.995 -161.675 ;
        RECT -76.325 -163.365 -75.995 -163.035 ;
        RECT -76.325 -164.725 -75.995 -164.395 ;
        RECT -76.325 -166.085 -75.995 -165.755 ;
        RECT -76.325 -167.445 -75.995 -167.115 ;
        RECT -76.325 -168.805 -75.995 -168.475 ;
        RECT -76.325 -170.165 -75.995 -169.835 ;
        RECT -76.325 -171.525 -75.995 -171.195 ;
        RECT -76.325 -172.885 -75.995 -172.555 ;
        RECT -76.325 -174.245 -75.995 -173.915 ;
        RECT -76.325 -175.605 -75.995 -175.275 ;
        RECT -76.325 -176.965 -75.995 -176.635 ;
        RECT -76.325 -178.325 -75.995 -177.995 ;
        RECT -76.325 -179.685 -75.995 -179.355 ;
        RECT -76.325 -181.045 -75.995 -180.715 ;
        RECT -76.325 -182.405 -75.995 -182.075 ;
        RECT -76.325 -183.765 -75.995 -183.435 ;
        RECT -76.325 -185.125 -75.995 -184.795 ;
        RECT -76.325 -186.485 -75.995 -186.155 ;
        RECT -76.325 -187.845 -75.995 -187.515 ;
        RECT -76.325 -189.205 -75.995 -188.875 ;
        RECT -76.325 -190.565 -75.995 -190.235 ;
        RECT -76.325 -191.925 -75.995 -191.595 ;
        RECT -76.325 -193.285 -75.995 -192.955 ;
        RECT -76.325 -194.645 -75.995 -194.315 ;
        RECT -76.325 -196.005 -75.995 -195.675 ;
        RECT -76.325 -197.365 -75.995 -197.035 ;
        RECT -76.325 -198.725 -75.995 -198.395 ;
        RECT -76.325 -200.085 -75.995 -199.755 ;
        RECT -76.325 -201.445 -75.995 -201.115 ;
        RECT -76.325 -202.805 -75.995 -202.475 ;
        RECT -76.325 -204.165 -75.995 -203.835 ;
        RECT -76.325 -205.525 -75.995 -205.195 ;
        RECT -76.325 -206.885 -75.995 -206.555 ;
        RECT -76.325 -208.245 -75.995 -207.915 ;
        RECT -76.325 -209.605 -75.995 -209.275 ;
        RECT -76.325 -210.965 -75.995 -210.635 ;
        RECT -76.325 -212.325 -75.995 -211.995 ;
        RECT -76.325 -213.685 -75.995 -213.355 ;
        RECT -76.325 -215.045 -75.995 -214.715 ;
        RECT -76.325 -216.405 -75.995 -216.075 ;
        RECT -76.325 -217.765 -75.995 -217.435 ;
        RECT -76.325 -219.125 -75.995 -218.795 ;
        RECT -76.325 -220.485 -75.995 -220.155 ;
        RECT -76.325 -221.845 -75.995 -221.515 ;
        RECT -76.325 -223.205 -75.995 -222.875 ;
        RECT -76.325 -224.565 -75.995 -224.235 ;
        RECT -76.325 -226.155 -75.995 -225.825 ;
        RECT -76.325 -227.285 -75.995 -226.955 ;
        RECT -76.325 -228.645 -75.995 -228.315 ;
        RECT -76.325 -231.365 -75.995 -231.035 ;
        RECT -76.325 -234.085 -75.995 -233.755 ;
        RECT -76.325 -235.445 -75.995 -235.115 ;
        RECT -76.325 -236.805 -75.995 -236.475 ;
        RECT -76.325 -238.165 -75.995 -237.835 ;
        RECT -76.325 -243.81 -75.995 -242.68 ;
        RECT -76.32 -243.925 -76 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.965 -137.525 -74.635 -137.195 ;
        RECT -74.965 -138.885 -74.635 -138.555 ;
        RECT -74.965 -140.245 -74.635 -139.915 ;
        RECT -74.965 -141.605 -74.635 -141.275 ;
        RECT -74.965 -142.965 -74.635 -142.635 ;
        RECT -74.965 -144.325 -74.635 -143.995 ;
        RECT -74.965 -145.685 -74.635 -145.355 ;
        RECT -74.965 -147.045 -74.635 -146.715 ;
        RECT -74.965 -148.405 -74.635 -148.075 ;
        RECT -74.965 -149.765 -74.635 -149.435 ;
        RECT -74.965 -151.125 -74.635 -150.795 ;
        RECT -74.965 -152.485 -74.635 -152.155 ;
        RECT -74.965 -153.845 -74.635 -153.515 ;
        RECT -74.965 -155.205 -74.635 -154.875 ;
        RECT -74.965 -156.565 -74.635 -156.235 ;
        RECT -74.965 -157.925 -74.635 -157.595 ;
        RECT -74.965 -159.285 -74.635 -158.955 ;
        RECT -74.965 -160.645 -74.635 -160.315 ;
        RECT -74.965 -162.005 -74.635 -161.675 ;
        RECT -74.965 -163.365 -74.635 -163.035 ;
        RECT -74.965 -164.725 -74.635 -164.395 ;
        RECT -74.965 -166.085 -74.635 -165.755 ;
        RECT -74.965 -167.445 -74.635 -167.115 ;
        RECT -74.965 -168.805 -74.635 -168.475 ;
        RECT -74.965 -170.165 -74.635 -169.835 ;
        RECT -74.965 -171.525 -74.635 -171.195 ;
        RECT -74.965 -172.885 -74.635 -172.555 ;
        RECT -74.965 -174.245 -74.635 -173.915 ;
        RECT -74.965 -175.605 -74.635 -175.275 ;
        RECT -74.965 -176.965 -74.635 -176.635 ;
        RECT -74.965 -178.325 -74.635 -177.995 ;
        RECT -74.965 -179.685 -74.635 -179.355 ;
        RECT -74.965 -181.045 -74.635 -180.715 ;
        RECT -74.965 -182.405 -74.635 -182.075 ;
        RECT -74.965 -183.765 -74.635 -183.435 ;
        RECT -74.965 -185.125 -74.635 -184.795 ;
        RECT -74.965 -186.485 -74.635 -186.155 ;
        RECT -74.965 -187.845 -74.635 -187.515 ;
        RECT -74.965 -189.205 -74.635 -188.875 ;
        RECT -74.965 -190.565 -74.635 -190.235 ;
        RECT -74.965 -191.925 -74.635 -191.595 ;
        RECT -74.965 -193.285 -74.635 -192.955 ;
        RECT -74.965 -194.645 -74.635 -194.315 ;
        RECT -74.965 -196.005 -74.635 -195.675 ;
        RECT -74.965 -197.365 -74.635 -197.035 ;
        RECT -74.965 -198.725 -74.635 -198.395 ;
        RECT -74.965 -200.085 -74.635 -199.755 ;
        RECT -74.965 -201.445 -74.635 -201.115 ;
        RECT -74.965 -202.805 -74.635 -202.475 ;
        RECT -74.965 -204.165 -74.635 -203.835 ;
        RECT -74.965 -205.525 -74.635 -205.195 ;
        RECT -74.965 -206.885 -74.635 -206.555 ;
        RECT -74.965 -208.245 -74.635 -207.915 ;
        RECT -74.965 -209.605 -74.635 -209.275 ;
        RECT -74.965 -210.965 -74.635 -210.635 ;
        RECT -74.965 -212.325 -74.635 -211.995 ;
        RECT -74.965 -213.685 -74.635 -213.355 ;
        RECT -74.965 -215.045 -74.635 -214.715 ;
        RECT -74.965 -216.405 -74.635 -216.075 ;
        RECT -74.965 -217.765 -74.635 -217.435 ;
        RECT -74.965 -219.125 -74.635 -218.795 ;
        RECT -74.965 -220.485 -74.635 -220.155 ;
        RECT -74.965 -221.845 -74.635 -221.515 ;
        RECT -74.965 -223.205 -74.635 -222.875 ;
        RECT -74.965 -224.565 -74.635 -224.235 ;
        RECT -74.965 -226.155 -74.635 -225.825 ;
        RECT -74.965 -227.285 -74.635 -226.955 ;
        RECT -74.965 -228.645 -74.635 -228.315 ;
        RECT -74.965 -230.005 -74.635 -229.675 ;
        RECT -74.965 -231.365 -74.635 -231.035 ;
        RECT -74.965 -234.085 -74.635 -233.755 ;
        RECT -74.965 -235.445 -74.635 -235.115 ;
        RECT -74.965 -236.805 -74.635 -236.475 ;
        RECT -74.965 -238.165 -74.635 -237.835 ;
        RECT -74.965 -243.81 -74.635 -242.68 ;
        RECT -74.96 -243.925 -74.64 248.005 ;
        RECT -74.965 246.76 -74.635 247.89 ;
        RECT -74.965 241.915 -74.635 242.245 ;
        RECT -74.965 240.555 -74.635 240.885 ;
        RECT -74.965 239.195 -74.635 239.525 ;
        RECT -74.965 237.835 -74.635 238.165 ;
        RECT -74.965 236.475 -74.635 236.805 ;
        RECT -74.965 235.115 -74.635 235.445 ;
        RECT -74.965 233.755 -74.635 234.085 ;
        RECT -74.965 232.395 -74.635 232.725 ;
        RECT -74.965 231.035 -74.635 231.365 ;
        RECT -74.965 229.675 -74.635 230.005 ;
        RECT -74.965 228.315 -74.635 228.645 ;
        RECT -74.965 226.955 -74.635 227.285 ;
        RECT -74.965 225.595 -74.635 225.925 ;
        RECT -74.965 224.235 -74.635 224.565 ;
        RECT -74.965 222.875 -74.635 223.205 ;
        RECT -74.965 221.515 -74.635 221.845 ;
        RECT -74.965 220.155 -74.635 220.485 ;
        RECT -74.965 218.795 -74.635 219.125 ;
        RECT -74.965 217.435 -74.635 217.765 ;
        RECT -74.965 216.075 -74.635 216.405 ;
        RECT -74.965 214.715 -74.635 215.045 ;
        RECT -74.965 213.355 -74.635 213.685 ;
        RECT -74.965 211.995 -74.635 212.325 ;
        RECT -74.965 210.635 -74.635 210.965 ;
        RECT -74.965 209.275 -74.635 209.605 ;
        RECT -74.965 207.915 -74.635 208.245 ;
        RECT -74.965 206.555 -74.635 206.885 ;
        RECT -74.965 205.195 -74.635 205.525 ;
        RECT -74.965 203.835 -74.635 204.165 ;
        RECT -74.965 202.475 -74.635 202.805 ;
        RECT -74.965 201.115 -74.635 201.445 ;
        RECT -74.965 199.755 -74.635 200.085 ;
        RECT -74.965 198.395 -74.635 198.725 ;
        RECT -74.965 197.035 -74.635 197.365 ;
        RECT -74.965 195.675 -74.635 196.005 ;
        RECT -74.965 194.315 -74.635 194.645 ;
        RECT -74.965 192.955 -74.635 193.285 ;
        RECT -74.965 191.595 -74.635 191.925 ;
        RECT -74.965 190.235 -74.635 190.565 ;
        RECT -74.965 188.875 -74.635 189.205 ;
        RECT -74.965 187.515 -74.635 187.845 ;
        RECT -74.965 186.155 -74.635 186.485 ;
        RECT -74.965 184.795 -74.635 185.125 ;
        RECT -74.965 183.435 -74.635 183.765 ;
        RECT -74.965 182.075 -74.635 182.405 ;
        RECT -74.965 180.715 -74.635 181.045 ;
        RECT -74.965 179.355 -74.635 179.685 ;
        RECT -74.965 177.995 -74.635 178.325 ;
        RECT -74.965 176.635 -74.635 176.965 ;
        RECT -74.965 175.275 -74.635 175.605 ;
        RECT -74.965 173.915 -74.635 174.245 ;
        RECT -74.965 172.555 -74.635 172.885 ;
        RECT -74.965 171.195 -74.635 171.525 ;
        RECT -74.965 169.835 -74.635 170.165 ;
        RECT -74.965 168.475 -74.635 168.805 ;
        RECT -74.965 167.115 -74.635 167.445 ;
        RECT -74.965 165.755 -74.635 166.085 ;
        RECT -74.965 164.395 -74.635 164.725 ;
        RECT -74.965 163.035 -74.635 163.365 ;
        RECT -74.965 161.675 -74.635 162.005 ;
        RECT -74.965 160.315 -74.635 160.645 ;
        RECT -74.965 158.955 -74.635 159.285 ;
        RECT -74.965 157.595 -74.635 157.925 ;
        RECT -74.965 156.235 -74.635 156.565 ;
        RECT -74.965 154.875 -74.635 155.205 ;
        RECT -74.965 153.515 -74.635 153.845 ;
        RECT -74.965 152.155 -74.635 152.485 ;
        RECT -74.965 150.795 -74.635 151.125 ;
        RECT -74.965 149.435 -74.635 149.765 ;
        RECT -74.965 148.075 -74.635 148.405 ;
        RECT -74.965 146.715 -74.635 147.045 ;
        RECT -74.965 145.355 -74.635 145.685 ;
        RECT -74.965 143.995 -74.635 144.325 ;
        RECT -74.965 142.635 -74.635 142.965 ;
        RECT -74.965 141.275 -74.635 141.605 ;
        RECT -74.965 139.915 -74.635 140.245 ;
        RECT -74.965 138.555 -74.635 138.885 ;
        RECT -74.965 137.195 -74.635 137.525 ;
        RECT -74.965 135.835 -74.635 136.165 ;
        RECT -74.965 134.475 -74.635 134.805 ;
        RECT -74.965 133.115 -74.635 133.445 ;
        RECT -74.965 131.755 -74.635 132.085 ;
        RECT -74.965 130.395 -74.635 130.725 ;
        RECT -74.965 129.035 -74.635 129.365 ;
        RECT -74.965 127.675 -74.635 128.005 ;
        RECT -74.965 126.315 -74.635 126.645 ;
        RECT -74.965 124.955 -74.635 125.285 ;
        RECT -74.965 123.595 -74.635 123.925 ;
        RECT -74.965 122.235 -74.635 122.565 ;
        RECT -74.965 120.875 -74.635 121.205 ;
        RECT -74.965 119.515 -74.635 119.845 ;
        RECT -74.965 118.155 -74.635 118.485 ;
        RECT -74.965 116.795 -74.635 117.125 ;
        RECT -74.965 115.435 -74.635 115.765 ;
        RECT -74.965 114.075 -74.635 114.405 ;
        RECT -74.965 112.715 -74.635 113.045 ;
        RECT -74.965 111.355 -74.635 111.685 ;
        RECT -74.965 109.995 -74.635 110.325 ;
        RECT -74.965 108.635 -74.635 108.965 ;
        RECT -74.965 107.275 -74.635 107.605 ;
        RECT -74.965 105.915 -74.635 106.245 ;
        RECT -74.965 104.555 -74.635 104.885 ;
        RECT -74.965 103.195 -74.635 103.525 ;
        RECT -74.965 101.835 -74.635 102.165 ;
        RECT -74.965 100.475 -74.635 100.805 ;
        RECT -74.965 99.115 -74.635 99.445 ;
        RECT -74.965 97.755 -74.635 98.085 ;
        RECT -74.965 96.395 -74.635 96.725 ;
        RECT -74.965 95.035 -74.635 95.365 ;
        RECT -74.965 93.675 -74.635 94.005 ;
        RECT -74.965 92.315 -74.635 92.645 ;
        RECT -74.965 90.955 -74.635 91.285 ;
        RECT -74.965 89.595 -74.635 89.925 ;
        RECT -74.965 88.235 -74.635 88.565 ;
        RECT -74.965 86.875 -74.635 87.205 ;
        RECT -74.965 85.515 -74.635 85.845 ;
        RECT -74.965 84.155 -74.635 84.485 ;
        RECT -74.965 82.795 -74.635 83.125 ;
        RECT -74.965 81.435 -74.635 81.765 ;
        RECT -74.965 80.075 -74.635 80.405 ;
        RECT -74.965 78.715 -74.635 79.045 ;
        RECT -74.965 77.355 -74.635 77.685 ;
        RECT -74.965 75.995 -74.635 76.325 ;
        RECT -74.965 74.635 -74.635 74.965 ;
        RECT -74.965 73.275 -74.635 73.605 ;
        RECT -74.965 71.915 -74.635 72.245 ;
        RECT -74.965 70.555 -74.635 70.885 ;
        RECT -74.965 69.195 -74.635 69.525 ;
        RECT -74.965 67.835 -74.635 68.165 ;
        RECT -74.965 66.475 -74.635 66.805 ;
        RECT -74.965 65.115 -74.635 65.445 ;
        RECT -74.965 63.755 -74.635 64.085 ;
        RECT -74.965 62.395 -74.635 62.725 ;
        RECT -74.965 61.035 -74.635 61.365 ;
        RECT -74.965 59.675 -74.635 60.005 ;
        RECT -74.965 58.315 -74.635 58.645 ;
        RECT -74.965 56.955 -74.635 57.285 ;
        RECT -74.965 55.595 -74.635 55.925 ;
        RECT -74.965 54.235 -74.635 54.565 ;
        RECT -74.965 52.875 -74.635 53.205 ;
        RECT -74.965 51.515 -74.635 51.845 ;
        RECT -74.965 50.155 -74.635 50.485 ;
        RECT -74.965 48.795 -74.635 49.125 ;
        RECT -74.965 47.435 -74.635 47.765 ;
        RECT -74.965 46.075 -74.635 46.405 ;
        RECT -74.965 44.715 -74.635 45.045 ;
        RECT -74.965 43.355 -74.635 43.685 ;
        RECT -74.965 41.995 -74.635 42.325 ;
        RECT -74.965 40.635 -74.635 40.965 ;
        RECT -74.965 39.275 -74.635 39.605 ;
        RECT -74.965 37.915 -74.635 38.245 ;
        RECT -74.965 36.555 -74.635 36.885 ;
        RECT -74.965 35.195 -74.635 35.525 ;
        RECT -74.965 33.835 -74.635 34.165 ;
        RECT -74.965 32.475 -74.635 32.805 ;
        RECT -74.965 31.115 -74.635 31.445 ;
        RECT -74.965 29.755 -74.635 30.085 ;
        RECT -74.965 28.395 -74.635 28.725 ;
        RECT -74.965 27.035 -74.635 27.365 ;
        RECT -74.965 25.675 -74.635 26.005 ;
        RECT -74.965 24.315 -74.635 24.645 ;
        RECT -74.965 22.955 -74.635 23.285 ;
        RECT -74.965 21.595 -74.635 21.925 ;
        RECT -74.965 20.235 -74.635 20.565 ;
        RECT -74.965 18.875 -74.635 19.205 ;
        RECT -74.965 17.515 -74.635 17.845 ;
        RECT -74.965 16.155 -74.635 16.485 ;
        RECT -74.965 14.795 -74.635 15.125 ;
        RECT -74.965 13.435 -74.635 13.765 ;
        RECT -74.965 12.075 -74.635 12.405 ;
        RECT -74.965 10.715 -74.635 11.045 ;
        RECT -74.965 9.355 -74.635 9.685 ;
        RECT -74.965 7.995 -74.635 8.325 ;
        RECT -74.965 6.635 -74.635 6.965 ;
        RECT -74.965 5.275 -74.635 5.605 ;
        RECT -74.965 3.915 -74.635 4.245 ;
        RECT -74.965 2.555 -74.635 2.885 ;
        RECT -74.965 1.195 -74.635 1.525 ;
        RECT -74.965 -0.165 -74.635 0.165 ;
        RECT -74.965 -1.525 -74.635 -1.195 ;
        RECT -74.965 -2.885 -74.635 -2.555 ;
        RECT -74.965 -4.245 -74.635 -3.915 ;
        RECT -74.965 -5.605 -74.635 -5.275 ;
        RECT -74.965 -6.965 -74.635 -6.635 ;
        RECT -74.965 -8.325 -74.635 -7.995 ;
        RECT -74.965 -9.685 -74.635 -9.355 ;
        RECT -74.965 -11.045 -74.635 -10.715 ;
        RECT -74.965 -12.405 -74.635 -12.075 ;
        RECT -74.965 -13.765 -74.635 -13.435 ;
        RECT -74.965 -15.125 -74.635 -14.795 ;
        RECT -74.965 -16.485 -74.635 -16.155 ;
        RECT -74.965 -17.845 -74.635 -17.515 ;
        RECT -74.965 -19.205 -74.635 -18.875 ;
        RECT -74.965 -20.565 -74.635 -20.235 ;
        RECT -74.965 -21.925 -74.635 -21.595 ;
        RECT -74.965 -23.285 -74.635 -22.955 ;
        RECT -74.965 -24.645 -74.635 -24.315 ;
        RECT -74.965 -26.005 -74.635 -25.675 ;
        RECT -74.965 -27.365 -74.635 -27.035 ;
        RECT -74.965 -28.725 -74.635 -28.395 ;
        RECT -74.965 -30.085 -74.635 -29.755 ;
        RECT -74.965 -31.445 -74.635 -31.115 ;
        RECT -74.965 -32.805 -74.635 -32.475 ;
        RECT -74.965 -34.165 -74.635 -33.835 ;
        RECT -74.965 -35.525 -74.635 -35.195 ;
        RECT -74.965 -36.885 -74.635 -36.555 ;
        RECT -74.965 -38.245 -74.635 -37.915 ;
        RECT -74.965 -39.605 -74.635 -39.275 ;
        RECT -74.965 -40.965 -74.635 -40.635 ;
        RECT -74.965 -42.325 -74.635 -41.995 ;
        RECT -74.965 -43.685 -74.635 -43.355 ;
        RECT -74.965 -45.045 -74.635 -44.715 ;
        RECT -74.965 -46.405 -74.635 -46.075 ;
        RECT -74.965 -47.765 -74.635 -47.435 ;
        RECT -74.965 -49.125 -74.635 -48.795 ;
        RECT -74.965 -50.485 -74.635 -50.155 ;
        RECT -74.965 -51.845 -74.635 -51.515 ;
        RECT -74.965 -53.205 -74.635 -52.875 ;
        RECT -74.965 -54.565 -74.635 -54.235 ;
        RECT -74.965 -55.925 -74.635 -55.595 ;
        RECT -74.965 -57.285 -74.635 -56.955 ;
        RECT -74.965 -58.645 -74.635 -58.315 ;
        RECT -74.965 -60.005 -74.635 -59.675 ;
        RECT -74.965 -61.365 -74.635 -61.035 ;
        RECT -74.965 -62.725 -74.635 -62.395 ;
        RECT -74.965 -64.085 -74.635 -63.755 ;
        RECT -74.965 -65.445 -74.635 -65.115 ;
        RECT -74.965 -66.805 -74.635 -66.475 ;
        RECT -74.965 -68.165 -74.635 -67.835 ;
        RECT -74.965 -69.525 -74.635 -69.195 ;
        RECT -74.965 -70.885 -74.635 -70.555 ;
        RECT -74.965 -72.245 -74.635 -71.915 ;
        RECT -74.965 -73.605 -74.635 -73.275 ;
        RECT -74.965 -74.965 -74.635 -74.635 ;
        RECT -74.965 -76.325 -74.635 -75.995 ;
        RECT -74.965 -77.685 -74.635 -77.355 ;
        RECT -74.965 -79.045 -74.635 -78.715 ;
        RECT -74.965 -80.405 -74.635 -80.075 ;
        RECT -74.965 -81.765 -74.635 -81.435 ;
        RECT -74.965 -83.125 -74.635 -82.795 ;
        RECT -74.965 -84.485 -74.635 -84.155 ;
        RECT -74.965 -85.845 -74.635 -85.515 ;
        RECT -74.965 -87.205 -74.635 -86.875 ;
        RECT -74.965 -88.565 -74.635 -88.235 ;
        RECT -74.965 -89.925 -74.635 -89.595 ;
        RECT -74.965 -91.285 -74.635 -90.955 ;
        RECT -74.965 -92.645 -74.635 -92.315 ;
        RECT -74.965 -94.005 -74.635 -93.675 ;
        RECT -74.965 -95.365 -74.635 -95.035 ;
        RECT -74.965 -96.725 -74.635 -96.395 ;
        RECT -74.965 -98.085 -74.635 -97.755 ;
        RECT -74.965 -99.445 -74.635 -99.115 ;
        RECT -74.965 -100.805 -74.635 -100.475 ;
        RECT -74.965 -102.165 -74.635 -101.835 ;
        RECT -74.965 -103.525 -74.635 -103.195 ;
        RECT -74.965 -104.885 -74.635 -104.555 ;
        RECT -74.965 -106.245 -74.635 -105.915 ;
        RECT -74.965 -107.605 -74.635 -107.275 ;
        RECT -74.965 -108.965 -74.635 -108.635 ;
        RECT -74.965 -110.325 -74.635 -109.995 ;
        RECT -74.965 -111.685 -74.635 -111.355 ;
        RECT -74.965 -113.045 -74.635 -112.715 ;
        RECT -74.965 -114.405 -74.635 -114.075 ;
        RECT -74.965 -115.765 -74.635 -115.435 ;
        RECT -74.965 -117.125 -74.635 -116.795 ;
        RECT -74.965 -118.485 -74.635 -118.155 ;
        RECT -74.965 -119.845 -74.635 -119.515 ;
        RECT -74.965 -121.205 -74.635 -120.875 ;
        RECT -74.965 -122.565 -74.635 -122.235 ;
        RECT -74.965 -123.925 -74.635 -123.595 ;
        RECT -74.965 -125.285 -74.635 -124.955 ;
        RECT -74.965 -126.645 -74.635 -126.315 ;
        RECT -74.965 -128.005 -74.635 -127.675 ;
        RECT -74.965 -129.365 -74.635 -129.035 ;
        RECT -74.965 -130.725 -74.635 -130.395 ;
        RECT -74.965 -132.085 -74.635 -131.755 ;
        RECT -74.965 -133.445 -74.635 -133.115 ;
        RECT -74.965 -134.805 -74.635 -134.475 ;
        RECT -74.965 -136.165 -74.635 -135.835 ;
    END
    PORT
      LAYER met3 ;
        RECT -81.765 246.76 -81.435 247.89 ;
        RECT -81.765 241.915 -81.435 242.245 ;
        RECT -81.765 240.555 -81.435 240.885 ;
        RECT -81.765 239.195 -81.435 239.525 ;
        RECT -81.765 237.835 -81.435 238.165 ;
        RECT -81.765 236.475 -81.435 236.805 ;
        RECT -81.765 235.115 -81.435 235.445 ;
        RECT -81.765 233.755 -81.435 234.085 ;
        RECT -81.765 232.395 -81.435 232.725 ;
        RECT -81.765 231.035 -81.435 231.365 ;
        RECT -81.765 229.675 -81.435 230.005 ;
        RECT -81.765 228.315 -81.435 228.645 ;
        RECT -81.765 226.955 -81.435 227.285 ;
        RECT -81.765 225.595 -81.435 225.925 ;
        RECT -81.765 224.235 -81.435 224.565 ;
        RECT -81.765 222.875 -81.435 223.205 ;
        RECT -81.765 221.515 -81.435 221.845 ;
        RECT -81.765 220.155 -81.435 220.485 ;
        RECT -81.765 218.795 -81.435 219.125 ;
        RECT -81.765 217.435 -81.435 217.765 ;
        RECT -81.765 216.075 -81.435 216.405 ;
        RECT -81.765 214.715 -81.435 215.045 ;
        RECT -81.765 213.355 -81.435 213.685 ;
        RECT -81.765 211.995 -81.435 212.325 ;
        RECT -81.765 210.635 -81.435 210.965 ;
        RECT -81.765 209.275 -81.435 209.605 ;
        RECT -81.765 207.915 -81.435 208.245 ;
        RECT -81.765 206.555 -81.435 206.885 ;
        RECT -81.765 205.195 -81.435 205.525 ;
        RECT -81.765 203.835 -81.435 204.165 ;
        RECT -81.765 202.475 -81.435 202.805 ;
        RECT -81.765 201.115 -81.435 201.445 ;
        RECT -81.765 199.755 -81.435 200.085 ;
        RECT -81.765 198.395 -81.435 198.725 ;
        RECT -81.765 197.035 -81.435 197.365 ;
        RECT -81.765 195.675 -81.435 196.005 ;
        RECT -81.765 194.315 -81.435 194.645 ;
        RECT -81.765 192.955 -81.435 193.285 ;
        RECT -81.765 191.595 -81.435 191.925 ;
        RECT -81.765 190.235 -81.435 190.565 ;
        RECT -81.765 188.875 -81.435 189.205 ;
        RECT -81.765 187.515 -81.435 187.845 ;
        RECT -81.765 186.155 -81.435 186.485 ;
        RECT -81.765 184.795 -81.435 185.125 ;
        RECT -81.765 183.435 -81.435 183.765 ;
        RECT -81.765 182.075 -81.435 182.405 ;
        RECT -81.765 180.715 -81.435 181.045 ;
        RECT -81.765 179.355 -81.435 179.685 ;
        RECT -81.765 177.995 -81.435 178.325 ;
        RECT -81.765 176.635 -81.435 176.965 ;
        RECT -81.765 175.275 -81.435 175.605 ;
        RECT -81.765 173.915 -81.435 174.245 ;
        RECT -81.765 172.555 -81.435 172.885 ;
        RECT -81.765 171.195 -81.435 171.525 ;
        RECT -81.765 169.835 -81.435 170.165 ;
        RECT -81.765 168.475 -81.435 168.805 ;
        RECT -81.765 167.115 -81.435 167.445 ;
        RECT -81.765 165.755 -81.435 166.085 ;
        RECT -81.765 164.395 -81.435 164.725 ;
        RECT -81.765 163.035 -81.435 163.365 ;
        RECT -81.765 161.675 -81.435 162.005 ;
        RECT -81.765 160.315 -81.435 160.645 ;
        RECT -81.765 158.955 -81.435 159.285 ;
        RECT -81.765 157.595 -81.435 157.925 ;
        RECT -81.765 156.235 -81.435 156.565 ;
        RECT -81.765 154.875 -81.435 155.205 ;
        RECT -81.765 153.515 -81.435 153.845 ;
        RECT -81.765 152.155 -81.435 152.485 ;
        RECT -81.765 150.795 -81.435 151.125 ;
        RECT -81.765 149.435 -81.435 149.765 ;
        RECT -81.765 148.075 -81.435 148.405 ;
        RECT -81.765 146.715 -81.435 147.045 ;
        RECT -81.765 145.355 -81.435 145.685 ;
        RECT -81.765 143.995 -81.435 144.325 ;
        RECT -81.765 142.635 -81.435 142.965 ;
        RECT -81.765 141.275 -81.435 141.605 ;
        RECT -81.765 139.915 -81.435 140.245 ;
        RECT -81.765 138.555 -81.435 138.885 ;
        RECT -81.765 137.195 -81.435 137.525 ;
        RECT -81.765 135.835 -81.435 136.165 ;
        RECT -81.765 134.475 -81.435 134.805 ;
        RECT -81.765 133.115 -81.435 133.445 ;
        RECT -81.765 131.755 -81.435 132.085 ;
        RECT -81.765 130.395 -81.435 130.725 ;
        RECT -81.765 129.035 -81.435 129.365 ;
        RECT -81.765 127.675 -81.435 128.005 ;
        RECT -81.765 126.315 -81.435 126.645 ;
        RECT -81.765 124.955 -81.435 125.285 ;
        RECT -81.765 123.595 -81.435 123.925 ;
        RECT -81.765 122.235 -81.435 122.565 ;
        RECT -81.765 120.875 -81.435 121.205 ;
        RECT -81.765 119.515 -81.435 119.845 ;
        RECT -81.765 118.155 -81.435 118.485 ;
        RECT -81.765 116.795 -81.435 117.125 ;
        RECT -81.765 115.435 -81.435 115.765 ;
        RECT -81.765 114.075 -81.435 114.405 ;
        RECT -81.765 112.715 -81.435 113.045 ;
        RECT -81.765 111.355 -81.435 111.685 ;
        RECT -81.765 109.995 -81.435 110.325 ;
        RECT -81.765 108.635 -81.435 108.965 ;
        RECT -81.765 107.275 -81.435 107.605 ;
        RECT -81.765 105.915 -81.435 106.245 ;
        RECT -81.765 104.555 -81.435 104.885 ;
        RECT -81.765 103.195 -81.435 103.525 ;
        RECT -81.765 101.835 -81.435 102.165 ;
        RECT -81.765 100.475 -81.435 100.805 ;
        RECT -81.765 99.115 -81.435 99.445 ;
        RECT -81.765 97.755 -81.435 98.085 ;
        RECT -81.765 96.395 -81.435 96.725 ;
        RECT -81.765 95.035 -81.435 95.365 ;
        RECT -81.765 93.675 -81.435 94.005 ;
        RECT -81.765 92.315 -81.435 92.645 ;
        RECT -81.765 90.955 -81.435 91.285 ;
        RECT -81.765 89.595 -81.435 89.925 ;
        RECT -81.765 88.235 -81.435 88.565 ;
        RECT -81.765 86.875 -81.435 87.205 ;
        RECT -81.765 85.515 -81.435 85.845 ;
        RECT -81.765 84.155 -81.435 84.485 ;
        RECT -81.765 82.795 -81.435 83.125 ;
        RECT -81.765 81.435 -81.435 81.765 ;
        RECT -81.765 80.075 -81.435 80.405 ;
        RECT -81.765 78.715 -81.435 79.045 ;
        RECT -81.765 77.355 -81.435 77.685 ;
        RECT -81.765 75.995 -81.435 76.325 ;
        RECT -81.765 74.635 -81.435 74.965 ;
        RECT -81.765 73.275 -81.435 73.605 ;
        RECT -81.765 71.915 -81.435 72.245 ;
        RECT -81.765 70.555 -81.435 70.885 ;
        RECT -81.765 69.195 -81.435 69.525 ;
        RECT -81.765 67.835 -81.435 68.165 ;
        RECT -81.765 66.475 -81.435 66.805 ;
        RECT -81.765 65.115 -81.435 65.445 ;
        RECT -81.765 63.755 -81.435 64.085 ;
        RECT -81.765 62.395 -81.435 62.725 ;
        RECT -81.765 61.035 -81.435 61.365 ;
        RECT -81.765 59.675 -81.435 60.005 ;
        RECT -81.765 58.315 -81.435 58.645 ;
        RECT -81.765 56.955 -81.435 57.285 ;
        RECT -81.765 55.595 -81.435 55.925 ;
        RECT -81.765 54.235 -81.435 54.565 ;
        RECT -81.765 52.875 -81.435 53.205 ;
        RECT -81.765 51.515 -81.435 51.845 ;
        RECT -81.765 50.155 -81.435 50.485 ;
        RECT -81.765 48.795 -81.435 49.125 ;
        RECT -81.765 47.435 -81.435 47.765 ;
        RECT -81.765 46.075 -81.435 46.405 ;
        RECT -81.765 44.715 -81.435 45.045 ;
        RECT -81.765 43.355 -81.435 43.685 ;
        RECT -81.765 41.995 -81.435 42.325 ;
        RECT -81.765 40.635 -81.435 40.965 ;
        RECT -81.765 39.275 -81.435 39.605 ;
        RECT -81.765 37.915 -81.435 38.245 ;
        RECT -81.765 36.555 -81.435 36.885 ;
        RECT -81.765 35.195 -81.435 35.525 ;
        RECT -81.765 33.835 -81.435 34.165 ;
        RECT -81.765 32.475 -81.435 32.805 ;
        RECT -81.765 31.115 -81.435 31.445 ;
        RECT -81.765 29.755 -81.435 30.085 ;
        RECT -81.765 28.395 -81.435 28.725 ;
        RECT -81.765 27.035 -81.435 27.365 ;
        RECT -81.765 25.675 -81.435 26.005 ;
        RECT -81.765 24.315 -81.435 24.645 ;
        RECT -81.765 22.955 -81.435 23.285 ;
        RECT -81.765 21.595 -81.435 21.925 ;
        RECT -81.765 20.235 -81.435 20.565 ;
        RECT -81.765 18.875 -81.435 19.205 ;
        RECT -81.765 17.515 -81.435 17.845 ;
        RECT -81.765 16.155 -81.435 16.485 ;
        RECT -81.765 14.795 -81.435 15.125 ;
        RECT -81.765 13.435 -81.435 13.765 ;
        RECT -81.765 12.075 -81.435 12.405 ;
        RECT -81.765 10.715 -81.435 11.045 ;
        RECT -81.765 9.355 -81.435 9.685 ;
        RECT -81.765 7.995 -81.435 8.325 ;
        RECT -81.765 6.635 -81.435 6.965 ;
        RECT -81.765 5.275 -81.435 5.605 ;
        RECT -81.765 3.915 -81.435 4.245 ;
        RECT -81.765 2.555 -81.435 2.885 ;
        RECT -81.765 1.195 -81.435 1.525 ;
        RECT -81.765 -0.165 -81.435 0.165 ;
        RECT -81.765 -1.525 -81.435 -1.195 ;
        RECT -81.765 -2.885 -81.435 -2.555 ;
        RECT -81.765 -4.245 -81.435 -3.915 ;
        RECT -81.765 -5.605 -81.435 -5.275 ;
        RECT -81.765 -6.965 -81.435 -6.635 ;
        RECT -81.765 -8.325 -81.435 -7.995 ;
        RECT -81.765 -9.685 -81.435 -9.355 ;
        RECT -81.765 -11.045 -81.435 -10.715 ;
        RECT -81.765 -12.405 -81.435 -12.075 ;
        RECT -81.765 -13.765 -81.435 -13.435 ;
        RECT -81.765 -15.125 -81.435 -14.795 ;
        RECT -81.765 -16.485 -81.435 -16.155 ;
        RECT -81.765 -17.845 -81.435 -17.515 ;
        RECT -81.765 -19.205 -81.435 -18.875 ;
        RECT -81.765 -20.565 -81.435 -20.235 ;
        RECT -81.765 -21.925 -81.435 -21.595 ;
        RECT -81.765 -23.285 -81.435 -22.955 ;
        RECT -81.765 -24.645 -81.435 -24.315 ;
        RECT -81.765 -26.005 -81.435 -25.675 ;
        RECT -81.765 -27.365 -81.435 -27.035 ;
        RECT -81.765 -28.725 -81.435 -28.395 ;
        RECT -81.765 -30.085 -81.435 -29.755 ;
        RECT -81.765 -31.445 -81.435 -31.115 ;
        RECT -81.765 -32.805 -81.435 -32.475 ;
        RECT -81.765 -34.165 -81.435 -33.835 ;
        RECT -81.765 -35.525 -81.435 -35.195 ;
        RECT -81.765 -36.885 -81.435 -36.555 ;
        RECT -81.765 -38.245 -81.435 -37.915 ;
        RECT -81.765 -39.605 -81.435 -39.275 ;
        RECT -81.765 -40.965 -81.435 -40.635 ;
        RECT -81.765 -42.325 -81.435 -41.995 ;
        RECT -81.765 -43.685 -81.435 -43.355 ;
        RECT -81.765 -45.045 -81.435 -44.715 ;
        RECT -81.765 -46.405 -81.435 -46.075 ;
        RECT -81.765 -47.765 -81.435 -47.435 ;
        RECT -81.765 -49.125 -81.435 -48.795 ;
        RECT -81.765 -50.485 -81.435 -50.155 ;
        RECT -81.765 -51.845 -81.435 -51.515 ;
        RECT -81.765 -53.205 -81.435 -52.875 ;
        RECT -81.765 -54.565 -81.435 -54.235 ;
        RECT -81.765 -55.925 -81.435 -55.595 ;
        RECT -81.765 -57.285 -81.435 -56.955 ;
        RECT -81.765 -58.645 -81.435 -58.315 ;
        RECT -81.765 -60.005 -81.435 -59.675 ;
        RECT -81.765 -61.365 -81.435 -61.035 ;
        RECT -81.765 -62.725 -81.435 -62.395 ;
        RECT -81.765 -64.085 -81.435 -63.755 ;
        RECT -81.765 -65.445 -81.435 -65.115 ;
        RECT -81.765 -66.805 -81.435 -66.475 ;
        RECT -81.765 -68.165 -81.435 -67.835 ;
        RECT -81.765 -69.525 -81.435 -69.195 ;
        RECT -81.765 -70.885 -81.435 -70.555 ;
        RECT -81.765 -72.245 -81.435 -71.915 ;
        RECT -81.765 -73.605 -81.435 -73.275 ;
        RECT -81.765 -74.965 -81.435 -74.635 ;
        RECT -81.765 -76.325 -81.435 -75.995 ;
        RECT -81.765 -77.685 -81.435 -77.355 ;
        RECT -81.765 -79.045 -81.435 -78.715 ;
        RECT -81.765 -80.405 -81.435 -80.075 ;
        RECT -81.765 -81.765 -81.435 -81.435 ;
        RECT -81.765 -83.125 -81.435 -82.795 ;
        RECT -81.765 -84.485 -81.435 -84.155 ;
        RECT -81.765 -85.845 -81.435 -85.515 ;
        RECT -81.765 -87.205 -81.435 -86.875 ;
        RECT -81.765 -88.565 -81.435 -88.235 ;
        RECT -81.765 -89.925 -81.435 -89.595 ;
        RECT -81.765 -91.285 -81.435 -90.955 ;
        RECT -81.765 -92.645 -81.435 -92.315 ;
        RECT -81.765 -94.005 -81.435 -93.675 ;
        RECT -81.765 -95.365 -81.435 -95.035 ;
        RECT -81.765 -96.725 -81.435 -96.395 ;
        RECT -81.765 -98.085 -81.435 -97.755 ;
        RECT -81.765 -99.445 -81.435 -99.115 ;
        RECT -81.765 -100.805 -81.435 -100.475 ;
        RECT -81.765 -102.165 -81.435 -101.835 ;
        RECT -81.765 -103.525 -81.435 -103.195 ;
        RECT -81.765 -104.885 -81.435 -104.555 ;
        RECT -81.765 -106.245 -81.435 -105.915 ;
        RECT -81.765 -107.605 -81.435 -107.275 ;
        RECT -81.765 -108.965 -81.435 -108.635 ;
        RECT -81.765 -110.325 -81.435 -109.995 ;
        RECT -81.765 -111.685 -81.435 -111.355 ;
        RECT -81.765 -113.045 -81.435 -112.715 ;
        RECT -81.765 -114.405 -81.435 -114.075 ;
        RECT -81.765 -115.765 -81.435 -115.435 ;
        RECT -81.765 -117.125 -81.435 -116.795 ;
        RECT -81.765 -118.485 -81.435 -118.155 ;
        RECT -81.765 -119.845 -81.435 -119.515 ;
        RECT -81.765 -121.205 -81.435 -120.875 ;
        RECT -81.765 -122.565 -81.435 -122.235 ;
        RECT -81.765 -123.925 -81.435 -123.595 ;
        RECT -81.765 -125.285 -81.435 -124.955 ;
        RECT -81.765 -126.645 -81.435 -126.315 ;
        RECT -81.765 -128.005 -81.435 -127.675 ;
        RECT -81.765 -129.365 -81.435 -129.035 ;
        RECT -81.765 -130.725 -81.435 -130.395 ;
        RECT -81.765 -132.085 -81.435 -131.755 ;
        RECT -81.765 -133.445 -81.435 -133.115 ;
        RECT -81.765 -134.805 -81.435 -134.475 ;
        RECT -81.765 -136.165 -81.435 -135.835 ;
        RECT -81.765 -137.525 -81.435 -137.195 ;
        RECT -81.765 -138.885 -81.435 -138.555 ;
        RECT -81.765 -140.245 -81.435 -139.915 ;
        RECT -81.765 -141.605 -81.435 -141.275 ;
        RECT -81.765 -142.965 -81.435 -142.635 ;
        RECT -81.765 -144.325 -81.435 -143.995 ;
        RECT -81.765 -145.685 -81.435 -145.355 ;
        RECT -81.765 -147.045 -81.435 -146.715 ;
        RECT -81.765 -148.405 -81.435 -148.075 ;
        RECT -81.765 -149.765 -81.435 -149.435 ;
        RECT -81.765 -151.125 -81.435 -150.795 ;
        RECT -81.765 -152.485 -81.435 -152.155 ;
        RECT -81.765 -153.845 -81.435 -153.515 ;
        RECT -81.765 -155.205 -81.435 -154.875 ;
        RECT -81.765 -156.565 -81.435 -156.235 ;
        RECT -81.765 -157.925 -81.435 -157.595 ;
        RECT -81.765 -159.285 -81.435 -158.955 ;
        RECT -81.765 -160.645 -81.435 -160.315 ;
        RECT -81.765 -162.005 -81.435 -161.675 ;
        RECT -81.765 -163.365 -81.435 -163.035 ;
        RECT -81.765 -164.725 -81.435 -164.395 ;
        RECT -81.765 -166.085 -81.435 -165.755 ;
        RECT -81.765 -167.445 -81.435 -167.115 ;
        RECT -81.765 -168.805 -81.435 -168.475 ;
        RECT -81.765 -170.165 -81.435 -169.835 ;
        RECT -81.765 -171.525 -81.435 -171.195 ;
        RECT -81.765 -172.885 -81.435 -172.555 ;
        RECT -81.765 -174.245 -81.435 -173.915 ;
        RECT -81.765 -175.605 -81.435 -175.275 ;
        RECT -81.765 -176.965 -81.435 -176.635 ;
        RECT -81.765 -178.325 -81.435 -177.995 ;
        RECT -81.765 -179.685 -81.435 -179.355 ;
        RECT -81.765 -181.045 -81.435 -180.715 ;
        RECT -81.765 -182.405 -81.435 -182.075 ;
        RECT -81.765 -183.765 -81.435 -183.435 ;
        RECT -81.765 -185.125 -81.435 -184.795 ;
        RECT -81.765 -186.485 -81.435 -186.155 ;
        RECT -81.765 -187.845 -81.435 -187.515 ;
        RECT -81.765 -189.205 -81.435 -188.875 ;
        RECT -81.765 -190.565 -81.435 -190.235 ;
        RECT -81.765 -191.925 -81.435 -191.595 ;
        RECT -81.765 -193.285 -81.435 -192.955 ;
        RECT -81.765 -194.645 -81.435 -194.315 ;
        RECT -81.765 -196.005 -81.435 -195.675 ;
        RECT -81.765 -197.365 -81.435 -197.035 ;
        RECT -81.765 -198.725 -81.435 -198.395 ;
        RECT -81.765 -200.085 -81.435 -199.755 ;
        RECT -81.765 -201.445 -81.435 -201.115 ;
        RECT -81.765 -202.805 -81.435 -202.475 ;
        RECT -81.765 -204.165 -81.435 -203.835 ;
        RECT -81.765 -205.525 -81.435 -205.195 ;
        RECT -81.765 -206.885 -81.435 -206.555 ;
        RECT -81.765 -208.245 -81.435 -207.915 ;
        RECT -81.765 -209.605 -81.435 -209.275 ;
        RECT -81.765 -210.965 -81.435 -210.635 ;
        RECT -81.765 -212.325 -81.435 -211.995 ;
        RECT -81.765 -213.685 -81.435 -213.355 ;
        RECT -81.765 -215.045 -81.435 -214.715 ;
        RECT -81.765 -216.405 -81.435 -216.075 ;
        RECT -81.765 -217.765 -81.435 -217.435 ;
        RECT -81.765 -219.125 -81.435 -218.795 ;
        RECT -81.765 -220.485 -81.435 -220.155 ;
        RECT -81.765 -221.845 -81.435 -221.515 ;
        RECT -81.765 -223.205 -81.435 -222.875 ;
        RECT -81.765 -224.565 -81.435 -224.235 ;
        RECT -81.765 -225.925 -81.435 -225.595 ;
        RECT -81.765 -227.285 -81.435 -226.955 ;
        RECT -81.765 -228.645 -81.435 -228.315 ;
        RECT -81.765 -230.005 -81.435 -229.675 ;
        RECT -81.765 -231.365 -81.435 -231.035 ;
        RECT -81.765 -232.725 -81.435 -232.395 ;
        RECT -81.765 -234.085 -81.435 -233.755 ;
        RECT -81.765 -235.445 -81.435 -235.115 ;
        RECT -81.765 -236.805 -81.435 -236.475 ;
        RECT -81.765 -238.165 -81.435 -237.835 ;
        RECT -81.765 -243.81 -81.435 -242.68 ;
        RECT -81.76 -243.925 -81.44 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -80.405 246.76 -80.075 247.89 ;
        RECT -80.405 241.915 -80.075 242.245 ;
        RECT -80.405 240.555 -80.075 240.885 ;
        RECT -80.405 239.195 -80.075 239.525 ;
        RECT -80.405 237.835 -80.075 238.165 ;
        RECT -80.405 236.475 -80.075 236.805 ;
        RECT -80.405 235.115 -80.075 235.445 ;
        RECT -80.405 233.755 -80.075 234.085 ;
        RECT -80.405 232.395 -80.075 232.725 ;
        RECT -80.405 231.035 -80.075 231.365 ;
        RECT -80.405 229.675 -80.075 230.005 ;
        RECT -80.405 228.315 -80.075 228.645 ;
        RECT -80.405 226.955 -80.075 227.285 ;
        RECT -80.405 225.595 -80.075 225.925 ;
        RECT -80.405 224.235 -80.075 224.565 ;
        RECT -80.405 222.875 -80.075 223.205 ;
        RECT -80.405 221.515 -80.075 221.845 ;
        RECT -80.405 220.155 -80.075 220.485 ;
        RECT -80.405 218.795 -80.075 219.125 ;
        RECT -80.405 217.435 -80.075 217.765 ;
        RECT -80.405 216.075 -80.075 216.405 ;
        RECT -80.405 214.715 -80.075 215.045 ;
        RECT -80.405 213.355 -80.075 213.685 ;
        RECT -80.405 211.995 -80.075 212.325 ;
        RECT -80.405 210.635 -80.075 210.965 ;
        RECT -80.405 209.275 -80.075 209.605 ;
        RECT -80.405 207.915 -80.075 208.245 ;
        RECT -80.405 206.555 -80.075 206.885 ;
        RECT -80.405 205.195 -80.075 205.525 ;
        RECT -80.405 203.835 -80.075 204.165 ;
        RECT -80.405 202.475 -80.075 202.805 ;
        RECT -80.405 201.115 -80.075 201.445 ;
        RECT -80.405 199.755 -80.075 200.085 ;
        RECT -80.405 198.395 -80.075 198.725 ;
        RECT -80.405 197.035 -80.075 197.365 ;
        RECT -80.405 195.675 -80.075 196.005 ;
        RECT -80.405 194.315 -80.075 194.645 ;
        RECT -80.405 192.955 -80.075 193.285 ;
        RECT -80.405 191.595 -80.075 191.925 ;
        RECT -80.405 190.235 -80.075 190.565 ;
        RECT -80.405 188.875 -80.075 189.205 ;
        RECT -80.405 187.515 -80.075 187.845 ;
        RECT -80.405 186.155 -80.075 186.485 ;
        RECT -80.405 184.795 -80.075 185.125 ;
        RECT -80.405 183.435 -80.075 183.765 ;
        RECT -80.405 182.075 -80.075 182.405 ;
        RECT -80.405 180.715 -80.075 181.045 ;
        RECT -80.405 179.355 -80.075 179.685 ;
        RECT -80.405 177.995 -80.075 178.325 ;
        RECT -80.405 176.635 -80.075 176.965 ;
        RECT -80.405 175.275 -80.075 175.605 ;
        RECT -80.405 173.915 -80.075 174.245 ;
        RECT -80.405 172.555 -80.075 172.885 ;
        RECT -80.405 171.195 -80.075 171.525 ;
        RECT -80.405 169.835 -80.075 170.165 ;
        RECT -80.405 168.475 -80.075 168.805 ;
        RECT -80.405 167.115 -80.075 167.445 ;
        RECT -80.405 165.755 -80.075 166.085 ;
        RECT -80.405 164.395 -80.075 164.725 ;
        RECT -80.405 163.035 -80.075 163.365 ;
        RECT -80.405 161.675 -80.075 162.005 ;
        RECT -80.405 160.315 -80.075 160.645 ;
        RECT -80.405 158.955 -80.075 159.285 ;
        RECT -80.405 157.595 -80.075 157.925 ;
        RECT -80.405 156.235 -80.075 156.565 ;
        RECT -80.405 154.875 -80.075 155.205 ;
        RECT -80.405 153.515 -80.075 153.845 ;
        RECT -80.405 152.155 -80.075 152.485 ;
        RECT -80.405 150.795 -80.075 151.125 ;
        RECT -80.405 149.435 -80.075 149.765 ;
        RECT -80.405 148.075 -80.075 148.405 ;
        RECT -80.405 146.715 -80.075 147.045 ;
        RECT -80.405 145.355 -80.075 145.685 ;
        RECT -80.405 143.995 -80.075 144.325 ;
        RECT -80.405 142.635 -80.075 142.965 ;
        RECT -80.405 141.275 -80.075 141.605 ;
        RECT -80.405 139.915 -80.075 140.245 ;
        RECT -80.405 138.555 -80.075 138.885 ;
        RECT -80.405 137.195 -80.075 137.525 ;
        RECT -80.405 135.835 -80.075 136.165 ;
        RECT -80.405 134.475 -80.075 134.805 ;
        RECT -80.405 133.115 -80.075 133.445 ;
        RECT -80.405 131.755 -80.075 132.085 ;
        RECT -80.405 130.395 -80.075 130.725 ;
        RECT -80.405 129.035 -80.075 129.365 ;
        RECT -80.405 127.675 -80.075 128.005 ;
        RECT -80.405 126.315 -80.075 126.645 ;
        RECT -80.405 124.955 -80.075 125.285 ;
        RECT -80.405 123.595 -80.075 123.925 ;
        RECT -80.405 122.235 -80.075 122.565 ;
        RECT -80.405 120.875 -80.075 121.205 ;
        RECT -80.405 119.515 -80.075 119.845 ;
        RECT -80.405 118.155 -80.075 118.485 ;
        RECT -80.405 116.795 -80.075 117.125 ;
        RECT -80.405 115.435 -80.075 115.765 ;
        RECT -80.405 114.075 -80.075 114.405 ;
        RECT -80.405 112.715 -80.075 113.045 ;
        RECT -80.405 111.355 -80.075 111.685 ;
        RECT -80.405 109.995 -80.075 110.325 ;
        RECT -80.405 108.635 -80.075 108.965 ;
        RECT -80.405 107.275 -80.075 107.605 ;
        RECT -80.405 105.915 -80.075 106.245 ;
        RECT -80.405 104.555 -80.075 104.885 ;
        RECT -80.405 103.195 -80.075 103.525 ;
        RECT -80.405 101.835 -80.075 102.165 ;
        RECT -80.405 100.475 -80.075 100.805 ;
        RECT -80.405 99.115 -80.075 99.445 ;
        RECT -80.405 97.755 -80.075 98.085 ;
        RECT -80.405 96.395 -80.075 96.725 ;
        RECT -80.405 95.035 -80.075 95.365 ;
        RECT -80.405 93.675 -80.075 94.005 ;
        RECT -80.405 92.315 -80.075 92.645 ;
        RECT -80.405 90.955 -80.075 91.285 ;
        RECT -80.405 89.595 -80.075 89.925 ;
        RECT -80.405 88.235 -80.075 88.565 ;
        RECT -80.405 86.875 -80.075 87.205 ;
        RECT -80.405 85.515 -80.075 85.845 ;
        RECT -80.405 84.155 -80.075 84.485 ;
        RECT -80.405 82.795 -80.075 83.125 ;
        RECT -80.405 81.435 -80.075 81.765 ;
        RECT -80.405 80.075 -80.075 80.405 ;
        RECT -80.405 78.715 -80.075 79.045 ;
        RECT -80.405 77.355 -80.075 77.685 ;
        RECT -80.405 75.995 -80.075 76.325 ;
        RECT -80.405 74.635 -80.075 74.965 ;
        RECT -80.405 73.275 -80.075 73.605 ;
        RECT -80.405 71.915 -80.075 72.245 ;
        RECT -80.405 70.555 -80.075 70.885 ;
        RECT -80.405 69.195 -80.075 69.525 ;
        RECT -80.405 67.835 -80.075 68.165 ;
        RECT -80.405 66.475 -80.075 66.805 ;
        RECT -80.405 65.115 -80.075 65.445 ;
        RECT -80.405 63.755 -80.075 64.085 ;
        RECT -80.405 62.395 -80.075 62.725 ;
        RECT -80.405 61.035 -80.075 61.365 ;
        RECT -80.405 59.675 -80.075 60.005 ;
        RECT -80.405 58.315 -80.075 58.645 ;
        RECT -80.405 56.955 -80.075 57.285 ;
        RECT -80.405 55.595 -80.075 55.925 ;
        RECT -80.405 54.235 -80.075 54.565 ;
        RECT -80.405 52.875 -80.075 53.205 ;
        RECT -80.405 51.515 -80.075 51.845 ;
        RECT -80.405 50.155 -80.075 50.485 ;
        RECT -80.405 48.795 -80.075 49.125 ;
        RECT -80.405 47.435 -80.075 47.765 ;
        RECT -80.405 46.075 -80.075 46.405 ;
        RECT -80.405 44.715 -80.075 45.045 ;
        RECT -80.405 43.355 -80.075 43.685 ;
        RECT -80.405 41.995 -80.075 42.325 ;
        RECT -80.405 40.635 -80.075 40.965 ;
        RECT -80.405 39.275 -80.075 39.605 ;
        RECT -80.405 37.915 -80.075 38.245 ;
        RECT -80.405 36.555 -80.075 36.885 ;
        RECT -80.405 35.195 -80.075 35.525 ;
        RECT -80.405 33.835 -80.075 34.165 ;
        RECT -80.405 32.475 -80.075 32.805 ;
        RECT -80.405 31.115 -80.075 31.445 ;
        RECT -80.405 29.755 -80.075 30.085 ;
        RECT -80.405 28.395 -80.075 28.725 ;
        RECT -80.405 27.035 -80.075 27.365 ;
        RECT -80.405 25.675 -80.075 26.005 ;
        RECT -80.405 24.315 -80.075 24.645 ;
        RECT -80.405 22.955 -80.075 23.285 ;
        RECT -80.405 21.595 -80.075 21.925 ;
        RECT -80.405 20.235 -80.075 20.565 ;
        RECT -80.405 18.875 -80.075 19.205 ;
        RECT -80.405 17.515 -80.075 17.845 ;
        RECT -80.405 16.155 -80.075 16.485 ;
        RECT -80.405 14.795 -80.075 15.125 ;
        RECT -80.405 13.435 -80.075 13.765 ;
        RECT -80.405 12.075 -80.075 12.405 ;
        RECT -80.405 10.715 -80.075 11.045 ;
        RECT -80.405 9.355 -80.075 9.685 ;
        RECT -80.405 7.995 -80.075 8.325 ;
        RECT -80.405 6.635 -80.075 6.965 ;
        RECT -80.405 5.275 -80.075 5.605 ;
        RECT -80.405 3.915 -80.075 4.245 ;
        RECT -80.405 2.555 -80.075 2.885 ;
        RECT -80.405 1.195 -80.075 1.525 ;
        RECT -80.405 -0.165 -80.075 0.165 ;
        RECT -80.405 -1.525 -80.075 -1.195 ;
        RECT -80.405 -2.885 -80.075 -2.555 ;
        RECT -80.405 -4.245 -80.075 -3.915 ;
        RECT -80.405 -5.605 -80.075 -5.275 ;
        RECT -80.405 -6.965 -80.075 -6.635 ;
        RECT -80.405 -8.325 -80.075 -7.995 ;
        RECT -80.405 -9.685 -80.075 -9.355 ;
        RECT -80.405 -11.045 -80.075 -10.715 ;
        RECT -80.405 -12.405 -80.075 -12.075 ;
        RECT -80.405 -13.765 -80.075 -13.435 ;
        RECT -80.405 -15.125 -80.075 -14.795 ;
        RECT -80.405 -16.485 -80.075 -16.155 ;
        RECT -80.405 -17.845 -80.075 -17.515 ;
        RECT -80.405 -19.205 -80.075 -18.875 ;
        RECT -80.405 -20.565 -80.075 -20.235 ;
        RECT -80.405 -21.925 -80.075 -21.595 ;
        RECT -80.405 -23.285 -80.075 -22.955 ;
        RECT -80.405 -24.645 -80.075 -24.315 ;
        RECT -80.405 -26.005 -80.075 -25.675 ;
        RECT -80.405 -27.365 -80.075 -27.035 ;
        RECT -80.405 -28.725 -80.075 -28.395 ;
        RECT -80.405 -30.085 -80.075 -29.755 ;
        RECT -80.405 -31.445 -80.075 -31.115 ;
        RECT -80.405 -32.805 -80.075 -32.475 ;
        RECT -80.405 -34.165 -80.075 -33.835 ;
        RECT -80.405 -35.525 -80.075 -35.195 ;
        RECT -80.405 -36.885 -80.075 -36.555 ;
        RECT -80.405 -38.245 -80.075 -37.915 ;
        RECT -80.405 -39.605 -80.075 -39.275 ;
        RECT -80.405 -40.965 -80.075 -40.635 ;
        RECT -80.405 -42.325 -80.075 -41.995 ;
        RECT -80.405 -43.685 -80.075 -43.355 ;
        RECT -80.405 -45.045 -80.075 -44.715 ;
        RECT -80.405 -46.405 -80.075 -46.075 ;
        RECT -80.405 -47.765 -80.075 -47.435 ;
        RECT -80.405 -49.125 -80.075 -48.795 ;
        RECT -80.405 -50.485 -80.075 -50.155 ;
        RECT -80.405 -51.845 -80.075 -51.515 ;
        RECT -80.405 -53.205 -80.075 -52.875 ;
        RECT -80.405 -54.565 -80.075 -54.235 ;
        RECT -80.405 -55.925 -80.075 -55.595 ;
        RECT -80.405 -57.285 -80.075 -56.955 ;
        RECT -80.405 -58.645 -80.075 -58.315 ;
        RECT -80.405 -60.005 -80.075 -59.675 ;
        RECT -80.405 -61.365 -80.075 -61.035 ;
        RECT -80.405 -62.725 -80.075 -62.395 ;
        RECT -80.405 -64.085 -80.075 -63.755 ;
        RECT -80.405 -65.445 -80.075 -65.115 ;
        RECT -80.405 -66.805 -80.075 -66.475 ;
        RECT -80.405 -68.165 -80.075 -67.835 ;
        RECT -80.405 -69.525 -80.075 -69.195 ;
        RECT -80.405 -70.885 -80.075 -70.555 ;
        RECT -80.405 -72.245 -80.075 -71.915 ;
        RECT -80.405 -73.605 -80.075 -73.275 ;
        RECT -80.405 -74.965 -80.075 -74.635 ;
        RECT -80.405 -76.325 -80.075 -75.995 ;
        RECT -80.405 -77.685 -80.075 -77.355 ;
        RECT -80.405 -79.045 -80.075 -78.715 ;
        RECT -80.405 -80.405 -80.075 -80.075 ;
        RECT -80.405 -81.765 -80.075 -81.435 ;
        RECT -80.405 -83.125 -80.075 -82.795 ;
        RECT -80.405 -84.485 -80.075 -84.155 ;
        RECT -80.405 -85.845 -80.075 -85.515 ;
        RECT -80.405 -87.205 -80.075 -86.875 ;
        RECT -80.405 -88.565 -80.075 -88.235 ;
        RECT -80.405 -89.925 -80.075 -89.595 ;
        RECT -80.405 -91.285 -80.075 -90.955 ;
        RECT -80.405 -92.645 -80.075 -92.315 ;
        RECT -80.405 -94.005 -80.075 -93.675 ;
        RECT -80.405 -95.365 -80.075 -95.035 ;
        RECT -80.405 -96.725 -80.075 -96.395 ;
        RECT -80.405 -98.085 -80.075 -97.755 ;
        RECT -80.405 -99.445 -80.075 -99.115 ;
        RECT -80.405 -100.805 -80.075 -100.475 ;
        RECT -80.405 -102.165 -80.075 -101.835 ;
        RECT -80.405 -103.525 -80.075 -103.195 ;
        RECT -80.405 -104.885 -80.075 -104.555 ;
        RECT -80.405 -106.245 -80.075 -105.915 ;
        RECT -80.405 -107.605 -80.075 -107.275 ;
        RECT -80.405 -108.965 -80.075 -108.635 ;
        RECT -80.405 -110.325 -80.075 -109.995 ;
        RECT -80.405 -111.685 -80.075 -111.355 ;
        RECT -80.405 -113.045 -80.075 -112.715 ;
        RECT -80.405 -114.405 -80.075 -114.075 ;
        RECT -80.405 -115.765 -80.075 -115.435 ;
        RECT -80.405 -117.125 -80.075 -116.795 ;
        RECT -80.405 -118.485 -80.075 -118.155 ;
        RECT -80.405 -119.845 -80.075 -119.515 ;
        RECT -80.405 -121.205 -80.075 -120.875 ;
        RECT -80.405 -122.565 -80.075 -122.235 ;
        RECT -80.405 -123.925 -80.075 -123.595 ;
        RECT -80.405 -125.285 -80.075 -124.955 ;
        RECT -80.405 -126.645 -80.075 -126.315 ;
        RECT -80.405 -128.005 -80.075 -127.675 ;
        RECT -80.405 -129.365 -80.075 -129.035 ;
        RECT -80.405 -130.725 -80.075 -130.395 ;
        RECT -80.405 -132.085 -80.075 -131.755 ;
        RECT -80.405 -133.445 -80.075 -133.115 ;
        RECT -80.405 -134.805 -80.075 -134.475 ;
        RECT -80.405 -136.165 -80.075 -135.835 ;
        RECT -80.405 -137.525 -80.075 -137.195 ;
        RECT -80.405 -138.885 -80.075 -138.555 ;
        RECT -80.405 -140.245 -80.075 -139.915 ;
        RECT -80.405 -141.605 -80.075 -141.275 ;
        RECT -80.405 -142.965 -80.075 -142.635 ;
        RECT -80.405 -144.325 -80.075 -143.995 ;
        RECT -80.405 -145.685 -80.075 -145.355 ;
        RECT -80.405 -147.045 -80.075 -146.715 ;
        RECT -80.405 -148.405 -80.075 -148.075 ;
        RECT -80.405 -149.765 -80.075 -149.435 ;
        RECT -80.405 -151.125 -80.075 -150.795 ;
        RECT -80.405 -152.485 -80.075 -152.155 ;
        RECT -80.405 -153.845 -80.075 -153.515 ;
        RECT -80.405 -155.205 -80.075 -154.875 ;
        RECT -80.405 -156.565 -80.075 -156.235 ;
        RECT -80.405 -157.925 -80.075 -157.595 ;
        RECT -80.405 -159.285 -80.075 -158.955 ;
        RECT -80.405 -160.645 -80.075 -160.315 ;
        RECT -80.405 -162.005 -80.075 -161.675 ;
        RECT -80.405 -163.365 -80.075 -163.035 ;
        RECT -80.405 -164.725 -80.075 -164.395 ;
        RECT -80.405 -166.085 -80.075 -165.755 ;
        RECT -80.405 -167.445 -80.075 -167.115 ;
        RECT -80.405 -168.805 -80.075 -168.475 ;
        RECT -80.405 -170.165 -80.075 -169.835 ;
        RECT -80.405 -171.525 -80.075 -171.195 ;
        RECT -80.405 -172.885 -80.075 -172.555 ;
        RECT -80.405 -174.245 -80.075 -173.915 ;
        RECT -80.405 -175.605 -80.075 -175.275 ;
        RECT -80.405 -176.965 -80.075 -176.635 ;
        RECT -80.405 -178.325 -80.075 -177.995 ;
        RECT -80.405 -179.685 -80.075 -179.355 ;
        RECT -80.405 -181.045 -80.075 -180.715 ;
        RECT -80.405 -182.405 -80.075 -182.075 ;
        RECT -80.405 -183.765 -80.075 -183.435 ;
        RECT -80.405 -185.125 -80.075 -184.795 ;
        RECT -80.405 -186.485 -80.075 -186.155 ;
        RECT -80.405 -187.845 -80.075 -187.515 ;
        RECT -80.405 -189.205 -80.075 -188.875 ;
        RECT -80.405 -190.565 -80.075 -190.235 ;
        RECT -80.405 -191.925 -80.075 -191.595 ;
        RECT -80.405 -193.285 -80.075 -192.955 ;
        RECT -80.405 -194.645 -80.075 -194.315 ;
        RECT -80.405 -196.005 -80.075 -195.675 ;
        RECT -80.405 -197.365 -80.075 -197.035 ;
        RECT -80.405 -198.725 -80.075 -198.395 ;
        RECT -80.405 -200.085 -80.075 -199.755 ;
        RECT -80.405 -201.445 -80.075 -201.115 ;
        RECT -80.405 -202.805 -80.075 -202.475 ;
        RECT -80.405 -204.165 -80.075 -203.835 ;
        RECT -80.405 -205.525 -80.075 -205.195 ;
        RECT -80.405 -206.885 -80.075 -206.555 ;
        RECT -80.405 -208.245 -80.075 -207.915 ;
        RECT -80.405 -209.605 -80.075 -209.275 ;
        RECT -80.405 -210.965 -80.075 -210.635 ;
        RECT -80.405 -212.325 -80.075 -211.995 ;
        RECT -80.405 -213.685 -80.075 -213.355 ;
        RECT -80.405 -215.045 -80.075 -214.715 ;
        RECT -80.405 -216.405 -80.075 -216.075 ;
        RECT -80.405 -217.765 -80.075 -217.435 ;
        RECT -80.405 -219.125 -80.075 -218.795 ;
        RECT -80.405 -220.485 -80.075 -220.155 ;
        RECT -80.405 -221.845 -80.075 -221.515 ;
        RECT -80.405 -223.205 -80.075 -222.875 ;
        RECT -80.405 -224.565 -80.075 -224.235 ;
        RECT -80.405 -225.925 -80.075 -225.595 ;
        RECT -80.405 -227.285 -80.075 -226.955 ;
        RECT -80.405 -228.645 -80.075 -228.315 ;
        RECT -80.405 -230.005 -80.075 -229.675 ;
        RECT -80.405 -231.365 -80.075 -231.035 ;
        RECT -80.405 -232.725 -80.075 -232.395 ;
        RECT -80.405 -234.085 -80.075 -233.755 ;
        RECT -80.405 -235.445 -80.075 -235.115 ;
        RECT -80.405 -236.805 -80.075 -236.475 ;
        RECT -80.405 -238.165 -80.075 -237.835 ;
        RECT -80.405 -243.81 -80.075 -242.68 ;
        RECT -80.4 -243.925 -80.08 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.045 -55.925 -78.715 -55.595 ;
        RECT -79.045 -57.285 -78.715 -56.955 ;
        RECT -79.045 -58.645 -78.715 -58.315 ;
        RECT -79.045 -60.005 -78.715 -59.675 ;
        RECT -79.045 -61.365 -78.715 -61.035 ;
        RECT -79.045 -62.725 -78.715 -62.395 ;
        RECT -79.045 -64.085 -78.715 -63.755 ;
        RECT -79.045 -65.445 -78.715 -65.115 ;
        RECT -79.045 -66.805 -78.715 -66.475 ;
        RECT -79.045 -68.165 -78.715 -67.835 ;
        RECT -79.045 -69.525 -78.715 -69.195 ;
        RECT -79.045 -70.885 -78.715 -70.555 ;
        RECT -79.045 -72.245 -78.715 -71.915 ;
        RECT -79.045 -73.605 -78.715 -73.275 ;
        RECT -79.045 -74.965 -78.715 -74.635 ;
        RECT -79.045 -76.325 -78.715 -75.995 ;
        RECT -79.045 -77.685 -78.715 -77.355 ;
        RECT -79.045 -79.045 -78.715 -78.715 ;
        RECT -79.045 -80.405 -78.715 -80.075 ;
        RECT -79.045 -81.765 -78.715 -81.435 ;
        RECT -79.045 -83.125 -78.715 -82.795 ;
        RECT -79.045 -84.485 -78.715 -84.155 ;
        RECT -79.045 -85.845 -78.715 -85.515 ;
        RECT -79.045 -87.205 -78.715 -86.875 ;
        RECT -79.045 -88.565 -78.715 -88.235 ;
        RECT -79.045 -89.925 -78.715 -89.595 ;
        RECT -79.045 -91.285 -78.715 -90.955 ;
        RECT -79.045 -92.645 -78.715 -92.315 ;
        RECT -79.045 -94.005 -78.715 -93.675 ;
        RECT -79.045 -95.365 -78.715 -95.035 ;
        RECT -79.045 -96.725 -78.715 -96.395 ;
        RECT -79.045 -98.085 -78.715 -97.755 ;
        RECT -79.045 -99.445 -78.715 -99.115 ;
        RECT -79.045 -100.805 -78.715 -100.475 ;
        RECT -79.045 -102.165 -78.715 -101.835 ;
        RECT -79.045 -103.525 -78.715 -103.195 ;
        RECT -79.045 -104.885 -78.715 -104.555 ;
        RECT -79.045 -106.245 -78.715 -105.915 ;
        RECT -79.045 -107.605 -78.715 -107.275 ;
        RECT -79.045 -108.965 -78.715 -108.635 ;
        RECT -79.045 -110.325 -78.715 -109.995 ;
        RECT -79.045 -111.685 -78.715 -111.355 ;
        RECT -79.045 -113.045 -78.715 -112.715 ;
        RECT -79.045 -114.405 -78.715 -114.075 ;
        RECT -79.045 -115.765 -78.715 -115.435 ;
        RECT -79.045 -117.125 -78.715 -116.795 ;
        RECT -79.045 -118.485 -78.715 -118.155 ;
        RECT -79.045 -119.845 -78.715 -119.515 ;
        RECT -79.045 -121.205 -78.715 -120.875 ;
        RECT -79.045 -122.565 -78.715 -122.235 ;
        RECT -79.045 -123.925 -78.715 -123.595 ;
        RECT -79.045 -125.285 -78.715 -124.955 ;
        RECT -79.045 -126.645 -78.715 -126.315 ;
        RECT -79.045 -128.005 -78.715 -127.675 ;
        RECT -79.045 -129.365 -78.715 -129.035 ;
        RECT -79.045 -130.725 -78.715 -130.395 ;
        RECT -79.045 -132.085 -78.715 -131.755 ;
        RECT -79.045 -133.445 -78.715 -133.115 ;
        RECT -79.045 -134.805 -78.715 -134.475 ;
        RECT -79.045 -136.165 -78.715 -135.835 ;
        RECT -79.045 -137.525 -78.715 -137.195 ;
        RECT -79.045 -138.885 -78.715 -138.555 ;
        RECT -79.045 -140.245 -78.715 -139.915 ;
        RECT -79.045 -141.605 -78.715 -141.275 ;
        RECT -79.045 -142.965 -78.715 -142.635 ;
        RECT -79.045 -144.325 -78.715 -143.995 ;
        RECT -79.045 -145.685 -78.715 -145.355 ;
        RECT -79.045 -147.045 -78.715 -146.715 ;
        RECT -79.045 -148.405 -78.715 -148.075 ;
        RECT -79.045 -149.765 -78.715 -149.435 ;
        RECT -79.045 -151.125 -78.715 -150.795 ;
        RECT -79.045 -152.485 -78.715 -152.155 ;
        RECT -79.045 -153.845 -78.715 -153.515 ;
        RECT -79.045 -155.205 -78.715 -154.875 ;
        RECT -79.045 -156.565 -78.715 -156.235 ;
        RECT -79.045 -157.925 -78.715 -157.595 ;
        RECT -79.045 -159.285 -78.715 -158.955 ;
        RECT -79.045 -160.645 -78.715 -160.315 ;
        RECT -79.045 -162.005 -78.715 -161.675 ;
        RECT -79.045 -163.365 -78.715 -163.035 ;
        RECT -79.045 -164.725 -78.715 -164.395 ;
        RECT -79.045 -166.085 -78.715 -165.755 ;
        RECT -79.045 -167.445 -78.715 -167.115 ;
        RECT -79.045 -168.805 -78.715 -168.475 ;
        RECT -79.045 -170.165 -78.715 -169.835 ;
        RECT -79.045 -171.525 -78.715 -171.195 ;
        RECT -79.045 -172.885 -78.715 -172.555 ;
        RECT -79.045 -174.245 -78.715 -173.915 ;
        RECT -79.045 -175.605 -78.715 -175.275 ;
        RECT -79.045 -176.965 -78.715 -176.635 ;
        RECT -79.045 -178.325 -78.715 -177.995 ;
        RECT -79.045 -179.685 -78.715 -179.355 ;
        RECT -79.045 -181.045 -78.715 -180.715 ;
        RECT -79.045 -182.405 -78.715 -182.075 ;
        RECT -79.045 -183.765 -78.715 -183.435 ;
        RECT -79.045 -185.125 -78.715 -184.795 ;
        RECT -79.045 -186.485 -78.715 -186.155 ;
        RECT -79.045 -187.845 -78.715 -187.515 ;
        RECT -79.045 -189.205 -78.715 -188.875 ;
        RECT -79.045 -190.565 -78.715 -190.235 ;
        RECT -79.045 -191.925 -78.715 -191.595 ;
        RECT -79.045 -193.285 -78.715 -192.955 ;
        RECT -79.045 -194.645 -78.715 -194.315 ;
        RECT -79.045 -196.005 -78.715 -195.675 ;
        RECT -79.045 -197.365 -78.715 -197.035 ;
        RECT -79.045 -198.725 -78.715 -198.395 ;
        RECT -79.045 -200.085 -78.715 -199.755 ;
        RECT -79.045 -201.445 -78.715 -201.115 ;
        RECT -79.045 -202.805 -78.715 -202.475 ;
        RECT -79.045 -204.165 -78.715 -203.835 ;
        RECT -79.045 -205.525 -78.715 -205.195 ;
        RECT -79.045 -206.885 -78.715 -206.555 ;
        RECT -79.045 -208.245 -78.715 -207.915 ;
        RECT -79.045 -209.605 -78.715 -209.275 ;
        RECT -79.045 -210.965 -78.715 -210.635 ;
        RECT -79.045 -212.325 -78.715 -211.995 ;
        RECT -79.045 -213.685 -78.715 -213.355 ;
        RECT -79.045 -215.045 -78.715 -214.715 ;
        RECT -79.045 -216.405 -78.715 -216.075 ;
        RECT -79.045 -217.765 -78.715 -217.435 ;
        RECT -79.045 -219.125 -78.715 -218.795 ;
        RECT -79.045 -220.485 -78.715 -220.155 ;
        RECT -79.045 -221.845 -78.715 -221.515 ;
        RECT -79.045 -223.205 -78.715 -222.875 ;
        RECT -79.045 -224.565 -78.715 -224.235 ;
        RECT -79.045 -225.925 -78.715 -225.595 ;
        RECT -79.045 -227.285 -78.715 -226.955 ;
        RECT -79.045 -228.645 -78.715 -228.315 ;
        RECT -79.045 -230.005 -78.715 -229.675 ;
        RECT -79.045 -231.365 -78.715 -231.035 ;
        RECT -79.045 -232.725 -78.715 -232.395 ;
        RECT -79.045 -234.085 -78.715 -233.755 ;
        RECT -79.045 -235.445 -78.715 -235.115 ;
        RECT -79.045 -236.805 -78.715 -236.475 ;
        RECT -79.045 -238.165 -78.715 -237.835 ;
        RECT -79.045 -243.81 -78.715 -242.68 ;
        RECT -79.04 -243.925 -78.72 248.005 ;
        RECT -79.045 246.76 -78.715 247.89 ;
        RECT -79.045 241.915 -78.715 242.245 ;
        RECT -79.045 240.555 -78.715 240.885 ;
        RECT -79.045 239.195 -78.715 239.525 ;
        RECT -79.045 237.835 -78.715 238.165 ;
        RECT -79.045 236.475 -78.715 236.805 ;
        RECT -79.045 235.115 -78.715 235.445 ;
        RECT -79.045 233.755 -78.715 234.085 ;
        RECT -79.045 232.395 -78.715 232.725 ;
        RECT -79.045 231.035 -78.715 231.365 ;
        RECT -79.045 229.675 -78.715 230.005 ;
        RECT -79.045 228.315 -78.715 228.645 ;
        RECT -79.045 226.955 -78.715 227.285 ;
        RECT -79.045 225.595 -78.715 225.925 ;
        RECT -79.045 224.235 -78.715 224.565 ;
        RECT -79.045 222.875 -78.715 223.205 ;
        RECT -79.045 221.515 -78.715 221.845 ;
        RECT -79.045 220.155 -78.715 220.485 ;
        RECT -79.045 218.795 -78.715 219.125 ;
        RECT -79.045 217.435 -78.715 217.765 ;
        RECT -79.045 216.075 -78.715 216.405 ;
        RECT -79.045 214.715 -78.715 215.045 ;
        RECT -79.045 213.355 -78.715 213.685 ;
        RECT -79.045 211.995 -78.715 212.325 ;
        RECT -79.045 210.635 -78.715 210.965 ;
        RECT -79.045 209.275 -78.715 209.605 ;
        RECT -79.045 207.915 -78.715 208.245 ;
        RECT -79.045 206.555 -78.715 206.885 ;
        RECT -79.045 205.195 -78.715 205.525 ;
        RECT -79.045 203.835 -78.715 204.165 ;
        RECT -79.045 202.475 -78.715 202.805 ;
        RECT -79.045 201.115 -78.715 201.445 ;
        RECT -79.045 199.755 -78.715 200.085 ;
        RECT -79.045 198.395 -78.715 198.725 ;
        RECT -79.045 197.035 -78.715 197.365 ;
        RECT -79.045 195.675 -78.715 196.005 ;
        RECT -79.045 194.315 -78.715 194.645 ;
        RECT -79.045 192.955 -78.715 193.285 ;
        RECT -79.045 191.595 -78.715 191.925 ;
        RECT -79.045 190.235 -78.715 190.565 ;
        RECT -79.045 188.875 -78.715 189.205 ;
        RECT -79.045 187.515 -78.715 187.845 ;
        RECT -79.045 186.155 -78.715 186.485 ;
        RECT -79.045 184.795 -78.715 185.125 ;
        RECT -79.045 183.435 -78.715 183.765 ;
        RECT -79.045 182.075 -78.715 182.405 ;
        RECT -79.045 180.715 -78.715 181.045 ;
        RECT -79.045 179.355 -78.715 179.685 ;
        RECT -79.045 177.995 -78.715 178.325 ;
        RECT -79.045 176.635 -78.715 176.965 ;
        RECT -79.045 175.275 -78.715 175.605 ;
        RECT -79.045 173.915 -78.715 174.245 ;
        RECT -79.045 172.555 -78.715 172.885 ;
        RECT -79.045 171.195 -78.715 171.525 ;
        RECT -79.045 169.835 -78.715 170.165 ;
        RECT -79.045 168.475 -78.715 168.805 ;
        RECT -79.045 167.115 -78.715 167.445 ;
        RECT -79.045 165.755 -78.715 166.085 ;
        RECT -79.045 164.395 -78.715 164.725 ;
        RECT -79.045 163.035 -78.715 163.365 ;
        RECT -79.045 161.675 -78.715 162.005 ;
        RECT -79.045 160.315 -78.715 160.645 ;
        RECT -79.045 158.955 -78.715 159.285 ;
        RECT -79.045 157.595 -78.715 157.925 ;
        RECT -79.045 156.235 -78.715 156.565 ;
        RECT -79.045 154.875 -78.715 155.205 ;
        RECT -79.045 153.515 -78.715 153.845 ;
        RECT -79.045 152.155 -78.715 152.485 ;
        RECT -79.045 150.795 -78.715 151.125 ;
        RECT -79.045 149.435 -78.715 149.765 ;
        RECT -79.045 148.075 -78.715 148.405 ;
        RECT -79.045 146.715 -78.715 147.045 ;
        RECT -79.045 145.355 -78.715 145.685 ;
        RECT -79.045 143.995 -78.715 144.325 ;
        RECT -79.045 142.635 -78.715 142.965 ;
        RECT -79.045 141.275 -78.715 141.605 ;
        RECT -79.045 139.915 -78.715 140.245 ;
        RECT -79.045 138.555 -78.715 138.885 ;
        RECT -79.045 137.195 -78.715 137.525 ;
        RECT -79.045 135.835 -78.715 136.165 ;
        RECT -79.045 134.475 -78.715 134.805 ;
        RECT -79.045 133.115 -78.715 133.445 ;
        RECT -79.045 131.755 -78.715 132.085 ;
        RECT -79.045 130.395 -78.715 130.725 ;
        RECT -79.045 129.035 -78.715 129.365 ;
        RECT -79.045 127.675 -78.715 128.005 ;
        RECT -79.045 126.315 -78.715 126.645 ;
        RECT -79.045 124.955 -78.715 125.285 ;
        RECT -79.045 123.595 -78.715 123.925 ;
        RECT -79.045 122.235 -78.715 122.565 ;
        RECT -79.045 120.875 -78.715 121.205 ;
        RECT -79.045 119.515 -78.715 119.845 ;
        RECT -79.045 118.155 -78.715 118.485 ;
        RECT -79.045 116.795 -78.715 117.125 ;
        RECT -79.045 115.435 -78.715 115.765 ;
        RECT -79.045 114.075 -78.715 114.405 ;
        RECT -79.045 112.715 -78.715 113.045 ;
        RECT -79.045 111.355 -78.715 111.685 ;
        RECT -79.045 109.995 -78.715 110.325 ;
        RECT -79.045 108.635 -78.715 108.965 ;
        RECT -79.045 107.275 -78.715 107.605 ;
        RECT -79.045 105.915 -78.715 106.245 ;
        RECT -79.045 104.555 -78.715 104.885 ;
        RECT -79.045 103.195 -78.715 103.525 ;
        RECT -79.045 101.835 -78.715 102.165 ;
        RECT -79.045 100.475 -78.715 100.805 ;
        RECT -79.045 99.115 -78.715 99.445 ;
        RECT -79.045 97.755 -78.715 98.085 ;
        RECT -79.045 96.395 -78.715 96.725 ;
        RECT -79.045 95.035 -78.715 95.365 ;
        RECT -79.045 93.675 -78.715 94.005 ;
        RECT -79.045 92.315 -78.715 92.645 ;
        RECT -79.045 90.955 -78.715 91.285 ;
        RECT -79.045 89.595 -78.715 89.925 ;
        RECT -79.045 88.235 -78.715 88.565 ;
        RECT -79.045 86.875 -78.715 87.205 ;
        RECT -79.045 85.515 -78.715 85.845 ;
        RECT -79.045 84.155 -78.715 84.485 ;
        RECT -79.045 82.795 -78.715 83.125 ;
        RECT -79.045 81.435 -78.715 81.765 ;
        RECT -79.045 80.075 -78.715 80.405 ;
        RECT -79.045 78.715 -78.715 79.045 ;
        RECT -79.045 77.355 -78.715 77.685 ;
        RECT -79.045 75.995 -78.715 76.325 ;
        RECT -79.045 74.635 -78.715 74.965 ;
        RECT -79.045 73.275 -78.715 73.605 ;
        RECT -79.045 71.915 -78.715 72.245 ;
        RECT -79.045 70.555 -78.715 70.885 ;
        RECT -79.045 69.195 -78.715 69.525 ;
        RECT -79.045 67.835 -78.715 68.165 ;
        RECT -79.045 66.475 -78.715 66.805 ;
        RECT -79.045 65.115 -78.715 65.445 ;
        RECT -79.045 63.755 -78.715 64.085 ;
        RECT -79.045 62.395 -78.715 62.725 ;
        RECT -79.045 61.035 -78.715 61.365 ;
        RECT -79.045 59.675 -78.715 60.005 ;
        RECT -79.045 58.315 -78.715 58.645 ;
        RECT -79.045 56.955 -78.715 57.285 ;
        RECT -79.045 55.595 -78.715 55.925 ;
        RECT -79.045 54.235 -78.715 54.565 ;
        RECT -79.045 52.875 -78.715 53.205 ;
        RECT -79.045 51.515 -78.715 51.845 ;
        RECT -79.045 50.155 -78.715 50.485 ;
        RECT -79.045 48.795 -78.715 49.125 ;
        RECT -79.045 47.435 -78.715 47.765 ;
        RECT -79.045 46.075 -78.715 46.405 ;
        RECT -79.045 44.715 -78.715 45.045 ;
        RECT -79.045 43.355 -78.715 43.685 ;
        RECT -79.045 41.995 -78.715 42.325 ;
        RECT -79.045 40.635 -78.715 40.965 ;
        RECT -79.045 39.275 -78.715 39.605 ;
        RECT -79.045 37.915 -78.715 38.245 ;
        RECT -79.045 36.555 -78.715 36.885 ;
        RECT -79.045 35.195 -78.715 35.525 ;
        RECT -79.045 33.835 -78.715 34.165 ;
        RECT -79.045 32.475 -78.715 32.805 ;
        RECT -79.045 31.115 -78.715 31.445 ;
        RECT -79.045 29.755 -78.715 30.085 ;
        RECT -79.045 28.395 -78.715 28.725 ;
        RECT -79.045 27.035 -78.715 27.365 ;
        RECT -79.045 25.675 -78.715 26.005 ;
        RECT -79.045 24.315 -78.715 24.645 ;
        RECT -79.045 22.955 -78.715 23.285 ;
        RECT -79.045 21.595 -78.715 21.925 ;
        RECT -79.045 20.235 -78.715 20.565 ;
        RECT -79.045 18.875 -78.715 19.205 ;
        RECT -79.045 17.515 -78.715 17.845 ;
        RECT -79.045 16.155 -78.715 16.485 ;
        RECT -79.045 14.795 -78.715 15.125 ;
        RECT -79.045 13.435 -78.715 13.765 ;
        RECT -79.045 12.075 -78.715 12.405 ;
        RECT -79.045 10.715 -78.715 11.045 ;
        RECT -79.045 9.355 -78.715 9.685 ;
        RECT -79.045 7.995 -78.715 8.325 ;
        RECT -79.045 6.635 -78.715 6.965 ;
        RECT -79.045 5.275 -78.715 5.605 ;
        RECT -79.045 3.915 -78.715 4.245 ;
        RECT -79.045 2.555 -78.715 2.885 ;
        RECT -79.045 1.195 -78.715 1.525 ;
        RECT -79.045 -0.165 -78.715 0.165 ;
        RECT -79.045 -1.525 -78.715 -1.195 ;
        RECT -79.045 -2.885 -78.715 -2.555 ;
        RECT -79.045 -4.245 -78.715 -3.915 ;
        RECT -79.045 -5.605 -78.715 -5.275 ;
        RECT -79.045 -6.965 -78.715 -6.635 ;
        RECT -79.045 -8.325 -78.715 -7.995 ;
        RECT -79.045 -9.685 -78.715 -9.355 ;
        RECT -79.045 -11.045 -78.715 -10.715 ;
        RECT -79.045 -12.405 -78.715 -12.075 ;
        RECT -79.045 -13.765 -78.715 -13.435 ;
        RECT -79.045 -15.125 -78.715 -14.795 ;
        RECT -79.045 -16.485 -78.715 -16.155 ;
        RECT -79.045 -17.845 -78.715 -17.515 ;
        RECT -79.045 -19.205 -78.715 -18.875 ;
        RECT -79.045 -20.565 -78.715 -20.235 ;
        RECT -79.045 -21.925 -78.715 -21.595 ;
        RECT -79.045 -23.285 -78.715 -22.955 ;
        RECT -79.045 -24.645 -78.715 -24.315 ;
        RECT -79.045 -26.005 -78.715 -25.675 ;
        RECT -79.045 -27.365 -78.715 -27.035 ;
        RECT -79.045 -28.725 -78.715 -28.395 ;
        RECT -79.045 -30.085 -78.715 -29.755 ;
        RECT -79.045 -31.445 -78.715 -31.115 ;
        RECT -79.045 -32.805 -78.715 -32.475 ;
        RECT -79.045 -34.165 -78.715 -33.835 ;
        RECT -79.045 -35.525 -78.715 -35.195 ;
        RECT -79.045 -36.885 -78.715 -36.555 ;
        RECT -79.045 -38.245 -78.715 -37.915 ;
        RECT -79.045 -39.605 -78.715 -39.275 ;
        RECT -79.045 -40.965 -78.715 -40.635 ;
        RECT -79.045 -42.325 -78.715 -41.995 ;
        RECT -79.045 -43.685 -78.715 -43.355 ;
        RECT -79.045 -45.045 -78.715 -44.715 ;
        RECT -79.045 -46.405 -78.715 -46.075 ;
        RECT -79.045 -47.765 -78.715 -47.435 ;
        RECT -79.045 -49.125 -78.715 -48.795 ;
        RECT -79.045 -50.485 -78.715 -50.155 ;
        RECT -79.045 -51.845 -78.715 -51.515 ;
        RECT -79.045 -53.205 -78.715 -52.875 ;
        RECT -79.045 -54.565 -78.715 -54.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -83.125 40.635 -82.795 40.965 ;
        RECT -83.125 39.275 -82.795 39.605 ;
        RECT -83.125 37.915 -82.795 38.245 ;
        RECT -83.125 36.555 -82.795 36.885 ;
        RECT -83.125 35.195 -82.795 35.525 ;
        RECT -83.125 33.835 -82.795 34.165 ;
        RECT -83.125 32.475 -82.795 32.805 ;
        RECT -83.125 31.115 -82.795 31.445 ;
        RECT -83.125 29.755 -82.795 30.085 ;
        RECT -83.125 28.395 -82.795 28.725 ;
        RECT -83.125 27.035 -82.795 27.365 ;
        RECT -83.125 25.675 -82.795 26.005 ;
        RECT -83.125 24.315 -82.795 24.645 ;
        RECT -83.125 22.955 -82.795 23.285 ;
        RECT -83.125 21.595 -82.795 21.925 ;
        RECT -83.125 20.235 -82.795 20.565 ;
        RECT -83.125 18.875 -82.795 19.205 ;
        RECT -83.125 17.515 -82.795 17.845 ;
        RECT -83.125 16.155 -82.795 16.485 ;
        RECT -83.125 14.795 -82.795 15.125 ;
        RECT -83.125 13.435 -82.795 13.765 ;
        RECT -83.125 12.075 -82.795 12.405 ;
        RECT -83.125 10.715 -82.795 11.045 ;
        RECT -83.125 9.355 -82.795 9.685 ;
        RECT -83.125 7.995 -82.795 8.325 ;
        RECT -83.125 6.635 -82.795 6.965 ;
        RECT -83.125 5.275 -82.795 5.605 ;
        RECT -83.125 3.915 -82.795 4.245 ;
        RECT -83.125 2.555 -82.795 2.885 ;
        RECT -83.125 1.195 -82.795 1.525 ;
        RECT -83.125 -0.165 -82.795 0.165 ;
        RECT -83.125 -1.525 -82.795 -1.195 ;
        RECT -83.125 -2.885 -82.795 -2.555 ;
        RECT -83.125 -4.245 -82.795 -3.915 ;
        RECT -83.125 -5.605 -82.795 -5.275 ;
        RECT -83.125 -6.965 -82.795 -6.635 ;
        RECT -83.125 -8.325 -82.795 -7.995 ;
        RECT -83.125 -9.685 -82.795 -9.355 ;
        RECT -83.125 -11.045 -82.795 -10.715 ;
        RECT -83.125 -12.405 -82.795 -12.075 ;
        RECT -83.125 -13.765 -82.795 -13.435 ;
        RECT -83.125 -15.125 -82.795 -14.795 ;
        RECT -83.125 -16.485 -82.795 -16.155 ;
        RECT -83.125 -17.845 -82.795 -17.515 ;
        RECT -83.125 -19.205 -82.795 -18.875 ;
        RECT -83.125 -20.565 -82.795 -20.235 ;
        RECT -83.125 -21.925 -82.795 -21.595 ;
        RECT -83.125 -23.285 -82.795 -22.955 ;
        RECT -83.125 -24.645 -82.795 -24.315 ;
        RECT -83.125 -26.005 -82.795 -25.675 ;
        RECT -83.125 -27.365 -82.795 -27.035 ;
        RECT -83.125 -28.725 -82.795 -28.395 ;
        RECT -83.125 -30.085 -82.795 -29.755 ;
        RECT -83.125 -31.445 -82.795 -31.115 ;
        RECT -83.125 -32.805 -82.795 -32.475 ;
        RECT -83.125 -34.165 -82.795 -33.835 ;
        RECT -83.125 -35.525 -82.795 -35.195 ;
        RECT -83.125 -36.885 -82.795 -36.555 ;
        RECT -83.125 -38.245 -82.795 -37.915 ;
        RECT -83.125 -39.605 -82.795 -39.275 ;
        RECT -83.125 -40.965 -82.795 -40.635 ;
        RECT -83.125 -42.325 -82.795 -41.995 ;
        RECT -83.125 -43.685 -82.795 -43.355 ;
        RECT -83.125 -45.045 -82.795 -44.715 ;
        RECT -83.125 -46.405 -82.795 -46.075 ;
        RECT -83.125 -47.765 -82.795 -47.435 ;
        RECT -83.125 -49.125 -82.795 -48.795 ;
        RECT -83.125 -50.485 -82.795 -50.155 ;
        RECT -83.125 -51.845 -82.795 -51.515 ;
        RECT -83.125 -53.205 -82.795 -52.875 ;
        RECT -83.125 -54.565 -82.795 -54.235 ;
        RECT -83.125 -55.925 -82.795 -55.595 ;
        RECT -83.125 -57.285 -82.795 -56.955 ;
        RECT -83.125 -58.645 -82.795 -58.315 ;
        RECT -83.125 -60.005 -82.795 -59.675 ;
        RECT -83.125 -61.365 -82.795 -61.035 ;
        RECT -83.125 -62.725 -82.795 -62.395 ;
        RECT -83.125 -64.085 -82.795 -63.755 ;
        RECT -83.125 -65.445 -82.795 -65.115 ;
        RECT -83.125 -66.805 -82.795 -66.475 ;
        RECT -83.125 -68.165 -82.795 -67.835 ;
        RECT -83.125 -69.525 -82.795 -69.195 ;
        RECT -83.125 -70.885 -82.795 -70.555 ;
        RECT -83.125 -72.245 -82.795 -71.915 ;
        RECT -83.125 -73.605 -82.795 -73.275 ;
        RECT -83.125 -74.965 -82.795 -74.635 ;
        RECT -83.125 -76.325 -82.795 -75.995 ;
        RECT -83.125 -77.685 -82.795 -77.355 ;
        RECT -83.125 -79.045 -82.795 -78.715 ;
        RECT -83.125 -80.405 -82.795 -80.075 ;
        RECT -83.125 -81.765 -82.795 -81.435 ;
        RECT -83.125 -83.125 -82.795 -82.795 ;
        RECT -83.125 -84.485 -82.795 -84.155 ;
        RECT -83.125 -85.845 -82.795 -85.515 ;
        RECT -83.125 -87.205 -82.795 -86.875 ;
        RECT -83.125 -88.565 -82.795 -88.235 ;
        RECT -83.125 -89.925 -82.795 -89.595 ;
        RECT -83.125 -91.285 -82.795 -90.955 ;
        RECT -83.125 -92.645 -82.795 -92.315 ;
        RECT -83.125 -94.005 -82.795 -93.675 ;
        RECT -83.125 -95.365 -82.795 -95.035 ;
        RECT -83.125 -96.725 -82.795 -96.395 ;
        RECT -83.125 -98.085 -82.795 -97.755 ;
        RECT -83.125 -99.445 -82.795 -99.115 ;
        RECT -83.125 -100.805 -82.795 -100.475 ;
        RECT -83.125 -102.165 -82.795 -101.835 ;
        RECT -83.125 -103.525 -82.795 -103.195 ;
        RECT -83.125 -104.885 -82.795 -104.555 ;
        RECT -83.125 -106.245 -82.795 -105.915 ;
        RECT -83.125 -107.605 -82.795 -107.275 ;
        RECT -83.125 -108.965 -82.795 -108.635 ;
        RECT -83.125 -110.325 -82.795 -109.995 ;
        RECT -83.125 -111.685 -82.795 -111.355 ;
        RECT -83.125 -113.045 -82.795 -112.715 ;
        RECT -83.125 -114.405 -82.795 -114.075 ;
        RECT -83.125 -115.765 -82.795 -115.435 ;
        RECT -83.125 -117.125 -82.795 -116.795 ;
        RECT -83.125 -118.485 -82.795 -118.155 ;
        RECT -83.125 -119.845 -82.795 -119.515 ;
        RECT -83.125 -121.205 -82.795 -120.875 ;
        RECT -83.125 -122.565 -82.795 -122.235 ;
        RECT -83.125 -123.925 -82.795 -123.595 ;
        RECT -83.125 -125.285 -82.795 -124.955 ;
        RECT -83.125 -126.645 -82.795 -126.315 ;
        RECT -83.125 -128.005 -82.795 -127.675 ;
        RECT -83.125 -129.365 -82.795 -129.035 ;
        RECT -83.125 -130.725 -82.795 -130.395 ;
        RECT -83.125 -132.085 -82.795 -131.755 ;
        RECT -83.125 -133.445 -82.795 -133.115 ;
        RECT -83.125 -134.805 -82.795 -134.475 ;
        RECT -83.125 -136.165 -82.795 -135.835 ;
        RECT -83.125 -137.525 -82.795 -137.195 ;
        RECT -83.125 -138.885 -82.795 -138.555 ;
        RECT -83.125 -140.245 -82.795 -139.915 ;
        RECT -83.125 -141.605 -82.795 -141.275 ;
        RECT -83.125 -142.965 -82.795 -142.635 ;
        RECT -83.125 -144.325 -82.795 -143.995 ;
        RECT -83.125 -145.685 -82.795 -145.355 ;
        RECT -83.125 -147.045 -82.795 -146.715 ;
        RECT -83.125 -148.405 -82.795 -148.075 ;
        RECT -83.125 -149.765 -82.795 -149.435 ;
        RECT -83.125 -151.125 -82.795 -150.795 ;
        RECT -83.125 -152.485 -82.795 -152.155 ;
        RECT -83.125 -153.845 -82.795 -153.515 ;
        RECT -83.125 -155.205 -82.795 -154.875 ;
        RECT -83.125 -156.565 -82.795 -156.235 ;
        RECT -83.125 -157.925 -82.795 -157.595 ;
        RECT -83.125 -159.285 -82.795 -158.955 ;
        RECT -83.125 -160.645 -82.795 -160.315 ;
        RECT -83.125 -162.005 -82.795 -161.675 ;
        RECT -83.125 -163.365 -82.795 -163.035 ;
        RECT -83.125 -164.725 -82.795 -164.395 ;
        RECT -83.125 -166.085 -82.795 -165.755 ;
        RECT -83.125 -167.445 -82.795 -167.115 ;
        RECT -83.125 -168.805 -82.795 -168.475 ;
        RECT -83.125 -170.165 -82.795 -169.835 ;
        RECT -83.125 -171.525 -82.795 -171.195 ;
        RECT -83.125 -172.885 -82.795 -172.555 ;
        RECT -83.125 -174.245 -82.795 -173.915 ;
        RECT -83.125 -175.605 -82.795 -175.275 ;
        RECT -83.125 -176.965 -82.795 -176.635 ;
        RECT -83.125 -178.325 -82.795 -177.995 ;
        RECT -83.125 -179.685 -82.795 -179.355 ;
        RECT -83.125 -181.045 -82.795 -180.715 ;
        RECT -83.125 -182.405 -82.795 -182.075 ;
        RECT -83.125 -183.765 -82.795 -183.435 ;
        RECT -83.125 -185.125 -82.795 -184.795 ;
        RECT -83.125 -186.485 -82.795 -186.155 ;
        RECT -83.125 -187.845 -82.795 -187.515 ;
        RECT -83.125 -189.205 -82.795 -188.875 ;
        RECT -83.125 -190.565 -82.795 -190.235 ;
        RECT -83.125 -191.925 -82.795 -191.595 ;
        RECT -83.125 -193.285 -82.795 -192.955 ;
        RECT -83.125 -194.645 -82.795 -194.315 ;
        RECT -83.125 -196.005 -82.795 -195.675 ;
        RECT -83.125 -197.365 -82.795 -197.035 ;
        RECT -83.125 -198.725 -82.795 -198.395 ;
        RECT -83.125 -200.085 -82.795 -199.755 ;
        RECT -83.125 -201.445 -82.795 -201.115 ;
        RECT -83.125 -202.805 -82.795 -202.475 ;
        RECT -83.125 -204.165 -82.795 -203.835 ;
        RECT -83.125 -205.525 -82.795 -205.195 ;
        RECT -83.125 -206.885 -82.795 -206.555 ;
        RECT -83.125 -208.245 -82.795 -207.915 ;
        RECT -83.125 -209.605 -82.795 -209.275 ;
        RECT -83.125 -210.965 -82.795 -210.635 ;
        RECT -83.125 -212.325 -82.795 -211.995 ;
        RECT -83.125 -213.685 -82.795 -213.355 ;
        RECT -83.125 -215.045 -82.795 -214.715 ;
        RECT -83.125 -216.405 -82.795 -216.075 ;
        RECT -83.125 -217.765 -82.795 -217.435 ;
        RECT -83.125 -219.125 -82.795 -218.795 ;
        RECT -83.125 -220.485 -82.795 -220.155 ;
        RECT -83.125 -221.845 -82.795 -221.515 ;
        RECT -83.125 -223.205 -82.795 -222.875 ;
        RECT -83.125 -224.565 -82.795 -224.235 ;
        RECT -83.125 -225.925 -82.795 -225.595 ;
        RECT -83.125 -227.285 -82.795 -226.955 ;
        RECT -83.125 -228.645 -82.795 -228.315 ;
        RECT -83.125 -230.005 -82.795 -229.675 ;
        RECT -83.125 -231.365 -82.795 -231.035 ;
        RECT -83.125 -232.725 -82.795 -232.395 ;
        RECT -83.125 -234.085 -82.795 -233.755 ;
        RECT -83.125 -235.445 -82.795 -235.115 ;
        RECT -83.125 -236.805 -82.795 -236.475 ;
        RECT -83.125 -238.165 -82.795 -237.835 ;
        RECT -83.125 -243.81 -82.795 -242.68 ;
        RECT -83.12 -243.925 -82.8 248.005 ;
        RECT -83.125 246.76 -82.795 247.89 ;
        RECT -83.125 241.915 -82.795 242.245 ;
        RECT -83.125 240.555 -82.795 240.885 ;
        RECT -83.125 239.195 -82.795 239.525 ;
        RECT -83.125 237.835 -82.795 238.165 ;
        RECT -83.125 236.475 -82.795 236.805 ;
        RECT -83.125 235.115 -82.795 235.445 ;
        RECT -83.125 233.755 -82.795 234.085 ;
        RECT -83.125 232.395 -82.795 232.725 ;
        RECT -83.125 231.035 -82.795 231.365 ;
        RECT -83.125 229.675 -82.795 230.005 ;
        RECT -83.125 228.315 -82.795 228.645 ;
        RECT -83.125 226.955 -82.795 227.285 ;
        RECT -83.125 225.595 -82.795 225.925 ;
        RECT -83.125 224.235 -82.795 224.565 ;
        RECT -83.125 222.875 -82.795 223.205 ;
        RECT -83.125 221.515 -82.795 221.845 ;
        RECT -83.125 220.155 -82.795 220.485 ;
        RECT -83.125 218.795 -82.795 219.125 ;
        RECT -83.125 217.435 -82.795 217.765 ;
        RECT -83.125 216.075 -82.795 216.405 ;
        RECT -83.125 214.715 -82.795 215.045 ;
        RECT -83.125 213.355 -82.795 213.685 ;
        RECT -83.125 211.995 -82.795 212.325 ;
        RECT -83.125 210.635 -82.795 210.965 ;
        RECT -83.125 209.275 -82.795 209.605 ;
        RECT -83.125 207.915 -82.795 208.245 ;
        RECT -83.125 206.555 -82.795 206.885 ;
        RECT -83.125 205.195 -82.795 205.525 ;
        RECT -83.125 203.835 -82.795 204.165 ;
        RECT -83.125 202.475 -82.795 202.805 ;
        RECT -83.125 201.115 -82.795 201.445 ;
        RECT -83.125 199.755 -82.795 200.085 ;
        RECT -83.125 198.395 -82.795 198.725 ;
        RECT -83.125 197.035 -82.795 197.365 ;
        RECT -83.125 195.675 -82.795 196.005 ;
        RECT -83.125 194.315 -82.795 194.645 ;
        RECT -83.125 192.955 -82.795 193.285 ;
        RECT -83.125 191.595 -82.795 191.925 ;
        RECT -83.125 190.235 -82.795 190.565 ;
        RECT -83.125 188.875 -82.795 189.205 ;
        RECT -83.125 187.515 -82.795 187.845 ;
        RECT -83.125 186.155 -82.795 186.485 ;
        RECT -83.125 184.795 -82.795 185.125 ;
        RECT -83.125 183.435 -82.795 183.765 ;
        RECT -83.125 182.075 -82.795 182.405 ;
        RECT -83.125 180.715 -82.795 181.045 ;
        RECT -83.125 179.355 -82.795 179.685 ;
        RECT -83.125 177.995 -82.795 178.325 ;
        RECT -83.125 176.635 -82.795 176.965 ;
        RECT -83.125 175.275 -82.795 175.605 ;
        RECT -83.125 173.915 -82.795 174.245 ;
        RECT -83.125 172.555 -82.795 172.885 ;
        RECT -83.125 171.195 -82.795 171.525 ;
        RECT -83.125 169.835 -82.795 170.165 ;
        RECT -83.125 168.475 -82.795 168.805 ;
        RECT -83.125 167.115 -82.795 167.445 ;
        RECT -83.125 165.755 -82.795 166.085 ;
        RECT -83.125 164.395 -82.795 164.725 ;
        RECT -83.125 163.035 -82.795 163.365 ;
        RECT -83.125 161.675 -82.795 162.005 ;
        RECT -83.125 160.315 -82.795 160.645 ;
        RECT -83.125 158.955 -82.795 159.285 ;
        RECT -83.125 157.595 -82.795 157.925 ;
        RECT -83.125 156.235 -82.795 156.565 ;
        RECT -83.125 154.875 -82.795 155.205 ;
        RECT -83.125 153.515 -82.795 153.845 ;
        RECT -83.125 152.155 -82.795 152.485 ;
        RECT -83.125 150.795 -82.795 151.125 ;
        RECT -83.125 149.435 -82.795 149.765 ;
        RECT -83.125 148.075 -82.795 148.405 ;
        RECT -83.125 146.715 -82.795 147.045 ;
        RECT -83.125 145.355 -82.795 145.685 ;
        RECT -83.125 143.995 -82.795 144.325 ;
        RECT -83.125 142.635 -82.795 142.965 ;
        RECT -83.125 141.275 -82.795 141.605 ;
        RECT -83.125 139.915 -82.795 140.245 ;
        RECT -83.125 138.555 -82.795 138.885 ;
        RECT -83.125 137.195 -82.795 137.525 ;
        RECT -83.125 135.835 -82.795 136.165 ;
        RECT -83.125 134.475 -82.795 134.805 ;
        RECT -83.125 133.115 -82.795 133.445 ;
        RECT -83.125 131.755 -82.795 132.085 ;
        RECT -83.125 130.395 -82.795 130.725 ;
        RECT -83.125 129.035 -82.795 129.365 ;
        RECT -83.125 127.675 -82.795 128.005 ;
        RECT -83.125 126.315 -82.795 126.645 ;
        RECT -83.125 124.955 -82.795 125.285 ;
        RECT -83.125 123.595 -82.795 123.925 ;
        RECT -83.125 122.235 -82.795 122.565 ;
        RECT -83.125 120.875 -82.795 121.205 ;
        RECT -83.125 119.515 -82.795 119.845 ;
        RECT -83.125 118.155 -82.795 118.485 ;
        RECT -83.125 116.795 -82.795 117.125 ;
        RECT -83.125 115.435 -82.795 115.765 ;
        RECT -83.125 114.075 -82.795 114.405 ;
        RECT -83.125 112.715 -82.795 113.045 ;
        RECT -83.125 111.355 -82.795 111.685 ;
        RECT -83.125 109.995 -82.795 110.325 ;
        RECT -83.125 108.635 -82.795 108.965 ;
        RECT -83.125 107.275 -82.795 107.605 ;
        RECT -83.125 105.915 -82.795 106.245 ;
        RECT -83.125 104.555 -82.795 104.885 ;
        RECT -83.125 103.195 -82.795 103.525 ;
        RECT -83.125 101.835 -82.795 102.165 ;
        RECT -83.125 100.475 -82.795 100.805 ;
        RECT -83.125 99.115 -82.795 99.445 ;
        RECT -83.125 97.755 -82.795 98.085 ;
        RECT -83.125 96.395 -82.795 96.725 ;
        RECT -83.125 95.035 -82.795 95.365 ;
        RECT -83.125 93.675 -82.795 94.005 ;
        RECT -83.125 92.315 -82.795 92.645 ;
        RECT -83.125 90.955 -82.795 91.285 ;
        RECT -83.125 89.595 -82.795 89.925 ;
        RECT -83.125 88.235 -82.795 88.565 ;
        RECT -83.125 86.875 -82.795 87.205 ;
        RECT -83.125 85.515 -82.795 85.845 ;
        RECT -83.125 84.155 -82.795 84.485 ;
        RECT -83.125 82.795 -82.795 83.125 ;
        RECT -83.125 81.435 -82.795 81.765 ;
        RECT -83.125 80.075 -82.795 80.405 ;
        RECT -83.125 78.715 -82.795 79.045 ;
        RECT -83.125 77.355 -82.795 77.685 ;
        RECT -83.125 75.995 -82.795 76.325 ;
        RECT -83.125 74.635 -82.795 74.965 ;
        RECT -83.125 73.275 -82.795 73.605 ;
        RECT -83.125 71.915 -82.795 72.245 ;
        RECT -83.125 70.555 -82.795 70.885 ;
        RECT -83.125 69.195 -82.795 69.525 ;
        RECT -83.125 67.835 -82.795 68.165 ;
        RECT -83.125 66.475 -82.795 66.805 ;
        RECT -83.125 65.115 -82.795 65.445 ;
        RECT -83.125 63.755 -82.795 64.085 ;
        RECT -83.125 62.395 -82.795 62.725 ;
        RECT -83.125 61.035 -82.795 61.365 ;
        RECT -83.125 59.675 -82.795 60.005 ;
        RECT -83.125 58.315 -82.795 58.645 ;
        RECT -83.125 56.955 -82.795 57.285 ;
        RECT -83.125 55.595 -82.795 55.925 ;
        RECT -83.125 54.235 -82.795 54.565 ;
        RECT -83.125 52.875 -82.795 53.205 ;
        RECT -83.125 51.515 -82.795 51.845 ;
        RECT -83.125 50.155 -82.795 50.485 ;
        RECT -83.125 48.795 -82.795 49.125 ;
        RECT -83.125 47.435 -82.795 47.765 ;
        RECT -83.125 46.075 -82.795 46.405 ;
        RECT -83.125 44.715 -82.795 45.045 ;
        RECT -83.125 43.355 -82.795 43.685 ;
        RECT -83.125 41.995 -82.795 42.325 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 360.915 244.04 361.245 245.17 ;
        RECT 360.915 242.595 361.245 242.925 ;
        RECT 360.915 241.235 361.245 241.565 ;
        RECT 360.915 239.875 361.245 240.205 ;
        RECT 360.915 238.515 361.245 238.845 ;
        RECT 360.915 237.155 361.245 237.485 ;
        RECT 360.915 -0.845 361.245 -0.515 ;
        RECT 360.915 -2.205 361.245 -1.875 ;
        RECT 360.915 -3.565 361.245 -3.235 ;
        RECT 360.915 -4.925 361.245 -4.595 ;
        RECT 360.915 -6.285 361.245 -5.955 ;
        RECT 360.915 -7.645 361.245 -7.315 ;
        RECT 360.915 -9.005 361.245 -8.675 ;
        RECT 360.915 -10.365 361.245 -10.035 ;
        RECT 360.915 -11.725 361.245 -11.395 ;
        RECT 360.915 -13.085 361.245 -12.755 ;
        RECT 360.915 -14.445 361.245 -14.115 ;
        RECT 360.915 -15.805 361.245 -15.475 ;
        RECT 360.915 -17.165 361.245 -16.835 ;
        RECT 360.915 -18.525 361.245 -18.195 ;
        RECT 360.915 -19.885 361.245 -19.555 ;
        RECT 360.915 -21.245 361.245 -20.915 ;
        RECT 360.915 -22.605 361.245 -22.275 ;
        RECT 360.915 -23.965 361.245 -23.635 ;
        RECT 360.915 -25.325 361.245 -24.995 ;
        RECT 360.915 -26.685 361.245 -26.355 ;
        RECT 360.915 -28.045 361.245 -27.715 ;
        RECT 360.915 -29.405 361.245 -29.075 ;
        RECT 360.915 -30.765 361.245 -30.435 ;
        RECT 360.915 -32.125 361.245 -31.795 ;
        RECT 360.915 -33.485 361.245 -33.155 ;
        RECT 360.915 -34.845 361.245 -34.515 ;
        RECT 360.915 -36.205 361.245 -35.875 ;
        RECT 360.915 -37.565 361.245 -37.235 ;
        RECT 360.915 -38.925 361.245 -38.595 ;
        RECT 360.915 -40.285 361.245 -39.955 ;
        RECT 360.915 -41.645 361.245 -41.315 ;
        RECT 360.915 -43.005 361.245 -42.675 ;
        RECT 360.915 -44.365 361.245 -44.035 ;
        RECT 360.915 -45.725 361.245 -45.395 ;
        RECT 360.915 -47.085 361.245 -46.755 ;
        RECT 360.915 -48.445 361.245 -48.115 ;
        RECT 360.915 -49.805 361.245 -49.475 ;
        RECT 360.915 -51.165 361.245 -50.835 ;
        RECT 360.915 -52.525 361.245 -52.195 ;
        RECT 360.915 -53.885 361.245 -53.555 ;
        RECT 360.915 -55.245 361.245 -54.915 ;
        RECT 360.915 -56.605 361.245 -56.275 ;
        RECT 360.915 -57.965 361.245 -57.635 ;
        RECT 360.915 -59.325 361.245 -58.995 ;
        RECT 360.915 -60.685 361.245 -60.355 ;
        RECT 360.915 -62.045 361.245 -61.715 ;
        RECT 360.915 -63.405 361.245 -63.075 ;
        RECT 360.915 -64.765 361.245 -64.435 ;
        RECT 360.915 -66.125 361.245 -65.795 ;
        RECT 360.915 -67.485 361.245 -67.155 ;
        RECT 360.915 -68.845 361.245 -68.515 ;
        RECT 360.915 -70.205 361.245 -69.875 ;
        RECT 360.915 -71.565 361.245 -71.235 ;
        RECT 360.915 -72.925 361.245 -72.595 ;
        RECT 360.915 -74.285 361.245 -73.955 ;
        RECT 360.915 -75.645 361.245 -75.315 ;
        RECT 360.915 -77.005 361.245 -76.675 ;
        RECT 360.915 -78.365 361.245 -78.035 ;
        RECT 360.915 -79.725 361.245 -79.395 ;
        RECT 360.915 -81.085 361.245 -80.755 ;
        RECT 360.915 -82.445 361.245 -82.115 ;
        RECT 360.915 -83.805 361.245 -83.475 ;
        RECT 360.915 -85.165 361.245 -84.835 ;
        RECT 360.915 -86.525 361.245 -86.195 ;
        RECT 360.915 -87.885 361.245 -87.555 ;
        RECT 360.915 -89.245 361.245 -88.915 ;
        RECT 360.915 -90.605 361.245 -90.275 ;
        RECT 360.915 -91.965 361.245 -91.635 ;
        RECT 360.915 -93.325 361.245 -92.995 ;
        RECT 360.915 -94.685 361.245 -94.355 ;
        RECT 360.915 -96.045 361.245 -95.715 ;
        RECT 360.915 -97.405 361.245 -97.075 ;
        RECT 360.915 -98.765 361.245 -98.435 ;
        RECT 360.915 -100.125 361.245 -99.795 ;
        RECT 360.915 -101.485 361.245 -101.155 ;
        RECT 360.915 -102.845 361.245 -102.515 ;
        RECT 360.915 -104.205 361.245 -103.875 ;
        RECT 360.915 -105.565 361.245 -105.235 ;
        RECT 360.915 -106.925 361.245 -106.595 ;
        RECT 360.915 -108.285 361.245 -107.955 ;
        RECT 360.915 -109.645 361.245 -109.315 ;
        RECT 360.915 -111.005 361.245 -110.675 ;
        RECT 360.915 -112.365 361.245 -112.035 ;
        RECT 360.915 -113.725 361.245 -113.395 ;
        RECT 360.915 -115.085 361.245 -114.755 ;
        RECT 360.915 -116.445 361.245 -116.115 ;
        RECT 360.915 -117.805 361.245 -117.475 ;
        RECT 360.915 -119.165 361.245 -118.835 ;
        RECT 360.915 -120.525 361.245 -120.195 ;
        RECT 360.915 -121.885 361.245 -121.555 ;
        RECT 360.915 -123.245 361.245 -122.915 ;
        RECT 360.915 -124.605 361.245 -124.275 ;
        RECT 360.915 -125.965 361.245 -125.635 ;
        RECT 360.915 -127.325 361.245 -126.995 ;
        RECT 360.915 -128.685 361.245 -128.355 ;
        RECT 360.915 -130.045 361.245 -129.715 ;
        RECT 360.915 -131.405 361.245 -131.075 ;
        RECT 360.915 -132.765 361.245 -132.435 ;
        RECT 360.915 -134.125 361.245 -133.795 ;
        RECT 360.915 -135.485 361.245 -135.155 ;
        RECT 360.915 -136.845 361.245 -136.515 ;
        RECT 360.915 -138.205 361.245 -137.875 ;
        RECT 360.915 -139.565 361.245 -139.235 ;
        RECT 360.915 -140.925 361.245 -140.595 ;
        RECT 360.915 -142.285 361.245 -141.955 ;
        RECT 360.915 -143.645 361.245 -143.315 ;
        RECT 360.915 -145.005 361.245 -144.675 ;
        RECT 360.915 -146.365 361.245 -146.035 ;
        RECT 360.915 -147.725 361.245 -147.395 ;
        RECT 360.915 -149.085 361.245 -148.755 ;
        RECT 360.915 -150.445 361.245 -150.115 ;
        RECT 360.915 -151.805 361.245 -151.475 ;
        RECT 360.915 -153.165 361.245 -152.835 ;
        RECT 360.915 -154.525 361.245 -154.195 ;
        RECT 360.915 -155.885 361.245 -155.555 ;
        RECT 360.915 -157.245 361.245 -156.915 ;
        RECT 360.915 -158.605 361.245 -158.275 ;
        RECT 360.915 -159.965 361.245 -159.635 ;
        RECT 360.915 -161.325 361.245 -160.995 ;
        RECT 360.915 -162.685 361.245 -162.355 ;
        RECT 360.915 -164.045 361.245 -163.715 ;
        RECT 360.915 -165.405 361.245 -165.075 ;
        RECT 360.915 -166.765 361.245 -166.435 ;
        RECT 360.915 -168.125 361.245 -167.795 ;
        RECT 360.915 -169.485 361.245 -169.155 ;
        RECT 360.915 -170.845 361.245 -170.515 ;
        RECT 360.915 -172.205 361.245 -171.875 ;
        RECT 360.915 -173.565 361.245 -173.235 ;
        RECT 360.915 -174.925 361.245 -174.595 ;
        RECT 360.915 -176.285 361.245 -175.955 ;
        RECT 360.915 -177.645 361.245 -177.315 ;
        RECT 360.915 -179.005 361.245 -178.675 ;
        RECT 360.915 -180.365 361.245 -180.035 ;
        RECT 360.915 -181.725 361.245 -181.395 ;
        RECT 360.915 -183.085 361.245 -182.755 ;
        RECT 360.915 -184.445 361.245 -184.115 ;
        RECT 360.915 -185.805 361.245 -185.475 ;
        RECT 360.915 -187.165 361.245 -186.835 ;
        RECT 360.915 -188.525 361.245 -188.195 ;
        RECT 360.915 -189.885 361.245 -189.555 ;
        RECT 360.915 -191.245 361.245 -190.915 ;
        RECT 360.915 -192.605 361.245 -192.275 ;
        RECT 360.915 -193.965 361.245 -193.635 ;
        RECT 360.915 -195.325 361.245 -194.995 ;
        RECT 360.915 -196.685 361.245 -196.355 ;
        RECT 360.915 -198.045 361.245 -197.715 ;
        RECT 360.915 -199.405 361.245 -199.075 ;
        RECT 360.915 -200.765 361.245 -200.435 ;
        RECT 360.915 -202.125 361.245 -201.795 ;
        RECT 360.915 -203.485 361.245 -203.155 ;
        RECT 360.915 -204.845 361.245 -204.515 ;
        RECT 360.915 -206.205 361.245 -205.875 ;
        RECT 360.915 -207.565 361.245 -207.235 ;
        RECT 360.915 -208.925 361.245 -208.595 ;
        RECT 360.915 -210.285 361.245 -209.955 ;
        RECT 360.915 -211.645 361.245 -211.315 ;
        RECT 360.915 -213.005 361.245 -212.675 ;
        RECT 360.915 -214.365 361.245 -214.035 ;
        RECT 360.915 -215.725 361.245 -215.395 ;
        RECT 360.915 -217.085 361.245 -216.755 ;
        RECT 360.915 -218.445 361.245 -218.115 ;
        RECT 360.915 -219.805 361.245 -219.475 ;
        RECT 360.915 -221.165 361.245 -220.835 ;
        RECT 360.915 -222.525 361.245 -222.195 ;
        RECT 360.915 -223.885 361.245 -223.555 ;
        RECT 360.915 -225.245 361.245 -224.915 ;
        RECT 360.915 -226.605 361.245 -226.275 ;
        RECT 360.915 -227.965 361.245 -227.635 ;
        RECT 360.915 -229.325 361.245 -228.995 ;
        RECT 360.915 -230.685 361.245 -230.355 ;
        RECT 360.915 -232.045 361.245 -231.715 ;
        RECT 360.915 -233.405 361.245 -233.075 ;
        RECT 360.915 -234.765 361.245 -234.435 ;
        RECT 360.915 -236.125 361.245 -235.795 ;
        RECT 360.915 -237.485 361.245 -237.155 ;
        RECT 360.915 -238.845 361.245 -238.515 ;
        RECT 360.915 -241.09 361.245 -239.96 ;
        RECT 360.92 -241.205 361.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.275 244.04 362.605 245.17 ;
        RECT 362.275 242.595 362.605 242.925 ;
        RECT 362.275 241.235 362.605 241.565 ;
        RECT 362.275 239.875 362.605 240.205 ;
        RECT 362.275 238.515 362.605 238.845 ;
        RECT 362.275 237.155 362.605 237.485 ;
        RECT 362.275 235.795 362.605 236.125 ;
        RECT 362.275 234.435 362.605 234.765 ;
        RECT 362.275 233.075 362.605 233.405 ;
        RECT 362.275 231.715 362.605 232.045 ;
        RECT 362.275 230.355 362.605 230.685 ;
        RECT 362.275 228.995 362.605 229.325 ;
        RECT 362.275 227.635 362.605 227.965 ;
        RECT 362.275 226.275 362.605 226.605 ;
        RECT 362.275 224.915 362.605 225.245 ;
        RECT 362.275 223.555 362.605 223.885 ;
        RECT 362.275 222.195 362.605 222.525 ;
        RECT 362.275 220.835 362.605 221.165 ;
        RECT 362.275 219.475 362.605 219.805 ;
        RECT 362.275 218.115 362.605 218.445 ;
        RECT 362.275 216.755 362.605 217.085 ;
        RECT 362.275 215.395 362.605 215.725 ;
        RECT 362.275 214.035 362.605 214.365 ;
        RECT 362.275 212.675 362.605 213.005 ;
        RECT 362.275 211.315 362.605 211.645 ;
        RECT 362.275 209.955 362.605 210.285 ;
        RECT 362.275 208.595 362.605 208.925 ;
        RECT 362.275 207.235 362.605 207.565 ;
        RECT 362.275 205.875 362.605 206.205 ;
        RECT 362.275 204.515 362.605 204.845 ;
        RECT 362.275 203.155 362.605 203.485 ;
        RECT 362.275 201.795 362.605 202.125 ;
        RECT 362.275 200.435 362.605 200.765 ;
        RECT 362.275 199.075 362.605 199.405 ;
        RECT 362.275 197.715 362.605 198.045 ;
        RECT 362.275 196.355 362.605 196.685 ;
        RECT 362.275 194.995 362.605 195.325 ;
        RECT 362.275 193.635 362.605 193.965 ;
        RECT 362.275 192.275 362.605 192.605 ;
        RECT 362.275 190.915 362.605 191.245 ;
        RECT 362.275 189.555 362.605 189.885 ;
        RECT 362.275 188.195 362.605 188.525 ;
        RECT 362.275 186.835 362.605 187.165 ;
        RECT 362.275 185.475 362.605 185.805 ;
        RECT 362.275 184.115 362.605 184.445 ;
        RECT 362.275 182.755 362.605 183.085 ;
        RECT 362.275 181.395 362.605 181.725 ;
        RECT 362.275 180.035 362.605 180.365 ;
        RECT 362.275 178.675 362.605 179.005 ;
        RECT 362.275 177.315 362.605 177.645 ;
        RECT 362.275 175.955 362.605 176.285 ;
        RECT 362.275 174.595 362.605 174.925 ;
        RECT 362.275 173.235 362.605 173.565 ;
        RECT 362.275 171.875 362.605 172.205 ;
        RECT 362.275 170.515 362.605 170.845 ;
        RECT 362.275 169.155 362.605 169.485 ;
        RECT 362.275 167.795 362.605 168.125 ;
        RECT 362.275 166.435 362.605 166.765 ;
        RECT 362.275 165.075 362.605 165.405 ;
        RECT 362.275 163.715 362.605 164.045 ;
        RECT 362.275 162.355 362.605 162.685 ;
        RECT 362.275 160.995 362.605 161.325 ;
        RECT 362.275 159.635 362.605 159.965 ;
        RECT 362.275 158.275 362.605 158.605 ;
        RECT 362.275 156.915 362.605 157.245 ;
        RECT 362.275 155.555 362.605 155.885 ;
        RECT 362.275 154.195 362.605 154.525 ;
        RECT 362.275 152.835 362.605 153.165 ;
        RECT 362.275 151.475 362.605 151.805 ;
        RECT 362.275 150.115 362.605 150.445 ;
        RECT 362.275 148.755 362.605 149.085 ;
        RECT 362.275 147.395 362.605 147.725 ;
        RECT 362.275 146.035 362.605 146.365 ;
        RECT 362.275 144.675 362.605 145.005 ;
        RECT 362.275 143.315 362.605 143.645 ;
        RECT 362.275 141.955 362.605 142.285 ;
        RECT 362.275 140.595 362.605 140.925 ;
        RECT 362.275 139.235 362.605 139.565 ;
        RECT 362.275 137.875 362.605 138.205 ;
        RECT 362.275 136.515 362.605 136.845 ;
        RECT 362.275 135.155 362.605 135.485 ;
        RECT 362.275 133.795 362.605 134.125 ;
        RECT 362.275 132.435 362.605 132.765 ;
        RECT 362.275 131.075 362.605 131.405 ;
        RECT 362.275 129.715 362.605 130.045 ;
        RECT 362.275 128.355 362.605 128.685 ;
        RECT 362.275 126.995 362.605 127.325 ;
        RECT 362.275 125.635 362.605 125.965 ;
        RECT 362.275 124.275 362.605 124.605 ;
        RECT 362.275 122.915 362.605 123.245 ;
        RECT 362.275 121.555 362.605 121.885 ;
        RECT 362.275 120.195 362.605 120.525 ;
        RECT 362.275 118.835 362.605 119.165 ;
        RECT 362.275 117.475 362.605 117.805 ;
        RECT 362.275 116.115 362.605 116.445 ;
        RECT 362.275 114.755 362.605 115.085 ;
        RECT 362.275 113.395 362.605 113.725 ;
        RECT 362.275 112.035 362.605 112.365 ;
        RECT 362.275 110.675 362.605 111.005 ;
        RECT 362.275 109.315 362.605 109.645 ;
        RECT 362.275 107.955 362.605 108.285 ;
        RECT 362.275 106.595 362.605 106.925 ;
        RECT 362.275 105.235 362.605 105.565 ;
        RECT 362.275 103.875 362.605 104.205 ;
        RECT 362.275 102.515 362.605 102.845 ;
        RECT 362.275 101.155 362.605 101.485 ;
        RECT 362.275 99.795 362.605 100.125 ;
        RECT 362.275 98.435 362.605 98.765 ;
        RECT 362.275 97.075 362.605 97.405 ;
        RECT 362.275 95.715 362.605 96.045 ;
        RECT 362.275 94.355 362.605 94.685 ;
        RECT 362.275 92.995 362.605 93.325 ;
        RECT 362.275 91.635 362.605 91.965 ;
        RECT 362.275 90.275 362.605 90.605 ;
        RECT 362.275 88.915 362.605 89.245 ;
        RECT 362.275 87.555 362.605 87.885 ;
        RECT 362.275 86.195 362.605 86.525 ;
        RECT 362.275 84.835 362.605 85.165 ;
        RECT 362.275 83.475 362.605 83.805 ;
        RECT 362.275 82.115 362.605 82.445 ;
        RECT 362.275 80.755 362.605 81.085 ;
        RECT 362.275 79.395 362.605 79.725 ;
        RECT 362.275 78.035 362.605 78.365 ;
        RECT 362.275 76.675 362.605 77.005 ;
        RECT 362.275 75.315 362.605 75.645 ;
        RECT 362.275 73.955 362.605 74.285 ;
        RECT 362.275 72.595 362.605 72.925 ;
        RECT 362.275 71.235 362.605 71.565 ;
        RECT 362.275 69.875 362.605 70.205 ;
        RECT 362.275 68.515 362.605 68.845 ;
        RECT 362.275 67.155 362.605 67.485 ;
        RECT 362.275 65.795 362.605 66.125 ;
        RECT 362.275 64.435 362.605 64.765 ;
        RECT 362.275 63.075 362.605 63.405 ;
        RECT 362.275 61.715 362.605 62.045 ;
        RECT 362.275 60.355 362.605 60.685 ;
        RECT 362.275 58.995 362.605 59.325 ;
        RECT 362.275 57.635 362.605 57.965 ;
        RECT 362.275 56.275 362.605 56.605 ;
        RECT 362.275 54.915 362.605 55.245 ;
        RECT 362.275 53.555 362.605 53.885 ;
        RECT 362.275 52.195 362.605 52.525 ;
        RECT 362.275 50.835 362.605 51.165 ;
        RECT 362.275 49.475 362.605 49.805 ;
        RECT 362.275 48.115 362.605 48.445 ;
        RECT 362.275 46.755 362.605 47.085 ;
        RECT 362.275 45.395 362.605 45.725 ;
        RECT 362.275 44.035 362.605 44.365 ;
        RECT 362.275 42.675 362.605 43.005 ;
        RECT 362.275 41.315 362.605 41.645 ;
        RECT 362.275 39.955 362.605 40.285 ;
        RECT 362.275 38.595 362.605 38.925 ;
        RECT 362.275 37.235 362.605 37.565 ;
        RECT 362.275 35.875 362.605 36.205 ;
        RECT 362.275 34.515 362.605 34.845 ;
        RECT 362.275 33.155 362.605 33.485 ;
        RECT 362.275 31.795 362.605 32.125 ;
        RECT 362.275 30.435 362.605 30.765 ;
        RECT 362.275 29.075 362.605 29.405 ;
        RECT 362.275 27.715 362.605 28.045 ;
        RECT 362.275 26.355 362.605 26.685 ;
        RECT 362.275 24.995 362.605 25.325 ;
        RECT 362.275 23.635 362.605 23.965 ;
        RECT 362.275 22.275 362.605 22.605 ;
        RECT 362.275 20.915 362.605 21.245 ;
        RECT 362.275 19.555 362.605 19.885 ;
        RECT 362.275 18.195 362.605 18.525 ;
        RECT 362.275 16.835 362.605 17.165 ;
        RECT 362.275 15.475 362.605 15.805 ;
        RECT 362.275 14.115 362.605 14.445 ;
        RECT 362.275 12.755 362.605 13.085 ;
        RECT 362.275 11.395 362.605 11.725 ;
        RECT 362.275 10.035 362.605 10.365 ;
        RECT 362.275 8.675 362.605 9.005 ;
        RECT 362.275 7.315 362.605 7.645 ;
        RECT 362.275 5.955 362.605 6.285 ;
        RECT 362.275 4.595 362.605 4.925 ;
        RECT 362.275 3.235 362.605 3.565 ;
        RECT 362.275 1.875 362.605 2.205 ;
        RECT 362.275 0.515 362.605 0.845 ;
        RECT 362.275 -0.845 362.605 -0.515 ;
        RECT 362.275 -2.205 362.605 -1.875 ;
        RECT 362.275 -3.565 362.605 -3.235 ;
        RECT 362.275 -4.925 362.605 -4.595 ;
        RECT 362.275 -6.285 362.605 -5.955 ;
        RECT 362.275 -7.645 362.605 -7.315 ;
        RECT 362.275 -9.005 362.605 -8.675 ;
        RECT 362.275 -10.365 362.605 -10.035 ;
        RECT 362.275 -11.725 362.605 -11.395 ;
        RECT 362.275 -13.085 362.605 -12.755 ;
        RECT 362.275 -14.445 362.605 -14.115 ;
        RECT 362.275 -15.805 362.605 -15.475 ;
        RECT 362.275 -17.165 362.605 -16.835 ;
        RECT 362.275 -18.525 362.605 -18.195 ;
        RECT 362.275 -19.885 362.605 -19.555 ;
        RECT 362.275 -21.245 362.605 -20.915 ;
        RECT 362.275 -22.605 362.605 -22.275 ;
        RECT 362.275 -23.965 362.605 -23.635 ;
        RECT 362.275 -25.325 362.605 -24.995 ;
        RECT 362.275 -26.685 362.605 -26.355 ;
        RECT 362.275 -28.045 362.605 -27.715 ;
        RECT 362.275 -29.405 362.605 -29.075 ;
        RECT 362.275 -30.765 362.605 -30.435 ;
        RECT 362.275 -32.125 362.605 -31.795 ;
        RECT 362.275 -33.485 362.605 -33.155 ;
        RECT 362.275 -34.845 362.605 -34.515 ;
        RECT 362.275 -36.205 362.605 -35.875 ;
        RECT 362.275 -37.565 362.605 -37.235 ;
        RECT 362.275 -38.925 362.605 -38.595 ;
        RECT 362.275 -40.285 362.605 -39.955 ;
        RECT 362.275 -41.645 362.605 -41.315 ;
        RECT 362.275 -43.005 362.605 -42.675 ;
        RECT 362.275 -44.365 362.605 -44.035 ;
        RECT 362.275 -45.725 362.605 -45.395 ;
        RECT 362.275 -47.085 362.605 -46.755 ;
        RECT 362.275 -48.445 362.605 -48.115 ;
        RECT 362.275 -49.805 362.605 -49.475 ;
        RECT 362.275 -51.165 362.605 -50.835 ;
        RECT 362.275 -52.525 362.605 -52.195 ;
        RECT 362.275 -53.885 362.605 -53.555 ;
        RECT 362.275 -55.245 362.605 -54.915 ;
        RECT 362.275 -56.605 362.605 -56.275 ;
        RECT 362.275 -57.965 362.605 -57.635 ;
        RECT 362.275 -59.325 362.605 -58.995 ;
        RECT 362.275 -60.685 362.605 -60.355 ;
        RECT 362.275 -62.045 362.605 -61.715 ;
        RECT 362.275 -63.405 362.605 -63.075 ;
        RECT 362.275 -64.765 362.605 -64.435 ;
        RECT 362.275 -66.125 362.605 -65.795 ;
        RECT 362.275 -67.485 362.605 -67.155 ;
        RECT 362.275 -68.845 362.605 -68.515 ;
        RECT 362.275 -70.205 362.605 -69.875 ;
        RECT 362.275 -71.565 362.605 -71.235 ;
        RECT 362.275 -72.925 362.605 -72.595 ;
        RECT 362.275 -74.285 362.605 -73.955 ;
        RECT 362.275 -75.645 362.605 -75.315 ;
        RECT 362.275 -77.005 362.605 -76.675 ;
        RECT 362.275 -78.365 362.605 -78.035 ;
        RECT 362.275 -79.725 362.605 -79.395 ;
        RECT 362.275 -81.085 362.605 -80.755 ;
        RECT 362.275 -82.445 362.605 -82.115 ;
        RECT 362.275 -83.805 362.605 -83.475 ;
        RECT 362.275 -85.165 362.605 -84.835 ;
        RECT 362.275 -86.525 362.605 -86.195 ;
        RECT 362.275 -87.885 362.605 -87.555 ;
        RECT 362.275 -89.245 362.605 -88.915 ;
        RECT 362.275 -90.605 362.605 -90.275 ;
        RECT 362.275 -91.965 362.605 -91.635 ;
        RECT 362.275 -93.325 362.605 -92.995 ;
        RECT 362.275 -94.685 362.605 -94.355 ;
        RECT 362.275 -96.045 362.605 -95.715 ;
        RECT 362.275 -97.405 362.605 -97.075 ;
        RECT 362.275 -98.765 362.605 -98.435 ;
        RECT 362.275 -100.125 362.605 -99.795 ;
        RECT 362.275 -101.485 362.605 -101.155 ;
        RECT 362.275 -102.845 362.605 -102.515 ;
        RECT 362.275 -104.205 362.605 -103.875 ;
        RECT 362.275 -105.565 362.605 -105.235 ;
        RECT 362.275 -106.925 362.605 -106.595 ;
        RECT 362.275 -108.285 362.605 -107.955 ;
        RECT 362.275 -109.645 362.605 -109.315 ;
        RECT 362.275 -111.005 362.605 -110.675 ;
        RECT 362.275 -112.365 362.605 -112.035 ;
        RECT 362.275 -113.725 362.605 -113.395 ;
        RECT 362.275 -115.085 362.605 -114.755 ;
        RECT 362.275 -116.445 362.605 -116.115 ;
        RECT 362.275 -117.805 362.605 -117.475 ;
        RECT 362.275 -119.165 362.605 -118.835 ;
        RECT 362.275 -120.525 362.605 -120.195 ;
        RECT 362.275 -121.885 362.605 -121.555 ;
        RECT 362.275 -123.245 362.605 -122.915 ;
        RECT 362.275 -124.605 362.605 -124.275 ;
        RECT 362.275 -125.965 362.605 -125.635 ;
        RECT 362.275 -127.325 362.605 -126.995 ;
        RECT 362.275 -128.685 362.605 -128.355 ;
        RECT 362.275 -130.045 362.605 -129.715 ;
        RECT 362.275 -131.405 362.605 -131.075 ;
        RECT 362.275 -132.765 362.605 -132.435 ;
        RECT 362.275 -134.125 362.605 -133.795 ;
        RECT 362.275 -135.485 362.605 -135.155 ;
        RECT 362.275 -136.845 362.605 -136.515 ;
        RECT 362.275 -138.205 362.605 -137.875 ;
        RECT 362.275 -139.565 362.605 -139.235 ;
        RECT 362.275 -140.925 362.605 -140.595 ;
        RECT 362.275 -142.285 362.605 -141.955 ;
        RECT 362.275 -143.645 362.605 -143.315 ;
        RECT 362.275 -145.005 362.605 -144.675 ;
        RECT 362.275 -146.365 362.605 -146.035 ;
        RECT 362.275 -147.725 362.605 -147.395 ;
        RECT 362.275 -149.085 362.605 -148.755 ;
        RECT 362.275 -150.445 362.605 -150.115 ;
        RECT 362.275 -151.805 362.605 -151.475 ;
        RECT 362.275 -153.165 362.605 -152.835 ;
        RECT 362.275 -154.525 362.605 -154.195 ;
        RECT 362.275 -155.885 362.605 -155.555 ;
        RECT 362.275 -157.245 362.605 -156.915 ;
        RECT 362.275 -158.605 362.605 -158.275 ;
        RECT 362.275 -159.965 362.605 -159.635 ;
        RECT 362.275 -161.325 362.605 -160.995 ;
        RECT 362.275 -162.685 362.605 -162.355 ;
        RECT 362.275 -164.045 362.605 -163.715 ;
        RECT 362.275 -165.405 362.605 -165.075 ;
        RECT 362.275 -166.765 362.605 -166.435 ;
        RECT 362.275 -168.125 362.605 -167.795 ;
        RECT 362.275 -169.485 362.605 -169.155 ;
        RECT 362.275 -170.845 362.605 -170.515 ;
        RECT 362.275 -172.205 362.605 -171.875 ;
        RECT 362.275 -173.565 362.605 -173.235 ;
        RECT 362.275 -174.925 362.605 -174.595 ;
        RECT 362.275 -176.285 362.605 -175.955 ;
        RECT 362.275 -177.645 362.605 -177.315 ;
        RECT 362.275 -179.005 362.605 -178.675 ;
        RECT 362.275 -180.365 362.605 -180.035 ;
        RECT 362.275 -181.725 362.605 -181.395 ;
        RECT 362.275 -183.085 362.605 -182.755 ;
        RECT 362.275 -184.445 362.605 -184.115 ;
        RECT 362.275 -185.805 362.605 -185.475 ;
        RECT 362.275 -187.165 362.605 -186.835 ;
        RECT 362.275 -188.525 362.605 -188.195 ;
        RECT 362.275 -189.885 362.605 -189.555 ;
        RECT 362.275 -191.245 362.605 -190.915 ;
        RECT 362.275 -192.605 362.605 -192.275 ;
        RECT 362.275 -193.965 362.605 -193.635 ;
        RECT 362.275 -195.325 362.605 -194.995 ;
        RECT 362.275 -196.685 362.605 -196.355 ;
        RECT 362.275 -198.045 362.605 -197.715 ;
        RECT 362.275 -199.405 362.605 -199.075 ;
        RECT 362.275 -200.765 362.605 -200.435 ;
        RECT 362.275 -202.125 362.605 -201.795 ;
        RECT 362.275 -203.485 362.605 -203.155 ;
        RECT 362.275 -204.845 362.605 -204.515 ;
        RECT 362.275 -206.205 362.605 -205.875 ;
        RECT 362.275 -207.565 362.605 -207.235 ;
        RECT 362.275 -208.925 362.605 -208.595 ;
        RECT 362.275 -210.285 362.605 -209.955 ;
        RECT 362.275 -211.645 362.605 -211.315 ;
        RECT 362.275 -213.005 362.605 -212.675 ;
        RECT 362.275 -214.365 362.605 -214.035 ;
        RECT 362.275 -215.725 362.605 -215.395 ;
        RECT 362.275 -217.085 362.605 -216.755 ;
        RECT 362.275 -218.445 362.605 -218.115 ;
        RECT 362.275 -219.805 362.605 -219.475 ;
        RECT 362.275 -221.165 362.605 -220.835 ;
        RECT 362.275 -222.525 362.605 -222.195 ;
        RECT 362.275 -223.885 362.605 -223.555 ;
        RECT 362.275 -225.245 362.605 -224.915 ;
        RECT 362.275 -226.605 362.605 -226.275 ;
        RECT 362.275 -227.965 362.605 -227.635 ;
        RECT 362.275 -229.325 362.605 -228.995 ;
        RECT 362.275 -230.685 362.605 -230.355 ;
        RECT 362.275 -232.045 362.605 -231.715 ;
        RECT 362.275 -233.405 362.605 -233.075 ;
        RECT 362.275 -234.765 362.605 -234.435 ;
        RECT 362.275 -236.125 362.605 -235.795 ;
        RECT 362.275 -237.485 362.605 -237.155 ;
        RECT 362.275 -238.845 362.605 -238.515 ;
        RECT 362.275 -241.09 362.605 -239.96 ;
        RECT 362.28 -241.205 362.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.635 244.04 363.965 245.17 ;
        RECT 363.635 242.595 363.965 242.925 ;
        RECT 363.635 241.235 363.965 241.565 ;
        RECT 363.635 239.875 363.965 240.205 ;
        RECT 363.635 238.515 363.965 238.845 ;
        RECT 363.635 237.155 363.965 237.485 ;
        RECT 363.635 235.795 363.965 236.125 ;
        RECT 363.635 234.435 363.965 234.765 ;
        RECT 363.635 233.075 363.965 233.405 ;
        RECT 363.635 231.715 363.965 232.045 ;
        RECT 363.635 230.355 363.965 230.685 ;
        RECT 363.635 228.995 363.965 229.325 ;
        RECT 363.635 227.635 363.965 227.965 ;
        RECT 363.635 226.275 363.965 226.605 ;
        RECT 363.635 224.915 363.965 225.245 ;
        RECT 363.635 223.555 363.965 223.885 ;
        RECT 363.635 222.195 363.965 222.525 ;
        RECT 363.635 220.835 363.965 221.165 ;
        RECT 363.635 219.475 363.965 219.805 ;
        RECT 363.635 218.115 363.965 218.445 ;
        RECT 363.635 216.755 363.965 217.085 ;
        RECT 363.635 215.395 363.965 215.725 ;
        RECT 363.635 214.035 363.965 214.365 ;
        RECT 363.635 212.675 363.965 213.005 ;
        RECT 363.635 211.315 363.965 211.645 ;
        RECT 363.635 209.955 363.965 210.285 ;
        RECT 363.635 208.595 363.965 208.925 ;
        RECT 363.635 207.235 363.965 207.565 ;
        RECT 363.635 205.875 363.965 206.205 ;
        RECT 363.635 204.515 363.965 204.845 ;
        RECT 363.635 203.155 363.965 203.485 ;
        RECT 363.635 201.795 363.965 202.125 ;
        RECT 363.635 200.435 363.965 200.765 ;
        RECT 363.635 199.075 363.965 199.405 ;
        RECT 363.635 197.715 363.965 198.045 ;
        RECT 363.635 196.355 363.965 196.685 ;
        RECT 363.635 194.995 363.965 195.325 ;
        RECT 363.635 193.635 363.965 193.965 ;
        RECT 363.635 192.275 363.965 192.605 ;
        RECT 363.635 190.915 363.965 191.245 ;
        RECT 363.635 189.555 363.965 189.885 ;
        RECT 363.635 188.195 363.965 188.525 ;
        RECT 363.635 186.835 363.965 187.165 ;
        RECT 363.635 185.475 363.965 185.805 ;
        RECT 363.635 184.115 363.965 184.445 ;
        RECT 363.635 182.755 363.965 183.085 ;
        RECT 363.635 181.395 363.965 181.725 ;
        RECT 363.635 180.035 363.965 180.365 ;
        RECT 363.635 178.675 363.965 179.005 ;
        RECT 363.635 177.315 363.965 177.645 ;
        RECT 363.635 175.955 363.965 176.285 ;
        RECT 363.635 174.595 363.965 174.925 ;
        RECT 363.635 173.235 363.965 173.565 ;
        RECT 363.635 171.875 363.965 172.205 ;
        RECT 363.635 170.515 363.965 170.845 ;
        RECT 363.635 169.155 363.965 169.485 ;
        RECT 363.635 167.795 363.965 168.125 ;
        RECT 363.635 166.435 363.965 166.765 ;
        RECT 363.635 165.075 363.965 165.405 ;
        RECT 363.635 163.715 363.965 164.045 ;
        RECT 363.635 162.355 363.965 162.685 ;
        RECT 363.635 160.995 363.965 161.325 ;
        RECT 363.635 159.635 363.965 159.965 ;
        RECT 363.635 158.275 363.965 158.605 ;
        RECT 363.635 156.915 363.965 157.245 ;
        RECT 363.635 155.555 363.965 155.885 ;
        RECT 363.635 154.195 363.965 154.525 ;
        RECT 363.635 152.835 363.965 153.165 ;
        RECT 363.635 151.475 363.965 151.805 ;
        RECT 363.635 150.115 363.965 150.445 ;
        RECT 363.635 148.755 363.965 149.085 ;
        RECT 363.635 147.395 363.965 147.725 ;
        RECT 363.635 146.035 363.965 146.365 ;
        RECT 363.635 144.675 363.965 145.005 ;
        RECT 363.635 143.315 363.965 143.645 ;
        RECT 363.635 141.955 363.965 142.285 ;
        RECT 363.635 140.595 363.965 140.925 ;
        RECT 363.635 139.235 363.965 139.565 ;
        RECT 363.635 137.875 363.965 138.205 ;
        RECT 363.635 136.515 363.965 136.845 ;
        RECT 363.635 135.155 363.965 135.485 ;
        RECT 363.635 133.795 363.965 134.125 ;
        RECT 363.635 132.435 363.965 132.765 ;
        RECT 363.635 131.075 363.965 131.405 ;
        RECT 363.635 129.715 363.965 130.045 ;
        RECT 363.635 128.355 363.965 128.685 ;
        RECT 363.635 126.995 363.965 127.325 ;
        RECT 363.635 125.635 363.965 125.965 ;
        RECT 363.635 124.275 363.965 124.605 ;
        RECT 363.635 122.915 363.965 123.245 ;
        RECT 363.635 121.555 363.965 121.885 ;
        RECT 363.635 120.195 363.965 120.525 ;
        RECT 363.635 118.835 363.965 119.165 ;
        RECT 363.635 117.475 363.965 117.805 ;
        RECT 363.635 116.115 363.965 116.445 ;
        RECT 363.635 114.755 363.965 115.085 ;
        RECT 363.635 113.395 363.965 113.725 ;
        RECT 363.635 112.035 363.965 112.365 ;
        RECT 363.635 110.675 363.965 111.005 ;
        RECT 363.635 109.315 363.965 109.645 ;
        RECT 363.635 107.955 363.965 108.285 ;
        RECT 363.635 106.595 363.965 106.925 ;
        RECT 363.635 105.235 363.965 105.565 ;
        RECT 363.635 103.875 363.965 104.205 ;
        RECT 363.635 102.515 363.965 102.845 ;
        RECT 363.635 101.155 363.965 101.485 ;
        RECT 363.635 99.795 363.965 100.125 ;
        RECT 363.635 98.435 363.965 98.765 ;
        RECT 363.635 97.075 363.965 97.405 ;
        RECT 363.635 95.715 363.965 96.045 ;
        RECT 363.635 94.355 363.965 94.685 ;
        RECT 363.635 92.995 363.965 93.325 ;
        RECT 363.635 91.635 363.965 91.965 ;
        RECT 363.635 90.275 363.965 90.605 ;
        RECT 363.635 88.915 363.965 89.245 ;
        RECT 363.635 87.555 363.965 87.885 ;
        RECT 363.635 86.195 363.965 86.525 ;
        RECT 363.635 84.835 363.965 85.165 ;
        RECT 363.635 83.475 363.965 83.805 ;
        RECT 363.635 82.115 363.965 82.445 ;
        RECT 363.635 80.755 363.965 81.085 ;
        RECT 363.635 79.395 363.965 79.725 ;
        RECT 363.635 78.035 363.965 78.365 ;
        RECT 363.635 76.675 363.965 77.005 ;
        RECT 363.635 75.315 363.965 75.645 ;
        RECT 363.635 73.955 363.965 74.285 ;
        RECT 363.635 72.595 363.965 72.925 ;
        RECT 363.635 71.235 363.965 71.565 ;
        RECT 363.635 69.875 363.965 70.205 ;
        RECT 363.635 68.515 363.965 68.845 ;
        RECT 363.635 67.155 363.965 67.485 ;
        RECT 363.635 65.795 363.965 66.125 ;
        RECT 363.635 64.435 363.965 64.765 ;
        RECT 363.635 63.075 363.965 63.405 ;
        RECT 363.635 61.715 363.965 62.045 ;
        RECT 363.635 60.355 363.965 60.685 ;
        RECT 363.635 58.995 363.965 59.325 ;
        RECT 363.635 57.635 363.965 57.965 ;
        RECT 363.635 56.275 363.965 56.605 ;
        RECT 363.635 54.915 363.965 55.245 ;
        RECT 363.635 53.555 363.965 53.885 ;
        RECT 363.635 52.195 363.965 52.525 ;
        RECT 363.635 50.835 363.965 51.165 ;
        RECT 363.635 49.475 363.965 49.805 ;
        RECT 363.635 48.115 363.965 48.445 ;
        RECT 363.635 46.755 363.965 47.085 ;
        RECT 363.635 45.395 363.965 45.725 ;
        RECT 363.635 44.035 363.965 44.365 ;
        RECT 363.635 42.675 363.965 43.005 ;
        RECT 363.635 41.315 363.965 41.645 ;
        RECT 363.635 39.955 363.965 40.285 ;
        RECT 363.635 38.595 363.965 38.925 ;
        RECT 363.635 37.235 363.965 37.565 ;
        RECT 363.635 35.875 363.965 36.205 ;
        RECT 363.635 34.515 363.965 34.845 ;
        RECT 363.635 33.155 363.965 33.485 ;
        RECT 363.635 31.795 363.965 32.125 ;
        RECT 363.635 30.435 363.965 30.765 ;
        RECT 363.635 29.075 363.965 29.405 ;
        RECT 363.635 27.715 363.965 28.045 ;
        RECT 363.635 26.355 363.965 26.685 ;
        RECT 363.635 24.995 363.965 25.325 ;
        RECT 363.635 23.635 363.965 23.965 ;
        RECT 363.635 22.275 363.965 22.605 ;
        RECT 363.635 20.915 363.965 21.245 ;
        RECT 363.635 19.555 363.965 19.885 ;
        RECT 363.635 18.195 363.965 18.525 ;
        RECT 363.635 16.835 363.965 17.165 ;
        RECT 363.635 15.475 363.965 15.805 ;
        RECT 363.635 14.115 363.965 14.445 ;
        RECT 363.635 12.755 363.965 13.085 ;
        RECT 363.635 11.395 363.965 11.725 ;
        RECT 363.635 10.035 363.965 10.365 ;
        RECT 363.635 8.675 363.965 9.005 ;
        RECT 363.635 7.315 363.965 7.645 ;
        RECT 363.635 5.955 363.965 6.285 ;
        RECT 363.635 4.595 363.965 4.925 ;
        RECT 363.635 3.235 363.965 3.565 ;
        RECT 363.635 1.875 363.965 2.205 ;
        RECT 363.635 0.515 363.965 0.845 ;
        RECT 363.635 -0.845 363.965 -0.515 ;
        RECT 363.635 -2.205 363.965 -1.875 ;
        RECT 363.635 -3.565 363.965 -3.235 ;
        RECT 363.635 -4.925 363.965 -4.595 ;
        RECT 363.635 -6.285 363.965 -5.955 ;
        RECT 363.635 -7.645 363.965 -7.315 ;
        RECT 363.635 -9.005 363.965 -8.675 ;
        RECT 363.635 -10.365 363.965 -10.035 ;
        RECT 363.635 -11.725 363.965 -11.395 ;
        RECT 363.635 -13.085 363.965 -12.755 ;
        RECT 363.635 -14.445 363.965 -14.115 ;
        RECT 363.635 -15.805 363.965 -15.475 ;
        RECT 363.635 -17.165 363.965 -16.835 ;
        RECT 363.635 -18.525 363.965 -18.195 ;
        RECT 363.635 -19.885 363.965 -19.555 ;
        RECT 363.635 -21.245 363.965 -20.915 ;
        RECT 363.635 -22.605 363.965 -22.275 ;
        RECT 363.635 -23.965 363.965 -23.635 ;
        RECT 363.635 -25.325 363.965 -24.995 ;
        RECT 363.635 -26.685 363.965 -26.355 ;
        RECT 363.635 -28.045 363.965 -27.715 ;
        RECT 363.635 -29.405 363.965 -29.075 ;
        RECT 363.635 -30.765 363.965 -30.435 ;
        RECT 363.635 -32.125 363.965 -31.795 ;
        RECT 363.635 -33.485 363.965 -33.155 ;
        RECT 363.635 -34.845 363.965 -34.515 ;
        RECT 363.635 -36.205 363.965 -35.875 ;
        RECT 363.635 -37.565 363.965 -37.235 ;
        RECT 363.635 -38.925 363.965 -38.595 ;
        RECT 363.635 -40.285 363.965 -39.955 ;
        RECT 363.635 -41.645 363.965 -41.315 ;
        RECT 363.635 -43.005 363.965 -42.675 ;
        RECT 363.635 -44.365 363.965 -44.035 ;
        RECT 363.635 -45.725 363.965 -45.395 ;
        RECT 363.635 -47.085 363.965 -46.755 ;
        RECT 363.635 -48.445 363.965 -48.115 ;
        RECT 363.635 -49.805 363.965 -49.475 ;
        RECT 363.635 -51.165 363.965 -50.835 ;
        RECT 363.635 -52.525 363.965 -52.195 ;
        RECT 363.635 -53.885 363.965 -53.555 ;
        RECT 363.635 -55.245 363.965 -54.915 ;
        RECT 363.635 -56.605 363.965 -56.275 ;
        RECT 363.635 -57.965 363.965 -57.635 ;
        RECT 363.635 -59.325 363.965 -58.995 ;
        RECT 363.635 -60.685 363.965 -60.355 ;
        RECT 363.635 -62.045 363.965 -61.715 ;
        RECT 363.635 -63.405 363.965 -63.075 ;
        RECT 363.635 -64.765 363.965 -64.435 ;
        RECT 363.635 -66.125 363.965 -65.795 ;
        RECT 363.635 -67.485 363.965 -67.155 ;
        RECT 363.635 -68.845 363.965 -68.515 ;
        RECT 363.635 -70.205 363.965 -69.875 ;
        RECT 363.635 -71.565 363.965 -71.235 ;
        RECT 363.635 -72.925 363.965 -72.595 ;
        RECT 363.635 -74.285 363.965 -73.955 ;
        RECT 363.635 -75.645 363.965 -75.315 ;
        RECT 363.635 -77.005 363.965 -76.675 ;
        RECT 363.635 -78.365 363.965 -78.035 ;
        RECT 363.635 -79.725 363.965 -79.395 ;
        RECT 363.635 -81.085 363.965 -80.755 ;
        RECT 363.635 -82.445 363.965 -82.115 ;
        RECT 363.635 -83.805 363.965 -83.475 ;
        RECT 363.635 -85.165 363.965 -84.835 ;
        RECT 363.635 -86.525 363.965 -86.195 ;
        RECT 363.635 -87.885 363.965 -87.555 ;
        RECT 363.635 -89.245 363.965 -88.915 ;
        RECT 363.635 -90.605 363.965 -90.275 ;
        RECT 363.635 -91.965 363.965 -91.635 ;
        RECT 363.635 -93.325 363.965 -92.995 ;
        RECT 363.635 -94.685 363.965 -94.355 ;
        RECT 363.635 -96.045 363.965 -95.715 ;
        RECT 363.635 -97.405 363.965 -97.075 ;
        RECT 363.635 -98.765 363.965 -98.435 ;
        RECT 363.635 -100.125 363.965 -99.795 ;
        RECT 363.635 -101.485 363.965 -101.155 ;
        RECT 363.635 -102.845 363.965 -102.515 ;
        RECT 363.635 -104.205 363.965 -103.875 ;
        RECT 363.635 -105.565 363.965 -105.235 ;
        RECT 363.635 -106.925 363.965 -106.595 ;
        RECT 363.635 -108.285 363.965 -107.955 ;
        RECT 363.635 -109.645 363.965 -109.315 ;
        RECT 363.635 -111.005 363.965 -110.675 ;
        RECT 363.635 -112.365 363.965 -112.035 ;
        RECT 363.635 -113.725 363.965 -113.395 ;
        RECT 363.635 -115.085 363.965 -114.755 ;
        RECT 363.635 -116.445 363.965 -116.115 ;
        RECT 363.635 -117.805 363.965 -117.475 ;
        RECT 363.635 -119.165 363.965 -118.835 ;
        RECT 363.635 -120.525 363.965 -120.195 ;
        RECT 363.635 -121.885 363.965 -121.555 ;
        RECT 363.635 -123.245 363.965 -122.915 ;
        RECT 363.635 -124.605 363.965 -124.275 ;
        RECT 363.635 -125.965 363.965 -125.635 ;
        RECT 363.635 -127.325 363.965 -126.995 ;
        RECT 363.635 -128.685 363.965 -128.355 ;
        RECT 363.635 -130.045 363.965 -129.715 ;
        RECT 363.635 -131.405 363.965 -131.075 ;
        RECT 363.635 -132.765 363.965 -132.435 ;
        RECT 363.635 -134.125 363.965 -133.795 ;
        RECT 363.635 -135.485 363.965 -135.155 ;
        RECT 363.635 -136.845 363.965 -136.515 ;
        RECT 363.635 -138.205 363.965 -137.875 ;
        RECT 363.635 -139.565 363.965 -139.235 ;
        RECT 363.635 -140.925 363.965 -140.595 ;
        RECT 363.635 -142.285 363.965 -141.955 ;
        RECT 363.635 -143.645 363.965 -143.315 ;
        RECT 363.635 -145.005 363.965 -144.675 ;
        RECT 363.635 -146.365 363.965 -146.035 ;
        RECT 363.635 -147.725 363.965 -147.395 ;
        RECT 363.635 -149.085 363.965 -148.755 ;
        RECT 363.635 -150.445 363.965 -150.115 ;
        RECT 363.635 -151.805 363.965 -151.475 ;
        RECT 363.635 -153.165 363.965 -152.835 ;
        RECT 363.635 -154.525 363.965 -154.195 ;
        RECT 363.635 -155.885 363.965 -155.555 ;
        RECT 363.635 -157.245 363.965 -156.915 ;
        RECT 363.635 -158.605 363.965 -158.275 ;
        RECT 363.635 -159.965 363.965 -159.635 ;
        RECT 363.635 -161.325 363.965 -160.995 ;
        RECT 363.635 -162.685 363.965 -162.355 ;
        RECT 363.635 -164.045 363.965 -163.715 ;
        RECT 363.635 -165.405 363.965 -165.075 ;
        RECT 363.635 -166.765 363.965 -166.435 ;
        RECT 363.635 -168.125 363.965 -167.795 ;
        RECT 363.635 -169.485 363.965 -169.155 ;
        RECT 363.635 -170.845 363.965 -170.515 ;
        RECT 363.635 -172.205 363.965 -171.875 ;
        RECT 363.635 -173.565 363.965 -173.235 ;
        RECT 363.635 -174.925 363.965 -174.595 ;
        RECT 363.635 -176.285 363.965 -175.955 ;
        RECT 363.635 -177.645 363.965 -177.315 ;
        RECT 363.635 -179.005 363.965 -178.675 ;
        RECT 363.635 -180.365 363.965 -180.035 ;
        RECT 363.635 -181.725 363.965 -181.395 ;
        RECT 363.635 -183.085 363.965 -182.755 ;
        RECT 363.635 -184.445 363.965 -184.115 ;
        RECT 363.635 -185.805 363.965 -185.475 ;
        RECT 363.635 -187.165 363.965 -186.835 ;
        RECT 363.635 -188.525 363.965 -188.195 ;
        RECT 363.635 -189.885 363.965 -189.555 ;
        RECT 363.635 -191.245 363.965 -190.915 ;
        RECT 363.635 -192.605 363.965 -192.275 ;
        RECT 363.635 -193.965 363.965 -193.635 ;
        RECT 363.635 -195.325 363.965 -194.995 ;
        RECT 363.635 -196.685 363.965 -196.355 ;
        RECT 363.635 -198.045 363.965 -197.715 ;
        RECT 363.635 -199.405 363.965 -199.075 ;
        RECT 363.635 -200.765 363.965 -200.435 ;
        RECT 363.635 -202.125 363.965 -201.795 ;
        RECT 363.635 -203.485 363.965 -203.155 ;
        RECT 363.635 -204.845 363.965 -204.515 ;
        RECT 363.635 -206.205 363.965 -205.875 ;
        RECT 363.635 -207.565 363.965 -207.235 ;
        RECT 363.635 -208.925 363.965 -208.595 ;
        RECT 363.635 -210.285 363.965 -209.955 ;
        RECT 363.635 -211.645 363.965 -211.315 ;
        RECT 363.635 -213.005 363.965 -212.675 ;
        RECT 363.635 -214.365 363.965 -214.035 ;
        RECT 363.635 -215.725 363.965 -215.395 ;
        RECT 363.635 -217.085 363.965 -216.755 ;
        RECT 363.635 -218.445 363.965 -218.115 ;
        RECT 363.635 -219.805 363.965 -219.475 ;
        RECT 363.635 -221.165 363.965 -220.835 ;
        RECT 363.635 -222.525 363.965 -222.195 ;
        RECT 363.635 -223.885 363.965 -223.555 ;
        RECT 363.635 -225.245 363.965 -224.915 ;
        RECT 363.635 -226.605 363.965 -226.275 ;
        RECT 363.635 -227.965 363.965 -227.635 ;
        RECT 363.635 -229.325 363.965 -228.995 ;
        RECT 363.635 -230.685 363.965 -230.355 ;
        RECT 363.635 -232.045 363.965 -231.715 ;
        RECT 363.635 -233.405 363.965 -233.075 ;
        RECT 363.635 -234.765 363.965 -234.435 ;
        RECT 363.635 -236.125 363.965 -235.795 ;
        RECT 363.635 -237.485 363.965 -237.155 ;
        RECT 363.635 -238.845 363.965 -238.515 ;
        RECT 363.635 -241.09 363.965 -239.96 ;
        RECT 363.64 -241.205 363.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.835 244.04 357.165 245.17 ;
        RECT 356.835 242.595 357.165 242.925 ;
        RECT 356.835 241.235 357.165 241.565 ;
        RECT 356.835 239.875 357.165 240.205 ;
        RECT 356.835 238.515 357.165 238.845 ;
        RECT 356.835 237.155 357.165 237.485 ;
        RECT 356.835 235.975 357.165 236.305 ;
        RECT 356.835 233.925 357.165 234.255 ;
        RECT 356.835 231.995 357.165 232.325 ;
        RECT 356.835 230.155 357.165 230.485 ;
        RECT 356.835 228.665 357.165 228.995 ;
        RECT 356.835 226.995 357.165 227.325 ;
        RECT 356.835 225.505 357.165 225.835 ;
        RECT 356.835 223.835 357.165 224.165 ;
        RECT 356.835 222.345 357.165 222.675 ;
        RECT 356.835 220.675 357.165 221.005 ;
        RECT 356.835 219.185 357.165 219.515 ;
        RECT 356.835 217.775 357.165 218.105 ;
        RECT 356.835 215.935 357.165 216.265 ;
        RECT 356.835 214.445 357.165 214.775 ;
        RECT 356.835 212.775 357.165 213.105 ;
        RECT 356.835 211.285 357.165 211.615 ;
        RECT 356.835 209.615 357.165 209.945 ;
        RECT 356.835 208.125 357.165 208.455 ;
        RECT 356.835 206.455 357.165 206.785 ;
        RECT 356.835 204.965 357.165 205.295 ;
        RECT 356.835 203.555 357.165 203.885 ;
        RECT 356.835 201.715 357.165 202.045 ;
        RECT 356.835 200.225 357.165 200.555 ;
        RECT 356.835 198.555 357.165 198.885 ;
        RECT 356.835 197.065 357.165 197.395 ;
        RECT 356.835 195.395 357.165 195.725 ;
        RECT 356.835 193.905 357.165 194.235 ;
        RECT 356.835 192.235 357.165 192.565 ;
        RECT 356.835 190.745 357.165 191.075 ;
        RECT 356.835 189.335 357.165 189.665 ;
        RECT 356.835 187.495 357.165 187.825 ;
        RECT 356.835 186.005 357.165 186.335 ;
        RECT 356.835 184.335 357.165 184.665 ;
        RECT 356.835 182.845 357.165 183.175 ;
        RECT 356.835 181.175 357.165 181.505 ;
        RECT 356.835 179.685 357.165 180.015 ;
        RECT 356.835 178.015 357.165 178.345 ;
        RECT 356.835 176.525 357.165 176.855 ;
        RECT 356.835 175.115 357.165 175.445 ;
        RECT 356.835 173.275 357.165 173.605 ;
        RECT 356.835 171.785 357.165 172.115 ;
        RECT 356.835 170.115 357.165 170.445 ;
        RECT 356.835 168.625 357.165 168.955 ;
        RECT 356.835 166.955 357.165 167.285 ;
        RECT 356.835 165.465 357.165 165.795 ;
        RECT 356.835 163.795 357.165 164.125 ;
        RECT 356.835 162.305 357.165 162.635 ;
        RECT 356.835 160.895 357.165 161.225 ;
        RECT 356.835 159.055 357.165 159.385 ;
        RECT 356.835 157.565 357.165 157.895 ;
        RECT 356.835 155.895 357.165 156.225 ;
        RECT 356.835 154.405 357.165 154.735 ;
        RECT 356.835 152.735 357.165 153.065 ;
        RECT 356.835 151.245 357.165 151.575 ;
        RECT 356.835 149.575 357.165 149.905 ;
        RECT 356.835 148.085 357.165 148.415 ;
        RECT 356.835 146.675 357.165 147.005 ;
        RECT 356.835 144.835 357.165 145.165 ;
        RECT 356.835 143.345 357.165 143.675 ;
        RECT 356.835 141.675 357.165 142.005 ;
        RECT 356.835 140.185 357.165 140.515 ;
        RECT 356.835 138.515 357.165 138.845 ;
        RECT 356.835 137.025 357.165 137.355 ;
        RECT 356.835 135.355 357.165 135.685 ;
        RECT 356.835 133.865 357.165 134.195 ;
        RECT 356.835 132.455 357.165 132.785 ;
        RECT 356.835 130.615 357.165 130.945 ;
        RECT 356.835 129.125 357.165 129.455 ;
        RECT 356.835 127.455 357.165 127.785 ;
        RECT 356.835 125.965 357.165 126.295 ;
        RECT 356.835 124.295 357.165 124.625 ;
        RECT 356.835 122.805 357.165 123.135 ;
        RECT 356.835 121.135 357.165 121.465 ;
        RECT 356.835 119.645 357.165 119.975 ;
        RECT 356.835 118.235 357.165 118.565 ;
        RECT 356.835 116.395 357.165 116.725 ;
        RECT 356.835 114.905 357.165 115.235 ;
        RECT 356.835 113.235 357.165 113.565 ;
        RECT 356.835 111.745 357.165 112.075 ;
        RECT 356.835 110.075 357.165 110.405 ;
        RECT 356.835 108.585 357.165 108.915 ;
        RECT 356.835 106.915 357.165 107.245 ;
        RECT 356.835 105.425 357.165 105.755 ;
        RECT 356.835 104.015 357.165 104.345 ;
        RECT 356.835 102.175 357.165 102.505 ;
        RECT 356.835 100.685 357.165 101.015 ;
        RECT 356.835 99.015 357.165 99.345 ;
        RECT 356.835 97.525 357.165 97.855 ;
        RECT 356.835 95.855 357.165 96.185 ;
        RECT 356.835 94.365 357.165 94.695 ;
        RECT 356.835 92.695 357.165 93.025 ;
        RECT 356.835 91.205 357.165 91.535 ;
        RECT 356.835 89.795 357.165 90.125 ;
        RECT 356.835 87.955 357.165 88.285 ;
        RECT 356.835 86.465 357.165 86.795 ;
        RECT 356.835 84.795 357.165 85.125 ;
        RECT 356.835 83.305 357.165 83.635 ;
        RECT 356.835 81.635 357.165 81.965 ;
        RECT 356.835 80.145 357.165 80.475 ;
        RECT 356.835 78.475 357.165 78.805 ;
        RECT 356.835 76.985 357.165 77.315 ;
        RECT 356.835 75.575 357.165 75.905 ;
        RECT 356.835 73.735 357.165 74.065 ;
        RECT 356.835 72.245 357.165 72.575 ;
        RECT 356.835 70.575 357.165 70.905 ;
        RECT 356.835 69.085 357.165 69.415 ;
        RECT 356.835 67.415 357.165 67.745 ;
        RECT 356.835 65.925 357.165 66.255 ;
        RECT 356.835 64.255 357.165 64.585 ;
        RECT 356.835 62.765 357.165 63.095 ;
        RECT 356.835 61.355 357.165 61.685 ;
        RECT 356.835 59.515 357.165 59.845 ;
        RECT 356.835 58.025 357.165 58.355 ;
        RECT 356.835 56.355 357.165 56.685 ;
        RECT 356.835 54.865 357.165 55.195 ;
        RECT 356.835 53.195 357.165 53.525 ;
        RECT 356.835 51.705 357.165 52.035 ;
        RECT 356.835 50.035 357.165 50.365 ;
        RECT 356.835 48.545 357.165 48.875 ;
        RECT 356.835 47.135 357.165 47.465 ;
        RECT 356.835 45.295 357.165 45.625 ;
        RECT 356.835 43.805 357.165 44.135 ;
        RECT 356.835 42.135 357.165 42.465 ;
        RECT 356.835 40.645 357.165 40.975 ;
        RECT 356.835 38.975 357.165 39.305 ;
        RECT 356.835 37.485 357.165 37.815 ;
        RECT 356.835 35.815 357.165 36.145 ;
        RECT 356.835 34.325 357.165 34.655 ;
        RECT 356.835 32.915 357.165 33.245 ;
        RECT 356.835 31.075 357.165 31.405 ;
        RECT 356.835 29.585 357.165 29.915 ;
        RECT 356.835 27.915 357.165 28.245 ;
        RECT 356.835 26.425 357.165 26.755 ;
        RECT 356.835 24.755 357.165 25.085 ;
        RECT 356.835 23.265 357.165 23.595 ;
        RECT 356.835 21.595 357.165 21.925 ;
        RECT 356.835 20.105 357.165 20.435 ;
        RECT 356.835 18.695 357.165 19.025 ;
        RECT 356.835 16.855 357.165 17.185 ;
        RECT 356.835 15.365 357.165 15.695 ;
        RECT 356.835 13.695 357.165 14.025 ;
        RECT 356.835 12.205 357.165 12.535 ;
        RECT 356.835 10.535 357.165 10.865 ;
        RECT 356.835 9.045 357.165 9.375 ;
        RECT 356.835 7.375 357.165 7.705 ;
        RECT 356.835 5.885 357.165 6.215 ;
        RECT 356.835 4.475 357.165 4.805 ;
        RECT 356.835 2.115 357.165 2.445 ;
        RECT 356.835 0.06 357.165 0.39 ;
        RECT 356.835 -0.845 357.165 -0.515 ;
        RECT 356.835 -2.205 357.165 -1.875 ;
        RECT 356.835 -3.565 357.165 -3.235 ;
        RECT 356.835 -4.925 357.165 -4.595 ;
        RECT 356.835 -6.285 357.165 -5.955 ;
        RECT 356.835 -7.645 357.165 -7.315 ;
        RECT 356.835 -9.005 357.165 -8.675 ;
        RECT 356.835 -10.365 357.165 -10.035 ;
        RECT 356.835 -11.725 357.165 -11.395 ;
        RECT 356.835 -13.085 357.165 -12.755 ;
        RECT 356.835 -14.445 357.165 -14.115 ;
        RECT 356.835 -15.805 357.165 -15.475 ;
        RECT 356.835 -17.165 357.165 -16.835 ;
        RECT 356.835 -18.525 357.165 -18.195 ;
        RECT 356.835 -19.885 357.165 -19.555 ;
        RECT 356.835 -21.245 357.165 -20.915 ;
        RECT 356.835 -22.605 357.165 -22.275 ;
        RECT 356.835 -23.965 357.165 -23.635 ;
        RECT 356.835 -25.325 357.165 -24.995 ;
        RECT 356.835 -26.685 357.165 -26.355 ;
        RECT 356.835 -28.045 357.165 -27.715 ;
        RECT 356.835 -29.405 357.165 -29.075 ;
        RECT 356.835 -30.765 357.165 -30.435 ;
        RECT 356.835 -32.125 357.165 -31.795 ;
        RECT 356.835 -33.485 357.165 -33.155 ;
        RECT 356.835 -34.845 357.165 -34.515 ;
        RECT 356.835 -36.205 357.165 -35.875 ;
        RECT 356.835 -37.565 357.165 -37.235 ;
        RECT 356.835 -38.925 357.165 -38.595 ;
        RECT 356.835 -40.285 357.165 -39.955 ;
        RECT 356.835 -41.645 357.165 -41.315 ;
        RECT 356.835 -43.005 357.165 -42.675 ;
        RECT 356.835 -44.365 357.165 -44.035 ;
        RECT 356.835 -45.725 357.165 -45.395 ;
        RECT 356.835 -47.085 357.165 -46.755 ;
        RECT 356.835 -48.445 357.165 -48.115 ;
        RECT 356.835 -49.805 357.165 -49.475 ;
        RECT 356.835 -51.165 357.165 -50.835 ;
        RECT 356.835 -52.525 357.165 -52.195 ;
        RECT 356.835 -53.885 357.165 -53.555 ;
        RECT 356.835 -55.245 357.165 -54.915 ;
        RECT 356.835 -56.605 357.165 -56.275 ;
        RECT 356.835 -57.965 357.165 -57.635 ;
        RECT 356.835 -59.325 357.165 -58.995 ;
        RECT 356.835 -60.685 357.165 -60.355 ;
        RECT 356.835 -62.045 357.165 -61.715 ;
        RECT 356.835 -63.405 357.165 -63.075 ;
        RECT 356.835 -64.765 357.165 -64.435 ;
        RECT 356.835 -66.125 357.165 -65.795 ;
        RECT 356.835 -67.485 357.165 -67.155 ;
        RECT 356.835 -68.845 357.165 -68.515 ;
        RECT 356.835 -70.205 357.165 -69.875 ;
        RECT 356.835 -71.565 357.165 -71.235 ;
        RECT 356.835 -72.925 357.165 -72.595 ;
        RECT 356.835 -74.285 357.165 -73.955 ;
        RECT 356.835 -75.645 357.165 -75.315 ;
        RECT 356.835 -77.005 357.165 -76.675 ;
        RECT 356.835 -78.365 357.165 -78.035 ;
        RECT 356.835 -79.725 357.165 -79.395 ;
        RECT 356.835 -81.085 357.165 -80.755 ;
        RECT 356.835 -82.445 357.165 -82.115 ;
        RECT 356.835 -83.805 357.165 -83.475 ;
        RECT 356.835 -85.165 357.165 -84.835 ;
        RECT 356.835 -86.525 357.165 -86.195 ;
        RECT 356.835 -87.885 357.165 -87.555 ;
        RECT 356.835 -89.245 357.165 -88.915 ;
        RECT 356.835 -90.605 357.165 -90.275 ;
        RECT 356.835 -91.965 357.165 -91.635 ;
        RECT 356.835 -93.325 357.165 -92.995 ;
        RECT 356.835 -94.685 357.165 -94.355 ;
        RECT 356.835 -96.045 357.165 -95.715 ;
        RECT 356.835 -97.405 357.165 -97.075 ;
        RECT 356.835 -98.765 357.165 -98.435 ;
        RECT 356.835 -100.125 357.165 -99.795 ;
        RECT 356.835 -101.485 357.165 -101.155 ;
        RECT 356.835 -102.845 357.165 -102.515 ;
        RECT 356.835 -104.205 357.165 -103.875 ;
        RECT 356.835 -105.565 357.165 -105.235 ;
        RECT 356.835 -106.925 357.165 -106.595 ;
        RECT 356.835 -108.285 357.165 -107.955 ;
        RECT 356.835 -109.645 357.165 -109.315 ;
        RECT 356.835 -111.005 357.165 -110.675 ;
        RECT 356.835 -112.365 357.165 -112.035 ;
        RECT 356.835 -113.725 357.165 -113.395 ;
        RECT 356.835 -115.085 357.165 -114.755 ;
        RECT 356.835 -116.445 357.165 -116.115 ;
        RECT 356.835 -117.805 357.165 -117.475 ;
        RECT 356.835 -119.165 357.165 -118.835 ;
        RECT 356.835 -120.525 357.165 -120.195 ;
        RECT 356.835 -121.885 357.165 -121.555 ;
        RECT 356.835 -123.245 357.165 -122.915 ;
        RECT 356.835 -124.605 357.165 -124.275 ;
        RECT 356.835 -125.965 357.165 -125.635 ;
        RECT 356.835 -127.325 357.165 -126.995 ;
        RECT 356.835 -128.685 357.165 -128.355 ;
        RECT 356.835 -130.045 357.165 -129.715 ;
        RECT 356.835 -131.405 357.165 -131.075 ;
        RECT 356.835 -132.765 357.165 -132.435 ;
        RECT 356.835 -134.125 357.165 -133.795 ;
        RECT 356.835 -135.485 357.165 -135.155 ;
        RECT 356.835 -136.845 357.165 -136.515 ;
        RECT 356.835 -138.205 357.165 -137.875 ;
        RECT 356.835 -139.565 357.165 -139.235 ;
        RECT 356.835 -140.925 357.165 -140.595 ;
        RECT 356.835 -142.285 357.165 -141.955 ;
        RECT 356.835 -143.645 357.165 -143.315 ;
        RECT 356.835 -145.005 357.165 -144.675 ;
        RECT 356.835 -146.365 357.165 -146.035 ;
        RECT 356.835 -147.725 357.165 -147.395 ;
        RECT 356.835 -149.085 357.165 -148.755 ;
        RECT 356.835 -150.445 357.165 -150.115 ;
        RECT 356.835 -151.805 357.165 -151.475 ;
        RECT 356.835 -153.165 357.165 -152.835 ;
        RECT 356.835 -154.525 357.165 -154.195 ;
        RECT 356.835 -155.885 357.165 -155.555 ;
        RECT 356.835 -157.245 357.165 -156.915 ;
        RECT 356.835 -158.605 357.165 -158.275 ;
        RECT 356.835 -159.965 357.165 -159.635 ;
        RECT 356.835 -161.325 357.165 -160.995 ;
        RECT 356.835 -162.685 357.165 -162.355 ;
        RECT 356.835 -164.045 357.165 -163.715 ;
        RECT 356.835 -165.405 357.165 -165.075 ;
        RECT 356.835 -166.765 357.165 -166.435 ;
        RECT 356.835 -168.125 357.165 -167.795 ;
        RECT 356.835 -169.485 357.165 -169.155 ;
        RECT 356.835 -170.845 357.165 -170.515 ;
        RECT 356.835 -172.205 357.165 -171.875 ;
        RECT 356.835 -173.565 357.165 -173.235 ;
        RECT 356.835 -174.925 357.165 -174.595 ;
        RECT 356.835 -176.285 357.165 -175.955 ;
        RECT 356.835 -177.645 357.165 -177.315 ;
        RECT 356.835 -179.005 357.165 -178.675 ;
        RECT 356.835 -180.365 357.165 -180.035 ;
        RECT 356.835 -181.725 357.165 -181.395 ;
        RECT 356.835 -183.085 357.165 -182.755 ;
        RECT 356.835 -184.445 357.165 -184.115 ;
        RECT 356.835 -185.805 357.165 -185.475 ;
        RECT 356.835 -187.165 357.165 -186.835 ;
        RECT 356.835 -188.525 357.165 -188.195 ;
        RECT 356.835 -189.885 357.165 -189.555 ;
        RECT 356.835 -191.245 357.165 -190.915 ;
        RECT 356.835 -192.605 357.165 -192.275 ;
        RECT 356.835 -193.965 357.165 -193.635 ;
        RECT 356.835 -195.325 357.165 -194.995 ;
        RECT 356.835 -196.685 357.165 -196.355 ;
        RECT 356.835 -198.045 357.165 -197.715 ;
        RECT 356.835 -199.405 357.165 -199.075 ;
        RECT 356.835 -200.765 357.165 -200.435 ;
        RECT 356.835 -202.125 357.165 -201.795 ;
        RECT 356.835 -203.485 357.165 -203.155 ;
        RECT 356.835 -204.845 357.165 -204.515 ;
        RECT 356.835 -206.205 357.165 -205.875 ;
        RECT 356.835 -207.565 357.165 -207.235 ;
        RECT 356.835 -208.925 357.165 -208.595 ;
        RECT 356.835 -210.285 357.165 -209.955 ;
        RECT 356.835 -211.645 357.165 -211.315 ;
        RECT 356.835 -213.005 357.165 -212.675 ;
        RECT 356.835 -214.365 357.165 -214.035 ;
        RECT 356.835 -215.725 357.165 -215.395 ;
        RECT 356.835 -217.085 357.165 -216.755 ;
        RECT 356.835 -218.445 357.165 -218.115 ;
        RECT 356.835 -219.805 357.165 -219.475 ;
        RECT 356.835 -221.165 357.165 -220.835 ;
        RECT 356.835 -222.525 357.165 -222.195 ;
        RECT 356.835 -223.885 357.165 -223.555 ;
        RECT 356.835 -225.245 357.165 -224.915 ;
        RECT 356.835 -226.605 357.165 -226.275 ;
        RECT 356.835 -227.965 357.165 -227.635 ;
        RECT 356.835 -229.325 357.165 -228.995 ;
        RECT 356.835 -230.685 357.165 -230.355 ;
        RECT 356.835 -232.045 357.165 -231.715 ;
        RECT 356.835 -233.405 357.165 -233.075 ;
        RECT 356.835 -234.765 357.165 -234.435 ;
        RECT 356.835 -236.125 357.165 -235.795 ;
        RECT 356.835 -237.485 357.165 -237.155 ;
        RECT 356.835 -238.845 357.165 -238.515 ;
        RECT 356.835 -241.09 357.165 -239.96 ;
        RECT 356.84 -241.205 357.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.195 244.04 358.525 245.17 ;
        RECT 358.195 242.595 358.525 242.925 ;
        RECT 358.195 241.235 358.525 241.565 ;
        RECT 358.195 239.875 358.525 240.205 ;
        RECT 358.195 238.515 358.525 238.845 ;
        RECT 358.195 237.155 358.525 237.485 ;
        RECT 358.195 235.975 358.525 236.305 ;
        RECT 358.195 233.925 358.525 234.255 ;
        RECT 358.195 231.995 358.525 232.325 ;
        RECT 358.195 230.155 358.525 230.485 ;
        RECT 358.195 228.665 358.525 228.995 ;
        RECT 358.195 226.995 358.525 227.325 ;
        RECT 358.195 225.505 358.525 225.835 ;
        RECT 358.195 223.835 358.525 224.165 ;
        RECT 358.195 222.345 358.525 222.675 ;
        RECT 358.195 220.675 358.525 221.005 ;
        RECT 358.195 219.185 358.525 219.515 ;
        RECT 358.195 217.775 358.525 218.105 ;
        RECT 358.195 215.935 358.525 216.265 ;
        RECT 358.195 214.445 358.525 214.775 ;
        RECT 358.195 212.775 358.525 213.105 ;
        RECT 358.195 211.285 358.525 211.615 ;
        RECT 358.195 209.615 358.525 209.945 ;
        RECT 358.195 208.125 358.525 208.455 ;
        RECT 358.195 206.455 358.525 206.785 ;
        RECT 358.195 204.965 358.525 205.295 ;
        RECT 358.195 203.555 358.525 203.885 ;
        RECT 358.195 201.715 358.525 202.045 ;
        RECT 358.195 200.225 358.525 200.555 ;
        RECT 358.195 198.555 358.525 198.885 ;
        RECT 358.195 197.065 358.525 197.395 ;
        RECT 358.195 195.395 358.525 195.725 ;
        RECT 358.195 193.905 358.525 194.235 ;
        RECT 358.195 192.235 358.525 192.565 ;
        RECT 358.195 190.745 358.525 191.075 ;
        RECT 358.195 189.335 358.525 189.665 ;
        RECT 358.195 187.495 358.525 187.825 ;
        RECT 358.195 186.005 358.525 186.335 ;
        RECT 358.195 184.335 358.525 184.665 ;
        RECT 358.195 182.845 358.525 183.175 ;
        RECT 358.195 181.175 358.525 181.505 ;
        RECT 358.195 179.685 358.525 180.015 ;
        RECT 358.195 178.015 358.525 178.345 ;
        RECT 358.195 176.525 358.525 176.855 ;
        RECT 358.195 175.115 358.525 175.445 ;
        RECT 358.195 173.275 358.525 173.605 ;
        RECT 358.195 171.785 358.525 172.115 ;
        RECT 358.195 170.115 358.525 170.445 ;
        RECT 358.195 168.625 358.525 168.955 ;
        RECT 358.195 166.955 358.525 167.285 ;
        RECT 358.195 165.465 358.525 165.795 ;
        RECT 358.195 163.795 358.525 164.125 ;
        RECT 358.195 162.305 358.525 162.635 ;
        RECT 358.195 160.895 358.525 161.225 ;
        RECT 358.195 159.055 358.525 159.385 ;
        RECT 358.195 157.565 358.525 157.895 ;
        RECT 358.195 155.895 358.525 156.225 ;
        RECT 358.195 154.405 358.525 154.735 ;
        RECT 358.195 152.735 358.525 153.065 ;
        RECT 358.195 151.245 358.525 151.575 ;
        RECT 358.195 149.575 358.525 149.905 ;
        RECT 358.195 148.085 358.525 148.415 ;
        RECT 358.195 146.675 358.525 147.005 ;
        RECT 358.195 144.835 358.525 145.165 ;
        RECT 358.195 143.345 358.525 143.675 ;
        RECT 358.195 141.675 358.525 142.005 ;
        RECT 358.195 140.185 358.525 140.515 ;
        RECT 358.195 138.515 358.525 138.845 ;
        RECT 358.195 137.025 358.525 137.355 ;
        RECT 358.195 135.355 358.525 135.685 ;
        RECT 358.195 133.865 358.525 134.195 ;
        RECT 358.195 132.455 358.525 132.785 ;
        RECT 358.195 130.615 358.525 130.945 ;
        RECT 358.195 129.125 358.525 129.455 ;
        RECT 358.195 127.455 358.525 127.785 ;
        RECT 358.195 125.965 358.525 126.295 ;
        RECT 358.195 124.295 358.525 124.625 ;
        RECT 358.195 122.805 358.525 123.135 ;
        RECT 358.195 121.135 358.525 121.465 ;
        RECT 358.195 119.645 358.525 119.975 ;
        RECT 358.195 118.235 358.525 118.565 ;
        RECT 358.195 116.395 358.525 116.725 ;
        RECT 358.195 114.905 358.525 115.235 ;
        RECT 358.195 113.235 358.525 113.565 ;
        RECT 358.195 111.745 358.525 112.075 ;
        RECT 358.195 110.075 358.525 110.405 ;
        RECT 358.195 108.585 358.525 108.915 ;
        RECT 358.195 106.915 358.525 107.245 ;
        RECT 358.195 105.425 358.525 105.755 ;
        RECT 358.195 104.015 358.525 104.345 ;
        RECT 358.195 102.175 358.525 102.505 ;
        RECT 358.195 100.685 358.525 101.015 ;
        RECT 358.195 99.015 358.525 99.345 ;
        RECT 358.195 97.525 358.525 97.855 ;
        RECT 358.195 95.855 358.525 96.185 ;
        RECT 358.195 94.365 358.525 94.695 ;
        RECT 358.195 92.695 358.525 93.025 ;
        RECT 358.195 91.205 358.525 91.535 ;
        RECT 358.195 89.795 358.525 90.125 ;
        RECT 358.195 87.955 358.525 88.285 ;
        RECT 358.195 86.465 358.525 86.795 ;
        RECT 358.195 84.795 358.525 85.125 ;
        RECT 358.195 83.305 358.525 83.635 ;
        RECT 358.195 81.635 358.525 81.965 ;
        RECT 358.195 80.145 358.525 80.475 ;
        RECT 358.195 78.475 358.525 78.805 ;
        RECT 358.195 76.985 358.525 77.315 ;
        RECT 358.195 75.575 358.525 75.905 ;
        RECT 358.195 73.735 358.525 74.065 ;
        RECT 358.195 72.245 358.525 72.575 ;
        RECT 358.195 70.575 358.525 70.905 ;
        RECT 358.195 69.085 358.525 69.415 ;
        RECT 358.195 67.415 358.525 67.745 ;
        RECT 358.195 65.925 358.525 66.255 ;
        RECT 358.195 64.255 358.525 64.585 ;
        RECT 358.195 62.765 358.525 63.095 ;
        RECT 358.195 61.355 358.525 61.685 ;
        RECT 358.195 59.515 358.525 59.845 ;
        RECT 358.195 58.025 358.525 58.355 ;
        RECT 358.195 56.355 358.525 56.685 ;
        RECT 358.195 54.865 358.525 55.195 ;
        RECT 358.195 53.195 358.525 53.525 ;
        RECT 358.195 51.705 358.525 52.035 ;
        RECT 358.195 50.035 358.525 50.365 ;
        RECT 358.195 48.545 358.525 48.875 ;
        RECT 358.195 47.135 358.525 47.465 ;
        RECT 358.195 45.295 358.525 45.625 ;
        RECT 358.195 43.805 358.525 44.135 ;
        RECT 358.195 42.135 358.525 42.465 ;
        RECT 358.195 40.645 358.525 40.975 ;
        RECT 358.195 38.975 358.525 39.305 ;
        RECT 358.195 37.485 358.525 37.815 ;
        RECT 358.195 35.815 358.525 36.145 ;
        RECT 358.195 34.325 358.525 34.655 ;
        RECT 358.195 32.915 358.525 33.245 ;
        RECT 358.195 31.075 358.525 31.405 ;
        RECT 358.195 29.585 358.525 29.915 ;
        RECT 358.195 27.915 358.525 28.245 ;
        RECT 358.195 26.425 358.525 26.755 ;
        RECT 358.195 24.755 358.525 25.085 ;
        RECT 358.195 23.265 358.525 23.595 ;
        RECT 358.195 21.595 358.525 21.925 ;
        RECT 358.195 20.105 358.525 20.435 ;
        RECT 358.195 18.695 358.525 19.025 ;
        RECT 358.195 16.855 358.525 17.185 ;
        RECT 358.195 15.365 358.525 15.695 ;
        RECT 358.195 13.695 358.525 14.025 ;
        RECT 358.195 12.205 358.525 12.535 ;
        RECT 358.195 10.535 358.525 10.865 ;
        RECT 358.195 9.045 358.525 9.375 ;
        RECT 358.195 7.375 358.525 7.705 ;
        RECT 358.195 5.885 358.525 6.215 ;
        RECT 358.195 4.475 358.525 4.805 ;
        RECT 358.195 2.115 358.525 2.445 ;
        RECT 358.195 0.06 358.525 0.39 ;
        RECT 358.195 -0.845 358.525 -0.515 ;
        RECT 358.195 -2.205 358.525 -1.875 ;
        RECT 358.195 -3.565 358.525 -3.235 ;
        RECT 358.195 -4.925 358.525 -4.595 ;
        RECT 358.195 -6.285 358.525 -5.955 ;
        RECT 358.195 -7.645 358.525 -7.315 ;
        RECT 358.195 -9.005 358.525 -8.675 ;
        RECT 358.195 -10.365 358.525 -10.035 ;
        RECT 358.195 -11.725 358.525 -11.395 ;
        RECT 358.195 -13.085 358.525 -12.755 ;
        RECT 358.195 -14.445 358.525 -14.115 ;
        RECT 358.195 -15.805 358.525 -15.475 ;
        RECT 358.195 -17.165 358.525 -16.835 ;
        RECT 358.195 -18.525 358.525 -18.195 ;
        RECT 358.195 -19.885 358.525 -19.555 ;
        RECT 358.195 -21.245 358.525 -20.915 ;
        RECT 358.195 -22.605 358.525 -22.275 ;
        RECT 358.195 -23.965 358.525 -23.635 ;
        RECT 358.195 -25.325 358.525 -24.995 ;
        RECT 358.195 -26.685 358.525 -26.355 ;
        RECT 358.195 -28.045 358.525 -27.715 ;
        RECT 358.195 -29.405 358.525 -29.075 ;
        RECT 358.195 -30.765 358.525 -30.435 ;
        RECT 358.195 -32.125 358.525 -31.795 ;
        RECT 358.195 -33.485 358.525 -33.155 ;
        RECT 358.195 -34.845 358.525 -34.515 ;
        RECT 358.195 -36.205 358.525 -35.875 ;
        RECT 358.195 -37.565 358.525 -37.235 ;
        RECT 358.195 -38.925 358.525 -38.595 ;
        RECT 358.195 -40.285 358.525 -39.955 ;
        RECT 358.195 -41.645 358.525 -41.315 ;
        RECT 358.195 -43.005 358.525 -42.675 ;
        RECT 358.195 -44.365 358.525 -44.035 ;
        RECT 358.195 -45.725 358.525 -45.395 ;
        RECT 358.195 -47.085 358.525 -46.755 ;
        RECT 358.195 -48.445 358.525 -48.115 ;
        RECT 358.195 -49.805 358.525 -49.475 ;
        RECT 358.195 -51.165 358.525 -50.835 ;
        RECT 358.195 -52.525 358.525 -52.195 ;
        RECT 358.195 -53.885 358.525 -53.555 ;
        RECT 358.195 -55.245 358.525 -54.915 ;
        RECT 358.195 -56.605 358.525 -56.275 ;
        RECT 358.195 -57.965 358.525 -57.635 ;
        RECT 358.195 -59.325 358.525 -58.995 ;
        RECT 358.195 -60.685 358.525 -60.355 ;
        RECT 358.195 -62.045 358.525 -61.715 ;
        RECT 358.195 -63.405 358.525 -63.075 ;
        RECT 358.195 -64.765 358.525 -64.435 ;
        RECT 358.195 -66.125 358.525 -65.795 ;
        RECT 358.195 -67.485 358.525 -67.155 ;
        RECT 358.195 -68.845 358.525 -68.515 ;
        RECT 358.195 -70.205 358.525 -69.875 ;
        RECT 358.195 -71.565 358.525 -71.235 ;
        RECT 358.195 -72.925 358.525 -72.595 ;
        RECT 358.195 -74.285 358.525 -73.955 ;
        RECT 358.195 -75.645 358.525 -75.315 ;
        RECT 358.195 -77.005 358.525 -76.675 ;
        RECT 358.195 -78.365 358.525 -78.035 ;
        RECT 358.195 -79.725 358.525 -79.395 ;
        RECT 358.195 -81.085 358.525 -80.755 ;
        RECT 358.195 -82.445 358.525 -82.115 ;
        RECT 358.195 -83.805 358.525 -83.475 ;
        RECT 358.195 -85.165 358.525 -84.835 ;
        RECT 358.195 -86.525 358.525 -86.195 ;
        RECT 358.195 -87.885 358.525 -87.555 ;
        RECT 358.195 -89.245 358.525 -88.915 ;
        RECT 358.195 -90.605 358.525 -90.275 ;
        RECT 358.195 -91.965 358.525 -91.635 ;
        RECT 358.195 -93.325 358.525 -92.995 ;
        RECT 358.195 -94.685 358.525 -94.355 ;
        RECT 358.195 -96.045 358.525 -95.715 ;
        RECT 358.195 -97.405 358.525 -97.075 ;
        RECT 358.195 -98.765 358.525 -98.435 ;
        RECT 358.195 -100.125 358.525 -99.795 ;
        RECT 358.195 -101.485 358.525 -101.155 ;
        RECT 358.195 -102.845 358.525 -102.515 ;
        RECT 358.195 -104.205 358.525 -103.875 ;
        RECT 358.195 -105.565 358.525 -105.235 ;
        RECT 358.195 -106.925 358.525 -106.595 ;
        RECT 358.195 -108.285 358.525 -107.955 ;
        RECT 358.195 -109.645 358.525 -109.315 ;
        RECT 358.195 -111.005 358.525 -110.675 ;
        RECT 358.195 -112.365 358.525 -112.035 ;
        RECT 358.195 -113.725 358.525 -113.395 ;
        RECT 358.195 -115.085 358.525 -114.755 ;
        RECT 358.195 -116.445 358.525 -116.115 ;
        RECT 358.195 -117.805 358.525 -117.475 ;
        RECT 358.195 -119.165 358.525 -118.835 ;
        RECT 358.195 -120.525 358.525 -120.195 ;
        RECT 358.195 -121.885 358.525 -121.555 ;
        RECT 358.195 -123.245 358.525 -122.915 ;
        RECT 358.195 -124.605 358.525 -124.275 ;
        RECT 358.195 -125.965 358.525 -125.635 ;
        RECT 358.195 -127.325 358.525 -126.995 ;
        RECT 358.195 -128.685 358.525 -128.355 ;
        RECT 358.195 -130.045 358.525 -129.715 ;
        RECT 358.195 -131.405 358.525 -131.075 ;
        RECT 358.195 -132.765 358.525 -132.435 ;
        RECT 358.195 -134.125 358.525 -133.795 ;
        RECT 358.195 -135.485 358.525 -135.155 ;
        RECT 358.195 -136.845 358.525 -136.515 ;
        RECT 358.195 -138.205 358.525 -137.875 ;
        RECT 358.195 -139.565 358.525 -139.235 ;
        RECT 358.195 -140.925 358.525 -140.595 ;
        RECT 358.195 -142.285 358.525 -141.955 ;
        RECT 358.195 -143.645 358.525 -143.315 ;
        RECT 358.195 -145.005 358.525 -144.675 ;
        RECT 358.195 -146.365 358.525 -146.035 ;
        RECT 358.195 -147.725 358.525 -147.395 ;
        RECT 358.195 -149.085 358.525 -148.755 ;
        RECT 358.195 -150.445 358.525 -150.115 ;
        RECT 358.195 -151.805 358.525 -151.475 ;
        RECT 358.195 -153.165 358.525 -152.835 ;
        RECT 358.195 -154.525 358.525 -154.195 ;
        RECT 358.195 -155.885 358.525 -155.555 ;
        RECT 358.195 -157.245 358.525 -156.915 ;
        RECT 358.195 -158.605 358.525 -158.275 ;
        RECT 358.195 -159.965 358.525 -159.635 ;
        RECT 358.195 -161.325 358.525 -160.995 ;
        RECT 358.195 -162.685 358.525 -162.355 ;
        RECT 358.195 -164.045 358.525 -163.715 ;
        RECT 358.195 -165.405 358.525 -165.075 ;
        RECT 358.195 -166.765 358.525 -166.435 ;
        RECT 358.195 -168.125 358.525 -167.795 ;
        RECT 358.195 -169.485 358.525 -169.155 ;
        RECT 358.195 -170.845 358.525 -170.515 ;
        RECT 358.195 -172.205 358.525 -171.875 ;
        RECT 358.195 -173.565 358.525 -173.235 ;
        RECT 358.195 -174.925 358.525 -174.595 ;
        RECT 358.195 -176.285 358.525 -175.955 ;
        RECT 358.195 -177.645 358.525 -177.315 ;
        RECT 358.195 -179.005 358.525 -178.675 ;
        RECT 358.195 -180.365 358.525 -180.035 ;
        RECT 358.195 -181.725 358.525 -181.395 ;
        RECT 358.195 -183.085 358.525 -182.755 ;
        RECT 358.195 -184.445 358.525 -184.115 ;
        RECT 358.195 -185.805 358.525 -185.475 ;
        RECT 358.195 -187.165 358.525 -186.835 ;
        RECT 358.195 -188.525 358.525 -188.195 ;
        RECT 358.195 -189.885 358.525 -189.555 ;
        RECT 358.195 -191.245 358.525 -190.915 ;
        RECT 358.195 -192.605 358.525 -192.275 ;
        RECT 358.195 -193.965 358.525 -193.635 ;
        RECT 358.195 -195.325 358.525 -194.995 ;
        RECT 358.195 -196.685 358.525 -196.355 ;
        RECT 358.195 -198.045 358.525 -197.715 ;
        RECT 358.195 -199.405 358.525 -199.075 ;
        RECT 358.195 -200.765 358.525 -200.435 ;
        RECT 358.195 -202.125 358.525 -201.795 ;
        RECT 358.195 -203.485 358.525 -203.155 ;
        RECT 358.195 -204.845 358.525 -204.515 ;
        RECT 358.195 -206.205 358.525 -205.875 ;
        RECT 358.195 -207.565 358.525 -207.235 ;
        RECT 358.195 -208.925 358.525 -208.595 ;
        RECT 358.195 -210.285 358.525 -209.955 ;
        RECT 358.195 -211.645 358.525 -211.315 ;
        RECT 358.195 -213.005 358.525 -212.675 ;
        RECT 358.195 -214.365 358.525 -214.035 ;
        RECT 358.195 -215.725 358.525 -215.395 ;
        RECT 358.195 -217.085 358.525 -216.755 ;
        RECT 358.195 -218.445 358.525 -218.115 ;
        RECT 358.195 -219.805 358.525 -219.475 ;
        RECT 358.195 -221.165 358.525 -220.835 ;
        RECT 358.195 -222.525 358.525 -222.195 ;
        RECT 358.195 -223.885 358.525 -223.555 ;
        RECT 358.195 -225.245 358.525 -224.915 ;
        RECT 358.195 -226.605 358.525 -226.275 ;
        RECT 358.195 -227.965 358.525 -227.635 ;
        RECT 358.195 -229.325 358.525 -228.995 ;
        RECT 358.195 -230.685 358.525 -230.355 ;
        RECT 358.195 -232.045 358.525 -231.715 ;
        RECT 358.195 -233.405 358.525 -233.075 ;
        RECT 358.195 -234.765 358.525 -234.435 ;
        RECT 358.195 -236.125 358.525 -235.795 ;
        RECT 358.195 -237.485 358.525 -237.155 ;
        RECT 358.195 -238.845 358.525 -238.515 ;
        RECT 358.195 -241.09 358.525 -239.96 ;
        RECT 358.2 -241.205 358.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.555 86.465 359.885 86.795 ;
        RECT 359.555 84.795 359.885 85.125 ;
        RECT 359.555 83.305 359.885 83.635 ;
        RECT 359.555 81.635 359.885 81.965 ;
        RECT 359.555 80.145 359.885 80.475 ;
        RECT 359.555 78.475 359.885 78.805 ;
        RECT 359.555 76.985 359.885 77.315 ;
        RECT 359.555 75.575 359.885 75.905 ;
        RECT 359.555 73.735 359.885 74.065 ;
        RECT 359.555 72.245 359.885 72.575 ;
        RECT 359.555 70.575 359.885 70.905 ;
        RECT 359.555 69.085 359.885 69.415 ;
        RECT 359.555 67.415 359.885 67.745 ;
        RECT 359.555 65.925 359.885 66.255 ;
        RECT 359.555 64.255 359.885 64.585 ;
        RECT 359.555 62.765 359.885 63.095 ;
        RECT 359.555 61.355 359.885 61.685 ;
        RECT 359.555 59.515 359.885 59.845 ;
        RECT 359.555 58.025 359.885 58.355 ;
        RECT 359.555 56.355 359.885 56.685 ;
        RECT 359.555 54.865 359.885 55.195 ;
        RECT 359.555 53.195 359.885 53.525 ;
        RECT 359.555 51.705 359.885 52.035 ;
        RECT 359.555 50.035 359.885 50.365 ;
        RECT 359.555 48.545 359.885 48.875 ;
        RECT 359.555 47.135 359.885 47.465 ;
        RECT 359.555 45.295 359.885 45.625 ;
        RECT 359.555 43.805 359.885 44.135 ;
        RECT 359.555 42.135 359.885 42.465 ;
        RECT 359.555 40.645 359.885 40.975 ;
        RECT 359.555 38.975 359.885 39.305 ;
        RECT 359.555 37.485 359.885 37.815 ;
        RECT 359.555 35.815 359.885 36.145 ;
        RECT 359.555 34.325 359.885 34.655 ;
        RECT 359.555 32.915 359.885 33.245 ;
        RECT 359.555 31.075 359.885 31.405 ;
        RECT 359.555 29.585 359.885 29.915 ;
        RECT 359.555 27.915 359.885 28.245 ;
        RECT 359.555 26.425 359.885 26.755 ;
        RECT 359.555 24.755 359.885 25.085 ;
        RECT 359.555 23.265 359.885 23.595 ;
        RECT 359.555 21.595 359.885 21.925 ;
        RECT 359.555 20.105 359.885 20.435 ;
        RECT 359.555 18.695 359.885 19.025 ;
        RECT 359.555 16.855 359.885 17.185 ;
        RECT 359.555 15.365 359.885 15.695 ;
        RECT 359.555 13.695 359.885 14.025 ;
        RECT 359.555 12.205 359.885 12.535 ;
        RECT 359.555 10.535 359.885 10.865 ;
        RECT 359.555 9.045 359.885 9.375 ;
        RECT 359.555 7.375 359.885 7.705 ;
        RECT 359.555 5.885 359.885 6.215 ;
        RECT 359.555 4.475 359.885 4.805 ;
        RECT 359.555 2.115 359.885 2.445 ;
        RECT 359.555 0.06 359.885 0.39 ;
        RECT 359.555 -0.845 359.885 -0.515 ;
        RECT 359.555 -2.205 359.885 -1.875 ;
        RECT 359.555 -3.565 359.885 -3.235 ;
        RECT 359.555 -4.925 359.885 -4.595 ;
        RECT 359.555 -6.285 359.885 -5.955 ;
        RECT 359.555 -7.645 359.885 -7.315 ;
        RECT 359.555 -9.005 359.885 -8.675 ;
        RECT 359.555 -10.365 359.885 -10.035 ;
        RECT 359.555 -11.725 359.885 -11.395 ;
        RECT 359.555 -13.085 359.885 -12.755 ;
        RECT 359.555 -14.445 359.885 -14.115 ;
        RECT 359.555 -15.805 359.885 -15.475 ;
        RECT 359.555 -17.165 359.885 -16.835 ;
        RECT 359.555 -18.525 359.885 -18.195 ;
        RECT 359.555 -19.885 359.885 -19.555 ;
        RECT 359.555 -21.245 359.885 -20.915 ;
        RECT 359.555 -22.605 359.885 -22.275 ;
        RECT 359.555 -23.965 359.885 -23.635 ;
        RECT 359.555 -25.325 359.885 -24.995 ;
        RECT 359.555 -26.685 359.885 -26.355 ;
        RECT 359.555 -28.045 359.885 -27.715 ;
        RECT 359.555 -29.405 359.885 -29.075 ;
        RECT 359.555 -30.765 359.885 -30.435 ;
        RECT 359.555 -32.125 359.885 -31.795 ;
        RECT 359.555 -33.485 359.885 -33.155 ;
        RECT 359.555 -34.845 359.885 -34.515 ;
        RECT 359.555 -36.205 359.885 -35.875 ;
        RECT 359.555 -37.565 359.885 -37.235 ;
        RECT 359.555 -38.925 359.885 -38.595 ;
        RECT 359.555 -40.285 359.885 -39.955 ;
        RECT 359.555 -41.645 359.885 -41.315 ;
        RECT 359.555 -43.005 359.885 -42.675 ;
        RECT 359.555 -44.365 359.885 -44.035 ;
        RECT 359.555 -45.725 359.885 -45.395 ;
        RECT 359.555 -47.085 359.885 -46.755 ;
        RECT 359.555 -48.445 359.885 -48.115 ;
        RECT 359.555 -49.805 359.885 -49.475 ;
        RECT 359.555 -51.165 359.885 -50.835 ;
        RECT 359.555 -52.525 359.885 -52.195 ;
        RECT 359.555 -53.885 359.885 -53.555 ;
        RECT 359.555 -55.245 359.885 -54.915 ;
        RECT 359.555 -56.605 359.885 -56.275 ;
        RECT 359.555 -57.965 359.885 -57.635 ;
        RECT 359.555 -59.325 359.885 -58.995 ;
        RECT 359.555 -60.685 359.885 -60.355 ;
        RECT 359.555 -62.045 359.885 -61.715 ;
        RECT 359.555 -63.405 359.885 -63.075 ;
        RECT 359.555 -64.765 359.885 -64.435 ;
        RECT 359.555 -66.125 359.885 -65.795 ;
        RECT 359.555 -67.485 359.885 -67.155 ;
        RECT 359.555 -68.845 359.885 -68.515 ;
        RECT 359.555 -70.205 359.885 -69.875 ;
        RECT 359.555 -71.565 359.885 -71.235 ;
        RECT 359.555 -72.925 359.885 -72.595 ;
        RECT 359.555 -74.285 359.885 -73.955 ;
        RECT 359.555 -75.645 359.885 -75.315 ;
        RECT 359.555 -77.005 359.885 -76.675 ;
        RECT 359.555 -78.365 359.885 -78.035 ;
        RECT 359.555 -79.725 359.885 -79.395 ;
        RECT 359.555 -81.085 359.885 -80.755 ;
        RECT 359.555 -82.445 359.885 -82.115 ;
        RECT 359.555 -83.805 359.885 -83.475 ;
        RECT 359.555 -85.165 359.885 -84.835 ;
        RECT 359.555 -86.525 359.885 -86.195 ;
        RECT 359.555 -87.885 359.885 -87.555 ;
        RECT 359.555 -89.245 359.885 -88.915 ;
        RECT 359.555 -90.605 359.885 -90.275 ;
        RECT 359.555 -91.965 359.885 -91.635 ;
        RECT 359.555 -93.325 359.885 -92.995 ;
        RECT 359.555 -94.685 359.885 -94.355 ;
        RECT 359.555 -96.045 359.885 -95.715 ;
        RECT 359.555 -97.405 359.885 -97.075 ;
        RECT 359.555 -98.765 359.885 -98.435 ;
        RECT 359.555 -100.125 359.885 -99.795 ;
        RECT 359.555 -101.485 359.885 -101.155 ;
        RECT 359.555 -102.845 359.885 -102.515 ;
        RECT 359.555 -104.205 359.885 -103.875 ;
        RECT 359.555 -105.565 359.885 -105.235 ;
        RECT 359.555 -106.925 359.885 -106.595 ;
        RECT 359.555 -108.285 359.885 -107.955 ;
        RECT 359.555 -109.645 359.885 -109.315 ;
        RECT 359.555 -111.005 359.885 -110.675 ;
        RECT 359.555 -112.365 359.885 -112.035 ;
        RECT 359.555 -113.725 359.885 -113.395 ;
        RECT 359.555 -115.085 359.885 -114.755 ;
        RECT 359.555 -116.445 359.885 -116.115 ;
        RECT 359.555 -117.805 359.885 -117.475 ;
        RECT 359.555 -119.165 359.885 -118.835 ;
        RECT 359.555 -120.525 359.885 -120.195 ;
        RECT 359.555 -121.885 359.885 -121.555 ;
        RECT 359.555 -123.245 359.885 -122.915 ;
        RECT 359.555 -124.605 359.885 -124.275 ;
        RECT 359.555 -125.965 359.885 -125.635 ;
        RECT 359.555 -127.325 359.885 -126.995 ;
        RECT 359.555 -128.685 359.885 -128.355 ;
        RECT 359.555 -130.045 359.885 -129.715 ;
        RECT 359.555 -131.405 359.885 -131.075 ;
        RECT 359.555 -132.765 359.885 -132.435 ;
        RECT 359.555 -134.125 359.885 -133.795 ;
        RECT 359.555 -135.485 359.885 -135.155 ;
        RECT 359.555 -136.845 359.885 -136.515 ;
        RECT 359.555 -138.205 359.885 -137.875 ;
        RECT 359.555 -139.565 359.885 -139.235 ;
        RECT 359.555 -140.925 359.885 -140.595 ;
        RECT 359.555 -142.285 359.885 -141.955 ;
        RECT 359.555 -143.645 359.885 -143.315 ;
        RECT 359.555 -145.005 359.885 -144.675 ;
        RECT 359.555 -146.365 359.885 -146.035 ;
        RECT 359.555 -147.725 359.885 -147.395 ;
        RECT 359.555 -149.085 359.885 -148.755 ;
        RECT 359.555 -150.445 359.885 -150.115 ;
        RECT 359.555 -151.805 359.885 -151.475 ;
        RECT 359.555 -153.165 359.885 -152.835 ;
        RECT 359.555 -154.525 359.885 -154.195 ;
        RECT 359.555 -155.885 359.885 -155.555 ;
        RECT 359.555 -157.245 359.885 -156.915 ;
        RECT 359.555 -158.605 359.885 -158.275 ;
        RECT 359.555 -159.965 359.885 -159.635 ;
        RECT 359.555 -161.325 359.885 -160.995 ;
        RECT 359.555 -162.685 359.885 -162.355 ;
        RECT 359.555 -164.045 359.885 -163.715 ;
        RECT 359.555 -165.405 359.885 -165.075 ;
        RECT 359.555 -166.765 359.885 -166.435 ;
        RECT 359.555 -168.125 359.885 -167.795 ;
        RECT 359.555 -169.485 359.885 -169.155 ;
        RECT 359.555 -170.845 359.885 -170.515 ;
        RECT 359.555 -172.205 359.885 -171.875 ;
        RECT 359.555 -173.565 359.885 -173.235 ;
        RECT 359.555 -174.925 359.885 -174.595 ;
        RECT 359.555 -176.285 359.885 -175.955 ;
        RECT 359.555 -177.645 359.885 -177.315 ;
        RECT 359.555 -179.005 359.885 -178.675 ;
        RECT 359.555 -180.365 359.885 -180.035 ;
        RECT 359.555 -181.725 359.885 -181.395 ;
        RECT 359.555 -183.085 359.885 -182.755 ;
        RECT 359.555 -184.445 359.885 -184.115 ;
        RECT 359.555 -185.805 359.885 -185.475 ;
        RECT 359.555 -187.165 359.885 -186.835 ;
        RECT 359.555 -188.525 359.885 -188.195 ;
        RECT 359.555 -189.885 359.885 -189.555 ;
        RECT 359.555 -191.245 359.885 -190.915 ;
        RECT 359.555 -192.605 359.885 -192.275 ;
        RECT 359.555 -193.965 359.885 -193.635 ;
        RECT 359.555 -195.325 359.885 -194.995 ;
        RECT 359.555 -196.685 359.885 -196.355 ;
        RECT 359.555 -198.045 359.885 -197.715 ;
        RECT 359.555 -199.405 359.885 -199.075 ;
        RECT 359.555 -200.765 359.885 -200.435 ;
        RECT 359.555 -202.125 359.885 -201.795 ;
        RECT 359.555 -203.485 359.885 -203.155 ;
        RECT 359.555 -204.845 359.885 -204.515 ;
        RECT 359.555 -206.205 359.885 -205.875 ;
        RECT 359.555 -207.565 359.885 -207.235 ;
        RECT 359.555 -208.925 359.885 -208.595 ;
        RECT 359.555 -210.285 359.885 -209.955 ;
        RECT 359.555 -211.645 359.885 -211.315 ;
        RECT 359.555 -213.005 359.885 -212.675 ;
        RECT 359.555 -214.365 359.885 -214.035 ;
        RECT 359.555 -215.725 359.885 -215.395 ;
        RECT 359.555 -217.085 359.885 -216.755 ;
        RECT 359.555 -218.445 359.885 -218.115 ;
        RECT 359.555 -219.805 359.885 -219.475 ;
        RECT 359.555 -221.165 359.885 -220.835 ;
        RECT 359.555 -222.525 359.885 -222.195 ;
        RECT 359.555 -223.885 359.885 -223.555 ;
        RECT 359.555 -225.245 359.885 -224.915 ;
        RECT 359.555 -226.605 359.885 -226.275 ;
        RECT 359.555 -227.965 359.885 -227.635 ;
        RECT 359.555 -229.325 359.885 -228.995 ;
        RECT 359.555 -230.685 359.885 -230.355 ;
        RECT 359.555 -232.045 359.885 -231.715 ;
        RECT 359.555 -233.405 359.885 -233.075 ;
        RECT 359.555 -234.765 359.885 -234.435 ;
        RECT 359.555 -236.125 359.885 -235.795 ;
        RECT 359.555 -237.485 359.885 -237.155 ;
        RECT 359.555 -238.845 359.885 -238.515 ;
        RECT 359.555 -241.09 359.885 -239.96 ;
        RECT 359.56 -241.205 359.88 245.285 ;
        RECT 359.555 244.04 359.885 245.17 ;
        RECT 359.555 242.595 359.885 242.925 ;
        RECT 359.555 241.235 359.885 241.565 ;
        RECT 359.555 239.875 359.885 240.205 ;
        RECT 359.555 238.515 359.885 238.845 ;
        RECT 359.555 237.155 359.885 237.485 ;
        RECT 359.555 235.975 359.885 236.305 ;
        RECT 359.555 233.925 359.885 234.255 ;
        RECT 359.555 231.995 359.885 232.325 ;
        RECT 359.555 230.155 359.885 230.485 ;
        RECT 359.555 228.665 359.885 228.995 ;
        RECT 359.555 226.995 359.885 227.325 ;
        RECT 359.555 225.505 359.885 225.835 ;
        RECT 359.555 223.835 359.885 224.165 ;
        RECT 359.555 222.345 359.885 222.675 ;
        RECT 359.555 220.675 359.885 221.005 ;
        RECT 359.555 219.185 359.885 219.515 ;
        RECT 359.555 217.775 359.885 218.105 ;
        RECT 359.555 215.935 359.885 216.265 ;
        RECT 359.555 214.445 359.885 214.775 ;
        RECT 359.555 212.775 359.885 213.105 ;
        RECT 359.555 211.285 359.885 211.615 ;
        RECT 359.555 209.615 359.885 209.945 ;
        RECT 359.555 208.125 359.885 208.455 ;
        RECT 359.555 206.455 359.885 206.785 ;
        RECT 359.555 204.965 359.885 205.295 ;
        RECT 359.555 203.555 359.885 203.885 ;
        RECT 359.555 201.715 359.885 202.045 ;
        RECT 359.555 200.225 359.885 200.555 ;
        RECT 359.555 198.555 359.885 198.885 ;
        RECT 359.555 197.065 359.885 197.395 ;
        RECT 359.555 195.395 359.885 195.725 ;
        RECT 359.555 193.905 359.885 194.235 ;
        RECT 359.555 192.235 359.885 192.565 ;
        RECT 359.555 190.745 359.885 191.075 ;
        RECT 359.555 189.335 359.885 189.665 ;
        RECT 359.555 187.495 359.885 187.825 ;
        RECT 359.555 186.005 359.885 186.335 ;
        RECT 359.555 184.335 359.885 184.665 ;
        RECT 359.555 182.845 359.885 183.175 ;
        RECT 359.555 181.175 359.885 181.505 ;
        RECT 359.555 179.685 359.885 180.015 ;
        RECT 359.555 178.015 359.885 178.345 ;
        RECT 359.555 176.525 359.885 176.855 ;
        RECT 359.555 175.115 359.885 175.445 ;
        RECT 359.555 173.275 359.885 173.605 ;
        RECT 359.555 171.785 359.885 172.115 ;
        RECT 359.555 170.115 359.885 170.445 ;
        RECT 359.555 168.625 359.885 168.955 ;
        RECT 359.555 166.955 359.885 167.285 ;
        RECT 359.555 165.465 359.885 165.795 ;
        RECT 359.555 163.795 359.885 164.125 ;
        RECT 359.555 162.305 359.885 162.635 ;
        RECT 359.555 160.895 359.885 161.225 ;
        RECT 359.555 159.055 359.885 159.385 ;
        RECT 359.555 157.565 359.885 157.895 ;
        RECT 359.555 155.895 359.885 156.225 ;
        RECT 359.555 154.405 359.885 154.735 ;
        RECT 359.555 152.735 359.885 153.065 ;
        RECT 359.555 151.245 359.885 151.575 ;
        RECT 359.555 149.575 359.885 149.905 ;
        RECT 359.555 148.085 359.885 148.415 ;
        RECT 359.555 146.675 359.885 147.005 ;
        RECT 359.555 144.835 359.885 145.165 ;
        RECT 359.555 143.345 359.885 143.675 ;
        RECT 359.555 141.675 359.885 142.005 ;
        RECT 359.555 140.185 359.885 140.515 ;
        RECT 359.555 138.515 359.885 138.845 ;
        RECT 359.555 137.025 359.885 137.355 ;
        RECT 359.555 135.355 359.885 135.685 ;
        RECT 359.555 133.865 359.885 134.195 ;
        RECT 359.555 132.455 359.885 132.785 ;
        RECT 359.555 130.615 359.885 130.945 ;
        RECT 359.555 129.125 359.885 129.455 ;
        RECT 359.555 127.455 359.885 127.785 ;
        RECT 359.555 125.965 359.885 126.295 ;
        RECT 359.555 124.295 359.885 124.625 ;
        RECT 359.555 122.805 359.885 123.135 ;
        RECT 359.555 121.135 359.885 121.465 ;
        RECT 359.555 119.645 359.885 119.975 ;
        RECT 359.555 118.235 359.885 118.565 ;
        RECT 359.555 116.395 359.885 116.725 ;
        RECT 359.555 114.905 359.885 115.235 ;
        RECT 359.555 113.235 359.885 113.565 ;
        RECT 359.555 111.745 359.885 112.075 ;
        RECT 359.555 110.075 359.885 110.405 ;
        RECT 359.555 108.585 359.885 108.915 ;
        RECT 359.555 106.915 359.885 107.245 ;
        RECT 359.555 105.425 359.885 105.755 ;
        RECT 359.555 104.015 359.885 104.345 ;
        RECT 359.555 102.175 359.885 102.505 ;
        RECT 359.555 100.685 359.885 101.015 ;
        RECT 359.555 99.015 359.885 99.345 ;
        RECT 359.555 97.525 359.885 97.855 ;
        RECT 359.555 95.855 359.885 96.185 ;
        RECT 359.555 94.365 359.885 94.695 ;
        RECT 359.555 92.695 359.885 93.025 ;
        RECT 359.555 91.205 359.885 91.535 ;
        RECT 359.555 89.795 359.885 90.125 ;
        RECT 359.555 87.955 359.885 88.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 -123.245 344.925 -122.915 ;
        RECT 344.595 -124.605 344.925 -124.275 ;
        RECT 344.595 -125.965 344.925 -125.635 ;
        RECT 344.595 -127.325 344.925 -126.995 ;
        RECT 344.595 -128.685 344.925 -128.355 ;
        RECT 344.595 -130.045 344.925 -129.715 ;
        RECT 344.595 -131.405 344.925 -131.075 ;
        RECT 344.595 -132.765 344.925 -132.435 ;
        RECT 344.595 -134.125 344.925 -133.795 ;
        RECT 344.595 -135.485 344.925 -135.155 ;
        RECT 344.595 -136.845 344.925 -136.515 ;
        RECT 344.595 -138.205 344.925 -137.875 ;
        RECT 344.595 -139.565 344.925 -139.235 ;
        RECT 344.595 -140.925 344.925 -140.595 ;
        RECT 344.595 -142.285 344.925 -141.955 ;
        RECT 344.595 -143.645 344.925 -143.315 ;
        RECT 344.595 -145.005 344.925 -144.675 ;
        RECT 344.595 -146.365 344.925 -146.035 ;
        RECT 344.595 -147.725 344.925 -147.395 ;
        RECT 344.595 -149.085 344.925 -148.755 ;
        RECT 344.595 -150.445 344.925 -150.115 ;
        RECT 344.595 -151.805 344.925 -151.475 ;
        RECT 344.595 -153.165 344.925 -152.835 ;
        RECT 344.595 -154.525 344.925 -154.195 ;
        RECT 344.595 -155.885 344.925 -155.555 ;
        RECT 344.595 -157.245 344.925 -156.915 ;
        RECT 344.595 -158.605 344.925 -158.275 ;
        RECT 344.595 -159.965 344.925 -159.635 ;
        RECT 344.595 -161.325 344.925 -160.995 ;
        RECT 344.595 -162.685 344.925 -162.355 ;
        RECT 344.595 -164.045 344.925 -163.715 ;
        RECT 344.595 -165.405 344.925 -165.075 ;
        RECT 344.595 -166.765 344.925 -166.435 ;
        RECT 344.595 -168.125 344.925 -167.795 ;
        RECT 344.595 -169.485 344.925 -169.155 ;
        RECT 344.595 -170.845 344.925 -170.515 ;
        RECT 344.595 -172.205 344.925 -171.875 ;
        RECT 344.595 -173.565 344.925 -173.235 ;
        RECT 344.595 -174.925 344.925 -174.595 ;
        RECT 344.595 -176.285 344.925 -175.955 ;
        RECT 344.595 -177.645 344.925 -177.315 ;
        RECT 344.595 -179.005 344.925 -178.675 ;
        RECT 344.595 -180.365 344.925 -180.035 ;
        RECT 344.595 -181.725 344.925 -181.395 ;
        RECT 344.595 -183.085 344.925 -182.755 ;
        RECT 344.595 -184.445 344.925 -184.115 ;
        RECT 344.595 -185.805 344.925 -185.475 ;
        RECT 344.595 -187.165 344.925 -186.835 ;
        RECT 344.595 -188.525 344.925 -188.195 ;
        RECT 344.595 -189.885 344.925 -189.555 ;
        RECT 344.595 -191.245 344.925 -190.915 ;
        RECT 344.595 -192.605 344.925 -192.275 ;
        RECT 344.595 -193.965 344.925 -193.635 ;
        RECT 344.595 -195.325 344.925 -194.995 ;
        RECT 344.595 -196.685 344.925 -196.355 ;
        RECT 344.595 -198.045 344.925 -197.715 ;
        RECT 344.595 -199.405 344.925 -199.075 ;
        RECT 344.595 -200.765 344.925 -200.435 ;
        RECT 344.595 -202.125 344.925 -201.795 ;
        RECT 344.595 -203.485 344.925 -203.155 ;
        RECT 344.595 -204.845 344.925 -204.515 ;
        RECT 344.595 -206.205 344.925 -205.875 ;
        RECT 344.595 -207.565 344.925 -207.235 ;
        RECT 344.595 -208.925 344.925 -208.595 ;
        RECT 344.595 -210.285 344.925 -209.955 ;
        RECT 344.595 -211.645 344.925 -211.315 ;
        RECT 344.595 -213.005 344.925 -212.675 ;
        RECT 344.595 -214.365 344.925 -214.035 ;
        RECT 344.595 -215.725 344.925 -215.395 ;
        RECT 344.595 -217.085 344.925 -216.755 ;
        RECT 344.595 -218.445 344.925 -218.115 ;
        RECT 344.595 -219.805 344.925 -219.475 ;
        RECT 344.595 -221.165 344.925 -220.835 ;
        RECT 344.595 -222.525 344.925 -222.195 ;
        RECT 344.595 -223.885 344.925 -223.555 ;
        RECT 344.595 -225.245 344.925 -224.915 ;
        RECT 344.595 -226.605 344.925 -226.275 ;
        RECT 344.595 -227.965 344.925 -227.635 ;
        RECT 344.595 -229.325 344.925 -228.995 ;
        RECT 344.595 -230.685 344.925 -230.355 ;
        RECT 344.595 -232.045 344.925 -231.715 ;
        RECT 344.595 -233.405 344.925 -233.075 ;
        RECT 344.595 -234.765 344.925 -234.435 ;
        RECT 344.595 -236.125 344.925 -235.795 ;
        RECT 344.595 -237.485 344.925 -237.155 ;
        RECT 344.595 -238.845 344.925 -238.515 ;
        RECT 344.595 -241.09 344.925 -239.96 ;
        RECT 344.6 -241.205 344.92 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 244.04 346.285 245.17 ;
        RECT 345.955 242.595 346.285 242.925 ;
        RECT 345.955 241.235 346.285 241.565 ;
        RECT 345.955 239.875 346.285 240.205 ;
        RECT 345.955 238.515 346.285 238.845 ;
        RECT 345.955 237.155 346.285 237.485 ;
        RECT 345.96 237.155 346.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 -0.845 346.285 -0.515 ;
        RECT 345.955 -2.205 346.285 -1.875 ;
        RECT 345.955 -3.565 346.285 -3.235 ;
        RECT 345.96 -3.565 346.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 -123.245 346.285 -122.915 ;
        RECT 345.955 -124.605 346.285 -124.275 ;
        RECT 345.955 -125.965 346.285 -125.635 ;
        RECT 345.955 -127.325 346.285 -126.995 ;
        RECT 345.955 -128.685 346.285 -128.355 ;
        RECT 345.955 -130.045 346.285 -129.715 ;
        RECT 345.955 -131.405 346.285 -131.075 ;
        RECT 345.955 -132.765 346.285 -132.435 ;
        RECT 345.955 -134.125 346.285 -133.795 ;
        RECT 345.955 -135.485 346.285 -135.155 ;
        RECT 345.955 -136.845 346.285 -136.515 ;
        RECT 345.955 -138.205 346.285 -137.875 ;
        RECT 345.955 -139.565 346.285 -139.235 ;
        RECT 345.955 -140.925 346.285 -140.595 ;
        RECT 345.955 -142.285 346.285 -141.955 ;
        RECT 345.955 -143.645 346.285 -143.315 ;
        RECT 345.955 -145.005 346.285 -144.675 ;
        RECT 345.955 -146.365 346.285 -146.035 ;
        RECT 345.955 -147.725 346.285 -147.395 ;
        RECT 345.955 -149.085 346.285 -148.755 ;
        RECT 345.955 -150.445 346.285 -150.115 ;
        RECT 345.955 -151.805 346.285 -151.475 ;
        RECT 345.955 -153.165 346.285 -152.835 ;
        RECT 345.955 -154.525 346.285 -154.195 ;
        RECT 345.955 -155.885 346.285 -155.555 ;
        RECT 345.955 -157.245 346.285 -156.915 ;
        RECT 345.955 -158.605 346.285 -158.275 ;
        RECT 345.955 -159.965 346.285 -159.635 ;
        RECT 345.955 -161.325 346.285 -160.995 ;
        RECT 345.955 -162.685 346.285 -162.355 ;
        RECT 345.955 -164.045 346.285 -163.715 ;
        RECT 345.955 -165.405 346.285 -165.075 ;
        RECT 345.955 -166.765 346.285 -166.435 ;
        RECT 345.955 -168.125 346.285 -167.795 ;
        RECT 345.955 -169.485 346.285 -169.155 ;
        RECT 345.955 -170.845 346.285 -170.515 ;
        RECT 345.955 -172.205 346.285 -171.875 ;
        RECT 345.955 -173.565 346.285 -173.235 ;
        RECT 345.955 -174.925 346.285 -174.595 ;
        RECT 345.955 -176.285 346.285 -175.955 ;
        RECT 345.955 -177.645 346.285 -177.315 ;
        RECT 345.955 -179.005 346.285 -178.675 ;
        RECT 345.955 -180.365 346.285 -180.035 ;
        RECT 345.955 -181.725 346.285 -181.395 ;
        RECT 345.955 -183.085 346.285 -182.755 ;
        RECT 345.955 -184.445 346.285 -184.115 ;
        RECT 345.955 -185.805 346.285 -185.475 ;
        RECT 345.955 -187.165 346.285 -186.835 ;
        RECT 345.955 -188.525 346.285 -188.195 ;
        RECT 345.955 -189.885 346.285 -189.555 ;
        RECT 345.955 -191.245 346.285 -190.915 ;
        RECT 345.955 -192.605 346.285 -192.275 ;
        RECT 345.955 -193.965 346.285 -193.635 ;
        RECT 345.955 -195.325 346.285 -194.995 ;
        RECT 345.955 -196.685 346.285 -196.355 ;
        RECT 345.955 -198.045 346.285 -197.715 ;
        RECT 345.955 -199.405 346.285 -199.075 ;
        RECT 345.955 -200.765 346.285 -200.435 ;
        RECT 345.955 -202.125 346.285 -201.795 ;
        RECT 345.955 -203.485 346.285 -203.155 ;
        RECT 345.955 -204.845 346.285 -204.515 ;
        RECT 345.955 -206.205 346.285 -205.875 ;
        RECT 345.955 -207.565 346.285 -207.235 ;
        RECT 345.955 -208.925 346.285 -208.595 ;
        RECT 345.955 -210.285 346.285 -209.955 ;
        RECT 345.955 -211.645 346.285 -211.315 ;
        RECT 345.955 -213.005 346.285 -212.675 ;
        RECT 345.955 -214.365 346.285 -214.035 ;
        RECT 345.955 -215.725 346.285 -215.395 ;
        RECT 345.955 -217.085 346.285 -216.755 ;
        RECT 345.955 -218.445 346.285 -218.115 ;
        RECT 345.955 -219.805 346.285 -219.475 ;
        RECT 345.955 -221.165 346.285 -220.835 ;
        RECT 345.955 -222.525 346.285 -222.195 ;
        RECT 345.955 -223.885 346.285 -223.555 ;
        RECT 345.955 -225.245 346.285 -224.915 ;
        RECT 345.955 -226.605 346.285 -226.275 ;
        RECT 345.955 -227.965 346.285 -227.635 ;
        RECT 345.955 -229.325 346.285 -228.995 ;
        RECT 345.955 -230.685 346.285 -230.355 ;
        RECT 345.955 -232.045 346.285 -231.715 ;
        RECT 345.955 -233.405 346.285 -233.075 ;
        RECT 345.955 -234.765 346.285 -234.435 ;
        RECT 345.955 -236.125 346.285 -235.795 ;
        RECT 345.955 -237.485 346.285 -237.155 ;
        RECT 345.955 -238.845 346.285 -238.515 ;
        RECT 345.955 -241.09 346.285 -239.96 ;
        RECT 345.96 -241.205 346.28 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 244.04 347.645 245.17 ;
        RECT 347.315 242.595 347.645 242.925 ;
        RECT 347.315 241.235 347.645 241.565 ;
        RECT 347.315 239.875 347.645 240.205 ;
        RECT 347.315 238.515 347.645 238.845 ;
        RECT 347.315 237.155 347.645 237.485 ;
        RECT 347.32 237.155 347.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 -0.845 347.645 -0.515 ;
        RECT 347.315 -2.205 347.645 -1.875 ;
        RECT 347.315 -3.565 347.645 -3.235 ;
        RECT 347.32 -3.565 347.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 -123.245 347.645 -122.915 ;
        RECT 347.315 -124.605 347.645 -124.275 ;
        RECT 347.315 -125.965 347.645 -125.635 ;
        RECT 347.315 -127.325 347.645 -126.995 ;
        RECT 347.315 -128.685 347.645 -128.355 ;
        RECT 347.315 -130.045 347.645 -129.715 ;
        RECT 347.315 -131.405 347.645 -131.075 ;
        RECT 347.315 -132.765 347.645 -132.435 ;
        RECT 347.315 -134.125 347.645 -133.795 ;
        RECT 347.315 -135.485 347.645 -135.155 ;
        RECT 347.315 -136.845 347.645 -136.515 ;
        RECT 347.315 -138.205 347.645 -137.875 ;
        RECT 347.315 -139.565 347.645 -139.235 ;
        RECT 347.315 -140.925 347.645 -140.595 ;
        RECT 347.315 -142.285 347.645 -141.955 ;
        RECT 347.315 -143.645 347.645 -143.315 ;
        RECT 347.315 -145.005 347.645 -144.675 ;
        RECT 347.315 -146.365 347.645 -146.035 ;
        RECT 347.315 -147.725 347.645 -147.395 ;
        RECT 347.315 -149.085 347.645 -148.755 ;
        RECT 347.315 -150.445 347.645 -150.115 ;
        RECT 347.315 -151.805 347.645 -151.475 ;
        RECT 347.315 -153.165 347.645 -152.835 ;
        RECT 347.315 -154.525 347.645 -154.195 ;
        RECT 347.315 -155.885 347.645 -155.555 ;
        RECT 347.315 -157.245 347.645 -156.915 ;
        RECT 347.315 -158.605 347.645 -158.275 ;
        RECT 347.315 -159.965 347.645 -159.635 ;
        RECT 347.315 -161.325 347.645 -160.995 ;
        RECT 347.315 -162.685 347.645 -162.355 ;
        RECT 347.315 -164.045 347.645 -163.715 ;
        RECT 347.315 -165.405 347.645 -165.075 ;
        RECT 347.315 -166.765 347.645 -166.435 ;
        RECT 347.315 -168.125 347.645 -167.795 ;
        RECT 347.315 -169.485 347.645 -169.155 ;
        RECT 347.315 -170.845 347.645 -170.515 ;
        RECT 347.315 -172.205 347.645 -171.875 ;
        RECT 347.315 -173.565 347.645 -173.235 ;
        RECT 347.315 -174.925 347.645 -174.595 ;
        RECT 347.315 -176.285 347.645 -175.955 ;
        RECT 347.315 -177.645 347.645 -177.315 ;
        RECT 347.315 -179.005 347.645 -178.675 ;
        RECT 347.315 -180.365 347.645 -180.035 ;
        RECT 347.315 -181.725 347.645 -181.395 ;
        RECT 347.315 -183.085 347.645 -182.755 ;
        RECT 347.315 -184.445 347.645 -184.115 ;
        RECT 347.315 -185.805 347.645 -185.475 ;
        RECT 347.315 -187.165 347.645 -186.835 ;
        RECT 347.315 -188.525 347.645 -188.195 ;
        RECT 347.315 -189.885 347.645 -189.555 ;
        RECT 347.315 -191.245 347.645 -190.915 ;
        RECT 347.315 -192.605 347.645 -192.275 ;
        RECT 347.315 -193.965 347.645 -193.635 ;
        RECT 347.315 -195.325 347.645 -194.995 ;
        RECT 347.315 -196.685 347.645 -196.355 ;
        RECT 347.315 -198.045 347.645 -197.715 ;
        RECT 347.315 -199.405 347.645 -199.075 ;
        RECT 347.315 -200.765 347.645 -200.435 ;
        RECT 347.315 -202.125 347.645 -201.795 ;
        RECT 347.315 -203.485 347.645 -203.155 ;
        RECT 347.315 -204.845 347.645 -204.515 ;
        RECT 347.315 -206.205 347.645 -205.875 ;
        RECT 347.315 -207.565 347.645 -207.235 ;
        RECT 347.315 -208.925 347.645 -208.595 ;
        RECT 347.315 -210.285 347.645 -209.955 ;
        RECT 347.315 -211.645 347.645 -211.315 ;
        RECT 347.315 -213.005 347.645 -212.675 ;
        RECT 347.315 -214.365 347.645 -214.035 ;
        RECT 347.315 -215.725 347.645 -215.395 ;
        RECT 347.315 -217.085 347.645 -216.755 ;
        RECT 347.315 -218.445 347.645 -218.115 ;
        RECT 347.315 -219.805 347.645 -219.475 ;
        RECT 347.315 -221.165 347.645 -220.835 ;
        RECT 347.315 -222.525 347.645 -222.195 ;
        RECT 347.315 -223.885 347.645 -223.555 ;
        RECT 347.315 -225.245 347.645 -224.915 ;
        RECT 347.315 -226.605 347.645 -226.275 ;
        RECT 347.315 -227.965 347.645 -227.635 ;
        RECT 347.315 -229.325 347.645 -228.995 ;
        RECT 347.315 -230.685 347.645 -230.355 ;
        RECT 347.315 -232.045 347.645 -231.715 ;
        RECT 347.315 -233.405 347.645 -233.075 ;
        RECT 347.315 -234.765 347.645 -234.435 ;
        RECT 347.315 -236.125 347.645 -235.795 ;
        RECT 347.315 -237.485 347.645 -237.155 ;
        RECT 347.315 -238.845 347.645 -238.515 ;
        RECT 347.315 -241.09 347.645 -239.96 ;
        RECT 347.32 -241.205 347.64 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 244.04 349.005 245.17 ;
        RECT 348.675 242.595 349.005 242.925 ;
        RECT 348.675 241.235 349.005 241.565 ;
        RECT 348.675 239.875 349.005 240.205 ;
        RECT 348.675 238.515 349.005 238.845 ;
        RECT 348.675 237.155 349.005 237.485 ;
        RECT 348.68 237.155 349 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 -0.845 349.005 -0.515 ;
        RECT 348.675 -2.205 349.005 -1.875 ;
        RECT 348.675 -3.565 349.005 -3.235 ;
        RECT 348.68 -3.565 349 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 -123.245 349.005 -122.915 ;
        RECT 348.675 -124.605 349.005 -124.275 ;
        RECT 348.675 -125.965 349.005 -125.635 ;
        RECT 348.675 -127.325 349.005 -126.995 ;
        RECT 348.675 -128.685 349.005 -128.355 ;
        RECT 348.675 -130.045 349.005 -129.715 ;
        RECT 348.675 -131.405 349.005 -131.075 ;
        RECT 348.675 -132.765 349.005 -132.435 ;
        RECT 348.675 -134.125 349.005 -133.795 ;
        RECT 348.675 -135.485 349.005 -135.155 ;
        RECT 348.675 -136.845 349.005 -136.515 ;
        RECT 348.675 -138.205 349.005 -137.875 ;
        RECT 348.675 -139.565 349.005 -139.235 ;
        RECT 348.675 -140.925 349.005 -140.595 ;
        RECT 348.675 -142.285 349.005 -141.955 ;
        RECT 348.675 -143.645 349.005 -143.315 ;
        RECT 348.675 -145.005 349.005 -144.675 ;
        RECT 348.675 -146.365 349.005 -146.035 ;
        RECT 348.675 -147.725 349.005 -147.395 ;
        RECT 348.675 -149.085 349.005 -148.755 ;
        RECT 348.675 -150.445 349.005 -150.115 ;
        RECT 348.675 -151.805 349.005 -151.475 ;
        RECT 348.675 -153.165 349.005 -152.835 ;
        RECT 348.675 -154.525 349.005 -154.195 ;
        RECT 348.675 -155.885 349.005 -155.555 ;
        RECT 348.675 -157.245 349.005 -156.915 ;
        RECT 348.675 -158.605 349.005 -158.275 ;
        RECT 348.675 -159.965 349.005 -159.635 ;
        RECT 348.675 -161.325 349.005 -160.995 ;
        RECT 348.675 -162.685 349.005 -162.355 ;
        RECT 348.675 -164.045 349.005 -163.715 ;
        RECT 348.675 -165.405 349.005 -165.075 ;
        RECT 348.675 -166.765 349.005 -166.435 ;
        RECT 348.675 -168.125 349.005 -167.795 ;
        RECT 348.675 -169.485 349.005 -169.155 ;
        RECT 348.675 -170.845 349.005 -170.515 ;
        RECT 348.675 -172.205 349.005 -171.875 ;
        RECT 348.675 -173.565 349.005 -173.235 ;
        RECT 348.675 -174.925 349.005 -174.595 ;
        RECT 348.675 -176.285 349.005 -175.955 ;
        RECT 348.675 -177.645 349.005 -177.315 ;
        RECT 348.675 -179.005 349.005 -178.675 ;
        RECT 348.675 -180.365 349.005 -180.035 ;
        RECT 348.675 -181.725 349.005 -181.395 ;
        RECT 348.675 -183.085 349.005 -182.755 ;
        RECT 348.675 -184.445 349.005 -184.115 ;
        RECT 348.675 -185.805 349.005 -185.475 ;
        RECT 348.675 -187.165 349.005 -186.835 ;
        RECT 348.675 -188.525 349.005 -188.195 ;
        RECT 348.675 -189.885 349.005 -189.555 ;
        RECT 348.675 -191.245 349.005 -190.915 ;
        RECT 348.675 -192.605 349.005 -192.275 ;
        RECT 348.675 -193.965 349.005 -193.635 ;
        RECT 348.675 -195.325 349.005 -194.995 ;
        RECT 348.675 -196.685 349.005 -196.355 ;
        RECT 348.675 -198.045 349.005 -197.715 ;
        RECT 348.675 -199.405 349.005 -199.075 ;
        RECT 348.675 -200.765 349.005 -200.435 ;
        RECT 348.675 -202.125 349.005 -201.795 ;
        RECT 348.675 -203.485 349.005 -203.155 ;
        RECT 348.675 -204.845 349.005 -204.515 ;
        RECT 348.675 -206.205 349.005 -205.875 ;
        RECT 348.675 -207.565 349.005 -207.235 ;
        RECT 348.675 -208.925 349.005 -208.595 ;
        RECT 348.675 -210.285 349.005 -209.955 ;
        RECT 348.675 -211.645 349.005 -211.315 ;
        RECT 348.675 -213.005 349.005 -212.675 ;
        RECT 348.675 -214.365 349.005 -214.035 ;
        RECT 348.675 -215.725 349.005 -215.395 ;
        RECT 348.675 -217.085 349.005 -216.755 ;
        RECT 348.675 -218.445 349.005 -218.115 ;
        RECT 348.675 -219.805 349.005 -219.475 ;
        RECT 348.675 -221.165 349.005 -220.835 ;
        RECT 348.675 -222.525 349.005 -222.195 ;
        RECT 348.675 -223.885 349.005 -223.555 ;
        RECT 348.675 -225.245 349.005 -224.915 ;
        RECT 348.675 -226.605 349.005 -226.275 ;
        RECT 348.675 -227.965 349.005 -227.635 ;
        RECT 348.675 -229.325 349.005 -228.995 ;
        RECT 348.675 -230.685 349.005 -230.355 ;
        RECT 348.675 -232.045 349.005 -231.715 ;
        RECT 348.675 -233.405 349.005 -233.075 ;
        RECT 348.675 -234.765 349.005 -234.435 ;
        RECT 348.675 -236.125 349.005 -235.795 ;
        RECT 348.675 -237.485 349.005 -237.155 ;
        RECT 348.675 -238.845 349.005 -238.515 ;
        RECT 348.675 -241.09 349.005 -239.96 ;
        RECT 348.68 -241.205 349 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 244.04 350.365 245.17 ;
        RECT 350.035 242.595 350.365 242.925 ;
        RECT 350.035 241.235 350.365 241.565 ;
        RECT 350.035 239.875 350.365 240.205 ;
        RECT 350.035 238.515 350.365 238.845 ;
        RECT 350.035 237.155 350.365 237.485 ;
        RECT 350.04 237.155 350.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 -0.845 350.365 -0.515 ;
        RECT 350.035 -2.205 350.365 -1.875 ;
        RECT 350.035 -3.565 350.365 -3.235 ;
        RECT 350.04 -3.565 350.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 -123.245 350.365 -122.915 ;
        RECT 350.035 -124.605 350.365 -124.275 ;
        RECT 350.035 -125.965 350.365 -125.635 ;
        RECT 350.035 -127.325 350.365 -126.995 ;
        RECT 350.035 -128.685 350.365 -128.355 ;
        RECT 350.035 -130.045 350.365 -129.715 ;
        RECT 350.035 -131.405 350.365 -131.075 ;
        RECT 350.035 -132.765 350.365 -132.435 ;
        RECT 350.035 -134.125 350.365 -133.795 ;
        RECT 350.035 -135.485 350.365 -135.155 ;
        RECT 350.035 -136.845 350.365 -136.515 ;
        RECT 350.035 -138.205 350.365 -137.875 ;
        RECT 350.035 -139.565 350.365 -139.235 ;
        RECT 350.035 -140.925 350.365 -140.595 ;
        RECT 350.035 -142.285 350.365 -141.955 ;
        RECT 350.035 -143.645 350.365 -143.315 ;
        RECT 350.035 -145.005 350.365 -144.675 ;
        RECT 350.035 -146.365 350.365 -146.035 ;
        RECT 350.035 -147.725 350.365 -147.395 ;
        RECT 350.035 -149.085 350.365 -148.755 ;
        RECT 350.035 -150.445 350.365 -150.115 ;
        RECT 350.035 -151.805 350.365 -151.475 ;
        RECT 350.035 -153.165 350.365 -152.835 ;
        RECT 350.035 -154.525 350.365 -154.195 ;
        RECT 350.035 -155.885 350.365 -155.555 ;
        RECT 350.035 -157.245 350.365 -156.915 ;
        RECT 350.035 -158.605 350.365 -158.275 ;
        RECT 350.035 -159.965 350.365 -159.635 ;
        RECT 350.035 -161.325 350.365 -160.995 ;
        RECT 350.035 -162.685 350.365 -162.355 ;
        RECT 350.035 -164.045 350.365 -163.715 ;
        RECT 350.035 -165.405 350.365 -165.075 ;
        RECT 350.035 -166.765 350.365 -166.435 ;
        RECT 350.035 -168.125 350.365 -167.795 ;
        RECT 350.035 -169.485 350.365 -169.155 ;
        RECT 350.035 -170.845 350.365 -170.515 ;
        RECT 350.035 -172.205 350.365 -171.875 ;
        RECT 350.035 -173.565 350.365 -173.235 ;
        RECT 350.035 -174.925 350.365 -174.595 ;
        RECT 350.035 -176.285 350.365 -175.955 ;
        RECT 350.035 -177.645 350.365 -177.315 ;
        RECT 350.035 -179.005 350.365 -178.675 ;
        RECT 350.035 -180.365 350.365 -180.035 ;
        RECT 350.035 -181.725 350.365 -181.395 ;
        RECT 350.035 -183.085 350.365 -182.755 ;
        RECT 350.035 -184.445 350.365 -184.115 ;
        RECT 350.035 -185.805 350.365 -185.475 ;
        RECT 350.035 -187.165 350.365 -186.835 ;
        RECT 350.035 -188.525 350.365 -188.195 ;
        RECT 350.035 -189.885 350.365 -189.555 ;
        RECT 350.035 -191.245 350.365 -190.915 ;
        RECT 350.035 -192.605 350.365 -192.275 ;
        RECT 350.035 -193.965 350.365 -193.635 ;
        RECT 350.035 -195.325 350.365 -194.995 ;
        RECT 350.035 -196.685 350.365 -196.355 ;
        RECT 350.035 -198.045 350.365 -197.715 ;
        RECT 350.035 -199.405 350.365 -199.075 ;
        RECT 350.035 -200.765 350.365 -200.435 ;
        RECT 350.035 -202.125 350.365 -201.795 ;
        RECT 350.035 -203.485 350.365 -203.155 ;
        RECT 350.035 -204.845 350.365 -204.515 ;
        RECT 350.035 -206.205 350.365 -205.875 ;
        RECT 350.035 -207.565 350.365 -207.235 ;
        RECT 350.035 -208.925 350.365 -208.595 ;
        RECT 350.035 -210.285 350.365 -209.955 ;
        RECT 350.035 -211.645 350.365 -211.315 ;
        RECT 350.035 -213.005 350.365 -212.675 ;
        RECT 350.035 -214.365 350.365 -214.035 ;
        RECT 350.035 -215.725 350.365 -215.395 ;
        RECT 350.035 -217.085 350.365 -216.755 ;
        RECT 350.035 -218.445 350.365 -218.115 ;
        RECT 350.035 -219.805 350.365 -219.475 ;
        RECT 350.035 -221.165 350.365 -220.835 ;
        RECT 350.035 -222.525 350.365 -222.195 ;
        RECT 350.035 -223.885 350.365 -223.555 ;
        RECT 350.035 -225.245 350.365 -224.915 ;
        RECT 350.035 -226.605 350.365 -226.275 ;
        RECT 350.035 -227.965 350.365 -227.635 ;
        RECT 350.035 -229.325 350.365 -228.995 ;
        RECT 350.035 -230.685 350.365 -230.355 ;
        RECT 350.035 -232.045 350.365 -231.715 ;
        RECT 350.035 -233.405 350.365 -233.075 ;
        RECT 350.035 -234.765 350.365 -234.435 ;
        RECT 350.035 -236.125 350.365 -235.795 ;
        RECT 350.035 -237.485 350.365 -237.155 ;
        RECT 350.035 -238.845 350.365 -238.515 ;
        RECT 350.035 -241.09 350.365 -239.96 ;
        RECT 350.04 -241.205 350.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.395 244.04 351.725 245.17 ;
        RECT 351.395 242.595 351.725 242.925 ;
        RECT 351.395 241.235 351.725 241.565 ;
        RECT 351.395 239.875 351.725 240.205 ;
        RECT 351.395 238.515 351.725 238.845 ;
        RECT 351.395 237.155 351.725 237.485 ;
        RECT 351.4 237.155 351.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.395 -127.325 351.725 -126.995 ;
        RECT 351.395 -128.685 351.725 -128.355 ;
        RECT 351.395 -130.045 351.725 -129.715 ;
        RECT 351.395 -131.405 351.725 -131.075 ;
        RECT 351.395 -132.765 351.725 -132.435 ;
        RECT 351.395 -134.125 351.725 -133.795 ;
        RECT 351.395 -135.485 351.725 -135.155 ;
        RECT 351.395 -136.845 351.725 -136.515 ;
        RECT 351.395 -138.205 351.725 -137.875 ;
        RECT 351.395 -139.565 351.725 -139.235 ;
        RECT 351.395 -140.925 351.725 -140.595 ;
        RECT 351.395 -142.285 351.725 -141.955 ;
        RECT 351.395 -143.645 351.725 -143.315 ;
        RECT 351.395 -145.005 351.725 -144.675 ;
        RECT 351.395 -146.365 351.725 -146.035 ;
        RECT 351.395 -147.725 351.725 -147.395 ;
        RECT 351.395 -149.085 351.725 -148.755 ;
        RECT 351.395 -150.445 351.725 -150.115 ;
        RECT 351.395 -151.805 351.725 -151.475 ;
        RECT 351.395 -153.165 351.725 -152.835 ;
        RECT 351.395 -154.525 351.725 -154.195 ;
        RECT 351.395 -155.885 351.725 -155.555 ;
        RECT 351.395 -157.245 351.725 -156.915 ;
        RECT 351.395 -158.605 351.725 -158.275 ;
        RECT 351.395 -159.965 351.725 -159.635 ;
        RECT 351.395 -161.325 351.725 -160.995 ;
        RECT 351.395 -162.685 351.725 -162.355 ;
        RECT 351.395 -164.045 351.725 -163.715 ;
        RECT 351.395 -165.405 351.725 -165.075 ;
        RECT 351.395 -166.765 351.725 -166.435 ;
        RECT 351.395 -168.125 351.725 -167.795 ;
        RECT 351.395 -169.485 351.725 -169.155 ;
        RECT 351.395 -170.845 351.725 -170.515 ;
        RECT 351.395 -172.205 351.725 -171.875 ;
        RECT 351.395 -173.565 351.725 -173.235 ;
        RECT 351.395 -174.925 351.725 -174.595 ;
        RECT 351.395 -176.285 351.725 -175.955 ;
        RECT 351.395 -177.645 351.725 -177.315 ;
        RECT 351.395 -179.005 351.725 -178.675 ;
        RECT 351.395 -180.365 351.725 -180.035 ;
        RECT 351.395 -181.725 351.725 -181.395 ;
        RECT 351.395 -183.085 351.725 -182.755 ;
        RECT 351.395 -184.445 351.725 -184.115 ;
        RECT 351.395 -185.805 351.725 -185.475 ;
        RECT 351.395 -187.165 351.725 -186.835 ;
        RECT 351.395 -188.525 351.725 -188.195 ;
        RECT 351.395 -189.885 351.725 -189.555 ;
        RECT 351.395 -191.245 351.725 -190.915 ;
        RECT 351.395 -192.605 351.725 -192.275 ;
        RECT 351.395 -193.965 351.725 -193.635 ;
        RECT 351.395 -195.325 351.725 -194.995 ;
        RECT 351.395 -196.685 351.725 -196.355 ;
        RECT 351.395 -198.045 351.725 -197.715 ;
        RECT 351.395 -199.405 351.725 -199.075 ;
        RECT 351.395 -200.765 351.725 -200.435 ;
        RECT 351.395 -202.125 351.725 -201.795 ;
        RECT 351.395 -203.485 351.725 -203.155 ;
        RECT 351.395 -204.845 351.725 -204.515 ;
        RECT 351.395 -206.205 351.725 -205.875 ;
        RECT 351.395 -207.565 351.725 -207.235 ;
        RECT 351.395 -208.925 351.725 -208.595 ;
        RECT 351.395 -210.285 351.725 -209.955 ;
        RECT 351.395 -211.645 351.725 -211.315 ;
        RECT 351.395 -213.005 351.725 -212.675 ;
        RECT 351.395 -214.365 351.725 -214.035 ;
        RECT 351.395 -215.725 351.725 -215.395 ;
        RECT 351.395 -217.085 351.725 -216.755 ;
        RECT 351.395 -218.445 351.725 -218.115 ;
        RECT 351.395 -219.805 351.725 -219.475 ;
        RECT 351.395 -221.165 351.725 -220.835 ;
        RECT 351.395 -222.525 351.725 -222.195 ;
        RECT 351.395 -223.885 351.725 -223.555 ;
        RECT 351.395 -225.245 351.725 -224.915 ;
        RECT 351.395 -226.605 351.725 -226.275 ;
        RECT 351.395 -227.965 351.725 -227.635 ;
        RECT 351.395 -229.325 351.725 -228.995 ;
        RECT 351.395 -230.685 351.725 -230.355 ;
        RECT 351.395 -232.045 351.725 -231.715 ;
        RECT 351.395 -233.405 351.725 -233.075 ;
        RECT 351.395 -234.765 351.725 -234.435 ;
        RECT 351.395 -236.125 351.725 -235.795 ;
        RECT 351.395 -237.485 351.725 -237.155 ;
        RECT 351.395 -238.845 351.725 -238.515 ;
        RECT 351.395 -241.09 351.725 -239.96 ;
        RECT 351.4 -241.205 351.72 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.46 -125.535 351.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 244.04 353.085 245.17 ;
        RECT 352.755 242.595 353.085 242.925 ;
        RECT 352.755 241.235 353.085 241.565 ;
        RECT 352.755 239.875 353.085 240.205 ;
        RECT 352.755 238.515 353.085 238.845 ;
        RECT 352.755 237.155 353.085 237.485 ;
        RECT 352.76 237.155 353.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 -127.325 353.085 -126.995 ;
        RECT 352.755 -128.685 353.085 -128.355 ;
        RECT 352.755 -130.045 353.085 -129.715 ;
        RECT 352.755 -131.405 353.085 -131.075 ;
        RECT 352.755 -132.765 353.085 -132.435 ;
        RECT 352.755 -134.125 353.085 -133.795 ;
        RECT 352.755 -135.485 353.085 -135.155 ;
        RECT 352.755 -136.845 353.085 -136.515 ;
        RECT 352.755 -138.205 353.085 -137.875 ;
        RECT 352.755 -139.565 353.085 -139.235 ;
        RECT 352.755 -140.925 353.085 -140.595 ;
        RECT 352.755 -142.285 353.085 -141.955 ;
        RECT 352.755 -143.645 353.085 -143.315 ;
        RECT 352.755 -145.005 353.085 -144.675 ;
        RECT 352.755 -146.365 353.085 -146.035 ;
        RECT 352.755 -147.725 353.085 -147.395 ;
        RECT 352.755 -149.085 353.085 -148.755 ;
        RECT 352.755 -150.445 353.085 -150.115 ;
        RECT 352.755 -151.805 353.085 -151.475 ;
        RECT 352.755 -153.165 353.085 -152.835 ;
        RECT 352.755 -154.525 353.085 -154.195 ;
        RECT 352.755 -155.885 353.085 -155.555 ;
        RECT 352.755 -157.245 353.085 -156.915 ;
        RECT 352.755 -158.605 353.085 -158.275 ;
        RECT 352.755 -159.965 353.085 -159.635 ;
        RECT 352.755 -161.325 353.085 -160.995 ;
        RECT 352.755 -162.685 353.085 -162.355 ;
        RECT 352.755 -164.045 353.085 -163.715 ;
        RECT 352.755 -165.405 353.085 -165.075 ;
        RECT 352.755 -166.765 353.085 -166.435 ;
        RECT 352.755 -168.125 353.085 -167.795 ;
        RECT 352.755 -169.485 353.085 -169.155 ;
        RECT 352.755 -170.845 353.085 -170.515 ;
        RECT 352.755 -172.205 353.085 -171.875 ;
        RECT 352.755 -173.565 353.085 -173.235 ;
        RECT 352.755 -174.925 353.085 -174.595 ;
        RECT 352.755 -176.285 353.085 -175.955 ;
        RECT 352.755 -177.645 353.085 -177.315 ;
        RECT 352.755 -179.005 353.085 -178.675 ;
        RECT 352.755 -180.365 353.085 -180.035 ;
        RECT 352.755 -181.725 353.085 -181.395 ;
        RECT 352.755 -183.085 353.085 -182.755 ;
        RECT 352.755 -184.445 353.085 -184.115 ;
        RECT 352.755 -185.805 353.085 -185.475 ;
        RECT 352.755 -187.165 353.085 -186.835 ;
        RECT 352.755 -188.525 353.085 -188.195 ;
        RECT 352.755 -189.885 353.085 -189.555 ;
        RECT 352.755 -191.245 353.085 -190.915 ;
        RECT 352.755 -192.605 353.085 -192.275 ;
        RECT 352.755 -193.965 353.085 -193.635 ;
        RECT 352.755 -195.325 353.085 -194.995 ;
        RECT 352.755 -196.685 353.085 -196.355 ;
        RECT 352.755 -198.045 353.085 -197.715 ;
        RECT 352.755 -199.405 353.085 -199.075 ;
        RECT 352.755 -200.765 353.085 -200.435 ;
        RECT 352.755 -202.125 353.085 -201.795 ;
        RECT 352.755 -203.485 353.085 -203.155 ;
        RECT 352.755 -204.845 353.085 -204.515 ;
        RECT 352.755 -206.205 353.085 -205.875 ;
        RECT 352.755 -207.565 353.085 -207.235 ;
        RECT 352.755 -208.925 353.085 -208.595 ;
        RECT 352.755 -210.285 353.085 -209.955 ;
        RECT 352.755 -211.645 353.085 -211.315 ;
        RECT 352.755 -213.005 353.085 -212.675 ;
        RECT 352.755 -214.365 353.085 -214.035 ;
        RECT 352.755 -215.725 353.085 -215.395 ;
        RECT 352.755 -217.085 353.085 -216.755 ;
        RECT 352.755 -218.445 353.085 -218.115 ;
        RECT 352.755 -219.805 353.085 -219.475 ;
        RECT 352.755 -221.165 353.085 -220.835 ;
        RECT 352.755 -222.525 353.085 -222.195 ;
        RECT 352.755 -223.885 353.085 -223.555 ;
        RECT 352.755 -225.245 353.085 -224.915 ;
        RECT 352.755 -226.605 353.085 -226.275 ;
        RECT 352.755 -227.965 353.085 -227.635 ;
        RECT 352.755 -229.325 353.085 -228.995 ;
        RECT 352.755 -230.685 353.085 -230.355 ;
        RECT 352.755 -232.045 353.085 -231.715 ;
        RECT 352.755 -233.405 353.085 -233.075 ;
        RECT 352.755 -234.765 353.085 -234.435 ;
        RECT 352.755 -236.125 353.085 -235.795 ;
        RECT 352.755 -237.485 353.085 -237.155 ;
        RECT 352.755 -238.845 353.085 -238.515 ;
        RECT 352.755 -241.09 353.085 -239.96 ;
        RECT 352.76 -241.205 353.08 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 244.04 354.445 245.17 ;
        RECT 354.115 242.595 354.445 242.925 ;
        RECT 354.115 241.235 354.445 241.565 ;
        RECT 354.115 239.875 354.445 240.205 ;
        RECT 354.115 238.515 354.445 238.845 ;
        RECT 354.115 237.155 354.445 237.485 ;
        RECT 354.12 237.155 354.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 -0.845 354.445 -0.515 ;
        RECT 354.115 -2.205 354.445 -1.875 ;
        RECT 354.115 -3.565 354.445 -3.235 ;
        RECT 354.12 -3.565 354.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 -123.245 354.445 -122.915 ;
        RECT 354.115 -124.605 354.445 -124.275 ;
        RECT 354.115 -125.965 354.445 -125.635 ;
        RECT 354.115 -127.325 354.445 -126.995 ;
        RECT 354.115 -128.685 354.445 -128.355 ;
        RECT 354.115 -130.045 354.445 -129.715 ;
        RECT 354.115 -131.405 354.445 -131.075 ;
        RECT 354.115 -132.765 354.445 -132.435 ;
        RECT 354.115 -134.125 354.445 -133.795 ;
        RECT 354.115 -135.485 354.445 -135.155 ;
        RECT 354.115 -136.845 354.445 -136.515 ;
        RECT 354.115 -138.205 354.445 -137.875 ;
        RECT 354.115 -139.565 354.445 -139.235 ;
        RECT 354.115 -140.925 354.445 -140.595 ;
        RECT 354.115 -142.285 354.445 -141.955 ;
        RECT 354.115 -143.645 354.445 -143.315 ;
        RECT 354.115 -145.005 354.445 -144.675 ;
        RECT 354.115 -146.365 354.445 -146.035 ;
        RECT 354.115 -147.725 354.445 -147.395 ;
        RECT 354.115 -149.085 354.445 -148.755 ;
        RECT 354.115 -150.445 354.445 -150.115 ;
        RECT 354.115 -151.805 354.445 -151.475 ;
        RECT 354.115 -153.165 354.445 -152.835 ;
        RECT 354.115 -154.525 354.445 -154.195 ;
        RECT 354.115 -155.885 354.445 -155.555 ;
        RECT 354.115 -157.245 354.445 -156.915 ;
        RECT 354.115 -158.605 354.445 -158.275 ;
        RECT 354.115 -159.965 354.445 -159.635 ;
        RECT 354.115 -161.325 354.445 -160.995 ;
        RECT 354.115 -162.685 354.445 -162.355 ;
        RECT 354.115 -164.045 354.445 -163.715 ;
        RECT 354.115 -165.405 354.445 -165.075 ;
        RECT 354.115 -166.765 354.445 -166.435 ;
        RECT 354.115 -168.125 354.445 -167.795 ;
        RECT 354.115 -169.485 354.445 -169.155 ;
        RECT 354.115 -170.845 354.445 -170.515 ;
        RECT 354.115 -172.205 354.445 -171.875 ;
        RECT 354.115 -173.565 354.445 -173.235 ;
        RECT 354.115 -174.925 354.445 -174.595 ;
        RECT 354.115 -176.285 354.445 -175.955 ;
        RECT 354.115 -177.645 354.445 -177.315 ;
        RECT 354.115 -179.005 354.445 -178.675 ;
        RECT 354.115 -180.365 354.445 -180.035 ;
        RECT 354.115 -181.725 354.445 -181.395 ;
        RECT 354.115 -183.085 354.445 -182.755 ;
        RECT 354.115 -184.445 354.445 -184.115 ;
        RECT 354.115 -185.805 354.445 -185.475 ;
        RECT 354.115 -187.165 354.445 -186.835 ;
        RECT 354.115 -188.525 354.445 -188.195 ;
        RECT 354.115 -189.885 354.445 -189.555 ;
        RECT 354.115 -191.245 354.445 -190.915 ;
        RECT 354.115 -192.605 354.445 -192.275 ;
        RECT 354.115 -193.965 354.445 -193.635 ;
        RECT 354.115 -195.325 354.445 -194.995 ;
        RECT 354.115 -196.685 354.445 -196.355 ;
        RECT 354.115 -198.045 354.445 -197.715 ;
        RECT 354.115 -199.405 354.445 -199.075 ;
        RECT 354.115 -200.765 354.445 -200.435 ;
        RECT 354.115 -202.125 354.445 -201.795 ;
        RECT 354.115 -203.485 354.445 -203.155 ;
        RECT 354.115 -204.845 354.445 -204.515 ;
        RECT 354.115 -206.205 354.445 -205.875 ;
        RECT 354.115 -207.565 354.445 -207.235 ;
        RECT 354.115 -208.925 354.445 -208.595 ;
        RECT 354.115 -210.285 354.445 -209.955 ;
        RECT 354.115 -211.645 354.445 -211.315 ;
        RECT 354.115 -213.005 354.445 -212.675 ;
        RECT 354.115 -214.365 354.445 -214.035 ;
        RECT 354.115 -215.725 354.445 -215.395 ;
        RECT 354.115 -217.085 354.445 -216.755 ;
        RECT 354.115 -218.445 354.445 -218.115 ;
        RECT 354.115 -219.805 354.445 -219.475 ;
        RECT 354.115 -221.165 354.445 -220.835 ;
        RECT 354.115 -222.525 354.445 -222.195 ;
        RECT 354.115 -223.885 354.445 -223.555 ;
        RECT 354.115 -225.245 354.445 -224.915 ;
        RECT 354.115 -226.605 354.445 -226.275 ;
        RECT 354.115 -227.965 354.445 -227.635 ;
        RECT 354.115 -229.325 354.445 -228.995 ;
        RECT 354.115 -230.685 354.445 -230.355 ;
        RECT 354.115 -232.045 354.445 -231.715 ;
        RECT 354.115 -233.405 354.445 -233.075 ;
        RECT 354.115 -234.765 354.445 -234.435 ;
        RECT 354.115 -236.125 354.445 -235.795 ;
        RECT 354.115 -237.485 354.445 -237.155 ;
        RECT 354.115 -238.845 354.445 -238.515 ;
        RECT 354.115 -241.09 354.445 -239.96 ;
        RECT 354.12 -241.205 354.44 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.475 84.795 355.805 85.125 ;
        RECT 355.475 83.305 355.805 83.635 ;
        RECT 355.475 81.635 355.805 81.965 ;
        RECT 355.475 80.145 355.805 80.475 ;
        RECT 355.475 78.475 355.805 78.805 ;
        RECT 355.475 76.985 355.805 77.315 ;
        RECT 355.475 75.575 355.805 75.905 ;
        RECT 355.475 73.735 355.805 74.065 ;
        RECT 355.475 72.245 355.805 72.575 ;
        RECT 355.475 70.575 355.805 70.905 ;
        RECT 355.475 69.085 355.805 69.415 ;
        RECT 355.475 67.415 355.805 67.745 ;
        RECT 355.475 65.925 355.805 66.255 ;
        RECT 355.475 64.255 355.805 64.585 ;
        RECT 355.475 62.765 355.805 63.095 ;
        RECT 355.475 61.355 355.805 61.685 ;
        RECT 355.475 59.515 355.805 59.845 ;
        RECT 355.475 58.025 355.805 58.355 ;
        RECT 355.475 56.355 355.805 56.685 ;
        RECT 355.475 54.865 355.805 55.195 ;
        RECT 355.475 53.195 355.805 53.525 ;
        RECT 355.475 51.705 355.805 52.035 ;
        RECT 355.475 50.035 355.805 50.365 ;
        RECT 355.475 48.545 355.805 48.875 ;
        RECT 355.475 47.135 355.805 47.465 ;
        RECT 355.475 45.295 355.805 45.625 ;
        RECT 355.475 43.805 355.805 44.135 ;
        RECT 355.475 42.135 355.805 42.465 ;
        RECT 355.475 40.645 355.805 40.975 ;
        RECT 355.475 38.975 355.805 39.305 ;
        RECT 355.475 37.485 355.805 37.815 ;
        RECT 355.475 35.815 355.805 36.145 ;
        RECT 355.475 34.325 355.805 34.655 ;
        RECT 355.475 32.915 355.805 33.245 ;
        RECT 355.475 31.075 355.805 31.405 ;
        RECT 355.475 29.585 355.805 29.915 ;
        RECT 355.475 27.915 355.805 28.245 ;
        RECT 355.475 26.425 355.805 26.755 ;
        RECT 355.475 24.755 355.805 25.085 ;
        RECT 355.475 23.265 355.805 23.595 ;
        RECT 355.475 21.595 355.805 21.925 ;
        RECT 355.475 20.105 355.805 20.435 ;
        RECT 355.475 18.695 355.805 19.025 ;
        RECT 355.475 16.855 355.805 17.185 ;
        RECT 355.475 15.365 355.805 15.695 ;
        RECT 355.475 13.695 355.805 14.025 ;
        RECT 355.475 12.205 355.805 12.535 ;
        RECT 355.475 10.535 355.805 10.865 ;
        RECT 355.475 9.045 355.805 9.375 ;
        RECT 355.475 7.375 355.805 7.705 ;
        RECT 355.475 5.885 355.805 6.215 ;
        RECT 355.475 4.475 355.805 4.805 ;
        RECT 355.475 2.115 355.805 2.445 ;
        RECT 355.475 0.06 355.805 0.39 ;
        RECT 355.475 -0.845 355.805 -0.515 ;
        RECT 355.475 -2.205 355.805 -1.875 ;
        RECT 355.475 -3.565 355.805 -3.235 ;
        RECT 355.475 -4.925 355.805 -4.595 ;
        RECT 355.475 -6.285 355.805 -5.955 ;
        RECT 355.475 -7.645 355.805 -7.315 ;
        RECT 355.475 -9.005 355.805 -8.675 ;
        RECT 355.475 -10.365 355.805 -10.035 ;
        RECT 355.475 -11.725 355.805 -11.395 ;
        RECT 355.475 -13.085 355.805 -12.755 ;
        RECT 355.475 -14.445 355.805 -14.115 ;
        RECT 355.475 -15.805 355.805 -15.475 ;
        RECT 355.475 -17.165 355.805 -16.835 ;
        RECT 355.475 -18.525 355.805 -18.195 ;
        RECT 355.475 -19.885 355.805 -19.555 ;
        RECT 355.475 -21.245 355.805 -20.915 ;
        RECT 355.475 -22.605 355.805 -22.275 ;
        RECT 355.475 -23.965 355.805 -23.635 ;
        RECT 355.475 -25.325 355.805 -24.995 ;
        RECT 355.475 -26.685 355.805 -26.355 ;
        RECT 355.475 -28.045 355.805 -27.715 ;
        RECT 355.475 -29.405 355.805 -29.075 ;
        RECT 355.475 -30.765 355.805 -30.435 ;
        RECT 355.475 -32.125 355.805 -31.795 ;
        RECT 355.475 -33.485 355.805 -33.155 ;
        RECT 355.475 -34.845 355.805 -34.515 ;
        RECT 355.475 -36.205 355.805 -35.875 ;
        RECT 355.475 -37.565 355.805 -37.235 ;
        RECT 355.475 -38.925 355.805 -38.595 ;
        RECT 355.475 -40.285 355.805 -39.955 ;
        RECT 355.475 -41.645 355.805 -41.315 ;
        RECT 355.475 -43.005 355.805 -42.675 ;
        RECT 355.475 -44.365 355.805 -44.035 ;
        RECT 355.475 -45.725 355.805 -45.395 ;
        RECT 355.475 -47.085 355.805 -46.755 ;
        RECT 355.475 -48.445 355.805 -48.115 ;
        RECT 355.475 -49.805 355.805 -49.475 ;
        RECT 355.475 -51.165 355.805 -50.835 ;
        RECT 355.475 -52.525 355.805 -52.195 ;
        RECT 355.475 -53.885 355.805 -53.555 ;
        RECT 355.475 -55.245 355.805 -54.915 ;
        RECT 355.475 -56.605 355.805 -56.275 ;
        RECT 355.475 -57.965 355.805 -57.635 ;
        RECT 355.475 -59.325 355.805 -58.995 ;
        RECT 355.475 -60.685 355.805 -60.355 ;
        RECT 355.475 -62.045 355.805 -61.715 ;
        RECT 355.475 -63.405 355.805 -63.075 ;
        RECT 355.475 -64.765 355.805 -64.435 ;
        RECT 355.475 -66.125 355.805 -65.795 ;
        RECT 355.475 -67.485 355.805 -67.155 ;
        RECT 355.475 -68.845 355.805 -68.515 ;
        RECT 355.475 -70.205 355.805 -69.875 ;
        RECT 355.475 -71.565 355.805 -71.235 ;
        RECT 355.475 -72.925 355.805 -72.595 ;
        RECT 355.475 -74.285 355.805 -73.955 ;
        RECT 355.475 -75.645 355.805 -75.315 ;
        RECT 355.475 -77.005 355.805 -76.675 ;
        RECT 355.475 -78.365 355.805 -78.035 ;
        RECT 355.475 -79.725 355.805 -79.395 ;
        RECT 355.475 -81.085 355.805 -80.755 ;
        RECT 355.475 -82.445 355.805 -82.115 ;
        RECT 355.475 -83.805 355.805 -83.475 ;
        RECT 355.475 -85.165 355.805 -84.835 ;
        RECT 355.475 -86.525 355.805 -86.195 ;
        RECT 355.475 -87.885 355.805 -87.555 ;
        RECT 355.475 -89.245 355.805 -88.915 ;
        RECT 355.475 -90.605 355.805 -90.275 ;
        RECT 355.475 -91.965 355.805 -91.635 ;
        RECT 355.475 -93.325 355.805 -92.995 ;
        RECT 355.475 -94.685 355.805 -94.355 ;
        RECT 355.475 -96.045 355.805 -95.715 ;
        RECT 355.475 -97.405 355.805 -97.075 ;
        RECT 355.475 -98.765 355.805 -98.435 ;
        RECT 355.475 -100.125 355.805 -99.795 ;
        RECT 355.475 -101.485 355.805 -101.155 ;
        RECT 355.475 -102.845 355.805 -102.515 ;
        RECT 355.475 -104.205 355.805 -103.875 ;
        RECT 355.475 -105.565 355.805 -105.235 ;
        RECT 355.475 -106.925 355.805 -106.595 ;
        RECT 355.475 -108.285 355.805 -107.955 ;
        RECT 355.475 -109.645 355.805 -109.315 ;
        RECT 355.475 -111.005 355.805 -110.675 ;
        RECT 355.475 -112.365 355.805 -112.035 ;
        RECT 355.475 -113.725 355.805 -113.395 ;
        RECT 355.475 -115.085 355.805 -114.755 ;
        RECT 355.475 -116.445 355.805 -116.115 ;
        RECT 355.475 -117.805 355.805 -117.475 ;
        RECT 355.475 -119.165 355.805 -118.835 ;
        RECT 355.475 -120.525 355.805 -120.195 ;
        RECT 355.475 -121.885 355.805 -121.555 ;
        RECT 355.475 -123.245 355.805 -122.915 ;
        RECT 355.475 -124.605 355.805 -124.275 ;
        RECT 355.475 -125.965 355.805 -125.635 ;
        RECT 355.475 -127.325 355.805 -126.995 ;
        RECT 355.475 -128.685 355.805 -128.355 ;
        RECT 355.475 -130.045 355.805 -129.715 ;
        RECT 355.475 -131.405 355.805 -131.075 ;
        RECT 355.475 -132.765 355.805 -132.435 ;
        RECT 355.475 -134.125 355.805 -133.795 ;
        RECT 355.475 -135.485 355.805 -135.155 ;
        RECT 355.475 -136.845 355.805 -136.515 ;
        RECT 355.475 -138.205 355.805 -137.875 ;
        RECT 355.475 -139.565 355.805 -139.235 ;
        RECT 355.475 -140.925 355.805 -140.595 ;
        RECT 355.475 -142.285 355.805 -141.955 ;
        RECT 355.475 -143.645 355.805 -143.315 ;
        RECT 355.475 -145.005 355.805 -144.675 ;
        RECT 355.475 -146.365 355.805 -146.035 ;
        RECT 355.475 -147.725 355.805 -147.395 ;
        RECT 355.475 -149.085 355.805 -148.755 ;
        RECT 355.475 -150.445 355.805 -150.115 ;
        RECT 355.475 -151.805 355.805 -151.475 ;
        RECT 355.475 -153.165 355.805 -152.835 ;
        RECT 355.475 -154.525 355.805 -154.195 ;
        RECT 355.475 -155.885 355.805 -155.555 ;
        RECT 355.475 -157.245 355.805 -156.915 ;
        RECT 355.475 -158.605 355.805 -158.275 ;
        RECT 355.475 -159.965 355.805 -159.635 ;
        RECT 355.475 -161.325 355.805 -160.995 ;
        RECT 355.475 -162.685 355.805 -162.355 ;
        RECT 355.475 -164.045 355.805 -163.715 ;
        RECT 355.475 -165.405 355.805 -165.075 ;
        RECT 355.475 -166.765 355.805 -166.435 ;
        RECT 355.475 -168.125 355.805 -167.795 ;
        RECT 355.475 -169.485 355.805 -169.155 ;
        RECT 355.475 -170.845 355.805 -170.515 ;
        RECT 355.475 -172.205 355.805 -171.875 ;
        RECT 355.475 -173.565 355.805 -173.235 ;
        RECT 355.475 -174.925 355.805 -174.595 ;
        RECT 355.475 -176.285 355.805 -175.955 ;
        RECT 355.475 -177.645 355.805 -177.315 ;
        RECT 355.475 -179.005 355.805 -178.675 ;
        RECT 355.475 -180.365 355.805 -180.035 ;
        RECT 355.475 -181.725 355.805 -181.395 ;
        RECT 355.475 -183.085 355.805 -182.755 ;
        RECT 355.475 -184.445 355.805 -184.115 ;
        RECT 355.475 -185.805 355.805 -185.475 ;
        RECT 355.475 -187.165 355.805 -186.835 ;
        RECT 355.475 -188.525 355.805 -188.195 ;
        RECT 355.475 -189.885 355.805 -189.555 ;
        RECT 355.475 -191.245 355.805 -190.915 ;
        RECT 355.475 -192.605 355.805 -192.275 ;
        RECT 355.475 -193.965 355.805 -193.635 ;
        RECT 355.475 -195.325 355.805 -194.995 ;
        RECT 355.475 -196.685 355.805 -196.355 ;
        RECT 355.475 -198.045 355.805 -197.715 ;
        RECT 355.475 -199.405 355.805 -199.075 ;
        RECT 355.475 -200.765 355.805 -200.435 ;
        RECT 355.475 -202.125 355.805 -201.795 ;
        RECT 355.475 -203.485 355.805 -203.155 ;
        RECT 355.475 -204.845 355.805 -204.515 ;
        RECT 355.475 -206.205 355.805 -205.875 ;
        RECT 355.475 -207.565 355.805 -207.235 ;
        RECT 355.475 -208.925 355.805 -208.595 ;
        RECT 355.475 -210.285 355.805 -209.955 ;
        RECT 355.475 -211.645 355.805 -211.315 ;
        RECT 355.475 -213.005 355.805 -212.675 ;
        RECT 355.475 -214.365 355.805 -214.035 ;
        RECT 355.475 -215.725 355.805 -215.395 ;
        RECT 355.475 -217.085 355.805 -216.755 ;
        RECT 355.475 -218.445 355.805 -218.115 ;
        RECT 355.475 -219.805 355.805 -219.475 ;
        RECT 355.475 -221.165 355.805 -220.835 ;
        RECT 355.475 -222.525 355.805 -222.195 ;
        RECT 355.475 -223.885 355.805 -223.555 ;
        RECT 355.475 -225.245 355.805 -224.915 ;
        RECT 355.475 -226.605 355.805 -226.275 ;
        RECT 355.475 -227.965 355.805 -227.635 ;
        RECT 355.475 -229.325 355.805 -228.995 ;
        RECT 355.475 -230.685 355.805 -230.355 ;
        RECT 355.475 -232.045 355.805 -231.715 ;
        RECT 355.475 -233.405 355.805 -233.075 ;
        RECT 355.475 -234.765 355.805 -234.435 ;
        RECT 355.475 -236.125 355.805 -235.795 ;
        RECT 355.475 -237.485 355.805 -237.155 ;
        RECT 355.475 -238.845 355.805 -238.515 ;
        RECT 355.475 -241.09 355.805 -239.96 ;
        RECT 355.48 -241.205 355.8 245.285 ;
        RECT 355.475 244.04 355.805 245.17 ;
        RECT 355.475 242.595 355.805 242.925 ;
        RECT 355.475 241.235 355.805 241.565 ;
        RECT 355.475 239.875 355.805 240.205 ;
        RECT 355.475 238.515 355.805 238.845 ;
        RECT 355.475 237.155 355.805 237.485 ;
        RECT 355.475 235.975 355.805 236.305 ;
        RECT 355.475 233.925 355.805 234.255 ;
        RECT 355.475 231.995 355.805 232.325 ;
        RECT 355.475 230.155 355.805 230.485 ;
        RECT 355.475 228.665 355.805 228.995 ;
        RECT 355.475 226.995 355.805 227.325 ;
        RECT 355.475 225.505 355.805 225.835 ;
        RECT 355.475 223.835 355.805 224.165 ;
        RECT 355.475 222.345 355.805 222.675 ;
        RECT 355.475 220.675 355.805 221.005 ;
        RECT 355.475 219.185 355.805 219.515 ;
        RECT 355.475 217.775 355.805 218.105 ;
        RECT 355.475 215.935 355.805 216.265 ;
        RECT 355.475 214.445 355.805 214.775 ;
        RECT 355.475 212.775 355.805 213.105 ;
        RECT 355.475 211.285 355.805 211.615 ;
        RECT 355.475 209.615 355.805 209.945 ;
        RECT 355.475 208.125 355.805 208.455 ;
        RECT 355.475 206.455 355.805 206.785 ;
        RECT 355.475 204.965 355.805 205.295 ;
        RECT 355.475 203.555 355.805 203.885 ;
        RECT 355.475 201.715 355.805 202.045 ;
        RECT 355.475 200.225 355.805 200.555 ;
        RECT 355.475 198.555 355.805 198.885 ;
        RECT 355.475 197.065 355.805 197.395 ;
        RECT 355.475 195.395 355.805 195.725 ;
        RECT 355.475 193.905 355.805 194.235 ;
        RECT 355.475 192.235 355.805 192.565 ;
        RECT 355.475 190.745 355.805 191.075 ;
        RECT 355.475 189.335 355.805 189.665 ;
        RECT 355.475 187.495 355.805 187.825 ;
        RECT 355.475 186.005 355.805 186.335 ;
        RECT 355.475 184.335 355.805 184.665 ;
        RECT 355.475 182.845 355.805 183.175 ;
        RECT 355.475 181.175 355.805 181.505 ;
        RECT 355.475 179.685 355.805 180.015 ;
        RECT 355.475 178.015 355.805 178.345 ;
        RECT 355.475 176.525 355.805 176.855 ;
        RECT 355.475 175.115 355.805 175.445 ;
        RECT 355.475 173.275 355.805 173.605 ;
        RECT 355.475 171.785 355.805 172.115 ;
        RECT 355.475 170.115 355.805 170.445 ;
        RECT 355.475 168.625 355.805 168.955 ;
        RECT 355.475 166.955 355.805 167.285 ;
        RECT 355.475 165.465 355.805 165.795 ;
        RECT 355.475 163.795 355.805 164.125 ;
        RECT 355.475 162.305 355.805 162.635 ;
        RECT 355.475 160.895 355.805 161.225 ;
        RECT 355.475 159.055 355.805 159.385 ;
        RECT 355.475 157.565 355.805 157.895 ;
        RECT 355.475 155.895 355.805 156.225 ;
        RECT 355.475 154.405 355.805 154.735 ;
        RECT 355.475 152.735 355.805 153.065 ;
        RECT 355.475 151.245 355.805 151.575 ;
        RECT 355.475 149.575 355.805 149.905 ;
        RECT 355.475 148.085 355.805 148.415 ;
        RECT 355.475 146.675 355.805 147.005 ;
        RECT 355.475 144.835 355.805 145.165 ;
        RECT 355.475 143.345 355.805 143.675 ;
        RECT 355.475 141.675 355.805 142.005 ;
        RECT 355.475 140.185 355.805 140.515 ;
        RECT 355.475 138.515 355.805 138.845 ;
        RECT 355.475 137.025 355.805 137.355 ;
        RECT 355.475 135.355 355.805 135.685 ;
        RECT 355.475 133.865 355.805 134.195 ;
        RECT 355.475 132.455 355.805 132.785 ;
        RECT 355.475 130.615 355.805 130.945 ;
        RECT 355.475 129.125 355.805 129.455 ;
        RECT 355.475 127.455 355.805 127.785 ;
        RECT 355.475 125.965 355.805 126.295 ;
        RECT 355.475 124.295 355.805 124.625 ;
        RECT 355.475 122.805 355.805 123.135 ;
        RECT 355.475 121.135 355.805 121.465 ;
        RECT 355.475 119.645 355.805 119.975 ;
        RECT 355.475 118.235 355.805 118.565 ;
        RECT 355.475 116.395 355.805 116.725 ;
        RECT 355.475 114.905 355.805 115.235 ;
        RECT 355.475 113.235 355.805 113.565 ;
        RECT 355.475 111.745 355.805 112.075 ;
        RECT 355.475 110.075 355.805 110.405 ;
        RECT 355.475 108.585 355.805 108.915 ;
        RECT 355.475 106.915 355.805 107.245 ;
        RECT 355.475 105.425 355.805 105.755 ;
        RECT 355.475 104.015 355.805 104.345 ;
        RECT 355.475 102.175 355.805 102.505 ;
        RECT 355.475 100.685 355.805 101.015 ;
        RECT 355.475 99.015 355.805 99.345 ;
        RECT 355.475 97.525 355.805 97.855 ;
        RECT 355.475 95.855 355.805 96.185 ;
        RECT 355.475 94.365 355.805 94.695 ;
        RECT 355.475 92.695 355.805 93.025 ;
        RECT 355.475 91.205 355.805 91.535 ;
        RECT 355.475 89.795 355.805 90.125 ;
        RECT 355.475 87.955 355.805 88.285 ;
        RECT 355.475 86.465 355.805 86.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 244.04 327.245 245.17 ;
        RECT 326.915 242.595 327.245 242.925 ;
        RECT 326.915 241.235 327.245 241.565 ;
        RECT 326.915 239.875 327.245 240.205 ;
        RECT 326.915 238.515 327.245 238.845 ;
        RECT 326.915 237.155 327.245 237.485 ;
        RECT 326.92 237.155 327.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 -0.845 327.245 -0.515 ;
        RECT 326.915 -2.205 327.245 -1.875 ;
        RECT 326.915 -3.565 327.245 -3.235 ;
        RECT 326.92 -3.565 327.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 -123.245 327.245 -122.915 ;
        RECT 326.915 -124.605 327.245 -124.275 ;
        RECT 326.915 -125.965 327.245 -125.635 ;
        RECT 326.915 -127.325 327.245 -126.995 ;
        RECT 326.915 -128.685 327.245 -128.355 ;
        RECT 326.915 -130.045 327.245 -129.715 ;
        RECT 326.915 -131.405 327.245 -131.075 ;
        RECT 326.915 -132.765 327.245 -132.435 ;
        RECT 326.915 -134.125 327.245 -133.795 ;
        RECT 326.915 -135.485 327.245 -135.155 ;
        RECT 326.915 -136.845 327.245 -136.515 ;
        RECT 326.915 -138.205 327.245 -137.875 ;
        RECT 326.915 -139.565 327.245 -139.235 ;
        RECT 326.915 -140.925 327.245 -140.595 ;
        RECT 326.915 -142.285 327.245 -141.955 ;
        RECT 326.915 -143.645 327.245 -143.315 ;
        RECT 326.915 -145.005 327.245 -144.675 ;
        RECT 326.915 -146.365 327.245 -146.035 ;
        RECT 326.915 -147.725 327.245 -147.395 ;
        RECT 326.915 -149.085 327.245 -148.755 ;
        RECT 326.915 -150.445 327.245 -150.115 ;
        RECT 326.915 -151.805 327.245 -151.475 ;
        RECT 326.915 -153.165 327.245 -152.835 ;
        RECT 326.915 -154.525 327.245 -154.195 ;
        RECT 326.915 -155.885 327.245 -155.555 ;
        RECT 326.915 -157.245 327.245 -156.915 ;
        RECT 326.915 -158.605 327.245 -158.275 ;
        RECT 326.915 -159.965 327.245 -159.635 ;
        RECT 326.915 -161.325 327.245 -160.995 ;
        RECT 326.915 -162.685 327.245 -162.355 ;
        RECT 326.915 -164.045 327.245 -163.715 ;
        RECT 326.915 -165.405 327.245 -165.075 ;
        RECT 326.915 -166.765 327.245 -166.435 ;
        RECT 326.915 -168.125 327.245 -167.795 ;
        RECT 326.915 -169.485 327.245 -169.155 ;
        RECT 326.915 -170.845 327.245 -170.515 ;
        RECT 326.915 -172.205 327.245 -171.875 ;
        RECT 326.915 -173.565 327.245 -173.235 ;
        RECT 326.915 -174.925 327.245 -174.595 ;
        RECT 326.915 -176.285 327.245 -175.955 ;
        RECT 326.915 -177.645 327.245 -177.315 ;
        RECT 326.915 -179.005 327.245 -178.675 ;
        RECT 326.915 -180.365 327.245 -180.035 ;
        RECT 326.915 -181.725 327.245 -181.395 ;
        RECT 326.915 -183.085 327.245 -182.755 ;
        RECT 326.915 -184.445 327.245 -184.115 ;
        RECT 326.915 -185.805 327.245 -185.475 ;
        RECT 326.915 -187.165 327.245 -186.835 ;
        RECT 326.915 -188.525 327.245 -188.195 ;
        RECT 326.915 -189.885 327.245 -189.555 ;
        RECT 326.915 -191.245 327.245 -190.915 ;
        RECT 326.915 -192.605 327.245 -192.275 ;
        RECT 326.915 -193.965 327.245 -193.635 ;
        RECT 326.915 -195.325 327.245 -194.995 ;
        RECT 326.915 -196.685 327.245 -196.355 ;
        RECT 326.915 -198.045 327.245 -197.715 ;
        RECT 326.915 -199.405 327.245 -199.075 ;
        RECT 326.915 -200.765 327.245 -200.435 ;
        RECT 326.915 -202.125 327.245 -201.795 ;
        RECT 326.915 -203.485 327.245 -203.155 ;
        RECT 326.915 -204.845 327.245 -204.515 ;
        RECT 326.915 -206.205 327.245 -205.875 ;
        RECT 326.915 -207.565 327.245 -207.235 ;
        RECT 326.915 -208.925 327.245 -208.595 ;
        RECT 326.915 -210.285 327.245 -209.955 ;
        RECT 326.915 -211.645 327.245 -211.315 ;
        RECT 326.915 -213.005 327.245 -212.675 ;
        RECT 326.915 -214.365 327.245 -214.035 ;
        RECT 326.915 -215.725 327.245 -215.395 ;
        RECT 326.915 -217.085 327.245 -216.755 ;
        RECT 326.915 -218.445 327.245 -218.115 ;
        RECT 326.915 -219.805 327.245 -219.475 ;
        RECT 326.915 -221.165 327.245 -220.835 ;
        RECT 326.915 -222.525 327.245 -222.195 ;
        RECT 326.915 -223.885 327.245 -223.555 ;
        RECT 326.915 -225.245 327.245 -224.915 ;
        RECT 326.915 -226.605 327.245 -226.275 ;
        RECT 326.915 -227.965 327.245 -227.635 ;
        RECT 326.915 -229.325 327.245 -228.995 ;
        RECT 326.915 -230.685 327.245 -230.355 ;
        RECT 326.915 -232.045 327.245 -231.715 ;
        RECT 326.915 -233.405 327.245 -233.075 ;
        RECT 326.915 -234.765 327.245 -234.435 ;
        RECT 326.915 -236.125 327.245 -235.795 ;
        RECT 326.915 -237.485 327.245 -237.155 ;
        RECT 326.915 -238.845 327.245 -238.515 ;
        RECT 326.915 -241.09 327.245 -239.96 ;
        RECT 326.92 -241.205 327.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 244.04 328.605 245.17 ;
        RECT 328.275 242.595 328.605 242.925 ;
        RECT 328.275 241.235 328.605 241.565 ;
        RECT 328.275 239.875 328.605 240.205 ;
        RECT 328.275 238.515 328.605 238.845 ;
        RECT 328.275 237.155 328.605 237.485 ;
        RECT 328.28 237.155 328.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 -0.845 328.605 -0.515 ;
        RECT 328.275 -2.205 328.605 -1.875 ;
        RECT 328.275 -3.565 328.605 -3.235 ;
        RECT 328.28 -3.565 328.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 -123.245 328.605 -122.915 ;
        RECT 328.275 -124.605 328.605 -124.275 ;
        RECT 328.275 -125.965 328.605 -125.635 ;
        RECT 328.275 -127.325 328.605 -126.995 ;
        RECT 328.275 -128.685 328.605 -128.355 ;
        RECT 328.275 -130.045 328.605 -129.715 ;
        RECT 328.275 -131.405 328.605 -131.075 ;
        RECT 328.275 -132.765 328.605 -132.435 ;
        RECT 328.275 -134.125 328.605 -133.795 ;
        RECT 328.275 -135.485 328.605 -135.155 ;
        RECT 328.275 -136.845 328.605 -136.515 ;
        RECT 328.275 -138.205 328.605 -137.875 ;
        RECT 328.275 -139.565 328.605 -139.235 ;
        RECT 328.275 -140.925 328.605 -140.595 ;
        RECT 328.275 -142.285 328.605 -141.955 ;
        RECT 328.275 -143.645 328.605 -143.315 ;
        RECT 328.275 -145.005 328.605 -144.675 ;
        RECT 328.275 -146.365 328.605 -146.035 ;
        RECT 328.275 -147.725 328.605 -147.395 ;
        RECT 328.275 -149.085 328.605 -148.755 ;
        RECT 328.275 -150.445 328.605 -150.115 ;
        RECT 328.275 -151.805 328.605 -151.475 ;
        RECT 328.275 -153.165 328.605 -152.835 ;
        RECT 328.275 -154.525 328.605 -154.195 ;
        RECT 328.275 -155.885 328.605 -155.555 ;
        RECT 328.275 -157.245 328.605 -156.915 ;
        RECT 328.275 -158.605 328.605 -158.275 ;
        RECT 328.275 -159.965 328.605 -159.635 ;
        RECT 328.275 -161.325 328.605 -160.995 ;
        RECT 328.275 -162.685 328.605 -162.355 ;
        RECT 328.275 -164.045 328.605 -163.715 ;
        RECT 328.275 -165.405 328.605 -165.075 ;
        RECT 328.275 -166.765 328.605 -166.435 ;
        RECT 328.275 -168.125 328.605 -167.795 ;
        RECT 328.275 -169.485 328.605 -169.155 ;
        RECT 328.275 -170.845 328.605 -170.515 ;
        RECT 328.275 -172.205 328.605 -171.875 ;
        RECT 328.275 -173.565 328.605 -173.235 ;
        RECT 328.275 -174.925 328.605 -174.595 ;
        RECT 328.275 -176.285 328.605 -175.955 ;
        RECT 328.275 -177.645 328.605 -177.315 ;
        RECT 328.275 -179.005 328.605 -178.675 ;
        RECT 328.275 -180.365 328.605 -180.035 ;
        RECT 328.275 -181.725 328.605 -181.395 ;
        RECT 328.275 -183.085 328.605 -182.755 ;
        RECT 328.275 -184.445 328.605 -184.115 ;
        RECT 328.275 -185.805 328.605 -185.475 ;
        RECT 328.275 -187.165 328.605 -186.835 ;
        RECT 328.275 -188.525 328.605 -188.195 ;
        RECT 328.275 -189.885 328.605 -189.555 ;
        RECT 328.275 -191.245 328.605 -190.915 ;
        RECT 328.275 -192.605 328.605 -192.275 ;
        RECT 328.275 -193.965 328.605 -193.635 ;
        RECT 328.275 -195.325 328.605 -194.995 ;
        RECT 328.275 -196.685 328.605 -196.355 ;
        RECT 328.275 -198.045 328.605 -197.715 ;
        RECT 328.275 -199.405 328.605 -199.075 ;
        RECT 328.275 -200.765 328.605 -200.435 ;
        RECT 328.275 -202.125 328.605 -201.795 ;
        RECT 328.275 -203.485 328.605 -203.155 ;
        RECT 328.275 -204.845 328.605 -204.515 ;
        RECT 328.275 -206.205 328.605 -205.875 ;
        RECT 328.275 -207.565 328.605 -207.235 ;
        RECT 328.275 -208.925 328.605 -208.595 ;
        RECT 328.275 -210.285 328.605 -209.955 ;
        RECT 328.275 -211.645 328.605 -211.315 ;
        RECT 328.275 -213.005 328.605 -212.675 ;
        RECT 328.275 -214.365 328.605 -214.035 ;
        RECT 328.275 -215.725 328.605 -215.395 ;
        RECT 328.275 -217.085 328.605 -216.755 ;
        RECT 328.275 -218.445 328.605 -218.115 ;
        RECT 328.275 -219.805 328.605 -219.475 ;
        RECT 328.275 -221.165 328.605 -220.835 ;
        RECT 328.275 -222.525 328.605 -222.195 ;
        RECT 328.275 -223.885 328.605 -223.555 ;
        RECT 328.275 -225.245 328.605 -224.915 ;
        RECT 328.275 -226.605 328.605 -226.275 ;
        RECT 328.275 -227.965 328.605 -227.635 ;
        RECT 328.275 -229.325 328.605 -228.995 ;
        RECT 328.275 -230.685 328.605 -230.355 ;
        RECT 328.275 -232.045 328.605 -231.715 ;
        RECT 328.275 -233.405 328.605 -233.075 ;
        RECT 328.275 -234.765 328.605 -234.435 ;
        RECT 328.275 -236.125 328.605 -235.795 ;
        RECT 328.275 -237.485 328.605 -237.155 ;
        RECT 328.275 -238.845 328.605 -238.515 ;
        RECT 328.275 -241.09 328.605 -239.96 ;
        RECT 328.28 -241.205 328.6 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 244.04 329.965 245.17 ;
        RECT 329.635 242.595 329.965 242.925 ;
        RECT 329.635 241.235 329.965 241.565 ;
        RECT 329.635 239.875 329.965 240.205 ;
        RECT 329.635 238.515 329.965 238.845 ;
        RECT 329.635 237.155 329.965 237.485 ;
        RECT 329.64 237.155 329.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 -127.325 329.965 -126.995 ;
        RECT 329.635 -128.685 329.965 -128.355 ;
        RECT 329.635 -130.045 329.965 -129.715 ;
        RECT 329.635 -131.405 329.965 -131.075 ;
        RECT 329.635 -132.765 329.965 -132.435 ;
        RECT 329.635 -134.125 329.965 -133.795 ;
        RECT 329.635 -135.485 329.965 -135.155 ;
        RECT 329.635 -136.845 329.965 -136.515 ;
        RECT 329.635 -138.205 329.965 -137.875 ;
        RECT 329.635 -139.565 329.965 -139.235 ;
        RECT 329.635 -140.925 329.965 -140.595 ;
        RECT 329.635 -142.285 329.965 -141.955 ;
        RECT 329.635 -143.645 329.965 -143.315 ;
        RECT 329.635 -145.005 329.965 -144.675 ;
        RECT 329.635 -146.365 329.965 -146.035 ;
        RECT 329.635 -147.725 329.965 -147.395 ;
        RECT 329.635 -149.085 329.965 -148.755 ;
        RECT 329.635 -150.445 329.965 -150.115 ;
        RECT 329.635 -151.805 329.965 -151.475 ;
        RECT 329.635 -153.165 329.965 -152.835 ;
        RECT 329.635 -154.525 329.965 -154.195 ;
        RECT 329.635 -155.885 329.965 -155.555 ;
        RECT 329.635 -157.245 329.965 -156.915 ;
        RECT 329.635 -158.605 329.965 -158.275 ;
        RECT 329.635 -159.965 329.965 -159.635 ;
        RECT 329.635 -161.325 329.965 -160.995 ;
        RECT 329.635 -162.685 329.965 -162.355 ;
        RECT 329.635 -164.045 329.965 -163.715 ;
        RECT 329.635 -165.405 329.965 -165.075 ;
        RECT 329.635 -166.765 329.965 -166.435 ;
        RECT 329.635 -168.125 329.965 -167.795 ;
        RECT 329.635 -169.485 329.965 -169.155 ;
        RECT 329.635 -170.845 329.965 -170.515 ;
        RECT 329.635 -172.205 329.965 -171.875 ;
        RECT 329.635 -173.565 329.965 -173.235 ;
        RECT 329.635 -174.925 329.965 -174.595 ;
        RECT 329.635 -176.285 329.965 -175.955 ;
        RECT 329.635 -177.645 329.965 -177.315 ;
        RECT 329.635 -179.005 329.965 -178.675 ;
        RECT 329.635 -180.365 329.965 -180.035 ;
        RECT 329.635 -181.725 329.965 -181.395 ;
        RECT 329.635 -183.085 329.965 -182.755 ;
        RECT 329.635 -184.445 329.965 -184.115 ;
        RECT 329.635 -185.805 329.965 -185.475 ;
        RECT 329.635 -187.165 329.965 -186.835 ;
        RECT 329.635 -188.525 329.965 -188.195 ;
        RECT 329.635 -189.885 329.965 -189.555 ;
        RECT 329.635 -191.245 329.965 -190.915 ;
        RECT 329.635 -192.605 329.965 -192.275 ;
        RECT 329.635 -193.965 329.965 -193.635 ;
        RECT 329.635 -195.325 329.965 -194.995 ;
        RECT 329.635 -196.685 329.965 -196.355 ;
        RECT 329.635 -198.045 329.965 -197.715 ;
        RECT 329.635 -199.405 329.965 -199.075 ;
        RECT 329.635 -200.765 329.965 -200.435 ;
        RECT 329.635 -202.125 329.965 -201.795 ;
        RECT 329.635 -203.485 329.965 -203.155 ;
        RECT 329.635 -204.845 329.965 -204.515 ;
        RECT 329.635 -206.205 329.965 -205.875 ;
        RECT 329.635 -207.565 329.965 -207.235 ;
        RECT 329.635 -208.925 329.965 -208.595 ;
        RECT 329.635 -210.285 329.965 -209.955 ;
        RECT 329.635 -211.645 329.965 -211.315 ;
        RECT 329.635 -213.005 329.965 -212.675 ;
        RECT 329.635 -214.365 329.965 -214.035 ;
        RECT 329.635 -215.725 329.965 -215.395 ;
        RECT 329.635 -217.085 329.965 -216.755 ;
        RECT 329.635 -218.445 329.965 -218.115 ;
        RECT 329.635 -219.805 329.965 -219.475 ;
        RECT 329.635 -221.165 329.965 -220.835 ;
        RECT 329.635 -222.525 329.965 -222.195 ;
        RECT 329.635 -223.885 329.965 -223.555 ;
        RECT 329.635 -225.245 329.965 -224.915 ;
        RECT 329.635 -226.605 329.965 -226.275 ;
        RECT 329.635 -227.965 329.965 -227.635 ;
        RECT 329.635 -229.325 329.965 -228.995 ;
        RECT 329.635 -230.685 329.965 -230.355 ;
        RECT 329.635 -232.045 329.965 -231.715 ;
        RECT 329.635 -233.405 329.965 -233.075 ;
        RECT 329.635 -234.765 329.965 -234.435 ;
        RECT 329.635 -236.125 329.965 -235.795 ;
        RECT 329.635 -237.485 329.965 -237.155 ;
        RECT 329.635 -238.845 329.965 -238.515 ;
        RECT 329.635 -241.09 329.965 -239.96 ;
        RECT 329.64 -241.205 329.96 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.31 -125.535 330.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 244.04 331.325 245.17 ;
        RECT 330.995 242.595 331.325 242.925 ;
        RECT 330.995 241.235 331.325 241.565 ;
        RECT 330.995 239.875 331.325 240.205 ;
        RECT 330.995 238.515 331.325 238.845 ;
        RECT 330.995 237.155 331.325 237.485 ;
        RECT 331 237.155 331.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 -0.845 331.325 -0.515 ;
        RECT 330.995 -2.205 331.325 -1.875 ;
        RECT 330.995 -3.565 331.325 -3.235 ;
        RECT 331 -3.565 331.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 244.04 332.685 245.17 ;
        RECT 332.355 242.595 332.685 242.925 ;
        RECT 332.355 241.235 332.685 241.565 ;
        RECT 332.355 239.875 332.685 240.205 ;
        RECT 332.355 238.515 332.685 238.845 ;
        RECT 332.355 237.155 332.685 237.485 ;
        RECT 332.36 237.155 332.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 -0.845 332.685 -0.515 ;
        RECT 332.355 -2.205 332.685 -1.875 ;
        RECT 332.355 -3.565 332.685 -3.235 ;
        RECT 332.36 -3.565 332.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 244.04 334.045 245.17 ;
        RECT 333.715 242.595 334.045 242.925 ;
        RECT 333.715 241.235 334.045 241.565 ;
        RECT 333.715 239.875 334.045 240.205 ;
        RECT 333.715 238.515 334.045 238.845 ;
        RECT 333.715 237.155 334.045 237.485 ;
        RECT 333.72 237.155 334.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 -0.845 334.045 -0.515 ;
        RECT 333.715 -2.205 334.045 -1.875 ;
        RECT 333.715 -3.565 334.045 -3.235 ;
        RECT 333.72 -3.565 334.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 -123.245 334.045 -122.915 ;
        RECT 333.715 -124.605 334.045 -124.275 ;
        RECT 333.715 -125.965 334.045 -125.635 ;
        RECT 333.715 -127.325 334.045 -126.995 ;
        RECT 333.715 -128.685 334.045 -128.355 ;
        RECT 333.715 -130.045 334.045 -129.715 ;
        RECT 333.715 -131.405 334.045 -131.075 ;
        RECT 333.715 -132.765 334.045 -132.435 ;
        RECT 333.715 -134.125 334.045 -133.795 ;
        RECT 333.715 -135.485 334.045 -135.155 ;
        RECT 333.715 -136.845 334.045 -136.515 ;
        RECT 333.715 -138.205 334.045 -137.875 ;
        RECT 333.715 -139.565 334.045 -139.235 ;
        RECT 333.715 -140.925 334.045 -140.595 ;
        RECT 333.715 -142.285 334.045 -141.955 ;
        RECT 333.715 -143.645 334.045 -143.315 ;
        RECT 333.715 -145.005 334.045 -144.675 ;
        RECT 333.715 -146.365 334.045 -146.035 ;
        RECT 333.715 -147.725 334.045 -147.395 ;
        RECT 333.715 -149.085 334.045 -148.755 ;
        RECT 333.715 -150.445 334.045 -150.115 ;
        RECT 333.715 -151.805 334.045 -151.475 ;
        RECT 333.715 -153.165 334.045 -152.835 ;
        RECT 333.715 -154.525 334.045 -154.195 ;
        RECT 333.715 -155.885 334.045 -155.555 ;
        RECT 333.715 -157.245 334.045 -156.915 ;
        RECT 333.715 -158.605 334.045 -158.275 ;
        RECT 333.715 -159.965 334.045 -159.635 ;
        RECT 333.715 -161.325 334.045 -160.995 ;
        RECT 333.715 -162.685 334.045 -162.355 ;
        RECT 333.715 -164.045 334.045 -163.715 ;
        RECT 333.715 -165.405 334.045 -165.075 ;
        RECT 333.715 -166.765 334.045 -166.435 ;
        RECT 333.715 -168.125 334.045 -167.795 ;
        RECT 333.715 -169.485 334.045 -169.155 ;
        RECT 333.715 -170.845 334.045 -170.515 ;
        RECT 333.715 -172.205 334.045 -171.875 ;
        RECT 333.715 -173.565 334.045 -173.235 ;
        RECT 333.715 -174.925 334.045 -174.595 ;
        RECT 333.715 -176.285 334.045 -175.955 ;
        RECT 333.715 -177.645 334.045 -177.315 ;
        RECT 333.715 -179.005 334.045 -178.675 ;
        RECT 333.715 -180.365 334.045 -180.035 ;
        RECT 333.715 -181.725 334.045 -181.395 ;
        RECT 333.715 -183.085 334.045 -182.755 ;
        RECT 333.715 -184.445 334.045 -184.115 ;
        RECT 333.715 -185.805 334.045 -185.475 ;
        RECT 333.715 -187.165 334.045 -186.835 ;
        RECT 333.715 -188.525 334.045 -188.195 ;
        RECT 333.715 -189.885 334.045 -189.555 ;
        RECT 333.715 -191.245 334.045 -190.915 ;
        RECT 333.715 -192.605 334.045 -192.275 ;
        RECT 333.715 -193.965 334.045 -193.635 ;
        RECT 333.715 -195.325 334.045 -194.995 ;
        RECT 333.715 -196.685 334.045 -196.355 ;
        RECT 333.715 -198.045 334.045 -197.715 ;
        RECT 333.715 -199.405 334.045 -199.075 ;
        RECT 333.715 -200.765 334.045 -200.435 ;
        RECT 333.715 -202.125 334.045 -201.795 ;
        RECT 333.715 -203.485 334.045 -203.155 ;
        RECT 333.715 -204.845 334.045 -204.515 ;
        RECT 333.715 -206.205 334.045 -205.875 ;
        RECT 333.715 -207.565 334.045 -207.235 ;
        RECT 333.715 -208.925 334.045 -208.595 ;
        RECT 333.715 -210.285 334.045 -209.955 ;
        RECT 333.715 -211.645 334.045 -211.315 ;
        RECT 333.715 -213.005 334.045 -212.675 ;
        RECT 333.715 -214.365 334.045 -214.035 ;
        RECT 333.715 -215.725 334.045 -215.395 ;
        RECT 333.715 -217.085 334.045 -216.755 ;
        RECT 333.715 -218.445 334.045 -218.115 ;
        RECT 333.715 -219.805 334.045 -219.475 ;
        RECT 333.715 -221.165 334.045 -220.835 ;
        RECT 333.715 -222.525 334.045 -222.195 ;
        RECT 333.715 -223.885 334.045 -223.555 ;
        RECT 333.715 -225.245 334.045 -224.915 ;
        RECT 333.715 -226.605 334.045 -226.275 ;
        RECT 333.715 -227.965 334.045 -227.635 ;
        RECT 333.715 -229.325 334.045 -228.995 ;
        RECT 333.715 -230.685 334.045 -230.355 ;
        RECT 333.715 -232.045 334.045 -231.715 ;
        RECT 333.715 -233.405 334.045 -233.075 ;
        RECT 333.715 -234.765 334.045 -234.435 ;
        RECT 333.715 -236.125 334.045 -235.795 ;
        RECT 333.715 -237.485 334.045 -237.155 ;
        RECT 333.715 -238.845 334.045 -238.515 ;
        RECT 333.715 -241.09 334.045 -239.96 ;
        RECT 333.72 -241.205 334.04 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 244.04 335.405 245.17 ;
        RECT 335.075 242.595 335.405 242.925 ;
        RECT 335.075 241.235 335.405 241.565 ;
        RECT 335.075 239.875 335.405 240.205 ;
        RECT 335.075 238.515 335.405 238.845 ;
        RECT 335.075 237.155 335.405 237.485 ;
        RECT 335.08 237.155 335.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 -0.845 335.405 -0.515 ;
        RECT 335.075 -2.205 335.405 -1.875 ;
        RECT 335.075 -3.565 335.405 -3.235 ;
        RECT 335.08 -3.565 335.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 -123.245 335.405 -122.915 ;
        RECT 335.075 -124.605 335.405 -124.275 ;
        RECT 335.075 -125.965 335.405 -125.635 ;
        RECT 335.075 -127.325 335.405 -126.995 ;
        RECT 335.075 -128.685 335.405 -128.355 ;
        RECT 335.075 -130.045 335.405 -129.715 ;
        RECT 335.075 -131.405 335.405 -131.075 ;
        RECT 335.075 -132.765 335.405 -132.435 ;
        RECT 335.075 -134.125 335.405 -133.795 ;
        RECT 335.075 -135.485 335.405 -135.155 ;
        RECT 335.075 -136.845 335.405 -136.515 ;
        RECT 335.075 -138.205 335.405 -137.875 ;
        RECT 335.075 -139.565 335.405 -139.235 ;
        RECT 335.075 -140.925 335.405 -140.595 ;
        RECT 335.075 -142.285 335.405 -141.955 ;
        RECT 335.075 -143.645 335.405 -143.315 ;
        RECT 335.075 -145.005 335.405 -144.675 ;
        RECT 335.075 -146.365 335.405 -146.035 ;
        RECT 335.075 -147.725 335.405 -147.395 ;
        RECT 335.075 -149.085 335.405 -148.755 ;
        RECT 335.075 -150.445 335.405 -150.115 ;
        RECT 335.075 -151.805 335.405 -151.475 ;
        RECT 335.075 -153.165 335.405 -152.835 ;
        RECT 335.075 -154.525 335.405 -154.195 ;
        RECT 335.075 -155.885 335.405 -155.555 ;
        RECT 335.075 -157.245 335.405 -156.915 ;
        RECT 335.075 -158.605 335.405 -158.275 ;
        RECT 335.075 -159.965 335.405 -159.635 ;
        RECT 335.075 -161.325 335.405 -160.995 ;
        RECT 335.075 -162.685 335.405 -162.355 ;
        RECT 335.075 -164.045 335.405 -163.715 ;
        RECT 335.075 -165.405 335.405 -165.075 ;
        RECT 335.075 -166.765 335.405 -166.435 ;
        RECT 335.075 -168.125 335.405 -167.795 ;
        RECT 335.075 -169.485 335.405 -169.155 ;
        RECT 335.075 -170.845 335.405 -170.515 ;
        RECT 335.075 -172.205 335.405 -171.875 ;
        RECT 335.075 -173.565 335.405 -173.235 ;
        RECT 335.075 -174.925 335.405 -174.595 ;
        RECT 335.075 -176.285 335.405 -175.955 ;
        RECT 335.075 -177.645 335.405 -177.315 ;
        RECT 335.075 -179.005 335.405 -178.675 ;
        RECT 335.075 -180.365 335.405 -180.035 ;
        RECT 335.075 -181.725 335.405 -181.395 ;
        RECT 335.075 -183.085 335.405 -182.755 ;
        RECT 335.075 -184.445 335.405 -184.115 ;
        RECT 335.075 -185.805 335.405 -185.475 ;
        RECT 335.075 -187.165 335.405 -186.835 ;
        RECT 335.075 -188.525 335.405 -188.195 ;
        RECT 335.075 -189.885 335.405 -189.555 ;
        RECT 335.075 -191.245 335.405 -190.915 ;
        RECT 335.075 -192.605 335.405 -192.275 ;
        RECT 335.075 -193.965 335.405 -193.635 ;
        RECT 335.075 -195.325 335.405 -194.995 ;
        RECT 335.075 -196.685 335.405 -196.355 ;
        RECT 335.075 -198.045 335.405 -197.715 ;
        RECT 335.075 -199.405 335.405 -199.075 ;
        RECT 335.075 -200.765 335.405 -200.435 ;
        RECT 335.075 -202.125 335.405 -201.795 ;
        RECT 335.075 -203.485 335.405 -203.155 ;
        RECT 335.075 -204.845 335.405 -204.515 ;
        RECT 335.075 -206.205 335.405 -205.875 ;
        RECT 335.075 -207.565 335.405 -207.235 ;
        RECT 335.075 -208.925 335.405 -208.595 ;
        RECT 335.075 -210.285 335.405 -209.955 ;
        RECT 335.075 -211.645 335.405 -211.315 ;
        RECT 335.075 -213.005 335.405 -212.675 ;
        RECT 335.075 -214.365 335.405 -214.035 ;
        RECT 335.075 -215.725 335.405 -215.395 ;
        RECT 335.075 -217.085 335.405 -216.755 ;
        RECT 335.075 -218.445 335.405 -218.115 ;
        RECT 335.075 -219.805 335.405 -219.475 ;
        RECT 335.075 -221.165 335.405 -220.835 ;
        RECT 335.075 -222.525 335.405 -222.195 ;
        RECT 335.075 -223.885 335.405 -223.555 ;
        RECT 335.075 -225.245 335.405 -224.915 ;
        RECT 335.075 -226.605 335.405 -226.275 ;
        RECT 335.075 -227.965 335.405 -227.635 ;
        RECT 335.075 -229.325 335.405 -228.995 ;
        RECT 335.075 -230.685 335.405 -230.355 ;
        RECT 335.075 -232.045 335.405 -231.715 ;
        RECT 335.075 -233.405 335.405 -233.075 ;
        RECT 335.075 -234.765 335.405 -234.435 ;
        RECT 335.075 -236.125 335.405 -235.795 ;
        RECT 335.075 -237.485 335.405 -237.155 ;
        RECT 335.075 -238.845 335.405 -238.515 ;
        RECT 335.075 -241.09 335.405 -239.96 ;
        RECT 335.08 -241.205 335.4 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 244.04 336.765 245.17 ;
        RECT 336.435 242.595 336.765 242.925 ;
        RECT 336.435 241.235 336.765 241.565 ;
        RECT 336.435 239.875 336.765 240.205 ;
        RECT 336.435 238.515 336.765 238.845 ;
        RECT 336.435 237.155 336.765 237.485 ;
        RECT 336.44 237.155 336.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 -0.845 336.765 -0.515 ;
        RECT 336.435 -2.205 336.765 -1.875 ;
        RECT 336.435 -3.565 336.765 -3.235 ;
        RECT 336.44 -3.565 336.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 -123.245 336.765 -122.915 ;
        RECT 336.435 -124.605 336.765 -124.275 ;
        RECT 336.435 -125.965 336.765 -125.635 ;
        RECT 336.435 -127.325 336.765 -126.995 ;
        RECT 336.435 -128.685 336.765 -128.355 ;
        RECT 336.435 -130.045 336.765 -129.715 ;
        RECT 336.435 -131.405 336.765 -131.075 ;
        RECT 336.435 -132.765 336.765 -132.435 ;
        RECT 336.435 -134.125 336.765 -133.795 ;
        RECT 336.435 -135.485 336.765 -135.155 ;
        RECT 336.435 -136.845 336.765 -136.515 ;
        RECT 336.435 -138.205 336.765 -137.875 ;
        RECT 336.435 -139.565 336.765 -139.235 ;
        RECT 336.435 -140.925 336.765 -140.595 ;
        RECT 336.435 -142.285 336.765 -141.955 ;
        RECT 336.435 -143.645 336.765 -143.315 ;
        RECT 336.435 -145.005 336.765 -144.675 ;
        RECT 336.435 -146.365 336.765 -146.035 ;
        RECT 336.435 -147.725 336.765 -147.395 ;
        RECT 336.435 -149.085 336.765 -148.755 ;
        RECT 336.435 -150.445 336.765 -150.115 ;
        RECT 336.435 -151.805 336.765 -151.475 ;
        RECT 336.435 -153.165 336.765 -152.835 ;
        RECT 336.435 -154.525 336.765 -154.195 ;
        RECT 336.435 -155.885 336.765 -155.555 ;
        RECT 336.435 -157.245 336.765 -156.915 ;
        RECT 336.435 -158.605 336.765 -158.275 ;
        RECT 336.435 -159.965 336.765 -159.635 ;
        RECT 336.435 -161.325 336.765 -160.995 ;
        RECT 336.435 -162.685 336.765 -162.355 ;
        RECT 336.435 -164.045 336.765 -163.715 ;
        RECT 336.435 -165.405 336.765 -165.075 ;
        RECT 336.435 -166.765 336.765 -166.435 ;
        RECT 336.435 -168.125 336.765 -167.795 ;
        RECT 336.435 -169.485 336.765 -169.155 ;
        RECT 336.435 -170.845 336.765 -170.515 ;
        RECT 336.435 -172.205 336.765 -171.875 ;
        RECT 336.435 -173.565 336.765 -173.235 ;
        RECT 336.435 -174.925 336.765 -174.595 ;
        RECT 336.435 -176.285 336.765 -175.955 ;
        RECT 336.435 -177.645 336.765 -177.315 ;
        RECT 336.435 -179.005 336.765 -178.675 ;
        RECT 336.435 -180.365 336.765 -180.035 ;
        RECT 336.435 -181.725 336.765 -181.395 ;
        RECT 336.435 -183.085 336.765 -182.755 ;
        RECT 336.435 -184.445 336.765 -184.115 ;
        RECT 336.435 -185.805 336.765 -185.475 ;
        RECT 336.435 -187.165 336.765 -186.835 ;
        RECT 336.435 -188.525 336.765 -188.195 ;
        RECT 336.435 -189.885 336.765 -189.555 ;
        RECT 336.435 -191.245 336.765 -190.915 ;
        RECT 336.435 -192.605 336.765 -192.275 ;
        RECT 336.435 -193.965 336.765 -193.635 ;
        RECT 336.435 -195.325 336.765 -194.995 ;
        RECT 336.435 -196.685 336.765 -196.355 ;
        RECT 336.435 -198.045 336.765 -197.715 ;
        RECT 336.435 -199.405 336.765 -199.075 ;
        RECT 336.435 -200.765 336.765 -200.435 ;
        RECT 336.435 -202.125 336.765 -201.795 ;
        RECT 336.435 -203.485 336.765 -203.155 ;
        RECT 336.435 -204.845 336.765 -204.515 ;
        RECT 336.435 -206.205 336.765 -205.875 ;
        RECT 336.435 -207.565 336.765 -207.235 ;
        RECT 336.435 -208.925 336.765 -208.595 ;
        RECT 336.435 -210.285 336.765 -209.955 ;
        RECT 336.435 -211.645 336.765 -211.315 ;
        RECT 336.435 -213.005 336.765 -212.675 ;
        RECT 336.435 -214.365 336.765 -214.035 ;
        RECT 336.435 -215.725 336.765 -215.395 ;
        RECT 336.435 -217.085 336.765 -216.755 ;
        RECT 336.435 -218.445 336.765 -218.115 ;
        RECT 336.435 -219.805 336.765 -219.475 ;
        RECT 336.435 -221.165 336.765 -220.835 ;
        RECT 336.435 -222.525 336.765 -222.195 ;
        RECT 336.435 -223.885 336.765 -223.555 ;
        RECT 336.435 -225.245 336.765 -224.915 ;
        RECT 336.435 -226.605 336.765 -226.275 ;
        RECT 336.435 -227.965 336.765 -227.635 ;
        RECT 336.435 -229.325 336.765 -228.995 ;
        RECT 336.435 -230.685 336.765 -230.355 ;
        RECT 336.435 -232.045 336.765 -231.715 ;
        RECT 336.435 -233.405 336.765 -233.075 ;
        RECT 336.435 -234.765 336.765 -234.435 ;
        RECT 336.435 -236.125 336.765 -235.795 ;
        RECT 336.435 -237.485 336.765 -237.155 ;
        RECT 336.435 -238.845 336.765 -238.515 ;
        RECT 336.435 -241.09 336.765 -239.96 ;
        RECT 336.44 -241.205 336.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 244.04 338.125 245.17 ;
        RECT 337.795 242.595 338.125 242.925 ;
        RECT 337.795 241.235 338.125 241.565 ;
        RECT 337.795 239.875 338.125 240.205 ;
        RECT 337.795 238.515 338.125 238.845 ;
        RECT 337.795 237.155 338.125 237.485 ;
        RECT 337.8 237.155 338.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 -0.845 338.125 -0.515 ;
        RECT 337.795 -2.205 338.125 -1.875 ;
        RECT 337.795 -3.565 338.125 -3.235 ;
        RECT 337.8 -3.565 338.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 -123.245 338.125 -122.915 ;
        RECT 337.795 -124.605 338.125 -124.275 ;
        RECT 337.795 -125.965 338.125 -125.635 ;
        RECT 337.795 -127.325 338.125 -126.995 ;
        RECT 337.795 -128.685 338.125 -128.355 ;
        RECT 337.795 -130.045 338.125 -129.715 ;
        RECT 337.795 -131.405 338.125 -131.075 ;
        RECT 337.795 -132.765 338.125 -132.435 ;
        RECT 337.795 -134.125 338.125 -133.795 ;
        RECT 337.795 -135.485 338.125 -135.155 ;
        RECT 337.795 -136.845 338.125 -136.515 ;
        RECT 337.795 -138.205 338.125 -137.875 ;
        RECT 337.795 -139.565 338.125 -139.235 ;
        RECT 337.795 -140.925 338.125 -140.595 ;
        RECT 337.795 -142.285 338.125 -141.955 ;
        RECT 337.795 -143.645 338.125 -143.315 ;
        RECT 337.795 -145.005 338.125 -144.675 ;
        RECT 337.795 -146.365 338.125 -146.035 ;
        RECT 337.795 -147.725 338.125 -147.395 ;
        RECT 337.795 -149.085 338.125 -148.755 ;
        RECT 337.795 -150.445 338.125 -150.115 ;
        RECT 337.795 -151.805 338.125 -151.475 ;
        RECT 337.795 -153.165 338.125 -152.835 ;
        RECT 337.795 -154.525 338.125 -154.195 ;
        RECT 337.795 -155.885 338.125 -155.555 ;
        RECT 337.795 -157.245 338.125 -156.915 ;
        RECT 337.795 -158.605 338.125 -158.275 ;
        RECT 337.795 -159.965 338.125 -159.635 ;
        RECT 337.795 -161.325 338.125 -160.995 ;
        RECT 337.795 -162.685 338.125 -162.355 ;
        RECT 337.795 -164.045 338.125 -163.715 ;
        RECT 337.795 -165.405 338.125 -165.075 ;
        RECT 337.795 -166.765 338.125 -166.435 ;
        RECT 337.795 -168.125 338.125 -167.795 ;
        RECT 337.795 -169.485 338.125 -169.155 ;
        RECT 337.795 -170.845 338.125 -170.515 ;
        RECT 337.795 -172.205 338.125 -171.875 ;
        RECT 337.795 -173.565 338.125 -173.235 ;
        RECT 337.795 -174.925 338.125 -174.595 ;
        RECT 337.795 -176.285 338.125 -175.955 ;
        RECT 337.795 -177.645 338.125 -177.315 ;
        RECT 337.795 -179.005 338.125 -178.675 ;
        RECT 337.795 -180.365 338.125 -180.035 ;
        RECT 337.795 -181.725 338.125 -181.395 ;
        RECT 337.795 -183.085 338.125 -182.755 ;
        RECT 337.795 -184.445 338.125 -184.115 ;
        RECT 337.795 -185.805 338.125 -185.475 ;
        RECT 337.795 -187.165 338.125 -186.835 ;
        RECT 337.795 -188.525 338.125 -188.195 ;
        RECT 337.795 -189.885 338.125 -189.555 ;
        RECT 337.795 -191.245 338.125 -190.915 ;
        RECT 337.795 -192.605 338.125 -192.275 ;
        RECT 337.795 -193.965 338.125 -193.635 ;
        RECT 337.795 -195.325 338.125 -194.995 ;
        RECT 337.795 -196.685 338.125 -196.355 ;
        RECT 337.795 -198.045 338.125 -197.715 ;
        RECT 337.795 -199.405 338.125 -199.075 ;
        RECT 337.795 -200.765 338.125 -200.435 ;
        RECT 337.795 -202.125 338.125 -201.795 ;
        RECT 337.795 -203.485 338.125 -203.155 ;
        RECT 337.795 -204.845 338.125 -204.515 ;
        RECT 337.795 -206.205 338.125 -205.875 ;
        RECT 337.795 -207.565 338.125 -207.235 ;
        RECT 337.795 -208.925 338.125 -208.595 ;
        RECT 337.795 -210.285 338.125 -209.955 ;
        RECT 337.795 -211.645 338.125 -211.315 ;
        RECT 337.795 -213.005 338.125 -212.675 ;
        RECT 337.795 -214.365 338.125 -214.035 ;
        RECT 337.795 -215.725 338.125 -215.395 ;
        RECT 337.795 -217.085 338.125 -216.755 ;
        RECT 337.795 -218.445 338.125 -218.115 ;
        RECT 337.795 -219.805 338.125 -219.475 ;
        RECT 337.795 -221.165 338.125 -220.835 ;
        RECT 337.795 -222.525 338.125 -222.195 ;
        RECT 337.795 -223.885 338.125 -223.555 ;
        RECT 337.795 -225.245 338.125 -224.915 ;
        RECT 337.795 -226.605 338.125 -226.275 ;
        RECT 337.795 -227.965 338.125 -227.635 ;
        RECT 337.795 -229.325 338.125 -228.995 ;
        RECT 337.795 -230.685 338.125 -230.355 ;
        RECT 337.795 -232.045 338.125 -231.715 ;
        RECT 337.795 -233.405 338.125 -233.075 ;
        RECT 337.795 -234.765 338.125 -234.435 ;
        RECT 337.795 -236.125 338.125 -235.795 ;
        RECT 337.795 -237.485 338.125 -237.155 ;
        RECT 337.795 -238.845 338.125 -238.515 ;
        RECT 337.795 -241.09 338.125 -239.96 ;
        RECT 337.8 -241.205 338.12 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 244.04 339.485 245.17 ;
        RECT 339.155 242.595 339.485 242.925 ;
        RECT 339.155 241.235 339.485 241.565 ;
        RECT 339.155 239.875 339.485 240.205 ;
        RECT 339.155 238.515 339.485 238.845 ;
        RECT 339.155 237.155 339.485 237.485 ;
        RECT 339.16 237.155 339.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 -0.845 339.485 -0.515 ;
        RECT 339.155 -2.205 339.485 -1.875 ;
        RECT 339.155 -3.565 339.485 -3.235 ;
        RECT 339.16 -3.565 339.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 -123.245 339.485 -122.915 ;
        RECT 339.155 -124.605 339.485 -124.275 ;
        RECT 339.155 -125.965 339.485 -125.635 ;
        RECT 339.155 -127.325 339.485 -126.995 ;
        RECT 339.155 -128.685 339.485 -128.355 ;
        RECT 339.155 -130.045 339.485 -129.715 ;
        RECT 339.155 -131.405 339.485 -131.075 ;
        RECT 339.155 -132.765 339.485 -132.435 ;
        RECT 339.155 -134.125 339.485 -133.795 ;
        RECT 339.155 -135.485 339.485 -135.155 ;
        RECT 339.155 -136.845 339.485 -136.515 ;
        RECT 339.155 -138.205 339.485 -137.875 ;
        RECT 339.155 -139.565 339.485 -139.235 ;
        RECT 339.155 -140.925 339.485 -140.595 ;
        RECT 339.155 -142.285 339.485 -141.955 ;
        RECT 339.155 -143.645 339.485 -143.315 ;
        RECT 339.155 -145.005 339.485 -144.675 ;
        RECT 339.155 -146.365 339.485 -146.035 ;
        RECT 339.155 -147.725 339.485 -147.395 ;
        RECT 339.155 -149.085 339.485 -148.755 ;
        RECT 339.155 -150.445 339.485 -150.115 ;
        RECT 339.155 -151.805 339.485 -151.475 ;
        RECT 339.155 -153.165 339.485 -152.835 ;
        RECT 339.155 -154.525 339.485 -154.195 ;
        RECT 339.155 -155.885 339.485 -155.555 ;
        RECT 339.155 -157.245 339.485 -156.915 ;
        RECT 339.155 -158.605 339.485 -158.275 ;
        RECT 339.155 -159.965 339.485 -159.635 ;
        RECT 339.155 -161.325 339.485 -160.995 ;
        RECT 339.155 -162.685 339.485 -162.355 ;
        RECT 339.155 -164.045 339.485 -163.715 ;
        RECT 339.155 -165.405 339.485 -165.075 ;
        RECT 339.155 -166.765 339.485 -166.435 ;
        RECT 339.155 -168.125 339.485 -167.795 ;
        RECT 339.155 -169.485 339.485 -169.155 ;
        RECT 339.155 -170.845 339.485 -170.515 ;
        RECT 339.155 -172.205 339.485 -171.875 ;
        RECT 339.155 -173.565 339.485 -173.235 ;
        RECT 339.155 -174.925 339.485 -174.595 ;
        RECT 339.155 -176.285 339.485 -175.955 ;
        RECT 339.155 -177.645 339.485 -177.315 ;
        RECT 339.155 -179.005 339.485 -178.675 ;
        RECT 339.155 -180.365 339.485 -180.035 ;
        RECT 339.155 -181.725 339.485 -181.395 ;
        RECT 339.155 -183.085 339.485 -182.755 ;
        RECT 339.155 -184.445 339.485 -184.115 ;
        RECT 339.155 -185.805 339.485 -185.475 ;
        RECT 339.155 -187.165 339.485 -186.835 ;
        RECT 339.155 -188.525 339.485 -188.195 ;
        RECT 339.155 -189.885 339.485 -189.555 ;
        RECT 339.155 -191.245 339.485 -190.915 ;
        RECT 339.155 -192.605 339.485 -192.275 ;
        RECT 339.155 -193.965 339.485 -193.635 ;
        RECT 339.155 -195.325 339.485 -194.995 ;
        RECT 339.155 -196.685 339.485 -196.355 ;
        RECT 339.155 -198.045 339.485 -197.715 ;
        RECT 339.155 -199.405 339.485 -199.075 ;
        RECT 339.155 -200.765 339.485 -200.435 ;
        RECT 339.155 -202.125 339.485 -201.795 ;
        RECT 339.155 -203.485 339.485 -203.155 ;
        RECT 339.155 -204.845 339.485 -204.515 ;
        RECT 339.155 -206.205 339.485 -205.875 ;
        RECT 339.155 -207.565 339.485 -207.235 ;
        RECT 339.155 -208.925 339.485 -208.595 ;
        RECT 339.155 -210.285 339.485 -209.955 ;
        RECT 339.155 -211.645 339.485 -211.315 ;
        RECT 339.155 -213.005 339.485 -212.675 ;
        RECT 339.155 -214.365 339.485 -214.035 ;
        RECT 339.155 -215.725 339.485 -215.395 ;
        RECT 339.155 -217.085 339.485 -216.755 ;
        RECT 339.155 -218.445 339.485 -218.115 ;
        RECT 339.155 -219.805 339.485 -219.475 ;
        RECT 339.155 -221.165 339.485 -220.835 ;
        RECT 339.155 -222.525 339.485 -222.195 ;
        RECT 339.155 -223.885 339.485 -223.555 ;
        RECT 339.155 -225.245 339.485 -224.915 ;
        RECT 339.155 -226.605 339.485 -226.275 ;
        RECT 339.155 -227.965 339.485 -227.635 ;
        RECT 339.155 -229.325 339.485 -228.995 ;
        RECT 339.155 -230.685 339.485 -230.355 ;
        RECT 339.155 -232.045 339.485 -231.715 ;
        RECT 339.155 -233.405 339.485 -233.075 ;
        RECT 339.155 -234.765 339.485 -234.435 ;
        RECT 339.155 -236.125 339.485 -235.795 ;
        RECT 339.155 -237.485 339.485 -237.155 ;
        RECT 339.155 -238.845 339.485 -238.515 ;
        RECT 339.155 -241.09 339.485 -239.96 ;
        RECT 339.16 -241.205 339.48 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 244.04 340.845 245.17 ;
        RECT 340.515 242.595 340.845 242.925 ;
        RECT 340.515 241.235 340.845 241.565 ;
        RECT 340.515 239.875 340.845 240.205 ;
        RECT 340.515 238.515 340.845 238.845 ;
        RECT 340.515 237.155 340.845 237.485 ;
        RECT 340.52 237.155 340.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 -127.325 340.845 -126.995 ;
        RECT 340.515 -128.685 340.845 -128.355 ;
        RECT 340.515 -130.045 340.845 -129.715 ;
        RECT 340.515 -131.405 340.845 -131.075 ;
        RECT 340.515 -132.765 340.845 -132.435 ;
        RECT 340.515 -134.125 340.845 -133.795 ;
        RECT 340.515 -135.485 340.845 -135.155 ;
        RECT 340.515 -136.845 340.845 -136.515 ;
        RECT 340.515 -138.205 340.845 -137.875 ;
        RECT 340.515 -139.565 340.845 -139.235 ;
        RECT 340.515 -140.925 340.845 -140.595 ;
        RECT 340.515 -142.285 340.845 -141.955 ;
        RECT 340.515 -143.645 340.845 -143.315 ;
        RECT 340.515 -145.005 340.845 -144.675 ;
        RECT 340.515 -146.365 340.845 -146.035 ;
        RECT 340.515 -147.725 340.845 -147.395 ;
        RECT 340.515 -149.085 340.845 -148.755 ;
        RECT 340.515 -150.445 340.845 -150.115 ;
        RECT 340.515 -151.805 340.845 -151.475 ;
        RECT 340.515 -153.165 340.845 -152.835 ;
        RECT 340.515 -154.525 340.845 -154.195 ;
        RECT 340.515 -155.885 340.845 -155.555 ;
        RECT 340.515 -157.245 340.845 -156.915 ;
        RECT 340.515 -158.605 340.845 -158.275 ;
        RECT 340.515 -159.965 340.845 -159.635 ;
        RECT 340.515 -161.325 340.845 -160.995 ;
        RECT 340.515 -162.685 340.845 -162.355 ;
        RECT 340.515 -164.045 340.845 -163.715 ;
        RECT 340.515 -165.405 340.845 -165.075 ;
        RECT 340.515 -166.765 340.845 -166.435 ;
        RECT 340.515 -168.125 340.845 -167.795 ;
        RECT 340.515 -169.485 340.845 -169.155 ;
        RECT 340.515 -170.845 340.845 -170.515 ;
        RECT 340.515 -172.205 340.845 -171.875 ;
        RECT 340.515 -173.565 340.845 -173.235 ;
        RECT 340.515 -174.925 340.845 -174.595 ;
        RECT 340.515 -176.285 340.845 -175.955 ;
        RECT 340.515 -177.645 340.845 -177.315 ;
        RECT 340.515 -179.005 340.845 -178.675 ;
        RECT 340.515 -180.365 340.845 -180.035 ;
        RECT 340.515 -181.725 340.845 -181.395 ;
        RECT 340.515 -183.085 340.845 -182.755 ;
        RECT 340.515 -184.445 340.845 -184.115 ;
        RECT 340.515 -185.805 340.845 -185.475 ;
        RECT 340.515 -187.165 340.845 -186.835 ;
        RECT 340.515 -188.525 340.845 -188.195 ;
        RECT 340.515 -189.885 340.845 -189.555 ;
        RECT 340.515 -191.245 340.845 -190.915 ;
        RECT 340.515 -192.605 340.845 -192.275 ;
        RECT 340.515 -193.965 340.845 -193.635 ;
        RECT 340.515 -195.325 340.845 -194.995 ;
        RECT 340.515 -196.685 340.845 -196.355 ;
        RECT 340.515 -198.045 340.845 -197.715 ;
        RECT 340.515 -199.405 340.845 -199.075 ;
        RECT 340.515 -200.765 340.845 -200.435 ;
        RECT 340.515 -202.125 340.845 -201.795 ;
        RECT 340.515 -203.485 340.845 -203.155 ;
        RECT 340.515 -204.845 340.845 -204.515 ;
        RECT 340.515 -206.205 340.845 -205.875 ;
        RECT 340.515 -207.565 340.845 -207.235 ;
        RECT 340.515 -208.925 340.845 -208.595 ;
        RECT 340.515 -210.285 340.845 -209.955 ;
        RECT 340.515 -211.645 340.845 -211.315 ;
        RECT 340.515 -213.005 340.845 -212.675 ;
        RECT 340.515 -214.365 340.845 -214.035 ;
        RECT 340.515 -215.725 340.845 -215.395 ;
        RECT 340.515 -217.085 340.845 -216.755 ;
        RECT 340.515 -218.445 340.845 -218.115 ;
        RECT 340.515 -219.805 340.845 -219.475 ;
        RECT 340.515 -221.165 340.845 -220.835 ;
        RECT 340.515 -222.525 340.845 -222.195 ;
        RECT 340.515 -223.885 340.845 -223.555 ;
        RECT 340.515 -225.245 340.845 -224.915 ;
        RECT 340.515 -226.605 340.845 -226.275 ;
        RECT 340.515 -227.965 340.845 -227.635 ;
        RECT 340.515 -229.325 340.845 -228.995 ;
        RECT 340.515 -230.685 340.845 -230.355 ;
        RECT 340.515 -232.045 340.845 -231.715 ;
        RECT 340.515 -233.405 340.845 -233.075 ;
        RECT 340.515 -234.765 340.845 -234.435 ;
        RECT 340.515 -236.125 340.845 -235.795 ;
        RECT 340.515 -237.485 340.845 -237.155 ;
        RECT 340.515 -238.845 340.845 -238.515 ;
        RECT 340.515 -241.09 340.845 -239.96 ;
        RECT 340.52 -241.205 340.84 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.21 -125.535 341.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.875 244.04 342.205 245.17 ;
        RECT 341.875 242.595 342.205 242.925 ;
        RECT 341.875 241.235 342.205 241.565 ;
        RECT 341.875 239.875 342.205 240.205 ;
        RECT 341.875 238.515 342.205 238.845 ;
        RECT 341.875 237.155 342.205 237.485 ;
        RECT 341.88 237.155 342.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 244.04 343.565 245.17 ;
        RECT 343.235 242.595 343.565 242.925 ;
        RECT 343.235 241.235 343.565 241.565 ;
        RECT 343.235 239.875 343.565 240.205 ;
        RECT 343.235 238.515 343.565 238.845 ;
        RECT 343.235 237.155 343.565 237.485 ;
        RECT 343.24 237.155 343.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 -0.845 343.565 -0.515 ;
        RECT 343.235 -2.205 343.565 -1.875 ;
        RECT 343.235 -3.565 343.565 -3.235 ;
        RECT 343.24 -3.565 343.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 244.04 344.925 245.17 ;
        RECT 344.595 242.595 344.925 242.925 ;
        RECT 344.595 241.235 344.925 241.565 ;
        RECT 344.595 239.875 344.925 240.205 ;
        RECT 344.595 238.515 344.925 238.845 ;
        RECT 344.595 237.155 344.925 237.485 ;
        RECT 344.6 237.155 344.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 -0.845 344.925 -0.515 ;
        RECT 344.595 -2.205 344.925 -1.875 ;
        RECT 344.595 -3.565 344.925 -3.235 ;
        RECT 344.6 -3.565 344.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 244.04 308.205 245.17 ;
        RECT 307.875 242.595 308.205 242.925 ;
        RECT 307.875 241.235 308.205 241.565 ;
        RECT 307.875 239.875 308.205 240.205 ;
        RECT 307.875 238.515 308.205 238.845 ;
        RECT 307.875 237.155 308.205 237.485 ;
        RECT 307.88 237.155 308.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 -127.325 308.205 -126.995 ;
        RECT 307.875 -128.685 308.205 -128.355 ;
        RECT 307.875 -130.045 308.205 -129.715 ;
        RECT 307.875 -131.405 308.205 -131.075 ;
        RECT 307.875 -132.765 308.205 -132.435 ;
        RECT 307.875 -134.125 308.205 -133.795 ;
        RECT 307.875 -135.485 308.205 -135.155 ;
        RECT 307.875 -136.845 308.205 -136.515 ;
        RECT 307.875 -138.205 308.205 -137.875 ;
        RECT 307.875 -139.565 308.205 -139.235 ;
        RECT 307.875 -140.925 308.205 -140.595 ;
        RECT 307.875 -142.285 308.205 -141.955 ;
        RECT 307.875 -143.645 308.205 -143.315 ;
        RECT 307.875 -145.005 308.205 -144.675 ;
        RECT 307.875 -146.365 308.205 -146.035 ;
        RECT 307.875 -147.725 308.205 -147.395 ;
        RECT 307.875 -149.085 308.205 -148.755 ;
        RECT 307.875 -150.445 308.205 -150.115 ;
        RECT 307.875 -151.805 308.205 -151.475 ;
        RECT 307.875 -153.165 308.205 -152.835 ;
        RECT 307.875 -154.525 308.205 -154.195 ;
        RECT 307.875 -155.885 308.205 -155.555 ;
        RECT 307.875 -157.245 308.205 -156.915 ;
        RECT 307.875 -158.605 308.205 -158.275 ;
        RECT 307.875 -159.965 308.205 -159.635 ;
        RECT 307.875 -161.325 308.205 -160.995 ;
        RECT 307.875 -162.685 308.205 -162.355 ;
        RECT 307.875 -164.045 308.205 -163.715 ;
        RECT 307.875 -165.405 308.205 -165.075 ;
        RECT 307.875 -166.765 308.205 -166.435 ;
        RECT 307.875 -168.125 308.205 -167.795 ;
        RECT 307.875 -169.485 308.205 -169.155 ;
        RECT 307.875 -170.845 308.205 -170.515 ;
        RECT 307.875 -172.205 308.205 -171.875 ;
        RECT 307.875 -173.565 308.205 -173.235 ;
        RECT 307.875 -174.925 308.205 -174.595 ;
        RECT 307.875 -176.285 308.205 -175.955 ;
        RECT 307.875 -177.645 308.205 -177.315 ;
        RECT 307.875 -179.005 308.205 -178.675 ;
        RECT 307.875 -180.365 308.205 -180.035 ;
        RECT 307.875 -181.725 308.205 -181.395 ;
        RECT 307.875 -183.085 308.205 -182.755 ;
        RECT 307.875 -184.445 308.205 -184.115 ;
        RECT 307.875 -185.805 308.205 -185.475 ;
        RECT 307.875 -187.165 308.205 -186.835 ;
        RECT 307.875 -188.525 308.205 -188.195 ;
        RECT 307.875 -189.885 308.205 -189.555 ;
        RECT 307.875 -191.245 308.205 -190.915 ;
        RECT 307.875 -192.605 308.205 -192.275 ;
        RECT 307.875 -193.965 308.205 -193.635 ;
        RECT 307.875 -195.325 308.205 -194.995 ;
        RECT 307.875 -196.685 308.205 -196.355 ;
        RECT 307.875 -198.045 308.205 -197.715 ;
        RECT 307.875 -199.405 308.205 -199.075 ;
        RECT 307.875 -200.765 308.205 -200.435 ;
        RECT 307.875 -202.125 308.205 -201.795 ;
        RECT 307.875 -203.485 308.205 -203.155 ;
        RECT 307.875 -204.845 308.205 -204.515 ;
        RECT 307.875 -206.205 308.205 -205.875 ;
        RECT 307.875 -207.565 308.205 -207.235 ;
        RECT 307.875 -208.925 308.205 -208.595 ;
        RECT 307.875 -210.285 308.205 -209.955 ;
        RECT 307.875 -211.645 308.205 -211.315 ;
        RECT 307.875 -213.005 308.205 -212.675 ;
        RECT 307.875 -214.365 308.205 -214.035 ;
        RECT 307.875 -215.725 308.205 -215.395 ;
        RECT 307.875 -217.085 308.205 -216.755 ;
        RECT 307.875 -218.445 308.205 -218.115 ;
        RECT 307.875 -219.805 308.205 -219.475 ;
        RECT 307.875 -221.165 308.205 -220.835 ;
        RECT 307.875 -222.525 308.205 -222.195 ;
        RECT 307.875 -223.885 308.205 -223.555 ;
        RECT 307.875 -225.245 308.205 -224.915 ;
        RECT 307.875 -226.605 308.205 -226.275 ;
        RECT 307.875 -227.965 308.205 -227.635 ;
        RECT 307.875 -229.325 308.205 -228.995 ;
        RECT 307.875 -230.685 308.205 -230.355 ;
        RECT 307.875 -232.045 308.205 -231.715 ;
        RECT 307.875 -233.405 308.205 -233.075 ;
        RECT 307.875 -234.765 308.205 -234.435 ;
        RECT 307.875 -236.125 308.205 -235.795 ;
        RECT 307.875 -237.485 308.205 -237.155 ;
        RECT 307.875 -238.845 308.205 -238.515 ;
        RECT 307.875 -241.09 308.205 -239.96 ;
        RECT 307.88 -241.205 308.2 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.51 -125.535 308.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 244.04 309.565 245.17 ;
        RECT 309.235 242.595 309.565 242.925 ;
        RECT 309.235 241.235 309.565 241.565 ;
        RECT 309.235 239.875 309.565 240.205 ;
        RECT 309.235 238.515 309.565 238.845 ;
        RECT 309.235 237.155 309.565 237.485 ;
        RECT 309.24 237.155 309.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 -0.845 309.565 -0.515 ;
        RECT 309.235 -2.205 309.565 -1.875 ;
        RECT 309.235 -3.565 309.565 -3.235 ;
        RECT 309.24 -3.565 309.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 244.04 310.925 245.17 ;
        RECT 310.595 242.595 310.925 242.925 ;
        RECT 310.595 241.235 310.925 241.565 ;
        RECT 310.595 239.875 310.925 240.205 ;
        RECT 310.595 238.515 310.925 238.845 ;
        RECT 310.595 237.155 310.925 237.485 ;
        RECT 310.6 237.155 310.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 -0.845 310.925 -0.515 ;
        RECT 310.595 -2.205 310.925 -1.875 ;
        RECT 310.595 -3.565 310.925 -3.235 ;
        RECT 310.6 -3.565 310.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 244.04 312.285 245.17 ;
        RECT 311.955 242.595 312.285 242.925 ;
        RECT 311.955 241.235 312.285 241.565 ;
        RECT 311.955 239.875 312.285 240.205 ;
        RECT 311.955 238.515 312.285 238.845 ;
        RECT 311.955 237.155 312.285 237.485 ;
        RECT 311.96 237.155 312.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 -0.845 312.285 -0.515 ;
        RECT 311.955 -2.205 312.285 -1.875 ;
        RECT 311.955 -3.565 312.285 -3.235 ;
        RECT 311.96 -3.565 312.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 -123.245 312.285 -122.915 ;
        RECT 311.955 -124.605 312.285 -124.275 ;
        RECT 311.955 -125.965 312.285 -125.635 ;
        RECT 311.955 -127.325 312.285 -126.995 ;
        RECT 311.955 -128.685 312.285 -128.355 ;
        RECT 311.955 -130.045 312.285 -129.715 ;
        RECT 311.955 -131.405 312.285 -131.075 ;
        RECT 311.955 -132.765 312.285 -132.435 ;
        RECT 311.955 -134.125 312.285 -133.795 ;
        RECT 311.955 -135.485 312.285 -135.155 ;
        RECT 311.955 -136.845 312.285 -136.515 ;
        RECT 311.955 -138.205 312.285 -137.875 ;
        RECT 311.955 -139.565 312.285 -139.235 ;
        RECT 311.955 -140.925 312.285 -140.595 ;
        RECT 311.955 -142.285 312.285 -141.955 ;
        RECT 311.955 -143.645 312.285 -143.315 ;
        RECT 311.955 -145.005 312.285 -144.675 ;
        RECT 311.955 -146.365 312.285 -146.035 ;
        RECT 311.955 -147.725 312.285 -147.395 ;
        RECT 311.955 -149.085 312.285 -148.755 ;
        RECT 311.955 -150.445 312.285 -150.115 ;
        RECT 311.955 -151.805 312.285 -151.475 ;
        RECT 311.955 -153.165 312.285 -152.835 ;
        RECT 311.955 -154.525 312.285 -154.195 ;
        RECT 311.955 -155.885 312.285 -155.555 ;
        RECT 311.955 -157.245 312.285 -156.915 ;
        RECT 311.955 -158.605 312.285 -158.275 ;
        RECT 311.955 -159.965 312.285 -159.635 ;
        RECT 311.955 -161.325 312.285 -160.995 ;
        RECT 311.955 -162.685 312.285 -162.355 ;
        RECT 311.955 -164.045 312.285 -163.715 ;
        RECT 311.955 -165.405 312.285 -165.075 ;
        RECT 311.955 -166.765 312.285 -166.435 ;
        RECT 311.955 -168.125 312.285 -167.795 ;
        RECT 311.955 -169.485 312.285 -169.155 ;
        RECT 311.955 -170.845 312.285 -170.515 ;
        RECT 311.955 -172.205 312.285 -171.875 ;
        RECT 311.955 -173.565 312.285 -173.235 ;
        RECT 311.955 -174.925 312.285 -174.595 ;
        RECT 311.955 -176.285 312.285 -175.955 ;
        RECT 311.955 -177.645 312.285 -177.315 ;
        RECT 311.955 -179.005 312.285 -178.675 ;
        RECT 311.955 -180.365 312.285 -180.035 ;
        RECT 311.955 -181.725 312.285 -181.395 ;
        RECT 311.955 -183.085 312.285 -182.755 ;
        RECT 311.955 -184.445 312.285 -184.115 ;
        RECT 311.955 -185.805 312.285 -185.475 ;
        RECT 311.955 -187.165 312.285 -186.835 ;
        RECT 311.955 -188.525 312.285 -188.195 ;
        RECT 311.955 -189.885 312.285 -189.555 ;
        RECT 311.955 -191.245 312.285 -190.915 ;
        RECT 311.955 -192.605 312.285 -192.275 ;
        RECT 311.955 -193.965 312.285 -193.635 ;
        RECT 311.955 -195.325 312.285 -194.995 ;
        RECT 311.955 -196.685 312.285 -196.355 ;
        RECT 311.955 -198.045 312.285 -197.715 ;
        RECT 311.955 -199.405 312.285 -199.075 ;
        RECT 311.955 -200.765 312.285 -200.435 ;
        RECT 311.955 -202.125 312.285 -201.795 ;
        RECT 311.955 -203.485 312.285 -203.155 ;
        RECT 311.955 -204.845 312.285 -204.515 ;
        RECT 311.955 -206.205 312.285 -205.875 ;
        RECT 311.955 -207.565 312.285 -207.235 ;
        RECT 311.955 -208.925 312.285 -208.595 ;
        RECT 311.955 -210.285 312.285 -209.955 ;
        RECT 311.955 -211.645 312.285 -211.315 ;
        RECT 311.955 -213.005 312.285 -212.675 ;
        RECT 311.955 -214.365 312.285 -214.035 ;
        RECT 311.955 -215.725 312.285 -215.395 ;
        RECT 311.955 -217.085 312.285 -216.755 ;
        RECT 311.955 -218.445 312.285 -218.115 ;
        RECT 311.955 -219.805 312.285 -219.475 ;
        RECT 311.955 -221.165 312.285 -220.835 ;
        RECT 311.955 -222.525 312.285 -222.195 ;
        RECT 311.955 -223.885 312.285 -223.555 ;
        RECT 311.955 -225.245 312.285 -224.915 ;
        RECT 311.955 -226.605 312.285 -226.275 ;
        RECT 311.955 -227.965 312.285 -227.635 ;
        RECT 311.955 -229.325 312.285 -228.995 ;
        RECT 311.955 -230.685 312.285 -230.355 ;
        RECT 311.955 -232.045 312.285 -231.715 ;
        RECT 311.955 -233.405 312.285 -233.075 ;
        RECT 311.955 -234.765 312.285 -234.435 ;
        RECT 311.955 -236.125 312.285 -235.795 ;
        RECT 311.955 -237.485 312.285 -237.155 ;
        RECT 311.955 -238.845 312.285 -238.515 ;
        RECT 311.955 -241.09 312.285 -239.96 ;
        RECT 311.96 -241.205 312.28 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 244.04 313.645 245.17 ;
        RECT 313.315 242.595 313.645 242.925 ;
        RECT 313.315 241.235 313.645 241.565 ;
        RECT 313.315 239.875 313.645 240.205 ;
        RECT 313.315 238.515 313.645 238.845 ;
        RECT 313.315 237.155 313.645 237.485 ;
        RECT 313.32 237.155 313.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 -0.845 313.645 -0.515 ;
        RECT 313.315 -2.205 313.645 -1.875 ;
        RECT 313.315 -3.565 313.645 -3.235 ;
        RECT 313.32 -3.565 313.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 -123.245 313.645 -122.915 ;
        RECT 313.315 -124.605 313.645 -124.275 ;
        RECT 313.315 -125.965 313.645 -125.635 ;
        RECT 313.315 -127.325 313.645 -126.995 ;
        RECT 313.315 -128.685 313.645 -128.355 ;
        RECT 313.315 -130.045 313.645 -129.715 ;
        RECT 313.315 -131.405 313.645 -131.075 ;
        RECT 313.315 -132.765 313.645 -132.435 ;
        RECT 313.315 -134.125 313.645 -133.795 ;
        RECT 313.315 -135.485 313.645 -135.155 ;
        RECT 313.315 -136.845 313.645 -136.515 ;
        RECT 313.315 -138.205 313.645 -137.875 ;
        RECT 313.315 -139.565 313.645 -139.235 ;
        RECT 313.315 -140.925 313.645 -140.595 ;
        RECT 313.315 -142.285 313.645 -141.955 ;
        RECT 313.315 -143.645 313.645 -143.315 ;
        RECT 313.315 -145.005 313.645 -144.675 ;
        RECT 313.315 -146.365 313.645 -146.035 ;
        RECT 313.315 -147.725 313.645 -147.395 ;
        RECT 313.315 -149.085 313.645 -148.755 ;
        RECT 313.315 -150.445 313.645 -150.115 ;
        RECT 313.315 -151.805 313.645 -151.475 ;
        RECT 313.315 -153.165 313.645 -152.835 ;
        RECT 313.315 -154.525 313.645 -154.195 ;
        RECT 313.315 -155.885 313.645 -155.555 ;
        RECT 313.315 -157.245 313.645 -156.915 ;
        RECT 313.315 -158.605 313.645 -158.275 ;
        RECT 313.315 -159.965 313.645 -159.635 ;
        RECT 313.315 -161.325 313.645 -160.995 ;
        RECT 313.315 -162.685 313.645 -162.355 ;
        RECT 313.315 -164.045 313.645 -163.715 ;
        RECT 313.315 -165.405 313.645 -165.075 ;
        RECT 313.315 -166.765 313.645 -166.435 ;
        RECT 313.315 -168.125 313.645 -167.795 ;
        RECT 313.315 -169.485 313.645 -169.155 ;
        RECT 313.315 -170.845 313.645 -170.515 ;
        RECT 313.315 -172.205 313.645 -171.875 ;
        RECT 313.315 -173.565 313.645 -173.235 ;
        RECT 313.315 -174.925 313.645 -174.595 ;
        RECT 313.315 -176.285 313.645 -175.955 ;
        RECT 313.315 -177.645 313.645 -177.315 ;
        RECT 313.315 -179.005 313.645 -178.675 ;
        RECT 313.315 -180.365 313.645 -180.035 ;
        RECT 313.315 -181.725 313.645 -181.395 ;
        RECT 313.315 -183.085 313.645 -182.755 ;
        RECT 313.315 -184.445 313.645 -184.115 ;
        RECT 313.315 -185.805 313.645 -185.475 ;
        RECT 313.315 -187.165 313.645 -186.835 ;
        RECT 313.315 -188.525 313.645 -188.195 ;
        RECT 313.315 -189.885 313.645 -189.555 ;
        RECT 313.315 -191.245 313.645 -190.915 ;
        RECT 313.315 -192.605 313.645 -192.275 ;
        RECT 313.315 -193.965 313.645 -193.635 ;
        RECT 313.315 -195.325 313.645 -194.995 ;
        RECT 313.315 -196.685 313.645 -196.355 ;
        RECT 313.315 -198.045 313.645 -197.715 ;
        RECT 313.315 -199.405 313.645 -199.075 ;
        RECT 313.315 -200.765 313.645 -200.435 ;
        RECT 313.315 -202.125 313.645 -201.795 ;
        RECT 313.315 -203.485 313.645 -203.155 ;
        RECT 313.315 -204.845 313.645 -204.515 ;
        RECT 313.315 -206.205 313.645 -205.875 ;
        RECT 313.315 -207.565 313.645 -207.235 ;
        RECT 313.315 -208.925 313.645 -208.595 ;
        RECT 313.315 -210.285 313.645 -209.955 ;
        RECT 313.315 -211.645 313.645 -211.315 ;
        RECT 313.315 -213.005 313.645 -212.675 ;
        RECT 313.315 -214.365 313.645 -214.035 ;
        RECT 313.315 -215.725 313.645 -215.395 ;
        RECT 313.315 -217.085 313.645 -216.755 ;
        RECT 313.315 -218.445 313.645 -218.115 ;
        RECT 313.315 -219.805 313.645 -219.475 ;
        RECT 313.315 -221.165 313.645 -220.835 ;
        RECT 313.315 -222.525 313.645 -222.195 ;
        RECT 313.315 -223.885 313.645 -223.555 ;
        RECT 313.315 -225.245 313.645 -224.915 ;
        RECT 313.315 -226.605 313.645 -226.275 ;
        RECT 313.315 -227.965 313.645 -227.635 ;
        RECT 313.315 -229.325 313.645 -228.995 ;
        RECT 313.315 -230.685 313.645 -230.355 ;
        RECT 313.315 -232.045 313.645 -231.715 ;
        RECT 313.315 -233.405 313.645 -233.075 ;
        RECT 313.315 -234.765 313.645 -234.435 ;
        RECT 313.315 -236.125 313.645 -235.795 ;
        RECT 313.315 -237.485 313.645 -237.155 ;
        RECT 313.315 -238.845 313.645 -238.515 ;
        RECT 313.315 -241.09 313.645 -239.96 ;
        RECT 313.32 -241.205 313.64 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 244.04 315.005 245.17 ;
        RECT 314.675 242.595 315.005 242.925 ;
        RECT 314.675 241.235 315.005 241.565 ;
        RECT 314.675 239.875 315.005 240.205 ;
        RECT 314.675 238.515 315.005 238.845 ;
        RECT 314.675 237.155 315.005 237.485 ;
        RECT 314.68 237.155 315 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 -0.845 315.005 -0.515 ;
        RECT 314.675 -2.205 315.005 -1.875 ;
        RECT 314.675 -3.565 315.005 -3.235 ;
        RECT 314.68 -3.565 315 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 -123.245 315.005 -122.915 ;
        RECT 314.675 -124.605 315.005 -124.275 ;
        RECT 314.675 -125.965 315.005 -125.635 ;
        RECT 314.675 -127.325 315.005 -126.995 ;
        RECT 314.675 -128.685 315.005 -128.355 ;
        RECT 314.675 -130.045 315.005 -129.715 ;
        RECT 314.675 -131.405 315.005 -131.075 ;
        RECT 314.675 -132.765 315.005 -132.435 ;
        RECT 314.675 -134.125 315.005 -133.795 ;
        RECT 314.675 -135.485 315.005 -135.155 ;
        RECT 314.675 -136.845 315.005 -136.515 ;
        RECT 314.675 -138.205 315.005 -137.875 ;
        RECT 314.675 -139.565 315.005 -139.235 ;
        RECT 314.675 -140.925 315.005 -140.595 ;
        RECT 314.675 -142.285 315.005 -141.955 ;
        RECT 314.675 -143.645 315.005 -143.315 ;
        RECT 314.675 -145.005 315.005 -144.675 ;
        RECT 314.675 -146.365 315.005 -146.035 ;
        RECT 314.675 -147.725 315.005 -147.395 ;
        RECT 314.675 -149.085 315.005 -148.755 ;
        RECT 314.675 -150.445 315.005 -150.115 ;
        RECT 314.675 -151.805 315.005 -151.475 ;
        RECT 314.675 -153.165 315.005 -152.835 ;
        RECT 314.675 -154.525 315.005 -154.195 ;
        RECT 314.675 -155.885 315.005 -155.555 ;
        RECT 314.675 -157.245 315.005 -156.915 ;
        RECT 314.675 -158.605 315.005 -158.275 ;
        RECT 314.675 -159.965 315.005 -159.635 ;
        RECT 314.675 -161.325 315.005 -160.995 ;
        RECT 314.675 -162.685 315.005 -162.355 ;
        RECT 314.675 -164.045 315.005 -163.715 ;
        RECT 314.675 -165.405 315.005 -165.075 ;
        RECT 314.675 -166.765 315.005 -166.435 ;
        RECT 314.675 -168.125 315.005 -167.795 ;
        RECT 314.675 -169.485 315.005 -169.155 ;
        RECT 314.675 -170.845 315.005 -170.515 ;
        RECT 314.675 -172.205 315.005 -171.875 ;
        RECT 314.675 -173.565 315.005 -173.235 ;
        RECT 314.675 -174.925 315.005 -174.595 ;
        RECT 314.675 -176.285 315.005 -175.955 ;
        RECT 314.675 -177.645 315.005 -177.315 ;
        RECT 314.675 -179.005 315.005 -178.675 ;
        RECT 314.675 -180.365 315.005 -180.035 ;
        RECT 314.675 -181.725 315.005 -181.395 ;
        RECT 314.675 -183.085 315.005 -182.755 ;
        RECT 314.675 -184.445 315.005 -184.115 ;
        RECT 314.675 -185.805 315.005 -185.475 ;
        RECT 314.675 -187.165 315.005 -186.835 ;
        RECT 314.675 -188.525 315.005 -188.195 ;
        RECT 314.675 -189.885 315.005 -189.555 ;
        RECT 314.675 -191.245 315.005 -190.915 ;
        RECT 314.675 -192.605 315.005 -192.275 ;
        RECT 314.675 -193.965 315.005 -193.635 ;
        RECT 314.675 -195.325 315.005 -194.995 ;
        RECT 314.675 -196.685 315.005 -196.355 ;
        RECT 314.675 -198.045 315.005 -197.715 ;
        RECT 314.675 -199.405 315.005 -199.075 ;
        RECT 314.675 -200.765 315.005 -200.435 ;
        RECT 314.675 -202.125 315.005 -201.795 ;
        RECT 314.675 -203.485 315.005 -203.155 ;
        RECT 314.675 -204.845 315.005 -204.515 ;
        RECT 314.675 -206.205 315.005 -205.875 ;
        RECT 314.675 -207.565 315.005 -207.235 ;
        RECT 314.675 -208.925 315.005 -208.595 ;
        RECT 314.675 -210.285 315.005 -209.955 ;
        RECT 314.675 -211.645 315.005 -211.315 ;
        RECT 314.675 -213.005 315.005 -212.675 ;
        RECT 314.675 -214.365 315.005 -214.035 ;
        RECT 314.675 -215.725 315.005 -215.395 ;
        RECT 314.675 -217.085 315.005 -216.755 ;
        RECT 314.675 -218.445 315.005 -218.115 ;
        RECT 314.675 -219.805 315.005 -219.475 ;
        RECT 314.675 -221.165 315.005 -220.835 ;
        RECT 314.675 -222.525 315.005 -222.195 ;
        RECT 314.675 -223.885 315.005 -223.555 ;
        RECT 314.675 -225.245 315.005 -224.915 ;
        RECT 314.675 -226.605 315.005 -226.275 ;
        RECT 314.675 -227.965 315.005 -227.635 ;
        RECT 314.675 -229.325 315.005 -228.995 ;
        RECT 314.675 -230.685 315.005 -230.355 ;
        RECT 314.675 -232.045 315.005 -231.715 ;
        RECT 314.675 -233.405 315.005 -233.075 ;
        RECT 314.675 -234.765 315.005 -234.435 ;
        RECT 314.675 -236.125 315.005 -235.795 ;
        RECT 314.675 -237.485 315.005 -237.155 ;
        RECT 314.675 -238.845 315.005 -238.515 ;
        RECT 314.675 -241.09 315.005 -239.96 ;
        RECT 314.68 -241.205 315 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 244.04 316.365 245.17 ;
        RECT 316.035 242.595 316.365 242.925 ;
        RECT 316.035 241.235 316.365 241.565 ;
        RECT 316.035 239.875 316.365 240.205 ;
        RECT 316.035 238.515 316.365 238.845 ;
        RECT 316.035 237.155 316.365 237.485 ;
        RECT 316.04 237.155 316.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 -0.845 316.365 -0.515 ;
        RECT 316.035 -2.205 316.365 -1.875 ;
        RECT 316.035 -3.565 316.365 -3.235 ;
        RECT 316.04 -3.565 316.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 -123.245 316.365 -122.915 ;
        RECT 316.035 -124.605 316.365 -124.275 ;
        RECT 316.035 -125.965 316.365 -125.635 ;
        RECT 316.035 -127.325 316.365 -126.995 ;
        RECT 316.035 -128.685 316.365 -128.355 ;
        RECT 316.035 -130.045 316.365 -129.715 ;
        RECT 316.035 -131.405 316.365 -131.075 ;
        RECT 316.035 -132.765 316.365 -132.435 ;
        RECT 316.035 -134.125 316.365 -133.795 ;
        RECT 316.035 -135.485 316.365 -135.155 ;
        RECT 316.035 -136.845 316.365 -136.515 ;
        RECT 316.035 -138.205 316.365 -137.875 ;
        RECT 316.035 -139.565 316.365 -139.235 ;
        RECT 316.035 -140.925 316.365 -140.595 ;
        RECT 316.035 -142.285 316.365 -141.955 ;
        RECT 316.035 -143.645 316.365 -143.315 ;
        RECT 316.035 -145.005 316.365 -144.675 ;
        RECT 316.035 -146.365 316.365 -146.035 ;
        RECT 316.035 -147.725 316.365 -147.395 ;
        RECT 316.035 -149.085 316.365 -148.755 ;
        RECT 316.035 -150.445 316.365 -150.115 ;
        RECT 316.035 -151.805 316.365 -151.475 ;
        RECT 316.035 -153.165 316.365 -152.835 ;
        RECT 316.035 -154.525 316.365 -154.195 ;
        RECT 316.035 -155.885 316.365 -155.555 ;
        RECT 316.035 -157.245 316.365 -156.915 ;
        RECT 316.035 -158.605 316.365 -158.275 ;
        RECT 316.035 -159.965 316.365 -159.635 ;
        RECT 316.035 -161.325 316.365 -160.995 ;
        RECT 316.035 -162.685 316.365 -162.355 ;
        RECT 316.035 -164.045 316.365 -163.715 ;
        RECT 316.035 -165.405 316.365 -165.075 ;
        RECT 316.035 -166.765 316.365 -166.435 ;
        RECT 316.035 -168.125 316.365 -167.795 ;
        RECT 316.035 -169.485 316.365 -169.155 ;
        RECT 316.035 -170.845 316.365 -170.515 ;
        RECT 316.035 -172.205 316.365 -171.875 ;
        RECT 316.035 -173.565 316.365 -173.235 ;
        RECT 316.035 -174.925 316.365 -174.595 ;
        RECT 316.035 -176.285 316.365 -175.955 ;
        RECT 316.035 -177.645 316.365 -177.315 ;
        RECT 316.035 -179.005 316.365 -178.675 ;
        RECT 316.035 -180.365 316.365 -180.035 ;
        RECT 316.035 -181.725 316.365 -181.395 ;
        RECT 316.035 -183.085 316.365 -182.755 ;
        RECT 316.035 -184.445 316.365 -184.115 ;
        RECT 316.035 -185.805 316.365 -185.475 ;
        RECT 316.035 -187.165 316.365 -186.835 ;
        RECT 316.035 -188.525 316.365 -188.195 ;
        RECT 316.035 -189.885 316.365 -189.555 ;
        RECT 316.035 -191.245 316.365 -190.915 ;
        RECT 316.035 -192.605 316.365 -192.275 ;
        RECT 316.035 -193.965 316.365 -193.635 ;
        RECT 316.035 -195.325 316.365 -194.995 ;
        RECT 316.035 -196.685 316.365 -196.355 ;
        RECT 316.035 -198.045 316.365 -197.715 ;
        RECT 316.035 -199.405 316.365 -199.075 ;
        RECT 316.035 -200.765 316.365 -200.435 ;
        RECT 316.035 -202.125 316.365 -201.795 ;
        RECT 316.035 -203.485 316.365 -203.155 ;
        RECT 316.035 -204.845 316.365 -204.515 ;
        RECT 316.035 -206.205 316.365 -205.875 ;
        RECT 316.035 -207.565 316.365 -207.235 ;
        RECT 316.035 -208.925 316.365 -208.595 ;
        RECT 316.035 -210.285 316.365 -209.955 ;
        RECT 316.035 -211.645 316.365 -211.315 ;
        RECT 316.035 -213.005 316.365 -212.675 ;
        RECT 316.035 -214.365 316.365 -214.035 ;
        RECT 316.035 -215.725 316.365 -215.395 ;
        RECT 316.035 -217.085 316.365 -216.755 ;
        RECT 316.035 -218.445 316.365 -218.115 ;
        RECT 316.035 -219.805 316.365 -219.475 ;
        RECT 316.035 -221.165 316.365 -220.835 ;
        RECT 316.035 -222.525 316.365 -222.195 ;
        RECT 316.035 -223.885 316.365 -223.555 ;
        RECT 316.035 -225.245 316.365 -224.915 ;
        RECT 316.035 -226.605 316.365 -226.275 ;
        RECT 316.035 -227.965 316.365 -227.635 ;
        RECT 316.035 -229.325 316.365 -228.995 ;
        RECT 316.035 -230.685 316.365 -230.355 ;
        RECT 316.035 -232.045 316.365 -231.715 ;
        RECT 316.035 -233.405 316.365 -233.075 ;
        RECT 316.035 -234.765 316.365 -234.435 ;
        RECT 316.035 -236.125 316.365 -235.795 ;
        RECT 316.035 -237.485 316.365 -237.155 ;
        RECT 316.035 -238.845 316.365 -238.515 ;
        RECT 316.035 -241.09 316.365 -239.96 ;
        RECT 316.04 -241.205 316.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 244.04 317.725 245.17 ;
        RECT 317.395 242.595 317.725 242.925 ;
        RECT 317.395 241.235 317.725 241.565 ;
        RECT 317.395 239.875 317.725 240.205 ;
        RECT 317.395 238.515 317.725 238.845 ;
        RECT 317.395 237.155 317.725 237.485 ;
        RECT 317.4 237.155 317.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 -0.845 317.725 -0.515 ;
        RECT 317.395 -2.205 317.725 -1.875 ;
        RECT 317.395 -3.565 317.725 -3.235 ;
        RECT 317.4 -3.565 317.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 -123.245 317.725 -122.915 ;
        RECT 317.395 -124.605 317.725 -124.275 ;
        RECT 317.395 -125.965 317.725 -125.635 ;
        RECT 317.395 -127.325 317.725 -126.995 ;
        RECT 317.395 -128.685 317.725 -128.355 ;
        RECT 317.395 -130.045 317.725 -129.715 ;
        RECT 317.395 -131.405 317.725 -131.075 ;
        RECT 317.395 -132.765 317.725 -132.435 ;
        RECT 317.395 -134.125 317.725 -133.795 ;
        RECT 317.395 -135.485 317.725 -135.155 ;
        RECT 317.395 -136.845 317.725 -136.515 ;
        RECT 317.395 -138.205 317.725 -137.875 ;
        RECT 317.395 -139.565 317.725 -139.235 ;
        RECT 317.395 -140.925 317.725 -140.595 ;
        RECT 317.395 -142.285 317.725 -141.955 ;
        RECT 317.395 -143.645 317.725 -143.315 ;
        RECT 317.395 -145.005 317.725 -144.675 ;
        RECT 317.395 -146.365 317.725 -146.035 ;
        RECT 317.395 -147.725 317.725 -147.395 ;
        RECT 317.395 -149.085 317.725 -148.755 ;
        RECT 317.395 -150.445 317.725 -150.115 ;
        RECT 317.395 -151.805 317.725 -151.475 ;
        RECT 317.395 -153.165 317.725 -152.835 ;
        RECT 317.395 -154.525 317.725 -154.195 ;
        RECT 317.395 -155.885 317.725 -155.555 ;
        RECT 317.395 -157.245 317.725 -156.915 ;
        RECT 317.395 -158.605 317.725 -158.275 ;
        RECT 317.395 -159.965 317.725 -159.635 ;
        RECT 317.395 -161.325 317.725 -160.995 ;
        RECT 317.395 -162.685 317.725 -162.355 ;
        RECT 317.395 -164.045 317.725 -163.715 ;
        RECT 317.395 -165.405 317.725 -165.075 ;
        RECT 317.395 -166.765 317.725 -166.435 ;
        RECT 317.395 -168.125 317.725 -167.795 ;
        RECT 317.395 -169.485 317.725 -169.155 ;
        RECT 317.395 -170.845 317.725 -170.515 ;
        RECT 317.395 -172.205 317.725 -171.875 ;
        RECT 317.395 -173.565 317.725 -173.235 ;
        RECT 317.395 -174.925 317.725 -174.595 ;
        RECT 317.395 -176.285 317.725 -175.955 ;
        RECT 317.395 -177.645 317.725 -177.315 ;
        RECT 317.395 -179.005 317.725 -178.675 ;
        RECT 317.395 -180.365 317.725 -180.035 ;
        RECT 317.395 -181.725 317.725 -181.395 ;
        RECT 317.395 -183.085 317.725 -182.755 ;
        RECT 317.395 -184.445 317.725 -184.115 ;
        RECT 317.395 -185.805 317.725 -185.475 ;
        RECT 317.395 -187.165 317.725 -186.835 ;
        RECT 317.395 -188.525 317.725 -188.195 ;
        RECT 317.395 -189.885 317.725 -189.555 ;
        RECT 317.395 -191.245 317.725 -190.915 ;
        RECT 317.395 -192.605 317.725 -192.275 ;
        RECT 317.395 -193.965 317.725 -193.635 ;
        RECT 317.395 -195.325 317.725 -194.995 ;
        RECT 317.395 -196.685 317.725 -196.355 ;
        RECT 317.395 -198.045 317.725 -197.715 ;
        RECT 317.395 -199.405 317.725 -199.075 ;
        RECT 317.395 -200.765 317.725 -200.435 ;
        RECT 317.395 -202.125 317.725 -201.795 ;
        RECT 317.395 -203.485 317.725 -203.155 ;
        RECT 317.395 -204.845 317.725 -204.515 ;
        RECT 317.395 -206.205 317.725 -205.875 ;
        RECT 317.395 -207.565 317.725 -207.235 ;
        RECT 317.395 -208.925 317.725 -208.595 ;
        RECT 317.395 -210.285 317.725 -209.955 ;
        RECT 317.395 -211.645 317.725 -211.315 ;
        RECT 317.395 -213.005 317.725 -212.675 ;
        RECT 317.395 -214.365 317.725 -214.035 ;
        RECT 317.395 -215.725 317.725 -215.395 ;
        RECT 317.395 -217.085 317.725 -216.755 ;
        RECT 317.395 -218.445 317.725 -218.115 ;
        RECT 317.395 -219.805 317.725 -219.475 ;
        RECT 317.395 -221.165 317.725 -220.835 ;
        RECT 317.395 -222.525 317.725 -222.195 ;
        RECT 317.395 -223.885 317.725 -223.555 ;
        RECT 317.395 -225.245 317.725 -224.915 ;
        RECT 317.395 -226.605 317.725 -226.275 ;
        RECT 317.395 -227.965 317.725 -227.635 ;
        RECT 317.395 -229.325 317.725 -228.995 ;
        RECT 317.395 -230.685 317.725 -230.355 ;
        RECT 317.395 -232.045 317.725 -231.715 ;
        RECT 317.395 -233.405 317.725 -233.075 ;
        RECT 317.395 -234.765 317.725 -234.435 ;
        RECT 317.395 -236.125 317.725 -235.795 ;
        RECT 317.395 -237.485 317.725 -237.155 ;
        RECT 317.395 -238.845 317.725 -238.515 ;
        RECT 317.395 -241.09 317.725 -239.96 ;
        RECT 317.4 -241.205 317.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 244.04 319.085 245.17 ;
        RECT 318.755 242.595 319.085 242.925 ;
        RECT 318.755 241.235 319.085 241.565 ;
        RECT 318.755 239.875 319.085 240.205 ;
        RECT 318.755 238.515 319.085 238.845 ;
        RECT 318.755 237.155 319.085 237.485 ;
        RECT 318.76 237.155 319.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 -127.325 319.085 -126.995 ;
        RECT 318.755 -128.685 319.085 -128.355 ;
        RECT 318.755 -130.045 319.085 -129.715 ;
        RECT 318.755 -131.405 319.085 -131.075 ;
        RECT 318.755 -132.765 319.085 -132.435 ;
        RECT 318.755 -134.125 319.085 -133.795 ;
        RECT 318.755 -135.485 319.085 -135.155 ;
        RECT 318.755 -136.845 319.085 -136.515 ;
        RECT 318.755 -138.205 319.085 -137.875 ;
        RECT 318.755 -139.565 319.085 -139.235 ;
        RECT 318.755 -140.925 319.085 -140.595 ;
        RECT 318.755 -142.285 319.085 -141.955 ;
        RECT 318.755 -143.645 319.085 -143.315 ;
        RECT 318.755 -145.005 319.085 -144.675 ;
        RECT 318.755 -146.365 319.085 -146.035 ;
        RECT 318.755 -147.725 319.085 -147.395 ;
        RECT 318.755 -149.085 319.085 -148.755 ;
        RECT 318.755 -150.445 319.085 -150.115 ;
        RECT 318.755 -151.805 319.085 -151.475 ;
        RECT 318.755 -153.165 319.085 -152.835 ;
        RECT 318.755 -154.525 319.085 -154.195 ;
        RECT 318.755 -155.885 319.085 -155.555 ;
        RECT 318.755 -157.245 319.085 -156.915 ;
        RECT 318.755 -158.605 319.085 -158.275 ;
        RECT 318.755 -159.965 319.085 -159.635 ;
        RECT 318.755 -161.325 319.085 -160.995 ;
        RECT 318.755 -162.685 319.085 -162.355 ;
        RECT 318.755 -164.045 319.085 -163.715 ;
        RECT 318.755 -165.405 319.085 -165.075 ;
        RECT 318.755 -166.765 319.085 -166.435 ;
        RECT 318.755 -168.125 319.085 -167.795 ;
        RECT 318.755 -169.485 319.085 -169.155 ;
        RECT 318.755 -170.845 319.085 -170.515 ;
        RECT 318.755 -172.205 319.085 -171.875 ;
        RECT 318.755 -173.565 319.085 -173.235 ;
        RECT 318.755 -174.925 319.085 -174.595 ;
        RECT 318.755 -176.285 319.085 -175.955 ;
        RECT 318.755 -177.645 319.085 -177.315 ;
        RECT 318.755 -179.005 319.085 -178.675 ;
        RECT 318.755 -180.365 319.085 -180.035 ;
        RECT 318.755 -181.725 319.085 -181.395 ;
        RECT 318.755 -183.085 319.085 -182.755 ;
        RECT 318.755 -184.445 319.085 -184.115 ;
        RECT 318.755 -185.805 319.085 -185.475 ;
        RECT 318.755 -187.165 319.085 -186.835 ;
        RECT 318.755 -188.525 319.085 -188.195 ;
        RECT 318.755 -189.885 319.085 -189.555 ;
        RECT 318.755 -191.245 319.085 -190.915 ;
        RECT 318.755 -192.605 319.085 -192.275 ;
        RECT 318.755 -193.965 319.085 -193.635 ;
        RECT 318.755 -195.325 319.085 -194.995 ;
        RECT 318.755 -196.685 319.085 -196.355 ;
        RECT 318.755 -198.045 319.085 -197.715 ;
        RECT 318.755 -199.405 319.085 -199.075 ;
        RECT 318.755 -200.765 319.085 -200.435 ;
        RECT 318.755 -202.125 319.085 -201.795 ;
        RECT 318.755 -203.485 319.085 -203.155 ;
        RECT 318.755 -204.845 319.085 -204.515 ;
        RECT 318.755 -206.205 319.085 -205.875 ;
        RECT 318.755 -207.565 319.085 -207.235 ;
        RECT 318.755 -208.925 319.085 -208.595 ;
        RECT 318.755 -210.285 319.085 -209.955 ;
        RECT 318.755 -211.645 319.085 -211.315 ;
        RECT 318.755 -213.005 319.085 -212.675 ;
        RECT 318.755 -214.365 319.085 -214.035 ;
        RECT 318.755 -215.725 319.085 -215.395 ;
        RECT 318.755 -217.085 319.085 -216.755 ;
        RECT 318.755 -218.445 319.085 -218.115 ;
        RECT 318.755 -219.805 319.085 -219.475 ;
        RECT 318.755 -221.165 319.085 -220.835 ;
        RECT 318.755 -222.525 319.085 -222.195 ;
        RECT 318.755 -223.885 319.085 -223.555 ;
        RECT 318.755 -225.245 319.085 -224.915 ;
        RECT 318.755 -226.605 319.085 -226.275 ;
        RECT 318.755 -227.965 319.085 -227.635 ;
        RECT 318.755 -229.325 319.085 -228.995 ;
        RECT 318.755 -230.685 319.085 -230.355 ;
        RECT 318.755 -232.045 319.085 -231.715 ;
        RECT 318.755 -233.405 319.085 -233.075 ;
        RECT 318.755 -234.765 319.085 -234.435 ;
        RECT 318.755 -236.125 319.085 -235.795 ;
        RECT 318.755 -237.485 319.085 -237.155 ;
        RECT 318.755 -238.845 319.085 -238.515 ;
        RECT 318.755 -241.09 319.085 -239.96 ;
        RECT 318.76 -241.205 319.08 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.41 -125.535 319.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 244.04 320.445 245.17 ;
        RECT 320.115 242.595 320.445 242.925 ;
        RECT 320.115 241.235 320.445 241.565 ;
        RECT 320.115 239.875 320.445 240.205 ;
        RECT 320.115 238.515 320.445 238.845 ;
        RECT 320.115 237.155 320.445 237.485 ;
        RECT 320.12 237.155 320.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 -0.845 320.445 -0.515 ;
        RECT 320.115 -2.205 320.445 -1.875 ;
        RECT 320.115 -3.565 320.445 -3.235 ;
        RECT 320.12 -3.565 320.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.475 244.04 321.805 245.17 ;
        RECT 321.475 242.595 321.805 242.925 ;
        RECT 321.475 241.235 321.805 241.565 ;
        RECT 321.475 239.875 321.805 240.205 ;
        RECT 321.475 238.515 321.805 238.845 ;
        RECT 321.475 237.155 321.805 237.485 ;
        RECT 321.48 237.155 321.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.475 -0.845 321.805 -0.515 ;
        RECT 321.475 -2.205 321.805 -1.875 ;
        RECT 321.475 -3.565 321.805 -3.235 ;
        RECT 321.48 -3.565 321.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 244.04 323.165 245.17 ;
        RECT 322.835 242.595 323.165 242.925 ;
        RECT 322.835 241.235 323.165 241.565 ;
        RECT 322.835 239.875 323.165 240.205 ;
        RECT 322.835 238.515 323.165 238.845 ;
        RECT 322.835 237.155 323.165 237.485 ;
        RECT 322.84 237.155 323.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 -0.845 323.165 -0.515 ;
        RECT 322.835 -2.205 323.165 -1.875 ;
        RECT 322.835 -3.565 323.165 -3.235 ;
        RECT 322.84 -3.565 323.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 -123.245 323.165 -122.915 ;
        RECT 322.835 -124.605 323.165 -124.275 ;
        RECT 322.835 -125.965 323.165 -125.635 ;
        RECT 322.835 -127.325 323.165 -126.995 ;
        RECT 322.835 -128.685 323.165 -128.355 ;
        RECT 322.835 -130.045 323.165 -129.715 ;
        RECT 322.835 -131.405 323.165 -131.075 ;
        RECT 322.835 -132.765 323.165 -132.435 ;
        RECT 322.835 -134.125 323.165 -133.795 ;
        RECT 322.835 -135.485 323.165 -135.155 ;
        RECT 322.835 -136.845 323.165 -136.515 ;
        RECT 322.835 -138.205 323.165 -137.875 ;
        RECT 322.835 -139.565 323.165 -139.235 ;
        RECT 322.835 -140.925 323.165 -140.595 ;
        RECT 322.835 -142.285 323.165 -141.955 ;
        RECT 322.835 -143.645 323.165 -143.315 ;
        RECT 322.835 -145.005 323.165 -144.675 ;
        RECT 322.835 -146.365 323.165 -146.035 ;
        RECT 322.835 -147.725 323.165 -147.395 ;
        RECT 322.835 -149.085 323.165 -148.755 ;
        RECT 322.835 -150.445 323.165 -150.115 ;
        RECT 322.835 -151.805 323.165 -151.475 ;
        RECT 322.835 -153.165 323.165 -152.835 ;
        RECT 322.835 -154.525 323.165 -154.195 ;
        RECT 322.835 -155.885 323.165 -155.555 ;
        RECT 322.835 -157.245 323.165 -156.915 ;
        RECT 322.835 -158.605 323.165 -158.275 ;
        RECT 322.835 -159.965 323.165 -159.635 ;
        RECT 322.835 -161.325 323.165 -160.995 ;
        RECT 322.835 -162.685 323.165 -162.355 ;
        RECT 322.835 -164.045 323.165 -163.715 ;
        RECT 322.835 -165.405 323.165 -165.075 ;
        RECT 322.835 -166.765 323.165 -166.435 ;
        RECT 322.835 -168.125 323.165 -167.795 ;
        RECT 322.835 -169.485 323.165 -169.155 ;
        RECT 322.835 -170.845 323.165 -170.515 ;
        RECT 322.835 -172.205 323.165 -171.875 ;
        RECT 322.835 -173.565 323.165 -173.235 ;
        RECT 322.835 -174.925 323.165 -174.595 ;
        RECT 322.835 -176.285 323.165 -175.955 ;
        RECT 322.835 -177.645 323.165 -177.315 ;
        RECT 322.835 -179.005 323.165 -178.675 ;
        RECT 322.835 -180.365 323.165 -180.035 ;
        RECT 322.835 -181.725 323.165 -181.395 ;
        RECT 322.835 -183.085 323.165 -182.755 ;
        RECT 322.835 -184.445 323.165 -184.115 ;
        RECT 322.835 -185.805 323.165 -185.475 ;
        RECT 322.835 -187.165 323.165 -186.835 ;
        RECT 322.835 -188.525 323.165 -188.195 ;
        RECT 322.835 -189.885 323.165 -189.555 ;
        RECT 322.835 -191.245 323.165 -190.915 ;
        RECT 322.835 -192.605 323.165 -192.275 ;
        RECT 322.835 -193.965 323.165 -193.635 ;
        RECT 322.835 -195.325 323.165 -194.995 ;
        RECT 322.835 -196.685 323.165 -196.355 ;
        RECT 322.835 -198.045 323.165 -197.715 ;
        RECT 322.835 -199.405 323.165 -199.075 ;
        RECT 322.835 -200.765 323.165 -200.435 ;
        RECT 322.835 -202.125 323.165 -201.795 ;
        RECT 322.835 -203.485 323.165 -203.155 ;
        RECT 322.835 -204.845 323.165 -204.515 ;
        RECT 322.835 -206.205 323.165 -205.875 ;
        RECT 322.835 -207.565 323.165 -207.235 ;
        RECT 322.835 -208.925 323.165 -208.595 ;
        RECT 322.835 -210.285 323.165 -209.955 ;
        RECT 322.835 -211.645 323.165 -211.315 ;
        RECT 322.835 -213.005 323.165 -212.675 ;
        RECT 322.835 -214.365 323.165 -214.035 ;
        RECT 322.835 -215.725 323.165 -215.395 ;
        RECT 322.835 -217.085 323.165 -216.755 ;
        RECT 322.835 -218.445 323.165 -218.115 ;
        RECT 322.835 -219.805 323.165 -219.475 ;
        RECT 322.835 -221.165 323.165 -220.835 ;
        RECT 322.835 -222.525 323.165 -222.195 ;
        RECT 322.835 -223.885 323.165 -223.555 ;
        RECT 322.835 -225.245 323.165 -224.915 ;
        RECT 322.835 -226.605 323.165 -226.275 ;
        RECT 322.835 -227.965 323.165 -227.635 ;
        RECT 322.835 -229.325 323.165 -228.995 ;
        RECT 322.835 -230.685 323.165 -230.355 ;
        RECT 322.835 -232.045 323.165 -231.715 ;
        RECT 322.835 -233.405 323.165 -233.075 ;
        RECT 322.835 -234.765 323.165 -234.435 ;
        RECT 322.835 -236.125 323.165 -235.795 ;
        RECT 322.835 -237.485 323.165 -237.155 ;
        RECT 322.835 -238.845 323.165 -238.515 ;
        RECT 322.835 -241.09 323.165 -239.96 ;
        RECT 322.84 -241.205 323.16 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 244.04 324.525 245.17 ;
        RECT 324.195 242.595 324.525 242.925 ;
        RECT 324.195 241.235 324.525 241.565 ;
        RECT 324.195 239.875 324.525 240.205 ;
        RECT 324.195 238.515 324.525 238.845 ;
        RECT 324.195 237.155 324.525 237.485 ;
        RECT 324.2 237.155 324.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 -0.845 324.525 -0.515 ;
        RECT 324.195 -2.205 324.525 -1.875 ;
        RECT 324.195 -3.565 324.525 -3.235 ;
        RECT 324.2 -3.565 324.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 -123.245 324.525 -122.915 ;
        RECT 324.195 -124.605 324.525 -124.275 ;
        RECT 324.195 -125.965 324.525 -125.635 ;
        RECT 324.195 -127.325 324.525 -126.995 ;
        RECT 324.195 -128.685 324.525 -128.355 ;
        RECT 324.195 -130.045 324.525 -129.715 ;
        RECT 324.195 -131.405 324.525 -131.075 ;
        RECT 324.195 -132.765 324.525 -132.435 ;
        RECT 324.195 -134.125 324.525 -133.795 ;
        RECT 324.195 -135.485 324.525 -135.155 ;
        RECT 324.195 -136.845 324.525 -136.515 ;
        RECT 324.195 -138.205 324.525 -137.875 ;
        RECT 324.195 -139.565 324.525 -139.235 ;
        RECT 324.195 -140.925 324.525 -140.595 ;
        RECT 324.195 -142.285 324.525 -141.955 ;
        RECT 324.195 -143.645 324.525 -143.315 ;
        RECT 324.195 -145.005 324.525 -144.675 ;
        RECT 324.195 -146.365 324.525 -146.035 ;
        RECT 324.195 -147.725 324.525 -147.395 ;
        RECT 324.195 -149.085 324.525 -148.755 ;
        RECT 324.195 -150.445 324.525 -150.115 ;
        RECT 324.195 -151.805 324.525 -151.475 ;
        RECT 324.195 -153.165 324.525 -152.835 ;
        RECT 324.195 -154.525 324.525 -154.195 ;
        RECT 324.195 -155.885 324.525 -155.555 ;
        RECT 324.195 -157.245 324.525 -156.915 ;
        RECT 324.195 -158.605 324.525 -158.275 ;
        RECT 324.195 -159.965 324.525 -159.635 ;
        RECT 324.195 -161.325 324.525 -160.995 ;
        RECT 324.195 -162.685 324.525 -162.355 ;
        RECT 324.195 -164.045 324.525 -163.715 ;
        RECT 324.195 -165.405 324.525 -165.075 ;
        RECT 324.195 -166.765 324.525 -166.435 ;
        RECT 324.195 -168.125 324.525 -167.795 ;
        RECT 324.195 -169.485 324.525 -169.155 ;
        RECT 324.195 -170.845 324.525 -170.515 ;
        RECT 324.195 -172.205 324.525 -171.875 ;
        RECT 324.195 -173.565 324.525 -173.235 ;
        RECT 324.195 -174.925 324.525 -174.595 ;
        RECT 324.195 -176.285 324.525 -175.955 ;
        RECT 324.195 -177.645 324.525 -177.315 ;
        RECT 324.195 -179.005 324.525 -178.675 ;
        RECT 324.195 -180.365 324.525 -180.035 ;
        RECT 324.195 -181.725 324.525 -181.395 ;
        RECT 324.195 -183.085 324.525 -182.755 ;
        RECT 324.195 -184.445 324.525 -184.115 ;
        RECT 324.195 -185.805 324.525 -185.475 ;
        RECT 324.195 -187.165 324.525 -186.835 ;
        RECT 324.195 -188.525 324.525 -188.195 ;
        RECT 324.195 -189.885 324.525 -189.555 ;
        RECT 324.195 -191.245 324.525 -190.915 ;
        RECT 324.195 -192.605 324.525 -192.275 ;
        RECT 324.195 -193.965 324.525 -193.635 ;
        RECT 324.195 -195.325 324.525 -194.995 ;
        RECT 324.195 -196.685 324.525 -196.355 ;
        RECT 324.195 -198.045 324.525 -197.715 ;
        RECT 324.195 -199.405 324.525 -199.075 ;
        RECT 324.195 -200.765 324.525 -200.435 ;
        RECT 324.195 -202.125 324.525 -201.795 ;
        RECT 324.195 -203.485 324.525 -203.155 ;
        RECT 324.195 -204.845 324.525 -204.515 ;
        RECT 324.195 -206.205 324.525 -205.875 ;
        RECT 324.195 -207.565 324.525 -207.235 ;
        RECT 324.195 -208.925 324.525 -208.595 ;
        RECT 324.195 -210.285 324.525 -209.955 ;
        RECT 324.195 -211.645 324.525 -211.315 ;
        RECT 324.195 -213.005 324.525 -212.675 ;
        RECT 324.195 -214.365 324.525 -214.035 ;
        RECT 324.195 -215.725 324.525 -215.395 ;
        RECT 324.195 -217.085 324.525 -216.755 ;
        RECT 324.195 -218.445 324.525 -218.115 ;
        RECT 324.195 -219.805 324.525 -219.475 ;
        RECT 324.195 -221.165 324.525 -220.835 ;
        RECT 324.195 -222.525 324.525 -222.195 ;
        RECT 324.195 -223.885 324.525 -223.555 ;
        RECT 324.195 -225.245 324.525 -224.915 ;
        RECT 324.195 -226.605 324.525 -226.275 ;
        RECT 324.195 -227.965 324.525 -227.635 ;
        RECT 324.195 -229.325 324.525 -228.995 ;
        RECT 324.195 -230.685 324.525 -230.355 ;
        RECT 324.195 -232.045 324.525 -231.715 ;
        RECT 324.195 -233.405 324.525 -233.075 ;
        RECT 324.195 -234.765 324.525 -234.435 ;
        RECT 324.195 -236.125 324.525 -235.795 ;
        RECT 324.195 -237.485 324.525 -237.155 ;
        RECT 324.195 -238.845 324.525 -238.515 ;
        RECT 324.195 -241.09 324.525 -239.96 ;
        RECT 324.2 -241.205 324.52 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 244.04 325.885 245.17 ;
        RECT 325.555 242.595 325.885 242.925 ;
        RECT 325.555 241.235 325.885 241.565 ;
        RECT 325.555 239.875 325.885 240.205 ;
        RECT 325.555 238.515 325.885 238.845 ;
        RECT 325.555 237.155 325.885 237.485 ;
        RECT 325.56 237.155 325.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 -0.845 325.885 -0.515 ;
        RECT 325.555 -2.205 325.885 -1.875 ;
        RECT 325.555 -3.565 325.885 -3.235 ;
        RECT 325.56 -3.565 325.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 -218.445 325.885 -218.115 ;
        RECT 325.555 -219.805 325.885 -219.475 ;
        RECT 325.555 -221.165 325.885 -220.835 ;
        RECT 325.555 -222.525 325.885 -222.195 ;
        RECT 325.555 -223.885 325.885 -223.555 ;
        RECT 325.555 -225.245 325.885 -224.915 ;
        RECT 325.555 -226.605 325.885 -226.275 ;
        RECT 325.555 -227.965 325.885 -227.635 ;
        RECT 325.555 -229.325 325.885 -228.995 ;
        RECT 325.555 -230.685 325.885 -230.355 ;
        RECT 325.555 -232.045 325.885 -231.715 ;
        RECT 325.555 -233.405 325.885 -233.075 ;
        RECT 325.555 -234.765 325.885 -234.435 ;
        RECT 325.555 -236.125 325.885 -235.795 ;
        RECT 325.555 -237.485 325.885 -237.155 ;
        RECT 325.555 -238.845 325.885 -238.515 ;
        RECT 325.555 -241.09 325.885 -239.96 ;
        RECT 325.56 -241.205 325.88 -122.24 ;
        RECT 325.555 -123.245 325.885 -122.915 ;
        RECT 325.555 -124.605 325.885 -124.275 ;
        RECT 325.555 -125.965 325.885 -125.635 ;
        RECT 325.555 -127.325 325.885 -126.995 ;
        RECT 325.555 -128.685 325.885 -128.355 ;
        RECT 325.555 -130.045 325.885 -129.715 ;
        RECT 325.555 -131.405 325.885 -131.075 ;
        RECT 325.555 -132.765 325.885 -132.435 ;
        RECT 325.555 -134.125 325.885 -133.795 ;
        RECT 325.555 -135.485 325.885 -135.155 ;
        RECT 325.555 -136.845 325.885 -136.515 ;
        RECT 325.555 -138.205 325.885 -137.875 ;
        RECT 325.555 -139.565 325.885 -139.235 ;
        RECT 325.555 -140.925 325.885 -140.595 ;
        RECT 325.555 -142.285 325.885 -141.955 ;
        RECT 325.555 -143.645 325.885 -143.315 ;
        RECT 325.555 -145.005 325.885 -144.675 ;
        RECT 325.555 -146.365 325.885 -146.035 ;
        RECT 325.555 -147.725 325.885 -147.395 ;
        RECT 325.555 -149.085 325.885 -148.755 ;
        RECT 325.555 -150.445 325.885 -150.115 ;
        RECT 325.555 -151.805 325.885 -151.475 ;
        RECT 325.555 -153.165 325.885 -152.835 ;
        RECT 325.555 -154.525 325.885 -154.195 ;
        RECT 325.555 -155.885 325.885 -155.555 ;
        RECT 325.555 -157.245 325.885 -156.915 ;
        RECT 325.555 -158.605 325.885 -158.275 ;
        RECT 325.555 -159.965 325.885 -159.635 ;
        RECT 325.555 -161.325 325.885 -160.995 ;
        RECT 325.555 -162.685 325.885 -162.355 ;
        RECT 325.555 -164.045 325.885 -163.715 ;
        RECT 325.555 -165.405 325.885 -165.075 ;
        RECT 325.555 -166.765 325.885 -166.435 ;
        RECT 325.555 -168.125 325.885 -167.795 ;
        RECT 325.555 -169.485 325.885 -169.155 ;
        RECT 325.555 -170.845 325.885 -170.515 ;
        RECT 325.555 -172.205 325.885 -171.875 ;
        RECT 325.555 -173.565 325.885 -173.235 ;
        RECT 325.555 -174.925 325.885 -174.595 ;
        RECT 325.555 -176.285 325.885 -175.955 ;
        RECT 325.555 -177.645 325.885 -177.315 ;
        RECT 325.555 -179.005 325.885 -178.675 ;
        RECT 325.555 -180.365 325.885 -180.035 ;
        RECT 325.555 -181.725 325.885 -181.395 ;
        RECT 325.555 -183.085 325.885 -182.755 ;
        RECT 325.555 -184.445 325.885 -184.115 ;
        RECT 325.555 -185.805 325.885 -185.475 ;
        RECT 325.555 -187.165 325.885 -186.835 ;
        RECT 325.555 -188.525 325.885 -188.195 ;
        RECT 325.555 -189.885 325.885 -189.555 ;
        RECT 325.555 -191.245 325.885 -190.915 ;
        RECT 325.555 -192.605 325.885 -192.275 ;
        RECT 325.555 -193.965 325.885 -193.635 ;
        RECT 325.555 -195.325 325.885 -194.995 ;
        RECT 325.555 -196.685 325.885 -196.355 ;
        RECT 325.555 -198.045 325.885 -197.715 ;
        RECT 325.555 -199.405 325.885 -199.075 ;
        RECT 325.555 -200.765 325.885 -200.435 ;
        RECT 325.555 -202.125 325.885 -201.795 ;
        RECT 325.555 -203.485 325.885 -203.155 ;
        RECT 325.555 -204.845 325.885 -204.515 ;
        RECT 325.555 -206.205 325.885 -205.875 ;
        RECT 325.555 -207.565 325.885 -207.235 ;
        RECT 325.555 -208.925 325.885 -208.595 ;
        RECT 325.555 -210.285 325.885 -209.955 ;
        RECT 325.555 -211.645 325.885 -211.315 ;
        RECT 325.555 -213.005 325.885 -212.675 ;
        RECT 325.555 -214.365 325.885 -214.035 ;
        RECT 325.555 -215.725 325.885 -215.395 ;
        RECT 325.555 -217.085 325.885 -216.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 244.04 291.885 245.17 ;
        RECT 291.555 242.595 291.885 242.925 ;
        RECT 291.555 241.235 291.885 241.565 ;
        RECT 291.555 239.875 291.885 240.205 ;
        RECT 291.555 238.515 291.885 238.845 ;
        RECT 291.555 237.155 291.885 237.485 ;
        RECT 291.56 237.155 291.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 -0.845 291.885 -0.515 ;
        RECT 291.555 -2.205 291.885 -1.875 ;
        RECT 291.555 -3.565 291.885 -3.235 ;
        RECT 291.56 -3.565 291.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 -123.245 291.885 -122.915 ;
        RECT 291.555 -124.605 291.885 -124.275 ;
        RECT 291.555 -125.965 291.885 -125.635 ;
        RECT 291.555 -127.325 291.885 -126.995 ;
        RECT 291.555 -128.685 291.885 -128.355 ;
        RECT 291.555 -130.045 291.885 -129.715 ;
        RECT 291.555 -131.405 291.885 -131.075 ;
        RECT 291.555 -132.765 291.885 -132.435 ;
        RECT 291.555 -134.125 291.885 -133.795 ;
        RECT 291.555 -135.485 291.885 -135.155 ;
        RECT 291.555 -136.845 291.885 -136.515 ;
        RECT 291.555 -138.205 291.885 -137.875 ;
        RECT 291.555 -139.565 291.885 -139.235 ;
        RECT 291.555 -140.925 291.885 -140.595 ;
        RECT 291.555 -142.285 291.885 -141.955 ;
        RECT 291.555 -143.645 291.885 -143.315 ;
        RECT 291.555 -145.005 291.885 -144.675 ;
        RECT 291.555 -146.365 291.885 -146.035 ;
        RECT 291.555 -147.725 291.885 -147.395 ;
        RECT 291.555 -149.085 291.885 -148.755 ;
        RECT 291.555 -150.445 291.885 -150.115 ;
        RECT 291.555 -151.805 291.885 -151.475 ;
        RECT 291.555 -153.165 291.885 -152.835 ;
        RECT 291.555 -154.525 291.885 -154.195 ;
        RECT 291.555 -155.885 291.885 -155.555 ;
        RECT 291.555 -157.245 291.885 -156.915 ;
        RECT 291.555 -158.605 291.885 -158.275 ;
        RECT 291.555 -159.965 291.885 -159.635 ;
        RECT 291.555 -161.325 291.885 -160.995 ;
        RECT 291.555 -162.685 291.885 -162.355 ;
        RECT 291.555 -164.045 291.885 -163.715 ;
        RECT 291.555 -165.405 291.885 -165.075 ;
        RECT 291.555 -166.765 291.885 -166.435 ;
        RECT 291.555 -168.125 291.885 -167.795 ;
        RECT 291.555 -169.485 291.885 -169.155 ;
        RECT 291.555 -170.845 291.885 -170.515 ;
        RECT 291.555 -172.205 291.885 -171.875 ;
        RECT 291.555 -173.565 291.885 -173.235 ;
        RECT 291.555 -174.925 291.885 -174.595 ;
        RECT 291.555 -176.285 291.885 -175.955 ;
        RECT 291.555 -177.645 291.885 -177.315 ;
        RECT 291.555 -179.005 291.885 -178.675 ;
        RECT 291.555 -180.365 291.885 -180.035 ;
        RECT 291.555 -181.725 291.885 -181.395 ;
        RECT 291.555 -183.085 291.885 -182.755 ;
        RECT 291.555 -184.445 291.885 -184.115 ;
        RECT 291.555 -185.805 291.885 -185.475 ;
        RECT 291.555 -187.165 291.885 -186.835 ;
        RECT 291.555 -188.525 291.885 -188.195 ;
        RECT 291.555 -189.885 291.885 -189.555 ;
        RECT 291.555 -191.245 291.885 -190.915 ;
        RECT 291.555 -192.605 291.885 -192.275 ;
        RECT 291.555 -193.965 291.885 -193.635 ;
        RECT 291.555 -195.325 291.885 -194.995 ;
        RECT 291.555 -196.685 291.885 -196.355 ;
        RECT 291.555 -198.045 291.885 -197.715 ;
        RECT 291.555 -199.405 291.885 -199.075 ;
        RECT 291.555 -200.765 291.885 -200.435 ;
        RECT 291.555 -202.125 291.885 -201.795 ;
        RECT 291.555 -203.485 291.885 -203.155 ;
        RECT 291.555 -204.845 291.885 -204.515 ;
        RECT 291.555 -206.205 291.885 -205.875 ;
        RECT 291.555 -207.565 291.885 -207.235 ;
        RECT 291.555 -208.925 291.885 -208.595 ;
        RECT 291.555 -210.285 291.885 -209.955 ;
        RECT 291.555 -211.645 291.885 -211.315 ;
        RECT 291.555 -213.005 291.885 -212.675 ;
        RECT 291.555 -214.365 291.885 -214.035 ;
        RECT 291.555 -215.725 291.885 -215.395 ;
        RECT 291.555 -217.085 291.885 -216.755 ;
        RECT 291.555 -218.445 291.885 -218.115 ;
        RECT 291.555 -219.805 291.885 -219.475 ;
        RECT 291.555 -221.165 291.885 -220.835 ;
        RECT 291.555 -222.525 291.885 -222.195 ;
        RECT 291.555 -223.885 291.885 -223.555 ;
        RECT 291.555 -225.245 291.885 -224.915 ;
        RECT 291.555 -226.605 291.885 -226.275 ;
        RECT 291.555 -227.965 291.885 -227.635 ;
        RECT 291.555 -229.325 291.885 -228.995 ;
        RECT 291.555 -230.685 291.885 -230.355 ;
        RECT 291.555 -232.045 291.885 -231.715 ;
        RECT 291.555 -233.405 291.885 -233.075 ;
        RECT 291.555 -234.765 291.885 -234.435 ;
        RECT 291.555 -236.125 291.885 -235.795 ;
        RECT 291.555 -237.485 291.885 -237.155 ;
        RECT 291.555 -238.845 291.885 -238.515 ;
        RECT 291.555 -241.09 291.885 -239.96 ;
        RECT 291.56 -241.205 291.88 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 244.04 293.245 245.17 ;
        RECT 292.915 242.595 293.245 242.925 ;
        RECT 292.915 241.235 293.245 241.565 ;
        RECT 292.915 239.875 293.245 240.205 ;
        RECT 292.915 238.515 293.245 238.845 ;
        RECT 292.915 237.155 293.245 237.485 ;
        RECT 292.92 237.155 293.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 -0.845 293.245 -0.515 ;
        RECT 292.915 -2.205 293.245 -1.875 ;
        RECT 292.915 -3.565 293.245 -3.235 ;
        RECT 292.92 -3.565 293.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 -123.245 293.245 -122.915 ;
        RECT 292.915 -124.605 293.245 -124.275 ;
        RECT 292.915 -125.965 293.245 -125.635 ;
        RECT 292.915 -127.325 293.245 -126.995 ;
        RECT 292.915 -128.685 293.245 -128.355 ;
        RECT 292.915 -130.045 293.245 -129.715 ;
        RECT 292.915 -131.405 293.245 -131.075 ;
        RECT 292.915 -132.765 293.245 -132.435 ;
        RECT 292.915 -134.125 293.245 -133.795 ;
        RECT 292.915 -135.485 293.245 -135.155 ;
        RECT 292.915 -136.845 293.245 -136.515 ;
        RECT 292.915 -138.205 293.245 -137.875 ;
        RECT 292.915 -139.565 293.245 -139.235 ;
        RECT 292.915 -140.925 293.245 -140.595 ;
        RECT 292.915 -142.285 293.245 -141.955 ;
        RECT 292.915 -143.645 293.245 -143.315 ;
        RECT 292.915 -145.005 293.245 -144.675 ;
        RECT 292.915 -146.365 293.245 -146.035 ;
        RECT 292.915 -147.725 293.245 -147.395 ;
        RECT 292.915 -149.085 293.245 -148.755 ;
        RECT 292.915 -150.445 293.245 -150.115 ;
        RECT 292.915 -151.805 293.245 -151.475 ;
        RECT 292.915 -153.165 293.245 -152.835 ;
        RECT 292.915 -154.525 293.245 -154.195 ;
        RECT 292.915 -155.885 293.245 -155.555 ;
        RECT 292.915 -157.245 293.245 -156.915 ;
        RECT 292.915 -158.605 293.245 -158.275 ;
        RECT 292.915 -159.965 293.245 -159.635 ;
        RECT 292.915 -161.325 293.245 -160.995 ;
        RECT 292.915 -162.685 293.245 -162.355 ;
        RECT 292.915 -164.045 293.245 -163.715 ;
        RECT 292.915 -165.405 293.245 -165.075 ;
        RECT 292.915 -166.765 293.245 -166.435 ;
        RECT 292.915 -168.125 293.245 -167.795 ;
        RECT 292.915 -169.485 293.245 -169.155 ;
        RECT 292.915 -170.845 293.245 -170.515 ;
        RECT 292.915 -172.205 293.245 -171.875 ;
        RECT 292.915 -173.565 293.245 -173.235 ;
        RECT 292.915 -174.925 293.245 -174.595 ;
        RECT 292.915 -176.285 293.245 -175.955 ;
        RECT 292.915 -177.645 293.245 -177.315 ;
        RECT 292.915 -179.005 293.245 -178.675 ;
        RECT 292.915 -180.365 293.245 -180.035 ;
        RECT 292.915 -181.725 293.245 -181.395 ;
        RECT 292.915 -183.085 293.245 -182.755 ;
        RECT 292.915 -184.445 293.245 -184.115 ;
        RECT 292.915 -185.805 293.245 -185.475 ;
        RECT 292.915 -187.165 293.245 -186.835 ;
        RECT 292.915 -188.525 293.245 -188.195 ;
        RECT 292.915 -189.885 293.245 -189.555 ;
        RECT 292.915 -191.245 293.245 -190.915 ;
        RECT 292.915 -192.605 293.245 -192.275 ;
        RECT 292.915 -193.965 293.245 -193.635 ;
        RECT 292.915 -195.325 293.245 -194.995 ;
        RECT 292.915 -196.685 293.245 -196.355 ;
        RECT 292.915 -198.045 293.245 -197.715 ;
        RECT 292.915 -199.405 293.245 -199.075 ;
        RECT 292.915 -200.765 293.245 -200.435 ;
        RECT 292.915 -202.125 293.245 -201.795 ;
        RECT 292.915 -203.485 293.245 -203.155 ;
        RECT 292.915 -204.845 293.245 -204.515 ;
        RECT 292.915 -206.205 293.245 -205.875 ;
        RECT 292.915 -207.565 293.245 -207.235 ;
        RECT 292.915 -208.925 293.245 -208.595 ;
        RECT 292.915 -210.285 293.245 -209.955 ;
        RECT 292.915 -211.645 293.245 -211.315 ;
        RECT 292.915 -213.005 293.245 -212.675 ;
        RECT 292.915 -214.365 293.245 -214.035 ;
        RECT 292.915 -215.725 293.245 -215.395 ;
        RECT 292.915 -217.085 293.245 -216.755 ;
        RECT 292.915 -218.445 293.245 -218.115 ;
        RECT 292.915 -219.805 293.245 -219.475 ;
        RECT 292.915 -221.165 293.245 -220.835 ;
        RECT 292.915 -222.525 293.245 -222.195 ;
        RECT 292.915 -223.885 293.245 -223.555 ;
        RECT 292.915 -225.245 293.245 -224.915 ;
        RECT 292.915 -226.605 293.245 -226.275 ;
        RECT 292.915 -227.965 293.245 -227.635 ;
        RECT 292.915 -229.325 293.245 -228.995 ;
        RECT 292.915 -230.685 293.245 -230.355 ;
        RECT 292.915 -232.045 293.245 -231.715 ;
        RECT 292.915 -233.405 293.245 -233.075 ;
        RECT 292.915 -234.765 293.245 -234.435 ;
        RECT 292.915 -236.125 293.245 -235.795 ;
        RECT 292.915 -237.485 293.245 -237.155 ;
        RECT 292.915 -238.845 293.245 -238.515 ;
        RECT 292.915 -241.09 293.245 -239.96 ;
        RECT 292.92 -241.205 293.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 244.04 294.605 245.17 ;
        RECT 294.275 242.595 294.605 242.925 ;
        RECT 294.275 241.235 294.605 241.565 ;
        RECT 294.275 239.875 294.605 240.205 ;
        RECT 294.275 238.515 294.605 238.845 ;
        RECT 294.275 237.155 294.605 237.485 ;
        RECT 294.28 237.155 294.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 -0.845 294.605 -0.515 ;
        RECT 294.275 -2.205 294.605 -1.875 ;
        RECT 294.275 -3.565 294.605 -3.235 ;
        RECT 294.28 -3.565 294.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 -123.245 294.605 -122.915 ;
        RECT 294.275 -124.605 294.605 -124.275 ;
        RECT 294.275 -125.965 294.605 -125.635 ;
        RECT 294.275 -127.325 294.605 -126.995 ;
        RECT 294.275 -128.685 294.605 -128.355 ;
        RECT 294.275 -130.045 294.605 -129.715 ;
        RECT 294.275 -131.405 294.605 -131.075 ;
        RECT 294.275 -132.765 294.605 -132.435 ;
        RECT 294.275 -134.125 294.605 -133.795 ;
        RECT 294.275 -135.485 294.605 -135.155 ;
        RECT 294.275 -136.845 294.605 -136.515 ;
        RECT 294.275 -138.205 294.605 -137.875 ;
        RECT 294.275 -139.565 294.605 -139.235 ;
        RECT 294.275 -140.925 294.605 -140.595 ;
        RECT 294.275 -142.285 294.605 -141.955 ;
        RECT 294.275 -143.645 294.605 -143.315 ;
        RECT 294.275 -145.005 294.605 -144.675 ;
        RECT 294.275 -146.365 294.605 -146.035 ;
        RECT 294.275 -147.725 294.605 -147.395 ;
        RECT 294.275 -149.085 294.605 -148.755 ;
        RECT 294.275 -150.445 294.605 -150.115 ;
        RECT 294.275 -151.805 294.605 -151.475 ;
        RECT 294.275 -153.165 294.605 -152.835 ;
        RECT 294.275 -154.525 294.605 -154.195 ;
        RECT 294.275 -155.885 294.605 -155.555 ;
        RECT 294.275 -157.245 294.605 -156.915 ;
        RECT 294.275 -158.605 294.605 -158.275 ;
        RECT 294.275 -159.965 294.605 -159.635 ;
        RECT 294.275 -161.325 294.605 -160.995 ;
        RECT 294.275 -162.685 294.605 -162.355 ;
        RECT 294.275 -164.045 294.605 -163.715 ;
        RECT 294.275 -165.405 294.605 -165.075 ;
        RECT 294.275 -166.765 294.605 -166.435 ;
        RECT 294.275 -168.125 294.605 -167.795 ;
        RECT 294.275 -169.485 294.605 -169.155 ;
        RECT 294.275 -170.845 294.605 -170.515 ;
        RECT 294.275 -172.205 294.605 -171.875 ;
        RECT 294.275 -173.565 294.605 -173.235 ;
        RECT 294.275 -174.925 294.605 -174.595 ;
        RECT 294.275 -176.285 294.605 -175.955 ;
        RECT 294.275 -177.645 294.605 -177.315 ;
        RECT 294.275 -179.005 294.605 -178.675 ;
        RECT 294.275 -180.365 294.605 -180.035 ;
        RECT 294.275 -181.725 294.605 -181.395 ;
        RECT 294.275 -183.085 294.605 -182.755 ;
        RECT 294.275 -184.445 294.605 -184.115 ;
        RECT 294.275 -185.805 294.605 -185.475 ;
        RECT 294.275 -187.165 294.605 -186.835 ;
        RECT 294.275 -188.525 294.605 -188.195 ;
        RECT 294.275 -189.885 294.605 -189.555 ;
        RECT 294.275 -191.245 294.605 -190.915 ;
        RECT 294.275 -192.605 294.605 -192.275 ;
        RECT 294.275 -193.965 294.605 -193.635 ;
        RECT 294.275 -195.325 294.605 -194.995 ;
        RECT 294.275 -196.685 294.605 -196.355 ;
        RECT 294.275 -198.045 294.605 -197.715 ;
        RECT 294.275 -199.405 294.605 -199.075 ;
        RECT 294.275 -200.765 294.605 -200.435 ;
        RECT 294.275 -202.125 294.605 -201.795 ;
        RECT 294.275 -203.485 294.605 -203.155 ;
        RECT 294.275 -204.845 294.605 -204.515 ;
        RECT 294.275 -206.205 294.605 -205.875 ;
        RECT 294.275 -207.565 294.605 -207.235 ;
        RECT 294.275 -208.925 294.605 -208.595 ;
        RECT 294.275 -210.285 294.605 -209.955 ;
        RECT 294.275 -211.645 294.605 -211.315 ;
        RECT 294.275 -213.005 294.605 -212.675 ;
        RECT 294.275 -214.365 294.605 -214.035 ;
        RECT 294.275 -215.725 294.605 -215.395 ;
        RECT 294.275 -217.085 294.605 -216.755 ;
        RECT 294.275 -218.445 294.605 -218.115 ;
        RECT 294.275 -219.805 294.605 -219.475 ;
        RECT 294.275 -221.165 294.605 -220.835 ;
        RECT 294.275 -222.525 294.605 -222.195 ;
        RECT 294.275 -223.885 294.605 -223.555 ;
        RECT 294.275 -225.245 294.605 -224.915 ;
        RECT 294.275 -226.605 294.605 -226.275 ;
        RECT 294.275 -227.965 294.605 -227.635 ;
        RECT 294.275 -229.325 294.605 -228.995 ;
        RECT 294.275 -230.685 294.605 -230.355 ;
        RECT 294.275 -232.045 294.605 -231.715 ;
        RECT 294.275 -233.405 294.605 -233.075 ;
        RECT 294.275 -234.765 294.605 -234.435 ;
        RECT 294.275 -236.125 294.605 -235.795 ;
        RECT 294.275 -237.485 294.605 -237.155 ;
        RECT 294.275 -238.845 294.605 -238.515 ;
        RECT 294.275 -241.09 294.605 -239.96 ;
        RECT 294.28 -241.205 294.6 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 244.04 295.965 245.17 ;
        RECT 295.635 242.595 295.965 242.925 ;
        RECT 295.635 241.235 295.965 241.565 ;
        RECT 295.635 239.875 295.965 240.205 ;
        RECT 295.635 238.515 295.965 238.845 ;
        RECT 295.635 237.155 295.965 237.485 ;
        RECT 295.64 237.155 295.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 -0.845 295.965 -0.515 ;
        RECT 295.635 -2.205 295.965 -1.875 ;
        RECT 295.635 -3.565 295.965 -3.235 ;
        RECT 295.64 -3.565 295.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 -123.245 295.965 -122.915 ;
        RECT 295.635 -124.605 295.965 -124.275 ;
        RECT 295.635 -125.965 295.965 -125.635 ;
        RECT 295.635 -127.325 295.965 -126.995 ;
        RECT 295.635 -128.685 295.965 -128.355 ;
        RECT 295.635 -130.045 295.965 -129.715 ;
        RECT 295.635 -131.405 295.965 -131.075 ;
        RECT 295.635 -132.765 295.965 -132.435 ;
        RECT 295.635 -134.125 295.965 -133.795 ;
        RECT 295.635 -135.485 295.965 -135.155 ;
        RECT 295.635 -136.845 295.965 -136.515 ;
        RECT 295.635 -138.205 295.965 -137.875 ;
        RECT 295.635 -139.565 295.965 -139.235 ;
        RECT 295.635 -140.925 295.965 -140.595 ;
        RECT 295.635 -142.285 295.965 -141.955 ;
        RECT 295.635 -143.645 295.965 -143.315 ;
        RECT 295.635 -145.005 295.965 -144.675 ;
        RECT 295.635 -146.365 295.965 -146.035 ;
        RECT 295.635 -147.725 295.965 -147.395 ;
        RECT 295.635 -149.085 295.965 -148.755 ;
        RECT 295.635 -150.445 295.965 -150.115 ;
        RECT 295.635 -151.805 295.965 -151.475 ;
        RECT 295.635 -153.165 295.965 -152.835 ;
        RECT 295.635 -154.525 295.965 -154.195 ;
        RECT 295.635 -155.885 295.965 -155.555 ;
        RECT 295.635 -157.245 295.965 -156.915 ;
        RECT 295.635 -158.605 295.965 -158.275 ;
        RECT 295.635 -159.965 295.965 -159.635 ;
        RECT 295.635 -161.325 295.965 -160.995 ;
        RECT 295.635 -162.685 295.965 -162.355 ;
        RECT 295.635 -164.045 295.965 -163.715 ;
        RECT 295.635 -165.405 295.965 -165.075 ;
        RECT 295.635 -166.765 295.965 -166.435 ;
        RECT 295.635 -168.125 295.965 -167.795 ;
        RECT 295.635 -169.485 295.965 -169.155 ;
        RECT 295.635 -170.845 295.965 -170.515 ;
        RECT 295.635 -172.205 295.965 -171.875 ;
        RECT 295.635 -173.565 295.965 -173.235 ;
        RECT 295.635 -174.925 295.965 -174.595 ;
        RECT 295.635 -176.285 295.965 -175.955 ;
        RECT 295.635 -177.645 295.965 -177.315 ;
        RECT 295.635 -179.005 295.965 -178.675 ;
        RECT 295.635 -180.365 295.965 -180.035 ;
        RECT 295.635 -181.725 295.965 -181.395 ;
        RECT 295.635 -183.085 295.965 -182.755 ;
        RECT 295.635 -184.445 295.965 -184.115 ;
        RECT 295.635 -185.805 295.965 -185.475 ;
        RECT 295.635 -187.165 295.965 -186.835 ;
        RECT 295.635 -188.525 295.965 -188.195 ;
        RECT 295.635 -189.885 295.965 -189.555 ;
        RECT 295.635 -191.245 295.965 -190.915 ;
        RECT 295.635 -192.605 295.965 -192.275 ;
        RECT 295.635 -193.965 295.965 -193.635 ;
        RECT 295.635 -195.325 295.965 -194.995 ;
        RECT 295.635 -196.685 295.965 -196.355 ;
        RECT 295.635 -198.045 295.965 -197.715 ;
        RECT 295.635 -199.405 295.965 -199.075 ;
        RECT 295.635 -200.765 295.965 -200.435 ;
        RECT 295.635 -202.125 295.965 -201.795 ;
        RECT 295.635 -203.485 295.965 -203.155 ;
        RECT 295.635 -204.845 295.965 -204.515 ;
        RECT 295.635 -206.205 295.965 -205.875 ;
        RECT 295.635 -207.565 295.965 -207.235 ;
        RECT 295.635 -208.925 295.965 -208.595 ;
        RECT 295.635 -210.285 295.965 -209.955 ;
        RECT 295.635 -211.645 295.965 -211.315 ;
        RECT 295.635 -213.005 295.965 -212.675 ;
        RECT 295.635 -214.365 295.965 -214.035 ;
        RECT 295.635 -215.725 295.965 -215.395 ;
        RECT 295.635 -217.085 295.965 -216.755 ;
        RECT 295.635 -218.445 295.965 -218.115 ;
        RECT 295.635 -219.805 295.965 -219.475 ;
        RECT 295.635 -221.165 295.965 -220.835 ;
        RECT 295.635 -222.525 295.965 -222.195 ;
        RECT 295.635 -223.885 295.965 -223.555 ;
        RECT 295.635 -225.245 295.965 -224.915 ;
        RECT 295.635 -226.605 295.965 -226.275 ;
        RECT 295.635 -227.965 295.965 -227.635 ;
        RECT 295.635 -229.325 295.965 -228.995 ;
        RECT 295.635 -230.685 295.965 -230.355 ;
        RECT 295.635 -232.045 295.965 -231.715 ;
        RECT 295.635 -233.405 295.965 -233.075 ;
        RECT 295.635 -234.765 295.965 -234.435 ;
        RECT 295.635 -236.125 295.965 -235.795 ;
        RECT 295.635 -237.485 295.965 -237.155 ;
        RECT 295.635 -238.845 295.965 -238.515 ;
        RECT 295.635 -241.09 295.965 -239.96 ;
        RECT 295.64 -241.205 295.96 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 244.04 297.325 245.17 ;
        RECT 296.995 242.595 297.325 242.925 ;
        RECT 296.995 241.235 297.325 241.565 ;
        RECT 296.995 239.875 297.325 240.205 ;
        RECT 296.995 238.515 297.325 238.845 ;
        RECT 296.995 237.155 297.325 237.485 ;
        RECT 297 237.155 297.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 -127.325 297.325 -126.995 ;
        RECT 296.995 -128.685 297.325 -128.355 ;
        RECT 296.995 -130.045 297.325 -129.715 ;
        RECT 296.995 -131.405 297.325 -131.075 ;
        RECT 296.995 -132.765 297.325 -132.435 ;
        RECT 296.995 -134.125 297.325 -133.795 ;
        RECT 296.995 -135.485 297.325 -135.155 ;
        RECT 296.995 -136.845 297.325 -136.515 ;
        RECT 296.995 -138.205 297.325 -137.875 ;
        RECT 296.995 -139.565 297.325 -139.235 ;
        RECT 296.995 -140.925 297.325 -140.595 ;
        RECT 296.995 -142.285 297.325 -141.955 ;
        RECT 296.995 -143.645 297.325 -143.315 ;
        RECT 296.995 -145.005 297.325 -144.675 ;
        RECT 296.995 -146.365 297.325 -146.035 ;
        RECT 296.995 -147.725 297.325 -147.395 ;
        RECT 296.995 -149.085 297.325 -148.755 ;
        RECT 296.995 -150.445 297.325 -150.115 ;
        RECT 296.995 -151.805 297.325 -151.475 ;
        RECT 296.995 -153.165 297.325 -152.835 ;
        RECT 296.995 -154.525 297.325 -154.195 ;
        RECT 296.995 -155.885 297.325 -155.555 ;
        RECT 296.995 -157.245 297.325 -156.915 ;
        RECT 296.995 -158.605 297.325 -158.275 ;
        RECT 296.995 -159.965 297.325 -159.635 ;
        RECT 296.995 -161.325 297.325 -160.995 ;
        RECT 296.995 -162.685 297.325 -162.355 ;
        RECT 296.995 -164.045 297.325 -163.715 ;
        RECT 296.995 -165.405 297.325 -165.075 ;
        RECT 296.995 -166.765 297.325 -166.435 ;
        RECT 296.995 -168.125 297.325 -167.795 ;
        RECT 296.995 -169.485 297.325 -169.155 ;
        RECT 296.995 -170.845 297.325 -170.515 ;
        RECT 296.995 -172.205 297.325 -171.875 ;
        RECT 296.995 -173.565 297.325 -173.235 ;
        RECT 296.995 -174.925 297.325 -174.595 ;
        RECT 296.995 -176.285 297.325 -175.955 ;
        RECT 296.995 -177.645 297.325 -177.315 ;
        RECT 296.995 -179.005 297.325 -178.675 ;
        RECT 296.995 -180.365 297.325 -180.035 ;
        RECT 296.995 -181.725 297.325 -181.395 ;
        RECT 296.995 -183.085 297.325 -182.755 ;
        RECT 296.995 -184.445 297.325 -184.115 ;
        RECT 296.995 -185.805 297.325 -185.475 ;
        RECT 296.995 -187.165 297.325 -186.835 ;
        RECT 296.995 -188.525 297.325 -188.195 ;
        RECT 296.995 -189.885 297.325 -189.555 ;
        RECT 296.995 -191.245 297.325 -190.915 ;
        RECT 296.995 -192.605 297.325 -192.275 ;
        RECT 296.995 -193.965 297.325 -193.635 ;
        RECT 296.995 -195.325 297.325 -194.995 ;
        RECT 296.995 -196.685 297.325 -196.355 ;
        RECT 296.995 -198.045 297.325 -197.715 ;
        RECT 296.995 -199.405 297.325 -199.075 ;
        RECT 296.995 -200.765 297.325 -200.435 ;
        RECT 296.995 -202.125 297.325 -201.795 ;
        RECT 296.995 -203.485 297.325 -203.155 ;
        RECT 296.995 -204.845 297.325 -204.515 ;
        RECT 296.995 -206.205 297.325 -205.875 ;
        RECT 296.995 -207.565 297.325 -207.235 ;
        RECT 296.995 -208.925 297.325 -208.595 ;
        RECT 296.995 -210.285 297.325 -209.955 ;
        RECT 296.995 -211.645 297.325 -211.315 ;
        RECT 296.995 -213.005 297.325 -212.675 ;
        RECT 296.995 -214.365 297.325 -214.035 ;
        RECT 296.995 -215.725 297.325 -215.395 ;
        RECT 296.995 -217.085 297.325 -216.755 ;
        RECT 296.995 -218.445 297.325 -218.115 ;
        RECT 296.995 -219.805 297.325 -219.475 ;
        RECT 296.995 -221.165 297.325 -220.835 ;
        RECT 296.995 -222.525 297.325 -222.195 ;
        RECT 296.995 -223.885 297.325 -223.555 ;
        RECT 296.995 -225.245 297.325 -224.915 ;
        RECT 296.995 -226.605 297.325 -226.275 ;
        RECT 296.995 -227.965 297.325 -227.635 ;
        RECT 296.995 -229.325 297.325 -228.995 ;
        RECT 296.995 -230.685 297.325 -230.355 ;
        RECT 296.995 -232.045 297.325 -231.715 ;
        RECT 296.995 -233.405 297.325 -233.075 ;
        RECT 296.995 -234.765 297.325 -234.435 ;
        RECT 296.995 -236.125 297.325 -235.795 ;
        RECT 296.995 -237.485 297.325 -237.155 ;
        RECT 296.995 -238.845 297.325 -238.515 ;
        RECT 296.995 -241.09 297.325 -239.96 ;
        RECT 297 -241.205 297.32 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.61 -125.535 297.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 244.04 298.685 245.17 ;
        RECT 298.355 242.595 298.685 242.925 ;
        RECT 298.355 241.235 298.685 241.565 ;
        RECT 298.355 239.875 298.685 240.205 ;
        RECT 298.355 238.515 298.685 238.845 ;
        RECT 298.355 237.155 298.685 237.485 ;
        RECT 298.36 237.155 298.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 -0.845 298.685 -0.515 ;
        RECT 298.355 -2.205 298.685 -1.875 ;
        RECT 298.355 -3.565 298.685 -3.235 ;
        RECT 298.36 -3.565 298.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 244.04 300.045 245.17 ;
        RECT 299.715 242.595 300.045 242.925 ;
        RECT 299.715 241.235 300.045 241.565 ;
        RECT 299.715 239.875 300.045 240.205 ;
        RECT 299.715 238.515 300.045 238.845 ;
        RECT 299.715 237.155 300.045 237.485 ;
        RECT 299.72 237.155 300.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 -0.845 300.045 -0.515 ;
        RECT 299.715 -2.205 300.045 -1.875 ;
        RECT 299.715 -3.565 300.045 -3.235 ;
        RECT 299.72 -3.565 300.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 244.04 301.405 245.17 ;
        RECT 301.075 242.595 301.405 242.925 ;
        RECT 301.075 241.235 301.405 241.565 ;
        RECT 301.075 239.875 301.405 240.205 ;
        RECT 301.075 238.515 301.405 238.845 ;
        RECT 301.075 237.155 301.405 237.485 ;
        RECT 301.08 237.155 301.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 -0.845 301.405 -0.515 ;
        RECT 301.075 -2.205 301.405 -1.875 ;
        RECT 301.075 -3.565 301.405 -3.235 ;
        RECT 301.08 -3.565 301.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 -123.245 301.405 -122.915 ;
        RECT 301.075 -124.605 301.405 -124.275 ;
        RECT 301.075 -125.965 301.405 -125.635 ;
        RECT 301.075 -127.325 301.405 -126.995 ;
        RECT 301.075 -128.685 301.405 -128.355 ;
        RECT 301.075 -130.045 301.405 -129.715 ;
        RECT 301.075 -131.405 301.405 -131.075 ;
        RECT 301.075 -132.765 301.405 -132.435 ;
        RECT 301.075 -134.125 301.405 -133.795 ;
        RECT 301.075 -135.485 301.405 -135.155 ;
        RECT 301.075 -136.845 301.405 -136.515 ;
        RECT 301.075 -138.205 301.405 -137.875 ;
        RECT 301.075 -139.565 301.405 -139.235 ;
        RECT 301.075 -140.925 301.405 -140.595 ;
        RECT 301.075 -142.285 301.405 -141.955 ;
        RECT 301.075 -143.645 301.405 -143.315 ;
        RECT 301.075 -145.005 301.405 -144.675 ;
        RECT 301.075 -146.365 301.405 -146.035 ;
        RECT 301.075 -147.725 301.405 -147.395 ;
        RECT 301.075 -149.085 301.405 -148.755 ;
        RECT 301.075 -150.445 301.405 -150.115 ;
        RECT 301.075 -151.805 301.405 -151.475 ;
        RECT 301.075 -153.165 301.405 -152.835 ;
        RECT 301.075 -154.525 301.405 -154.195 ;
        RECT 301.075 -155.885 301.405 -155.555 ;
        RECT 301.075 -157.245 301.405 -156.915 ;
        RECT 301.075 -158.605 301.405 -158.275 ;
        RECT 301.075 -159.965 301.405 -159.635 ;
        RECT 301.075 -161.325 301.405 -160.995 ;
        RECT 301.075 -162.685 301.405 -162.355 ;
        RECT 301.075 -164.045 301.405 -163.715 ;
        RECT 301.075 -165.405 301.405 -165.075 ;
        RECT 301.075 -166.765 301.405 -166.435 ;
        RECT 301.075 -168.125 301.405 -167.795 ;
        RECT 301.075 -169.485 301.405 -169.155 ;
        RECT 301.075 -170.845 301.405 -170.515 ;
        RECT 301.075 -172.205 301.405 -171.875 ;
        RECT 301.075 -173.565 301.405 -173.235 ;
        RECT 301.075 -174.925 301.405 -174.595 ;
        RECT 301.075 -176.285 301.405 -175.955 ;
        RECT 301.075 -177.645 301.405 -177.315 ;
        RECT 301.075 -179.005 301.405 -178.675 ;
        RECT 301.075 -180.365 301.405 -180.035 ;
        RECT 301.075 -181.725 301.405 -181.395 ;
        RECT 301.075 -183.085 301.405 -182.755 ;
        RECT 301.075 -184.445 301.405 -184.115 ;
        RECT 301.075 -185.805 301.405 -185.475 ;
        RECT 301.075 -187.165 301.405 -186.835 ;
        RECT 301.075 -188.525 301.405 -188.195 ;
        RECT 301.075 -189.885 301.405 -189.555 ;
        RECT 301.075 -191.245 301.405 -190.915 ;
        RECT 301.075 -192.605 301.405 -192.275 ;
        RECT 301.075 -193.965 301.405 -193.635 ;
        RECT 301.075 -195.325 301.405 -194.995 ;
        RECT 301.075 -196.685 301.405 -196.355 ;
        RECT 301.075 -198.045 301.405 -197.715 ;
        RECT 301.075 -199.405 301.405 -199.075 ;
        RECT 301.075 -200.765 301.405 -200.435 ;
        RECT 301.075 -202.125 301.405 -201.795 ;
        RECT 301.075 -203.485 301.405 -203.155 ;
        RECT 301.075 -204.845 301.405 -204.515 ;
        RECT 301.075 -206.205 301.405 -205.875 ;
        RECT 301.075 -207.565 301.405 -207.235 ;
        RECT 301.075 -208.925 301.405 -208.595 ;
        RECT 301.075 -210.285 301.405 -209.955 ;
        RECT 301.075 -211.645 301.405 -211.315 ;
        RECT 301.075 -213.005 301.405 -212.675 ;
        RECT 301.075 -214.365 301.405 -214.035 ;
        RECT 301.075 -215.725 301.405 -215.395 ;
        RECT 301.075 -217.085 301.405 -216.755 ;
        RECT 301.075 -218.445 301.405 -218.115 ;
        RECT 301.075 -219.805 301.405 -219.475 ;
        RECT 301.075 -221.165 301.405 -220.835 ;
        RECT 301.075 -222.525 301.405 -222.195 ;
        RECT 301.075 -223.885 301.405 -223.555 ;
        RECT 301.075 -225.245 301.405 -224.915 ;
        RECT 301.075 -226.605 301.405 -226.275 ;
        RECT 301.075 -227.965 301.405 -227.635 ;
        RECT 301.075 -229.325 301.405 -228.995 ;
        RECT 301.075 -230.685 301.405 -230.355 ;
        RECT 301.075 -232.045 301.405 -231.715 ;
        RECT 301.075 -233.405 301.405 -233.075 ;
        RECT 301.075 -234.765 301.405 -234.435 ;
        RECT 301.075 -236.125 301.405 -235.795 ;
        RECT 301.075 -237.485 301.405 -237.155 ;
        RECT 301.075 -238.845 301.405 -238.515 ;
        RECT 301.075 -241.09 301.405 -239.96 ;
        RECT 301.08 -241.205 301.4 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 244.04 302.765 245.17 ;
        RECT 302.435 242.595 302.765 242.925 ;
        RECT 302.435 241.235 302.765 241.565 ;
        RECT 302.435 239.875 302.765 240.205 ;
        RECT 302.435 238.515 302.765 238.845 ;
        RECT 302.435 237.155 302.765 237.485 ;
        RECT 302.44 237.155 302.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 -0.845 302.765 -0.515 ;
        RECT 302.435 -2.205 302.765 -1.875 ;
        RECT 302.435 -3.565 302.765 -3.235 ;
        RECT 302.44 -3.565 302.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 -123.245 302.765 -122.915 ;
        RECT 302.435 -124.605 302.765 -124.275 ;
        RECT 302.435 -125.965 302.765 -125.635 ;
        RECT 302.435 -127.325 302.765 -126.995 ;
        RECT 302.435 -128.685 302.765 -128.355 ;
        RECT 302.435 -130.045 302.765 -129.715 ;
        RECT 302.435 -131.405 302.765 -131.075 ;
        RECT 302.435 -132.765 302.765 -132.435 ;
        RECT 302.435 -134.125 302.765 -133.795 ;
        RECT 302.435 -135.485 302.765 -135.155 ;
        RECT 302.435 -136.845 302.765 -136.515 ;
        RECT 302.435 -138.205 302.765 -137.875 ;
        RECT 302.435 -139.565 302.765 -139.235 ;
        RECT 302.435 -140.925 302.765 -140.595 ;
        RECT 302.435 -142.285 302.765 -141.955 ;
        RECT 302.435 -143.645 302.765 -143.315 ;
        RECT 302.435 -145.005 302.765 -144.675 ;
        RECT 302.435 -146.365 302.765 -146.035 ;
        RECT 302.435 -147.725 302.765 -147.395 ;
        RECT 302.435 -149.085 302.765 -148.755 ;
        RECT 302.435 -150.445 302.765 -150.115 ;
        RECT 302.435 -151.805 302.765 -151.475 ;
        RECT 302.435 -153.165 302.765 -152.835 ;
        RECT 302.435 -154.525 302.765 -154.195 ;
        RECT 302.435 -155.885 302.765 -155.555 ;
        RECT 302.435 -157.245 302.765 -156.915 ;
        RECT 302.435 -158.605 302.765 -158.275 ;
        RECT 302.435 -159.965 302.765 -159.635 ;
        RECT 302.435 -161.325 302.765 -160.995 ;
        RECT 302.435 -162.685 302.765 -162.355 ;
        RECT 302.435 -164.045 302.765 -163.715 ;
        RECT 302.435 -165.405 302.765 -165.075 ;
        RECT 302.435 -166.765 302.765 -166.435 ;
        RECT 302.435 -168.125 302.765 -167.795 ;
        RECT 302.435 -169.485 302.765 -169.155 ;
        RECT 302.435 -170.845 302.765 -170.515 ;
        RECT 302.435 -172.205 302.765 -171.875 ;
        RECT 302.435 -173.565 302.765 -173.235 ;
        RECT 302.435 -174.925 302.765 -174.595 ;
        RECT 302.435 -176.285 302.765 -175.955 ;
        RECT 302.435 -177.645 302.765 -177.315 ;
        RECT 302.435 -179.005 302.765 -178.675 ;
        RECT 302.435 -180.365 302.765 -180.035 ;
        RECT 302.435 -181.725 302.765 -181.395 ;
        RECT 302.435 -183.085 302.765 -182.755 ;
        RECT 302.435 -184.445 302.765 -184.115 ;
        RECT 302.435 -185.805 302.765 -185.475 ;
        RECT 302.435 -187.165 302.765 -186.835 ;
        RECT 302.435 -188.525 302.765 -188.195 ;
        RECT 302.435 -189.885 302.765 -189.555 ;
        RECT 302.435 -191.245 302.765 -190.915 ;
        RECT 302.435 -192.605 302.765 -192.275 ;
        RECT 302.435 -193.965 302.765 -193.635 ;
        RECT 302.435 -195.325 302.765 -194.995 ;
        RECT 302.435 -196.685 302.765 -196.355 ;
        RECT 302.435 -198.045 302.765 -197.715 ;
        RECT 302.435 -199.405 302.765 -199.075 ;
        RECT 302.435 -200.765 302.765 -200.435 ;
        RECT 302.435 -202.125 302.765 -201.795 ;
        RECT 302.435 -203.485 302.765 -203.155 ;
        RECT 302.435 -204.845 302.765 -204.515 ;
        RECT 302.435 -206.205 302.765 -205.875 ;
        RECT 302.435 -207.565 302.765 -207.235 ;
        RECT 302.435 -208.925 302.765 -208.595 ;
        RECT 302.435 -210.285 302.765 -209.955 ;
        RECT 302.435 -211.645 302.765 -211.315 ;
        RECT 302.435 -213.005 302.765 -212.675 ;
        RECT 302.435 -214.365 302.765 -214.035 ;
        RECT 302.435 -215.725 302.765 -215.395 ;
        RECT 302.435 -217.085 302.765 -216.755 ;
        RECT 302.435 -218.445 302.765 -218.115 ;
        RECT 302.435 -219.805 302.765 -219.475 ;
        RECT 302.435 -221.165 302.765 -220.835 ;
        RECT 302.435 -222.525 302.765 -222.195 ;
        RECT 302.435 -223.885 302.765 -223.555 ;
        RECT 302.435 -225.245 302.765 -224.915 ;
        RECT 302.435 -226.605 302.765 -226.275 ;
        RECT 302.435 -227.965 302.765 -227.635 ;
        RECT 302.435 -229.325 302.765 -228.995 ;
        RECT 302.435 -230.685 302.765 -230.355 ;
        RECT 302.435 -232.045 302.765 -231.715 ;
        RECT 302.435 -233.405 302.765 -233.075 ;
        RECT 302.435 -234.765 302.765 -234.435 ;
        RECT 302.435 -236.125 302.765 -235.795 ;
        RECT 302.435 -237.485 302.765 -237.155 ;
        RECT 302.435 -238.845 302.765 -238.515 ;
        RECT 302.435 -241.09 302.765 -239.96 ;
        RECT 302.44 -241.205 302.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 244.04 304.125 245.17 ;
        RECT 303.795 242.595 304.125 242.925 ;
        RECT 303.795 241.235 304.125 241.565 ;
        RECT 303.795 239.875 304.125 240.205 ;
        RECT 303.795 238.515 304.125 238.845 ;
        RECT 303.795 237.155 304.125 237.485 ;
        RECT 303.8 237.155 304.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 -0.845 304.125 -0.515 ;
        RECT 303.795 -2.205 304.125 -1.875 ;
        RECT 303.795 -3.565 304.125 -3.235 ;
        RECT 303.8 -3.565 304.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 -123.245 304.125 -122.915 ;
        RECT 303.795 -124.605 304.125 -124.275 ;
        RECT 303.795 -125.965 304.125 -125.635 ;
        RECT 303.795 -127.325 304.125 -126.995 ;
        RECT 303.795 -128.685 304.125 -128.355 ;
        RECT 303.795 -130.045 304.125 -129.715 ;
        RECT 303.795 -131.405 304.125 -131.075 ;
        RECT 303.795 -132.765 304.125 -132.435 ;
        RECT 303.795 -134.125 304.125 -133.795 ;
        RECT 303.795 -135.485 304.125 -135.155 ;
        RECT 303.795 -136.845 304.125 -136.515 ;
        RECT 303.795 -138.205 304.125 -137.875 ;
        RECT 303.795 -139.565 304.125 -139.235 ;
        RECT 303.795 -140.925 304.125 -140.595 ;
        RECT 303.795 -142.285 304.125 -141.955 ;
        RECT 303.795 -143.645 304.125 -143.315 ;
        RECT 303.795 -145.005 304.125 -144.675 ;
        RECT 303.795 -146.365 304.125 -146.035 ;
        RECT 303.795 -147.725 304.125 -147.395 ;
        RECT 303.795 -149.085 304.125 -148.755 ;
        RECT 303.795 -150.445 304.125 -150.115 ;
        RECT 303.795 -151.805 304.125 -151.475 ;
        RECT 303.795 -153.165 304.125 -152.835 ;
        RECT 303.795 -154.525 304.125 -154.195 ;
        RECT 303.795 -155.885 304.125 -155.555 ;
        RECT 303.795 -157.245 304.125 -156.915 ;
        RECT 303.795 -158.605 304.125 -158.275 ;
        RECT 303.795 -159.965 304.125 -159.635 ;
        RECT 303.795 -161.325 304.125 -160.995 ;
        RECT 303.795 -162.685 304.125 -162.355 ;
        RECT 303.795 -164.045 304.125 -163.715 ;
        RECT 303.795 -165.405 304.125 -165.075 ;
        RECT 303.795 -166.765 304.125 -166.435 ;
        RECT 303.795 -168.125 304.125 -167.795 ;
        RECT 303.795 -169.485 304.125 -169.155 ;
        RECT 303.795 -170.845 304.125 -170.515 ;
        RECT 303.795 -172.205 304.125 -171.875 ;
        RECT 303.795 -173.565 304.125 -173.235 ;
        RECT 303.795 -174.925 304.125 -174.595 ;
        RECT 303.795 -176.285 304.125 -175.955 ;
        RECT 303.795 -177.645 304.125 -177.315 ;
        RECT 303.795 -179.005 304.125 -178.675 ;
        RECT 303.795 -180.365 304.125 -180.035 ;
        RECT 303.795 -181.725 304.125 -181.395 ;
        RECT 303.795 -183.085 304.125 -182.755 ;
        RECT 303.795 -184.445 304.125 -184.115 ;
        RECT 303.795 -185.805 304.125 -185.475 ;
        RECT 303.795 -187.165 304.125 -186.835 ;
        RECT 303.795 -188.525 304.125 -188.195 ;
        RECT 303.795 -189.885 304.125 -189.555 ;
        RECT 303.795 -191.245 304.125 -190.915 ;
        RECT 303.795 -192.605 304.125 -192.275 ;
        RECT 303.795 -193.965 304.125 -193.635 ;
        RECT 303.795 -195.325 304.125 -194.995 ;
        RECT 303.795 -196.685 304.125 -196.355 ;
        RECT 303.795 -198.045 304.125 -197.715 ;
        RECT 303.795 -199.405 304.125 -199.075 ;
        RECT 303.795 -200.765 304.125 -200.435 ;
        RECT 303.795 -202.125 304.125 -201.795 ;
        RECT 303.795 -203.485 304.125 -203.155 ;
        RECT 303.795 -204.845 304.125 -204.515 ;
        RECT 303.795 -206.205 304.125 -205.875 ;
        RECT 303.795 -207.565 304.125 -207.235 ;
        RECT 303.795 -208.925 304.125 -208.595 ;
        RECT 303.795 -210.285 304.125 -209.955 ;
        RECT 303.795 -211.645 304.125 -211.315 ;
        RECT 303.795 -213.005 304.125 -212.675 ;
        RECT 303.795 -214.365 304.125 -214.035 ;
        RECT 303.795 -215.725 304.125 -215.395 ;
        RECT 303.795 -217.085 304.125 -216.755 ;
        RECT 303.795 -218.445 304.125 -218.115 ;
        RECT 303.795 -219.805 304.125 -219.475 ;
        RECT 303.795 -221.165 304.125 -220.835 ;
        RECT 303.795 -222.525 304.125 -222.195 ;
        RECT 303.795 -223.885 304.125 -223.555 ;
        RECT 303.795 -225.245 304.125 -224.915 ;
        RECT 303.795 -226.605 304.125 -226.275 ;
        RECT 303.795 -227.965 304.125 -227.635 ;
        RECT 303.795 -229.325 304.125 -228.995 ;
        RECT 303.795 -230.685 304.125 -230.355 ;
        RECT 303.795 -232.045 304.125 -231.715 ;
        RECT 303.795 -233.405 304.125 -233.075 ;
        RECT 303.795 -234.765 304.125 -234.435 ;
        RECT 303.795 -236.125 304.125 -235.795 ;
        RECT 303.795 -237.485 304.125 -237.155 ;
        RECT 303.795 -238.845 304.125 -238.515 ;
        RECT 303.795 -241.09 304.125 -239.96 ;
        RECT 303.8 -241.205 304.12 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 244.04 305.485 245.17 ;
        RECT 305.155 242.595 305.485 242.925 ;
        RECT 305.155 241.235 305.485 241.565 ;
        RECT 305.155 239.875 305.485 240.205 ;
        RECT 305.155 238.515 305.485 238.845 ;
        RECT 305.155 237.155 305.485 237.485 ;
        RECT 305.16 237.155 305.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 -0.845 305.485 -0.515 ;
        RECT 305.155 -2.205 305.485 -1.875 ;
        RECT 305.155 -3.565 305.485 -3.235 ;
        RECT 305.16 -3.565 305.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 -123.245 305.485 -122.915 ;
        RECT 305.155 -124.605 305.485 -124.275 ;
        RECT 305.155 -125.965 305.485 -125.635 ;
        RECT 305.155 -127.325 305.485 -126.995 ;
        RECT 305.155 -128.685 305.485 -128.355 ;
        RECT 305.155 -130.045 305.485 -129.715 ;
        RECT 305.155 -131.405 305.485 -131.075 ;
        RECT 305.155 -132.765 305.485 -132.435 ;
        RECT 305.155 -134.125 305.485 -133.795 ;
        RECT 305.155 -135.485 305.485 -135.155 ;
        RECT 305.155 -136.845 305.485 -136.515 ;
        RECT 305.155 -138.205 305.485 -137.875 ;
        RECT 305.155 -139.565 305.485 -139.235 ;
        RECT 305.155 -140.925 305.485 -140.595 ;
        RECT 305.155 -142.285 305.485 -141.955 ;
        RECT 305.155 -143.645 305.485 -143.315 ;
        RECT 305.155 -145.005 305.485 -144.675 ;
        RECT 305.155 -146.365 305.485 -146.035 ;
        RECT 305.155 -147.725 305.485 -147.395 ;
        RECT 305.155 -149.085 305.485 -148.755 ;
        RECT 305.155 -150.445 305.485 -150.115 ;
        RECT 305.155 -151.805 305.485 -151.475 ;
        RECT 305.155 -153.165 305.485 -152.835 ;
        RECT 305.155 -154.525 305.485 -154.195 ;
        RECT 305.155 -155.885 305.485 -155.555 ;
        RECT 305.155 -157.245 305.485 -156.915 ;
        RECT 305.155 -158.605 305.485 -158.275 ;
        RECT 305.155 -159.965 305.485 -159.635 ;
        RECT 305.155 -161.325 305.485 -160.995 ;
        RECT 305.155 -162.685 305.485 -162.355 ;
        RECT 305.155 -164.045 305.485 -163.715 ;
        RECT 305.155 -165.405 305.485 -165.075 ;
        RECT 305.155 -166.765 305.485 -166.435 ;
        RECT 305.155 -168.125 305.485 -167.795 ;
        RECT 305.155 -169.485 305.485 -169.155 ;
        RECT 305.155 -170.845 305.485 -170.515 ;
        RECT 305.155 -172.205 305.485 -171.875 ;
        RECT 305.155 -173.565 305.485 -173.235 ;
        RECT 305.155 -174.925 305.485 -174.595 ;
        RECT 305.155 -176.285 305.485 -175.955 ;
        RECT 305.155 -177.645 305.485 -177.315 ;
        RECT 305.155 -179.005 305.485 -178.675 ;
        RECT 305.155 -180.365 305.485 -180.035 ;
        RECT 305.155 -181.725 305.485 -181.395 ;
        RECT 305.155 -183.085 305.485 -182.755 ;
        RECT 305.155 -184.445 305.485 -184.115 ;
        RECT 305.155 -185.805 305.485 -185.475 ;
        RECT 305.155 -187.165 305.485 -186.835 ;
        RECT 305.155 -188.525 305.485 -188.195 ;
        RECT 305.155 -189.885 305.485 -189.555 ;
        RECT 305.155 -191.245 305.485 -190.915 ;
        RECT 305.155 -192.605 305.485 -192.275 ;
        RECT 305.155 -193.965 305.485 -193.635 ;
        RECT 305.155 -195.325 305.485 -194.995 ;
        RECT 305.155 -196.685 305.485 -196.355 ;
        RECT 305.155 -198.045 305.485 -197.715 ;
        RECT 305.155 -199.405 305.485 -199.075 ;
        RECT 305.155 -200.765 305.485 -200.435 ;
        RECT 305.155 -202.125 305.485 -201.795 ;
        RECT 305.155 -203.485 305.485 -203.155 ;
        RECT 305.155 -204.845 305.485 -204.515 ;
        RECT 305.155 -206.205 305.485 -205.875 ;
        RECT 305.155 -207.565 305.485 -207.235 ;
        RECT 305.155 -208.925 305.485 -208.595 ;
        RECT 305.155 -210.285 305.485 -209.955 ;
        RECT 305.155 -211.645 305.485 -211.315 ;
        RECT 305.155 -213.005 305.485 -212.675 ;
        RECT 305.155 -214.365 305.485 -214.035 ;
        RECT 305.155 -215.725 305.485 -215.395 ;
        RECT 305.155 -217.085 305.485 -216.755 ;
        RECT 305.155 -218.445 305.485 -218.115 ;
        RECT 305.155 -219.805 305.485 -219.475 ;
        RECT 305.155 -221.165 305.485 -220.835 ;
        RECT 305.155 -222.525 305.485 -222.195 ;
        RECT 305.155 -223.885 305.485 -223.555 ;
        RECT 305.155 -225.245 305.485 -224.915 ;
        RECT 305.155 -226.605 305.485 -226.275 ;
        RECT 305.155 -227.965 305.485 -227.635 ;
        RECT 305.155 -229.325 305.485 -228.995 ;
        RECT 305.155 -230.685 305.485 -230.355 ;
        RECT 305.155 -232.045 305.485 -231.715 ;
        RECT 305.155 -233.405 305.485 -233.075 ;
        RECT 305.155 -234.765 305.485 -234.435 ;
        RECT 305.155 -236.125 305.485 -235.795 ;
        RECT 305.155 -237.485 305.485 -237.155 ;
        RECT 305.155 -238.845 305.485 -238.515 ;
        RECT 305.155 -241.09 305.485 -239.96 ;
        RECT 305.16 -241.205 305.48 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 244.04 306.845 245.17 ;
        RECT 306.515 242.595 306.845 242.925 ;
        RECT 306.515 241.235 306.845 241.565 ;
        RECT 306.515 239.875 306.845 240.205 ;
        RECT 306.515 238.515 306.845 238.845 ;
        RECT 306.515 237.155 306.845 237.485 ;
        RECT 306.52 237.155 306.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 -0.845 306.845 -0.515 ;
        RECT 306.515 -2.205 306.845 -1.875 ;
        RECT 306.515 -3.565 306.845 -3.235 ;
        RECT 306.52 -3.565 306.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 -188.525 306.845 -188.195 ;
        RECT 306.515 -189.885 306.845 -189.555 ;
        RECT 306.515 -191.245 306.845 -190.915 ;
        RECT 306.515 -192.605 306.845 -192.275 ;
        RECT 306.515 -193.965 306.845 -193.635 ;
        RECT 306.515 -195.325 306.845 -194.995 ;
        RECT 306.515 -196.685 306.845 -196.355 ;
        RECT 306.515 -198.045 306.845 -197.715 ;
        RECT 306.515 -199.405 306.845 -199.075 ;
        RECT 306.515 -200.765 306.845 -200.435 ;
        RECT 306.515 -202.125 306.845 -201.795 ;
        RECT 306.515 -203.485 306.845 -203.155 ;
        RECT 306.515 -204.845 306.845 -204.515 ;
        RECT 306.515 -206.205 306.845 -205.875 ;
        RECT 306.515 -207.565 306.845 -207.235 ;
        RECT 306.515 -208.925 306.845 -208.595 ;
        RECT 306.515 -210.285 306.845 -209.955 ;
        RECT 306.515 -211.645 306.845 -211.315 ;
        RECT 306.515 -213.005 306.845 -212.675 ;
        RECT 306.515 -214.365 306.845 -214.035 ;
        RECT 306.515 -215.725 306.845 -215.395 ;
        RECT 306.515 -217.085 306.845 -216.755 ;
        RECT 306.515 -218.445 306.845 -218.115 ;
        RECT 306.515 -219.805 306.845 -219.475 ;
        RECT 306.515 -221.165 306.845 -220.835 ;
        RECT 306.515 -222.525 306.845 -222.195 ;
        RECT 306.515 -223.885 306.845 -223.555 ;
        RECT 306.515 -225.245 306.845 -224.915 ;
        RECT 306.515 -226.605 306.845 -226.275 ;
        RECT 306.515 -227.965 306.845 -227.635 ;
        RECT 306.515 -229.325 306.845 -228.995 ;
        RECT 306.515 -230.685 306.845 -230.355 ;
        RECT 306.515 -232.045 306.845 -231.715 ;
        RECT 306.515 -233.405 306.845 -233.075 ;
        RECT 306.515 -234.765 306.845 -234.435 ;
        RECT 306.515 -236.125 306.845 -235.795 ;
        RECT 306.515 -237.485 306.845 -237.155 ;
        RECT 306.515 -238.845 306.845 -238.515 ;
        RECT 306.515 -241.09 306.845 -239.96 ;
        RECT 306.52 -241.205 306.84 -122.24 ;
        RECT 306.515 -123.245 306.845 -122.915 ;
        RECT 306.515 -124.605 306.845 -124.275 ;
        RECT 306.515 -125.965 306.845 -125.635 ;
        RECT 306.515 -127.325 306.845 -126.995 ;
        RECT 306.515 -128.685 306.845 -128.355 ;
        RECT 306.515 -130.045 306.845 -129.715 ;
        RECT 306.515 -131.405 306.845 -131.075 ;
        RECT 306.515 -132.765 306.845 -132.435 ;
        RECT 306.515 -134.125 306.845 -133.795 ;
        RECT 306.515 -135.485 306.845 -135.155 ;
        RECT 306.515 -136.845 306.845 -136.515 ;
        RECT 306.515 -138.205 306.845 -137.875 ;
        RECT 306.515 -139.565 306.845 -139.235 ;
        RECT 306.515 -140.925 306.845 -140.595 ;
        RECT 306.515 -142.285 306.845 -141.955 ;
        RECT 306.515 -143.645 306.845 -143.315 ;
        RECT 306.515 -145.005 306.845 -144.675 ;
        RECT 306.515 -146.365 306.845 -146.035 ;
        RECT 306.515 -147.725 306.845 -147.395 ;
        RECT 306.515 -149.085 306.845 -148.755 ;
        RECT 306.515 -150.445 306.845 -150.115 ;
        RECT 306.515 -151.805 306.845 -151.475 ;
        RECT 306.515 -153.165 306.845 -152.835 ;
        RECT 306.515 -154.525 306.845 -154.195 ;
        RECT 306.515 -155.885 306.845 -155.555 ;
        RECT 306.515 -157.245 306.845 -156.915 ;
        RECT 306.515 -158.605 306.845 -158.275 ;
        RECT 306.515 -159.965 306.845 -159.635 ;
        RECT 306.515 -161.325 306.845 -160.995 ;
        RECT 306.515 -162.685 306.845 -162.355 ;
        RECT 306.515 -164.045 306.845 -163.715 ;
        RECT 306.515 -165.405 306.845 -165.075 ;
        RECT 306.515 -166.765 306.845 -166.435 ;
        RECT 306.515 -168.125 306.845 -167.795 ;
        RECT 306.515 -169.485 306.845 -169.155 ;
        RECT 306.515 -170.845 306.845 -170.515 ;
        RECT 306.515 -172.205 306.845 -171.875 ;
        RECT 306.515 -173.565 306.845 -173.235 ;
        RECT 306.515 -174.925 306.845 -174.595 ;
        RECT 306.515 -176.285 306.845 -175.955 ;
        RECT 306.515 -177.645 306.845 -177.315 ;
        RECT 306.515 -179.005 306.845 -178.675 ;
        RECT 306.515 -180.365 306.845 -180.035 ;
        RECT 306.515 -181.725 306.845 -181.395 ;
        RECT 306.515 -183.085 306.845 -182.755 ;
        RECT 306.515 -184.445 306.845 -184.115 ;
        RECT 306.515 -185.805 306.845 -185.475 ;
        RECT 306.515 -187.165 306.845 -186.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 244.04 272.845 245.17 ;
        RECT 272.515 242.595 272.845 242.925 ;
        RECT 272.515 241.235 272.845 241.565 ;
        RECT 272.515 239.875 272.845 240.205 ;
        RECT 272.515 238.515 272.845 238.845 ;
        RECT 272.515 237.155 272.845 237.485 ;
        RECT 272.52 237.155 272.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 -0.845 272.845 -0.515 ;
        RECT 272.515 -2.205 272.845 -1.875 ;
        RECT 272.515 -3.565 272.845 -3.235 ;
        RECT 272.52 -3.565 272.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 -123.245 272.845 -122.915 ;
        RECT 272.515 -124.605 272.845 -124.275 ;
        RECT 272.515 -125.965 272.845 -125.635 ;
        RECT 272.515 -127.325 272.845 -126.995 ;
        RECT 272.515 -128.685 272.845 -128.355 ;
        RECT 272.515 -130.045 272.845 -129.715 ;
        RECT 272.515 -131.405 272.845 -131.075 ;
        RECT 272.515 -132.765 272.845 -132.435 ;
        RECT 272.515 -134.125 272.845 -133.795 ;
        RECT 272.515 -135.485 272.845 -135.155 ;
        RECT 272.515 -136.845 272.845 -136.515 ;
        RECT 272.515 -138.205 272.845 -137.875 ;
        RECT 272.515 -139.565 272.845 -139.235 ;
        RECT 272.515 -140.925 272.845 -140.595 ;
        RECT 272.515 -142.285 272.845 -141.955 ;
        RECT 272.515 -143.645 272.845 -143.315 ;
        RECT 272.515 -145.005 272.845 -144.675 ;
        RECT 272.515 -146.365 272.845 -146.035 ;
        RECT 272.515 -147.725 272.845 -147.395 ;
        RECT 272.515 -149.085 272.845 -148.755 ;
        RECT 272.515 -150.445 272.845 -150.115 ;
        RECT 272.515 -151.805 272.845 -151.475 ;
        RECT 272.515 -153.165 272.845 -152.835 ;
        RECT 272.515 -154.525 272.845 -154.195 ;
        RECT 272.515 -155.885 272.845 -155.555 ;
        RECT 272.515 -157.245 272.845 -156.915 ;
        RECT 272.515 -158.605 272.845 -158.275 ;
        RECT 272.515 -159.965 272.845 -159.635 ;
        RECT 272.515 -161.325 272.845 -160.995 ;
        RECT 272.515 -162.685 272.845 -162.355 ;
        RECT 272.515 -164.045 272.845 -163.715 ;
        RECT 272.515 -165.405 272.845 -165.075 ;
        RECT 272.515 -166.765 272.845 -166.435 ;
        RECT 272.515 -168.125 272.845 -167.795 ;
        RECT 272.515 -169.485 272.845 -169.155 ;
        RECT 272.515 -170.845 272.845 -170.515 ;
        RECT 272.515 -172.205 272.845 -171.875 ;
        RECT 272.515 -173.565 272.845 -173.235 ;
        RECT 272.515 -174.925 272.845 -174.595 ;
        RECT 272.515 -176.285 272.845 -175.955 ;
        RECT 272.515 -177.645 272.845 -177.315 ;
        RECT 272.515 -179.005 272.845 -178.675 ;
        RECT 272.515 -180.365 272.845 -180.035 ;
        RECT 272.515 -181.725 272.845 -181.395 ;
        RECT 272.515 -183.085 272.845 -182.755 ;
        RECT 272.515 -184.445 272.845 -184.115 ;
        RECT 272.515 -185.805 272.845 -185.475 ;
        RECT 272.515 -187.165 272.845 -186.835 ;
        RECT 272.515 -188.525 272.845 -188.195 ;
        RECT 272.515 -189.885 272.845 -189.555 ;
        RECT 272.515 -191.245 272.845 -190.915 ;
        RECT 272.515 -192.605 272.845 -192.275 ;
        RECT 272.515 -193.965 272.845 -193.635 ;
        RECT 272.515 -195.325 272.845 -194.995 ;
        RECT 272.515 -196.685 272.845 -196.355 ;
        RECT 272.515 -198.045 272.845 -197.715 ;
        RECT 272.515 -199.405 272.845 -199.075 ;
        RECT 272.515 -200.765 272.845 -200.435 ;
        RECT 272.515 -202.125 272.845 -201.795 ;
        RECT 272.515 -203.485 272.845 -203.155 ;
        RECT 272.515 -204.845 272.845 -204.515 ;
        RECT 272.515 -206.205 272.845 -205.875 ;
        RECT 272.515 -207.565 272.845 -207.235 ;
        RECT 272.515 -208.925 272.845 -208.595 ;
        RECT 272.515 -210.285 272.845 -209.955 ;
        RECT 272.515 -211.645 272.845 -211.315 ;
        RECT 272.515 -213.005 272.845 -212.675 ;
        RECT 272.515 -214.365 272.845 -214.035 ;
        RECT 272.515 -215.725 272.845 -215.395 ;
        RECT 272.515 -217.085 272.845 -216.755 ;
        RECT 272.515 -218.445 272.845 -218.115 ;
        RECT 272.515 -219.805 272.845 -219.475 ;
        RECT 272.515 -221.165 272.845 -220.835 ;
        RECT 272.515 -222.525 272.845 -222.195 ;
        RECT 272.515 -223.885 272.845 -223.555 ;
        RECT 272.515 -225.245 272.845 -224.915 ;
        RECT 272.515 -226.605 272.845 -226.275 ;
        RECT 272.515 -227.965 272.845 -227.635 ;
        RECT 272.515 -229.325 272.845 -228.995 ;
        RECT 272.515 -230.685 272.845 -230.355 ;
        RECT 272.515 -232.045 272.845 -231.715 ;
        RECT 272.515 -233.405 272.845 -233.075 ;
        RECT 272.515 -234.765 272.845 -234.435 ;
        RECT 272.515 -236.125 272.845 -235.795 ;
        RECT 272.515 -237.485 272.845 -237.155 ;
        RECT 272.515 -238.845 272.845 -238.515 ;
        RECT 272.515 -241.09 272.845 -239.96 ;
        RECT 272.52 -241.205 272.84 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 244.04 274.205 245.17 ;
        RECT 273.875 242.595 274.205 242.925 ;
        RECT 273.875 241.235 274.205 241.565 ;
        RECT 273.875 239.875 274.205 240.205 ;
        RECT 273.875 238.515 274.205 238.845 ;
        RECT 273.875 237.155 274.205 237.485 ;
        RECT 273.88 237.155 274.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 -0.845 274.205 -0.515 ;
        RECT 273.875 -2.205 274.205 -1.875 ;
        RECT 273.875 -3.565 274.205 -3.235 ;
        RECT 273.88 -3.565 274.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 -123.245 274.205 -122.915 ;
        RECT 273.875 -124.605 274.205 -124.275 ;
        RECT 273.875 -125.965 274.205 -125.635 ;
        RECT 273.875 -127.325 274.205 -126.995 ;
        RECT 273.875 -128.685 274.205 -128.355 ;
        RECT 273.875 -130.045 274.205 -129.715 ;
        RECT 273.875 -131.405 274.205 -131.075 ;
        RECT 273.875 -132.765 274.205 -132.435 ;
        RECT 273.875 -134.125 274.205 -133.795 ;
        RECT 273.875 -135.485 274.205 -135.155 ;
        RECT 273.875 -136.845 274.205 -136.515 ;
        RECT 273.875 -138.205 274.205 -137.875 ;
        RECT 273.875 -139.565 274.205 -139.235 ;
        RECT 273.875 -140.925 274.205 -140.595 ;
        RECT 273.875 -142.285 274.205 -141.955 ;
        RECT 273.875 -143.645 274.205 -143.315 ;
        RECT 273.875 -145.005 274.205 -144.675 ;
        RECT 273.875 -146.365 274.205 -146.035 ;
        RECT 273.875 -147.725 274.205 -147.395 ;
        RECT 273.875 -149.085 274.205 -148.755 ;
        RECT 273.875 -150.445 274.205 -150.115 ;
        RECT 273.875 -151.805 274.205 -151.475 ;
        RECT 273.875 -153.165 274.205 -152.835 ;
        RECT 273.875 -154.525 274.205 -154.195 ;
        RECT 273.875 -155.885 274.205 -155.555 ;
        RECT 273.875 -157.245 274.205 -156.915 ;
        RECT 273.875 -158.605 274.205 -158.275 ;
        RECT 273.875 -159.965 274.205 -159.635 ;
        RECT 273.875 -161.325 274.205 -160.995 ;
        RECT 273.875 -162.685 274.205 -162.355 ;
        RECT 273.875 -164.045 274.205 -163.715 ;
        RECT 273.875 -165.405 274.205 -165.075 ;
        RECT 273.875 -166.765 274.205 -166.435 ;
        RECT 273.875 -168.125 274.205 -167.795 ;
        RECT 273.875 -169.485 274.205 -169.155 ;
        RECT 273.875 -170.845 274.205 -170.515 ;
        RECT 273.875 -172.205 274.205 -171.875 ;
        RECT 273.875 -173.565 274.205 -173.235 ;
        RECT 273.875 -174.925 274.205 -174.595 ;
        RECT 273.875 -176.285 274.205 -175.955 ;
        RECT 273.875 -177.645 274.205 -177.315 ;
        RECT 273.875 -179.005 274.205 -178.675 ;
        RECT 273.875 -180.365 274.205 -180.035 ;
        RECT 273.875 -181.725 274.205 -181.395 ;
        RECT 273.875 -183.085 274.205 -182.755 ;
        RECT 273.875 -184.445 274.205 -184.115 ;
        RECT 273.875 -185.805 274.205 -185.475 ;
        RECT 273.875 -187.165 274.205 -186.835 ;
        RECT 273.875 -188.525 274.205 -188.195 ;
        RECT 273.875 -189.885 274.205 -189.555 ;
        RECT 273.875 -191.245 274.205 -190.915 ;
        RECT 273.875 -192.605 274.205 -192.275 ;
        RECT 273.875 -193.965 274.205 -193.635 ;
        RECT 273.875 -195.325 274.205 -194.995 ;
        RECT 273.875 -196.685 274.205 -196.355 ;
        RECT 273.875 -198.045 274.205 -197.715 ;
        RECT 273.875 -199.405 274.205 -199.075 ;
        RECT 273.875 -200.765 274.205 -200.435 ;
        RECT 273.875 -202.125 274.205 -201.795 ;
        RECT 273.875 -203.485 274.205 -203.155 ;
        RECT 273.875 -204.845 274.205 -204.515 ;
        RECT 273.875 -206.205 274.205 -205.875 ;
        RECT 273.875 -207.565 274.205 -207.235 ;
        RECT 273.875 -208.925 274.205 -208.595 ;
        RECT 273.875 -210.285 274.205 -209.955 ;
        RECT 273.875 -211.645 274.205 -211.315 ;
        RECT 273.875 -213.005 274.205 -212.675 ;
        RECT 273.875 -214.365 274.205 -214.035 ;
        RECT 273.875 -215.725 274.205 -215.395 ;
        RECT 273.875 -217.085 274.205 -216.755 ;
        RECT 273.875 -218.445 274.205 -218.115 ;
        RECT 273.875 -219.805 274.205 -219.475 ;
        RECT 273.875 -221.165 274.205 -220.835 ;
        RECT 273.875 -222.525 274.205 -222.195 ;
        RECT 273.875 -223.885 274.205 -223.555 ;
        RECT 273.875 -225.245 274.205 -224.915 ;
        RECT 273.875 -226.605 274.205 -226.275 ;
        RECT 273.875 -227.965 274.205 -227.635 ;
        RECT 273.875 -229.325 274.205 -228.995 ;
        RECT 273.875 -230.685 274.205 -230.355 ;
        RECT 273.875 -232.045 274.205 -231.715 ;
        RECT 273.875 -233.405 274.205 -233.075 ;
        RECT 273.875 -234.765 274.205 -234.435 ;
        RECT 273.875 -236.125 274.205 -235.795 ;
        RECT 273.875 -237.485 274.205 -237.155 ;
        RECT 273.875 -238.845 274.205 -238.515 ;
        RECT 273.875 -241.09 274.205 -239.96 ;
        RECT 273.88 -241.205 274.2 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 244.04 275.565 245.17 ;
        RECT 275.235 242.595 275.565 242.925 ;
        RECT 275.235 241.235 275.565 241.565 ;
        RECT 275.235 239.875 275.565 240.205 ;
        RECT 275.235 238.515 275.565 238.845 ;
        RECT 275.235 237.155 275.565 237.485 ;
        RECT 275.24 237.155 275.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 -127.325 275.565 -126.995 ;
        RECT 275.235 -128.685 275.565 -128.355 ;
        RECT 275.235 -130.045 275.565 -129.715 ;
        RECT 275.235 -131.405 275.565 -131.075 ;
        RECT 275.235 -132.765 275.565 -132.435 ;
        RECT 275.235 -134.125 275.565 -133.795 ;
        RECT 275.235 -135.485 275.565 -135.155 ;
        RECT 275.235 -136.845 275.565 -136.515 ;
        RECT 275.235 -138.205 275.565 -137.875 ;
        RECT 275.235 -139.565 275.565 -139.235 ;
        RECT 275.235 -140.925 275.565 -140.595 ;
        RECT 275.235 -142.285 275.565 -141.955 ;
        RECT 275.235 -143.645 275.565 -143.315 ;
        RECT 275.235 -145.005 275.565 -144.675 ;
        RECT 275.235 -146.365 275.565 -146.035 ;
        RECT 275.235 -147.725 275.565 -147.395 ;
        RECT 275.235 -149.085 275.565 -148.755 ;
        RECT 275.235 -150.445 275.565 -150.115 ;
        RECT 275.235 -151.805 275.565 -151.475 ;
        RECT 275.235 -153.165 275.565 -152.835 ;
        RECT 275.235 -154.525 275.565 -154.195 ;
        RECT 275.235 -155.885 275.565 -155.555 ;
        RECT 275.235 -157.245 275.565 -156.915 ;
        RECT 275.235 -158.605 275.565 -158.275 ;
        RECT 275.235 -159.965 275.565 -159.635 ;
        RECT 275.235 -161.325 275.565 -160.995 ;
        RECT 275.235 -162.685 275.565 -162.355 ;
        RECT 275.235 -164.045 275.565 -163.715 ;
        RECT 275.235 -165.405 275.565 -165.075 ;
        RECT 275.235 -166.765 275.565 -166.435 ;
        RECT 275.235 -168.125 275.565 -167.795 ;
        RECT 275.235 -169.485 275.565 -169.155 ;
        RECT 275.235 -170.845 275.565 -170.515 ;
        RECT 275.235 -172.205 275.565 -171.875 ;
        RECT 275.235 -173.565 275.565 -173.235 ;
        RECT 275.235 -174.925 275.565 -174.595 ;
        RECT 275.235 -176.285 275.565 -175.955 ;
        RECT 275.235 -177.645 275.565 -177.315 ;
        RECT 275.235 -179.005 275.565 -178.675 ;
        RECT 275.235 -180.365 275.565 -180.035 ;
        RECT 275.235 -181.725 275.565 -181.395 ;
        RECT 275.235 -183.085 275.565 -182.755 ;
        RECT 275.235 -184.445 275.565 -184.115 ;
        RECT 275.235 -185.805 275.565 -185.475 ;
        RECT 275.235 -187.165 275.565 -186.835 ;
        RECT 275.235 -188.525 275.565 -188.195 ;
        RECT 275.235 -189.885 275.565 -189.555 ;
        RECT 275.235 -191.245 275.565 -190.915 ;
        RECT 275.235 -192.605 275.565 -192.275 ;
        RECT 275.235 -193.965 275.565 -193.635 ;
        RECT 275.235 -195.325 275.565 -194.995 ;
        RECT 275.235 -196.685 275.565 -196.355 ;
        RECT 275.235 -198.045 275.565 -197.715 ;
        RECT 275.235 -199.405 275.565 -199.075 ;
        RECT 275.235 -200.765 275.565 -200.435 ;
        RECT 275.235 -202.125 275.565 -201.795 ;
        RECT 275.235 -203.485 275.565 -203.155 ;
        RECT 275.235 -204.845 275.565 -204.515 ;
        RECT 275.235 -206.205 275.565 -205.875 ;
        RECT 275.235 -207.565 275.565 -207.235 ;
        RECT 275.235 -208.925 275.565 -208.595 ;
        RECT 275.235 -210.285 275.565 -209.955 ;
        RECT 275.235 -211.645 275.565 -211.315 ;
        RECT 275.235 -213.005 275.565 -212.675 ;
        RECT 275.235 -214.365 275.565 -214.035 ;
        RECT 275.235 -215.725 275.565 -215.395 ;
        RECT 275.235 -217.085 275.565 -216.755 ;
        RECT 275.235 -218.445 275.565 -218.115 ;
        RECT 275.235 -219.805 275.565 -219.475 ;
        RECT 275.235 -221.165 275.565 -220.835 ;
        RECT 275.235 -222.525 275.565 -222.195 ;
        RECT 275.235 -223.885 275.565 -223.555 ;
        RECT 275.235 -225.245 275.565 -224.915 ;
        RECT 275.235 -226.605 275.565 -226.275 ;
        RECT 275.235 -227.965 275.565 -227.635 ;
        RECT 275.235 -229.325 275.565 -228.995 ;
        RECT 275.235 -230.685 275.565 -230.355 ;
        RECT 275.235 -232.045 275.565 -231.715 ;
        RECT 275.235 -233.405 275.565 -233.075 ;
        RECT 275.235 -234.765 275.565 -234.435 ;
        RECT 275.235 -236.125 275.565 -235.795 ;
        RECT 275.235 -237.485 275.565 -237.155 ;
        RECT 275.235 -238.845 275.565 -238.515 ;
        RECT 275.235 -241.09 275.565 -239.96 ;
        RECT 275.24 -241.205 275.56 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.81 -125.535 276.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 244.04 276.925 245.17 ;
        RECT 276.595 242.595 276.925 242.925 ;
        RECT 276.595 241.235 276.925 241.565 ;
        RECT 276.595 239.875 276.925 240.205 ;
        RECT 276.595 238.515 276.925 238.845 ;
        RECT 276.595 237.155 276.925 237.485 ;
        RECT 276.6 237.155 276.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 -0.845 276.925 -0.515 ;
        RECT 276.595 -2.205 276.925 -1.875 ;
        RECT 276.595 -3.565 276.925 -3.235 ;
        RECT 276.6 -3.565 276.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.955 244.04 278.285 245.17 ;
        RECT 277.955 242.595 278.285 242.925 ;
        RECT 277.955 241.235 278.285 241.565 ;
        RECT 277.955 239.875 278.285 240.205 ;
        RECT 277.955 238.515 278.285 238.845 ;
        RECT 277.955 237.155 278.285 237.485 ;
        RECT 277.96 237.155 278.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.955 -0.845 278.285 -0.515 ;
        RECT 277.955 -2.205 278.285 -1.875 ;
        RECT 277.955 -3.565 278.285 -3.235 ;
        RECT 277.96 -3.565 278.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 244.04 279.645 245.17 ;
        RECT 279.315 242.595 279.645 242.925 ;
        RECT 279.315 241.235 279.645 241.565 ;
        RECT 279.315 239.875 279.645 240.205 ;
        RECT 279.315 238.515 279.645 238.845 ;
        RECT 279.315 237.155 279.645 237.485 ;
        RECT 279.32 237.155 279.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 -0.845 279.645 -0.515 ;
        RECT 279.315 -2.205 279.645 -1.875 ;
        RECT 279.315 -3.565 279.645 -3.235 ;
        RECT 279.32 -3.565 279.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 -123.245 279.645 -122.915 ;
        RECT 279.315 -124.605 279.645 -124.275 ;
        RECT 279.315 -125.965 279.645 -125.635 ;
        RECT 279.315 -127.325 279.645 -126.995 ;
        RECT 279.315 -128.685 279.645 -128.355 ;
        RECT 279.315 -130.045 279.645 -129.715 ;
        RECT 279.315 -131.405 279.645 -131.075 ;
        RECT 279.315 -132.765 279.645 -132.435 ;
        RECT 279.315 -134.125 279.645 -133.795 ;
        RECT 279.315 -135.485 279.645 -135.155 ;
        RECT 279.315 -136.845 279.645 -136.515 ;
        RECT 279.315 -138.205 279.645 -137.875 ;
        RECT 279.315 -139.565 279.645 -139.235 ;
        RECT 279.315 -140.925 279.645 -140.595 ;
        RECT 279.315 -142.285 279.645 -141.955 ;
        RECT 279.315 -143.645 279.645 -143.315 ;
        RECT 279.315 -145.005 279.645 -144.675 ;
        RECT 279.315 -146.365 279.645 -146.035 ;
        RECT 279.315 -147.725 279.645 -147.395 ;
        RECT 279.315 -149.085 279.645 -148.755 ;
        RECT 279.315 -150.445 279.645 -150.115 ;
        RECT 279.315 -151.805 279.645 -151.475 ;
        RECT 279.315 -153.165 279.645 -152.835 ;
        RECT 279.315 -154.525 279.645 -154.195 ;
        RECT 279.315 -155.885 279.645 -155.555 ;
        RECT 279.315 -157.245 279.645 -156.915 ;
        RECT 279.315 -158.605 279.645 -158.275 ;
        RECT 279.315 -159.965 279.645 -159.635 ;
        RECT 279.315 -161.325 279.645 -160.995 ;
        RECT 279.315 -162.685 279.645 -162.355 ;
        RECT 279.315 -164.045 279.645 -163.715 ;
        RECT 279.315 -165.405 279.645 -165.075 ;
        RECT 279.315 -166.765 279.645 -166.435 ;
        RECT 279.315 -168.125 279.645 -167.795 ;
        RECT 279.315 -169.485 279.645 -169.155 ;
        RECT 279.315 -170.845 279.645 -170.515 ;
        RECT 279.315 -172.205 279.645 -171.875 ;
        RECT 279.315 -173.565 279.645 -173.235 ;
        RECT 279.315 -174.925 279.645 -174.595 ;
        RECT 279.315 -176.285 279.645 -175.955 ;
        RECT 279.315 -177.645 279.645 -177.315 ;
        RECT 279.315 -179.005 279.645 -178.675 ;
        RECT 279.315 -180.365 279.645 -180.035 ;
        RECT 279.315 -181.725 279.645 -181.395 ;
        RECT 279.315 -183.085 279.645 -182.755 ;
        RECT 279.315 -184.445 279.645 -184.115 ;
        RECT 279.315 -185.805 279.645 -185.475 ;
        RECT 279.315 -187.165 279.645 -186.835 ;
        RECT 279.315 -188.525 279.645 -188.195 ;
        RECT 279.315 -189.885 279.645 -189.555 ;
        RECT 279.315 -191.245 279.645 -190.915 ;
        RECT 279.315 -192.605 279.645 -192.275 ;
        RECT 279.315 -193.965 279.645 -193.635 ;
        RECT 279.315 -195.325 279.645 -194.995 ;
        RECT 279.315 -196.685 279.645 -196.355 ;
        RECT 279.315 -198.045 279.645 -197.715 ;
        RECT 279.315 -199.405 279.645 -199.075 ;
        RECT 279.315 -200.765 279.645 -200.435 ;
        RECT 279.315 -202.125 279.645 -201.795 ;
        RECT 279.315 -203.485 279.645 -203.155 ;
        RECT 279.315 -204.845 279.645 -204.515 ;
        RECT 279.315 -206.205 279.645 -205.875 ;
        RECT 279.315 -207.565 279.645 -207.235 ;
        RECT 279.315 -208.925 279.645 -208.595 ;
        RECT 279.315 -210.285 279.645 -209.955 ;
        RECT 279.315 -211.645 279.645 -211.315 ;
        RECT 279.315 -213.005 279.645 -212.675 ;
        RECT 279.315 -214.365 279.645 -214.035 ;
        RECT 279.315 -215.725 279.645 -215.395 ;
        RECT 279.315 -217.085 279.645 -216.755 ;
        RECT 279.315 -218.445 279.645 -218.115 ;
        RECT 279.315 -219.805 279.645 -219.475 ;
        RECT 279.315 -221.165 279.645 -220.835 ;
        RECT 279.315 -222.525 279.645 -222.195 ;
        RECT 279.315 -223.885 279.645 -223.555 ;
        RECT 279.315 -225.245 279.645 -224.915 ;
        RECT 279.315 -226.605 279.645 -226.275 ;
        RECT 279.315 -227.965 279.645 -227.635 ;
        RECT 279.315 -229.325 279.645 -228.995 ;
        RECT 279.315 -230.685 279.645 -230.355 ;
        RECT 279.315 -232.045 279.645 -231.715 ;
        RECT 279.315 -233.405 279.645 -233.075 ;
        RECT 279.315 -234.765 279.645 -234.435 ;
        RECT 279.315 -236.125 279.645 -235.795 ;
        RECT 279.315 -237.485 279.645 -237.155 ;
        RECT 279.315 -238.845 279.645 -238.515 ;
        RECT 279.315 -241.09 279.645 -239.96 ;
        RECT 279.32 -241.205 279.64 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 244.04 281.005 245.17 ;
        RECT 280.675 242.595 281.005 242.925 ;
        RECT 280.675 241.235 281.005 241.565 ;
        RECT 280.675 239.875 281.005 240.205 ;
        RECT 280.675 238.515 281.005 238.845 ;
        RECT 280.675 237.155 281.005 237.485 ;
        RECT 280.68 237.155 281 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 -0.845 281.005 -0.515 ;
        RECT 280.675 -2.205 281.005 -1.875 ;
        RECT 280.675 -3.565 281.005 -3.235 ;
        RECT 280.68 -3.565 281 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 -123.245 281.005 -122.915 ;
        RECT 280.675 -124.605 281.005 -124.275 ;
        RECT 280.675 -125.965 281.005 -125.635 ;
        RECT 280.675 -127.325 281.005 -126.995 ;
        RECT 280.675 -128.685 281.005 -128.355 ;
        RECT 280.675 -130.045 281.005 -129.715 ;
        RECT 280.675 -131.405 281.005 -131.075 ;
        RECT 280.675 -132.765 281.005 -132.435 ;
        RECT 280.675 -134.125 281.005 -133.795 ;
        RECT 280.675 -135.485 281.005 -135.155 ;
        RECT 280.675 -136.845 281.005 -136.515 ;
        RECT 280.675 -138.205 281.005 -137.875 ;
        RECT 280.675 -139.565 281.005 -139.235 ;
        RECT 280.675 -140.925 281.005 -140.595 ;
        RECT 280.675 -142.285 281.005 -141.955 ;
        RECT 280.675 -143.645 281.005 -143.315 ;
        RECT 280.675 -145.005 281.005 -144.675 ;
        RECT 280.675 -146.365 281.005 -146.035 ;
        RECT 280.675 -147.725 281.005 -147.395 ;
        RECT 280.675 -149.085 281.005 -148.755 ;
        RECT 280.675 -150.445 281.005 -150.115 ;
        RECT 280.675 -151.805 281.005 -151.475 ;
        RECT 280.675 -153.165 281.005 -152.835 ;
        RECT 280.675 -154.525 281.005 -154.195 ;
        RECT 280.675 -155.885 281.005 -155.555 ;
        RECT 280.675 -157.245 281.005 -156.915 ;
        RECT 280.675 -158.605 281.005 -158.275 ;
        RECT 280.675 -159.965 281.005 -159.635 ;
        RECT 280.675 -161.325 281.005 -160.995 ;
        RECT 280.675 -162.685 281.005 -162.355 ;
        RECT 280.675 -164.045 281.005 -163.715 ;
        RECT 280.675 -165.405 281.005 -165.075 ;
        RECT 280.675 -166.765 281.005 -166.435 ;
        RECT 280.675 -168.125 281.005 -167.795 ;
        RECT 280.675 -169.485 281.005 -169.155 ;
        RECT 280.675 -170.845 281.005 -170.515 ;
        RECT 280.675 -172.205 281.005 -171.875 ;
        RECT 280.675 -173.565 281.005 -173.235 ;
        RECT 280.675 -174.925 281.005 -174.595 ;
        RECT 280.675 -176.285 281.005 -175.955 ;
        RECT 280.675 -177.645 281.005 -177.315 ;
        RECT 280.675 -179.005 281.005 -178.675 ;
        RECT 280.675 -180.365 281.005 -180.035 ;
        RECT 280.675 -181.725 281.005 -181.395 ;
        RECT 280.675 -183.085 281.005 -182.755 ;
        RECT 280.675 -184.445 281.005 -184.115 ;
        RECT 280.675 -185.805 281.005 -185.475 ;
        RECT 280.675 -187.165 281.005 -186.835 ;
        RECT 280.675 -188.525 281.005 -188.195 ;
        RECT 280.675 -189.885 281.005 -189.555 ;
        RECT 280.675 -191.245 281.005 -190.915 ;
        RECT 280.675 -192.605 281.005 -192.275 ;
        RECT 280.675 -193.965 281.005 -193.635 ;
        RECT 280.675 -195.325 281.005 -194.995 ;
        RECT 280.675 -196.685 281.005 -196.355 ;
        RECT 280.675 -198.045 281.005 -197.715 ;
        RECT 280.675 -199.405 281.005 -199.075 ;
        RECT 280.675 -200.765 281.005 -200.435 ;
        RECT 280.675 -202.125 281.005 -201.795 ;
        RECT 280.675 -203.485 281.005 -203.155 ;
        RECT 280.675 -204.845 281.005 -204.515 ;
        RECT 280.675 -206.205 281.005 -205.875 ;
        RECT 280.675 -207.565 281.005 -207.235 ;
        RECT 280.675 -208.925 281.005 -208.595 ;
        RECT 280.675 -210.285 281.005 -209.955 ;
        RECT 280.675 -211.645 281.005 -211.315 ;
        RECT 280.675 -213.005 281.005 -212.675 ;
        RECT 280.675 -214.365 281.005 -214.035 ;
        RECT 280.675 -215.725 281.005 -215.395 ;
        RECT 280.675 -217.085 281.005 -216.755 ;
        RECT 280.675 -218.445 281.005 -218.115 ;
        RECT 280.675 -219.805 281.005 -219.475 ;
        RECT 280.675 -221.165 281.005 -220.835 ;
        RECT 280.675 -222.525 281.005 -222.195 ;
        RECT 280.675 -223.885 281.005 -223.555 ;
        RECT 280.675 -225.245 281.005 -224.915 ;
        RECT 280.675 -226.605 281.005 -226.275 ;
        RECT 280.675 -227.965 281.005 -227.635 ;
        RECT 280.675 -229.325 281.005 -228.995 ;
        RECT 280.675 -230.685 281.005 -230.355 ;
        RECT 280.675 -232.045 281.005 -231.715 ;
        RECT 280.675 -233.405 281.005 -233.075 ;
        RECT 280.675 -234.765 281.005 -234.435 ;
        RECT 280.675 -236.125 281.005 -235.795 ;
        RECT 280.675 -237.485 281.005 -237.155 ;
        RECT 280.675 -238.845 281.005 -238.515 ;
        RECT 280.675 -241.09 281.005 -239.96 ;
        RECT 280.68 -241.205 281 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 244.04 282.365 245.17 ;
        RECT 282.035 242.595 282.365 242.925 ;
        RECT 282.035 241.235 282.365 241.565 ;
        RECT 282.035 239.875 282.365 240.205 ;
        RECT 282.035 238.515 282.365 238.845 ;
        RECT 282.035 237.155 282.365 237.485 ;
        RECT 282.04 237.155 282.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 -0.845 282.365 -0.515 ;
        RECT 282.035 -2.205 282.365 -1.875 ;
        RECT 282.035 -3.565 282.365 -3.235 ;
        RECT 282.04 -3.565 282.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 -123.245 282.365 -122.915 ;
        RECT 282.035 -124.605 282.365 -124.275 ;
        RECT 282.035 -125.965 282.365 -125.635 ;
        RECT 282.035 -127.325 282.365 -126.995 ;
        RECT 282.035 -128.685 282.365 -128.355 ;
        RECT 282.035 -130.045 282.365 -129.715 ;
        RECT 282.035 -131.405 282.365 -131.075 ;
        RECT 282.035 -132.765 282.365 -132.435 ;
        RECT 282.035 -134.125 282.365 -133.795 ;
        RECT 282.035 -135.485 282.365 -135.155 ;
        RECT 282.035 -136.845 282.365 -136.515 ;
        RECT 282.035 -138.205 282.365 -137.875 ;
        RECT 282.035 -139.565 282.365 -139.235 ;
        RECT 282.035 -140.925 282.365 -140.595 ;
        RECT 282.035 -142.285 282.365 -141.955 ;
        RECT 282.035 -143.645 282.365 -143.315 ;
        RECT 282.035 -145.005 282.365 -144.675 ;
        RECT 282.035 -146.365 282.365 -146.035 ;
        RECT 282.035 -147.725 282.365 -147.395 ;
        RECT 282.035 -149.085 282.365 -148.755 ;
        RECT 282.035 -150.445 282.365 -150.115 ;
        RECT 282.035 -151.805 282.365 -151.475 ;
        RECT 282.035 -153.165 282.365 -152.835 ;
        RECT 282.035 -154.525 282.365 -154.195 ;
        RECT 282.035 -155.885 282.365 -155.555 ;
        RECT 282.035 -157.245 282.365 -156.915 ;
        RECT 282.035 -158.605 282.365 -158.275 ;
        RECT 282.035 -159.965 282.365 -159.635 ;
        RECT 282.035 -161.325 282.365 -160.995 ;
        RECT 282.035 -162.685 282.365 -162.355 ;
        RECT 282.035 -164.045 282.365 -163.715 ;
        RECT 282.035 -165.405 282.365 -165.075 ;
        RECT 282.035 -166.765 282.365 -166.435 ;
        RECT 282.035 -168.125 282.365 -167.795 ;
        RECT 282.035 -169.485 282.365 -169.155 ;
        RECT 282.035 -170.845 282.365 -170.515 ;
        RECT 282.035 -172.205 282.365 -171.875 ;
        RECT 282.035 -173.565 282.365 -173.235 ;
        RECT 282.035 -174.925 282.365 -174.595 ;
        RECT 282.035 -176.285 282.365 -175.955 ;
        RECT 282.035 -177.645 282.365 -177.315 ;
        RECT 282.035 -179.005 282.365 -178.675 ;
        RECT 282.035 -180.365 282.365 -180.035 ;
        RECT 282.035 -181.725 282.365 -181.395 ;
        RECT 282.035 -183.085 282.365 -182.755 ;
        RECT 282.035 -184.445 282.365 -184.115 ;
        RECT 282.035 -185.805 282.365 -185.475 ;
        RECT 282.035 -187.165 282.365 -186.835 ;
        RECT 282.035 -188.525 282.365 -188.195 ;
        RECT 282.035 -189.885 282.365 -189.555 ;
        RECT 282.035 -191.245 282.365 -190.915 ;
        RECT 282.035 -192.605 282.365 -192.275 ;
        RECT 282.035 -193.965 282.365 -193.635 ;
        RECT 282.035 -195.325 282.365 -194.995 ;
        RECT 282.035 -196.685 282.365 -196.355 ;
        RECT 282.035 -198.045 282.365 -197.715 ;
        RECT 282.035 -199.405 282.365 -199.075 ;
        RECT 282.035 -200.765 282.365 -200.435 ;
        RECT 282.035 -202.125 282.365 -201.795 ;
        RECT 282.035 -203.485 282.365 -203.155 ;
        RECT 282.035 -204.845 282.365 -204.515 ;
        RECT 282.035 -206.205 282.365 -205.875 ;
        RECT 282.035 -207.565 282.365 -207.235 ;
        RECT 282.035 -208.925 282.365 -208.595 ;
        RECT 282.035 -210.285 282.365 -209.955 ;
        RECT 282.035 -211.645 282.365 -211.315 ;
        RECT 282.035 -213.005 282.365 -212.675 ;
        RECT 282.035 -214.365 282.365 -214.035 ;
        RECT 282.035 -215.725 282.365 -215.395 ;
        RECT 282.035 -217.085 282.365 -216.755 ;
        RECT 282.035 -218.445 282.365 -218.115 ;
        RECT 282.035 -219.805 282.365 -219.475 ;
        RECT 282.035 -221.165 282.365 -220.835 ;
        RECT 282.035 -222.525 282.365 -222.195 ;
        RECT 282.035 -223.885 282.365 -223.555 ;
        RECT 282.035 -225.245 282.365 -224.915 ;
        RECT 282.035 -226.605 282.365 -226.275 ;
        RECT 282.035 -227.965 282.365 -227.635 ;
        RECT 282.035 -229.325 282.365 -228.995 ;
        RECT 282.035 -230.685 282.365 -230.355 ;
        RECT 282.035 -232.045 282.365 -231.715 ;
        RECT 282.035 -233.405 282.365 -233.075 ;
        RECT 282.035 -234.765 282.365 -234.435 ;
        RECT 282.035 -236.125 282.365 -235.795 ;
        RECT 282.035 -237.485 282.365 -237.155 ;
        RECT 282.035 -238.845 282.365 -238.515 ;
        RECT 282.035 -241.09 282.365 -239.96 ;
        RECT 282.04 -241.205 282.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 244.04 283.725 245.17 ;
        RECT 283.395 242.595 283.725 242.925 ;
        RECT 283.395 241.235 283.725 241.565 ;
        RECT 283.395 239.875 283.725 240.205 ;
        RECT 283.395 238.515 283.725 238.845 ;
        RECT 283.395 237.155 283.725 237.485 ;
        RECT 283.4 237.155 283.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 -0.845 283.725 -0.515 ;
        RECT 283.395 -2.205 283.725 -1.875 ;
        RECT 283.395 -3.565 283.725 -3.235 ;
        RECT 283.4 -3.565 283.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 -123.245 283.725 -122.915 ;
        RECT 283.395 -124.605 283.725 -124.275 ;
        RECT 283.395 -125.965 283.725 -125.635 ;
        RECT 283.395 -127.325 283.725 -126.995 ;
        RECT 283.395 -128.685 283.725 -128.355 ;
        RECT 283.395 -130.045 283.725 -129.715 ;
        RECT 283.395 -131.405 283.725 -131.075 ;
        RECT 283.395 -132.765 283.725 -132.435 ;
        RECT 283.395 -134.125 283.725 -133.795 ;
        RECT 283.395 -135.485 283.725 -135.155 ;
        RECT 283.395 -136.845 283.725 -136.515 ;
        RECT 283.395 -138.205 283.725 -137.875 ;
        RECT 283.395 -139.565 283.725 -139.235 ;
        RECT 283.395 -140.925 283.725 -140.595 ;
        RECT 283.395 -142.285 283.725 -141.955 ;
        RECT 283.395 -143.645 283.725 -143.315 ;
        RECT 283.395 -145.005 283.725 -144.675 ;
        RECT 283.395 -146.365 283.725 -146.035 ;
        RECT 283.395 -147.725 283.725 -147.395 ;
        RECT 283.395 -149.085 283.725 -148.755 ;
        RECT 283.395 -150.445 283.725 -150.115 ;
        RECT 283.395 -151.805 283.725 -151.475 ;
        RECT 283.395 -153.165 283.725 -152.835 ;
        RECT 283.395 -154.525 283.725 -154.195 ;
        RECT 283.395 -155.885 283.725 -155.555 ;
        RECT 283.395 -157.245 283.725 -156.915 ;
        RECT 283.395 -158.605 283.725 -158.275 ;
        RECT 283.395 -159.965 283.725 -159.635 ;
        RECT 283.395 -161.325 283.725 -160.995 ;
        RECT 283.395 -162.685 283.725 -162.355 ;
        RECT 283.395 -164.045 283.725 -163.715 ;
        RECT 283.395 -165.405 283.725 -165.075 ;
        RECT 283.395 -166.765 283.725 -166.435 ;
        RECT 283.395 -168.125 283.725 -167.795 ;
        RECT 283.395 -169.485 283.725 -169.155 ;
        RECT 283.395 -170.845 283.725 -170.515 ;
        RECT 283.395 -172.205 283.725 -171.875 ;
        RECT 283.395 -173.565 283.725 -173.235 ;
        RECT 283.395 -174.925 283.725 -174.595 ;
        RECT 283.395 -176.285 283.725 -175.955 ;
        RECT 283.395 -177.645 283.725 -177.315 ;
        RECT 283.395 -179.005 283.725 -178.675 ;
        RECT 283.395 -180.365 283.725 -180.035 ;
        RECT 283.395 -181.725 283.725 -181.395 ;
        RECT 283.395 -183.085 283.725 -182.755 ;
        RECT 283.395 -184.445 283.725 -184.115 ;
        RECT 283.395 -185.805 283.725 -185.475 ;
        RECT 283.395 -187.165 283.725 -186.835 ;
        RECT 283.395 -188.525 283.725 -188.195 ;
        RECT 283.395 -189.885 283.725 -189.555 ;
        RECT 283.395 -191.245 283.725 -190.915 ;
        RECT 283.395 -192.605 283.725 -192.275 ;
        RECT 283.395 -193.965 283.725 -193.635 ;
        RECT 283.395 -195.325 283.725 -194.995 ;
        RECT 283.395 -196.685 283.725 -196.355 ;
        RECT 283.395 -198.045 283.725 -197.715 ;
        RECT 283.395 -199.405 283.725 -199.075 ;
        RECT 283.395 -200.765 283.725 -200.435 ;
        RECT 283.395 -202.125 283.725 -201.795 ;
        RECT 283.395 -203.485 283.725 -203.155 ;
        RECT 283.395 -204.845 283.725 -204.515 ;
        RECT 283.395 -206.205 283.725 -205.875 ;
        RECT 283.395 -207.565 283.725 -207.235 ;
        RECT 283.395 -208.925 283.725 -208.595 ;
        RECT 283.395 -210.285 283.725 -209.955 ;
        RECT 283.395 -211.645 283.725 -211.315 ;
        RECT 283.395 -213.005 283.725 -212.675 ;
        RECT 283.395 -214.365 283.725 -214.035 ;
        RECT 283.395 -215.725 283.725 -215.395 ;
        RECT 283.395 -217.085 283.725 -216.755 ;
        RECT 283.395 -218.445 283.725 -218.115 ;
        RECT 283.395 -219.805 283.725 -219.475 ;
        RECT 283.395 -221.165 283.725 -220.835 ;
        RECT 283.395 -222.525 283.725 -222.195 ;
        RECT 283.395 -223.885 283.725 -223.555 ;
        RECT 283.395 -225.245 283.725 -224.915 ;
        RECT 283.395 -226.605 283.725 -226.275 ;
        RECT 283.395 -227.965 283.725 -227.635 ;
        RECT 283.395 -229.325 283.725 -228.995 ;
        RECT 283.395 -230.685 283.725 -230.355 ;
        RECT 283.395 -232.045 283.725 -231.715 ;
        RECT 283.395 -233.405 283.725 -233.075 ;
        RECT 283.395 -234.765 283.725 -234.435 ;
        RECT 283.395 -236.125 283.725 -235.795 ;
        RECT 283.395 -237.485 283.725 -237.155 ;
        RECT 283.395 -238.845 283.725 -238.515 ;
        RECT 283.395 -241.09 283.725 -239.96 ;
        RECT 283.4 -241.205 283.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 244.04 285.085 245.17 ;
        RECT 284.755 242.595 285.085 242.925 ;
        RECT 284.755 241.235 285.085 241.565 ;
        RECT 284.755 239.875 285.085 240.205 ;
        RECT 284.755 238.515 285.085 238.845 ;
        RECT 284.755 237.155 285.085 237.485 ;
        RECT 284.76 237.155 285.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 -0.845 285.085 -0.515 ;
        RECT 284.755 -2.205 285.085 -1.875 ;
        RECT 284.755 -3.565 285.085 -3.235 ;
        RECT 284.76 -3.565 285.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 -123.245 285.085 -122.915 ;
        RECT 284.755 -124.605 285.085 -124.275 ;
        RECT 284.755 -125.965 285.085 -125.635 ;
        RECT 284.755 -127.325 285.085 -126.995 ;
        RECT 284.755 -128.685 285.085 -128.355 ;
        RECT 284.755 -130.045 285.085 -129.715 ;
        RECT 284.755 -131.405 285.085 -131.075 ;
        RECT 284.755 -132.765 285.085 -132.435 ;
        RECT 284.755 -134.125 285.085 -133.795 ;
        RECT 284.755 -135.485 285.085 -135.155 ;
        RECT 284.755 -136.845 285.085 -136.515 ;
        RECT 284.755 -138.205 285.085 -137.875 ;
        RECT 284.755 -139.565 285.085 -139.235 ;
        RECT 284.755 -140.925 285.085 -140.595 ;
        RECT 284.755 -142.285 285.085 -141.955 ;
        RECT 284.755 -143.645 285.085 -143.315 ;
        RECT 284.755 -145.005 285.085 -144.675 ;
        RECT 284.755 -146.365 285.085 -146.035 ;
        RECT 284.755 -147.725 285.085 -147.395 ;
        RECT 284.755 -149.085 285.085 -148.755 ;
        RECT 284.755 -150.445 285.085 -150.115 ;
        RECT 284.755 -151.805 285.085 -151.475 ;
        RECT 284.755 -153.165 285.085 -152.835 ;
        RECT 284.755 -154.525 285.085 -154.195 ;
        RECT 284.755 -155.885 285.085 -155.555 ;
        RECT 284.755 -157.245 285.085 -156.915 ;
        RECT 284.755 -158.605 285.085 -158.275 ;
        RECT 284.755 -159.965 285.085 -159.635 ;
        RECT 284.755 -161.325 285.085 -160.995 ;
        RECT 284.755 -162.685 285.085 -162.355 ;
        RECT 284.755 -164.045 285.085 -163.715 ;
        RECT 284.755 -165.405 285.085 -165.075 ;
        RECT 284.755 -166.765 285.085 -166.435 ;
        RECT 284.755 -168.125 285.085 -167.795 ;
        RECT 284.755 -169.485 285.085 -169.155 ;
        RECT 284.755 -170.845 285.085 -170.515 ;
        RECT 284.755 -172.205 285.085 -171.875 ;
        RECT 284.755 -173.565 285.085 -173.235 ;
        RECT 284.755 -174.925 285.085 -174.595 ;
        RECT 284.755 -176.285 285.085 -175.955 ;
        RECT 284.755 -177.645 285.085 -177.315 ;
        RECT 284.755 -179.005 285.085 -178.675 ;
        RECT 284.755 -180.365 285.085 -180.035 ;
        RECT 284.755 -181.725 285.085 -181.395 ;
        RECT 284.755 -183.085 285.085 -182.755 ;
        RECT 284.755 -184.445 285.085 -184.115 ;
        RECT 284.755 -185.805 285.085 -185.475 ;
        RECT 284.755 -187.165 285.085 -186.835 ;
        RECT 284.755 -188.525 285.085 -188.195 ;
        RECT 284.755 -189.885 285.085 -189.555 ;
        RECT 284.755 -191.245 285.085 -190.915 ;
        RECT 284.755 -192.605 285.085 -192.275 ;
        RECT 284.755 -193.965 285.085 -193.635 ;
        RECT 284.755 -195.325 285.085 -194.995 ;
        RECT 284.755 -196.685 285.085 -196.355 ;
        RECT 284.755 -198.045 285.085 -197.715 ;
        RECT 284.755 -199.405 285.085 -199.075 ;
        RECT 284.755 -200.765 285.085 -200.435 ;
        RECT 284.755 -202.125 285.085 -201.795 ;
        RECT 284.755 -203.485 285.085 -203.155 ;
        RECT 284.755 -204.845 285.085 -204.515 ;
        RECT 284.755 -206.205 285.085 -205.875 ;
        RECT 284.755 -207.565 285.085 -207.235 ;
        RECT 284.755 -208.925 285.085 -208.595 ;
        RECT 284.755 -210.285 285.085 -209.955 ;
        RECT 284.755 -211.645 285.085 -211.315 ;
        RECT 284.755 -213.005 285.085 -212.675 ;
        RECT 284.755 -214.365 285.085 -214.035 ;
        RECT 284.755 -215.725 285.085 -215.395 ;
        RECT 284.755 -217.085 285.085 -216.755 ;
        RECT 284.755 -218.445 285.085 -218.115 ;
        RECT 284.755 -219.805 285.085 -219.475 ;
        RECT 284.755 -221.165 285.085 -220.835 ;
        RECT 284.755 -222.525 285.085 -222.195 ;
        RECT 284.755 -223.885 285.085 -223.555 ;
        RECT 284.755 -225.245 285.085 -224.915 ;
        RECT 284.755 -226.605 285.085 -226.275 ;
        RECT 284.755 -227.965 285.085 -227.635 ;
        RECT 284.755 -229.325 285.085 -228.995 ;
        RECT 284.755 -230.685 285.085 -230.355 ;
        RECT 284.755 -232.045 285.085 -231.715 ;
        RECT 284.755 -233.405 285.085 -233.075 ;
        RECT 284.755 -234.765 285.085 -234.435 ;
        RECT 284.755 -236.125 285.085 -235.795 ;
        RECT 284.755 -237.485 285.085 -237.155 ;
        RECT 284.755 -238.845 285.085 -238.515 ;
        RECT 284.755 -241.09 285.085 -239.96 ;
        RECT 284.76 -241.205 285.08 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 244.04 286.445 245.17 ;
        RECT 286.115 242.595 286.445 242.925 ;
        RECT 286.115 241.235 286.445 241.565 ;
        RECT 286.115 239.875 286.445 240.205 ;
        RECT 286.115 238.515 286.445 238.845 ;
        RECT 286.115 237.155 286.445 237.485 ;
        RECT 286.12 237.155 286.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 -127.325 286.445 -126.995 ;
        RECT 286.115 -128.685 286.445 -128.355 ;
        RECT 286.115 -130.045 286.445 -129.715 ;
        RECT 286.115 -131.405 286.445 -131.075 ;
        RECT 286.115 -132.765 286.445 -132.435 ;
        RECT 286.115 -134.125 286.445 -133.795 ;
        RECT 286.115 -135.485 286.445 -135.155 ;
        RECT 286.115 -136.845 286.445 -136.515 ;
        RECT 286.115 -138.205 286.445 -137.875 ;
        RECT 286.115 -139.565 286.445 -139.235 ;
        RECT 286.115 -140.925 286.445 -140.595 ;
        RECT 286.115 -142.285 286.445 -141.955 ;
        RECT 286.115 -143.645 286.445 -143.315 ;
        RECT 286.115 -145.005 286.445 -144.675 ;
        RECT 286.115 -146.365 286.445 -146.035 ;
        RECT 286.115 -147.725 286.445 -147.395 ;
        RECT 286.115 -149.085 286.445 -148.755 ;
        RECT 286.115 -150.445 286.445 -150.115 ;
        RECT 286.115 -151.805 286.445 -151.475 ;
        RECT 286.115 -153.165 286.445 -152.835 ;
        RECT 286.115 -154.525 286.445 -154.195 ;
        RECT 286.115 -155.885 286.445 -155.555 ;
        RECT 286.115 -157.245 286.445 -156.915 ;
        RECT 286.115 -158.605 286.445 -158.275 ;
        RECT 286.115 -159.965 286.445 -159.635 ;
        RECT 286.115 -161.325 286.445 -160.995 ;
        RECT 286.115 -162.685 286.445 -162.355 ;
        RECT 286.115 -164.045 286.445 -163.715 ;
        RECT 286.115 -165.405 286.445 -165.075 ;
        RECT 286.115 -166.765 286.445 -166.435 ;
        RECT 286.115 -168.125 286.445 -167.795 ;
        RECT 286.115 -169.485 286.445 -169.155 ;
        RECT 286.115 -170.845 286.445 -170.515 ;
        RECT 286.115 -172.205 286.445 -171.875 ;
        RECT 286.115 -173.565 286.445 -173.235 ;
        RECT 286.115 -174.925 286.445 -174.595 ;
        RECT 286.115 -176.285 286.445 -175.955 ;
        RECT 286.115 -177.645 286.445 -177.315 ;
        RECT 286.115 -179.005 286.445 -178.675 ;
        RECT 286.115 -180.365 286.445 -180.035 ;
        RECT 286.115 -181.725 286.445 -181.395 ;
        RECT 286.115 -183.085 286.445 -182.755 ;
        RECT 286.115 -184.445 286.445 -184.115 ;
        RECT 286.115 -185.805 286.445 -185.475 ;
        RECT 286.115 -187.165 286.445 -186.835 ;
        RECT 286.115 -188.525 286.445 -188.195 ;
        RECT 286.115 -189.885 286.445 -189.555 ;
        RECT 286.115 -191.245 286.445 -190.915 ;
        RECT 286.115 -192.605 286.445 -192.275 ;
        RECT 286.115 -193.965 286.445 -193.635 ;
        RECT 286.115 -195.325 286.445 -194.995 ;
        RECT 286.115 -196.685 286.445 -196.355 ;
        RECT 286.115 -198.045 286.445 -197.715 ;
        RECT 286.115 -199.405 286.445 -199.075 ;
        RECT 286.115 -200.765 286.445 -200.435 ;
        RECT 286.115 -202.125 286.445 -201.795 ;
        RECT 286.115 -203.485 286.445 -203.155 ;
        RECT 286.115 -204.845 286.445 -204.515 ;
        RECT 286.115 -206.205 286.445 -205.875 ;
        RECT 286.115 -207.565 286.445 -207.235 ;
        RECT 286.115 -208.925 286.445 -208.595 ;
        RECT 286.115 -210.285 286.445 -209.955 ;
        RECT 286.115 -211.645 286.445 -211.315 ;
        RECT 286.115 -213.005 286.445 -212.675 ;
        RECT 286.115 -214.365 286.445 -214.035 ;
        RECT 286.115 -215.725 286.445 -215.395 ;
        RECT 286.115 -217.085 286.445 -216.755 ;
        RECT 286.115 -218.445 286.445 -218.115 ;
        RECT 286.115 -219.805 286.445 -219.475 ;
        RECT 286.115 -221.165 286.445 -220.835 ;
        RECT 286.115 -222.525 286.445 -222.195 ;
        RECT 286.115 -223.885 286.445 -223.555 ;
        RECT 286.115 -225.245 286.445 -224.915 ;
        RECT 286.115 -226.605 286.445 -226.275 ;
        RECT 286.115 -227.965 286.445 -227.635 ;
        RECT 286.115 -229.325 286.445 -228.995 ;
        RECT 286.115 -230.685 286.445 -230.355 ;
        RECT 286.115 -232.045 286.445 -231.715 ;
        RECT 286.115 -233.405 286.445 -233.075 ;
        RECT 286.115 -234.765 286.445 -234.435 ;
        RECT 286.115 -236.125 286.445 -235.795 ;
        RECT 286.115 -237.485 286.445 -237.155 ;
        RECT 286.115 -238.845 286.445 -238.515 ;
        RECT 286.115 -241.09 286.445 -239.96 ;
        RECT 286.12 -241.205 286.44 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.71 -125.535 287.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 244.04 287.805 245.17 ;
        RECT 287.475 242.595 287.805 242.925 ;
        RECT 287.475 241.235 287.805 241.565 ;
        RECT 287.475 239.875 287.805 240.205 ;
        RECT 287.475 238.515 287.805 238.845 ;
        RECT 287.475 237.155 287.805 237.485 ;
        RECT 287.48 237.155 287.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 -0.845 287.805 -0.515 ;
        RECT 287.475 -2.205 287.805 -1.875 ;
        RECT 287.475 -3.565 287.805 -3.235 ;
        RECT 287.48 -3.565 287.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 244.04 289.165 245.17 ;
        RECT 288.835 242.595 289.165 242.925 ;
        RECT 288.835 241.235 289.165 241.565 ;
        RECT 288.835 239.875 289.165 240.205 ;
        RECT 288.835 238.515 289.165 238.845 ;
        RECT 288.835 237.155 289.165 237.485 ;
        RECT 288.84 237.155 289.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 -0.845 289.165 -0.515 ;
        RECT 288.835 -2.205 289.165 -1.875 ;
        RECT 288.835 -3.565 289.165 -3.235 ;
        RECT 288.84 -3.565 289.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 244.04 290.525 245.17 ;
        RECT 290.195 242.595 290.525 242.925 ;
        RECT 290.195 241.235 290.525 241.565 ;
        RECT 290.195 239.875 290.525 240.205 ;
        RECT 290.195 238.515 290.525 238.845 ;
        RECT 290.195 237.155 290.525 237.485 ;
        RECT 290.2 237.155 290.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 -0.845 290.525 -0.515 ;
        RECT 290.195 -2.205 290.525 -1.875 ;
        RECT 290.195 -3.565 290.525 -3.235 ;
        RECT 290.2 -3.565 290.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 -180.365 290.525 -180.035 ;
        RECT 290.195 -181.725 290.525 -181.395 ;
        RECT 290.195 -183.085 290.525 -182.755 ;
        RECT 290.195 -184.445 290.525 -184.115 ;
        RECT 290.195 -185.805 290.525 -185.475 ;
        RECT 290.195 -187.165 290.525 -186.835 ;
        RECT 290.195 -188.525 290.525 -188.195 ;
        RECT 290.195 -189.885 290.525 -189.555 ;
        RECT 290.195 -191.245 290.525 -190.915 ;
        RECT 290.195 -192.605 290.525 -192.275 ;
        RECT 290.195 -193.965 290.525 -193.635 ;
        RECT 290.195 -195.325 290.525 -194.995 ;
        RECT 290.195 -196.685 290.525 -196.355 ;
        RECT 290.195 -198.045 290.525 -197.715 ;
        RECT 290.195 -199.405 290.525 -199.075 ;
        RECT 290.195 -200.765 290.525 -200.435 ;
        RECT 290.195 -202.125 290.525 -201.795 ;
        RECT 290.195 -203.485 290.525 -203.155 ;
        RECT 290.195 -204.845 290.525 -204.515 ;
        RECT 290.195 -206.205 290.525 -205.875 ;
        RECT 290.195 -207.565 290.525 -207.235 ;
        RECT 290.195 -208.925 290.525 -208.595 ;
        RECT 290.195 -210.285 290.525 -209.955 ;
        RECT 290.195 -211.645 290.525 -211.315 ;
        RECT 290.195 -213.005 290.525 -212.675 ;
        RECT 290.195 -214.365 290.525 -214.035 ;
        RECT 290.195 -215.725 290.525 -215.395 ;
        RECT 290.195 -217.085 290.525 -216.755 ;
        RECT 290.195 -218.445 290.525 -218.115 ;
        RECT 290.195 -219.805 290.525 -219.475 ;
        RECT 290.195 -221.165 290.525 -220.835 ;
        RECT 290.195 -222.525 290.525 -222.195 ;
        RECT 290.195 -223.885 290.525 -223.555 ;
        RECT 290.195 -225.245 290.525 -224.915 ;
        RECT 290.195 -226.605 290.525 -226.275 ;
        RECT 290.195 -227.965 290.525 -227.635 ;
        RECT 290.195 -229.325 290.525 -228.995 ;
        RECT 290.195 -230.685 290.525 -230.355 ;
        RECT 290.195 -232.045 290.525 -231.715 ;
        RECT 290.195 -233.405 290.525 -233.075 ;
        RECT 290.195 -234.765 290.525 -234.435 ;
        RECT 290.195 -236.125 290.525 -235.795 ;
        RECT 290.195 -237.485 290.525 -237.155 ;
        RECT 290.195 -238.845 290.525 -238.515 ;
        RECT 290.195 -241.09 290.525 -239.96 ;
        RECT 290.2 -241.205 290.52 -122.24 ;
        RECT 290.195 -123.245 290.525 -122.915 ;
        RECT 290.195 -124.605 290.525 -124.275 ;
        RECT 290.195 -125.965 290.525 -125.635 ;
        RECT 290.195 -127.325 290.525 -126.995 ;
        RECT 290.195 -128.685 290.525 -128.355 ;
        RECT 290.195 -130.045 290.525 -129.715 ;
        RECT 290.195 -131.405 290.525 -131.075 ;
        RECT 290.195 -132.765 290.525 -132.435 ;
        RECT 290.195 -134.125 290.525 -133.795 ;
        RECT 290.195 -135.485 290.525 -135.155 ;
        RECT 290.195 -136.845 290.525 -136.515 ;
        RECT 290.195 -138.205 290.525 -137.875 ;
        RECT 290.195 -139.565 290.525 -139.235 ;
        RECT 290.195 -140.925 290.525 -140.595 ;
        RECT 290.195 -142.285 290.525 -141.955 ;
        RECT 290.195 -143.645 290.525 -143.315 ;
        RECT 290.195 -145.005 290.525 -144.675 ;
        RECT 290.195 -146.365 290.525 -146.035 ;
        RECT 290.195 -147.725 290.525 -147.395 ;
        RECT 290.195 -149.085 290.525 -148.755 ;
        RECT 290.195 -150.445 290.525 -150.115 ;
        RECT 290.195 -151.805 290.525 -151.475 ;
        RECT 290.195 -153.165 290.525 -152.835 ;
        RECT 290.195 -154.525 290.525 -154.195 ;
        RECT 290.195 -155.885 290.525 -155.555 ;
        RECT 290.195 -157.245 290.525 -156.915 ;
        RECT 290.195 -158.605 290.525 -158.275 ;
        RECT 290.195 -159.965 290.525 -159.635 ;
        RECT 290.195 -161.325 290.525 -160.995 ;
        RECT 290.195 -162.685 290.525 -162.355 ;
        RECT 290.195 -164.045 290.525 -163.715 ;
        RECT 290.195 -165.405 290.525 -165.075 ;
        RECT 290.195 -166.765 290.525 -166.435 ;
        RECT 290.195 -168.125 290.525 -167.795 ;
        RECT 290.195 -169.485 290.525 -169.155 ;
        RECT 290.195 -170.845 290.525 -170.515 ;
        RECT 290.195 -172.205 290.525 -171.875 ;
        RECT 290.195 -173.565 290.525 -173.235 ;
        RECT 290.195 -174.925 290.525 -174.595 ;
        RECT 290.195 -176.285 290.525 -175.955 ;
        RECT 290.195 -177.645 290.525 -177.315 ;
        RECT 290.195 -179.005 290.525 -178.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.475 -127.325 253.805 -126.995 ;
        RECT 253.475 -128.685 253.805 -128.355 ;
        RECT 253.475 -130.045 253.805 -129.715 ;
        RECT 253.475 -131.405 253.805 -131.075 ;
        RECT 253.475 -132.765 253.805 -132.435 ;
        RECT 253.475 -134.125 253.805 -133.795 ;
        RECT 253.475 -135.485 253.805 -135.155 ;
        RECT 253.475 -136.845 253.805 -136.515 ;
        RECT 253.475 -138.205 253.805 -137.875 ;
        RECT 253.475 -139.565 253.805 -139.235 ;
        RECT 253.475 -140.925 253.805 -140.595 ;
        RECT 253.475 -142.285 253.805 -141.955 ;
        RECT 253.475 -143.645 253.805 -143.315 ;
        RECT 253.475 -145.005 253.805 -144.675 ;
        RECT 253.475 -146.365 253.805 -146.035 ;
        RECT 253.475 -147.725 253.805 -147.395 ;
        RECT 253.475 -149.085 253.805 -148.755 ;
        RECT 253.475 -150.445 253.805 -150.115 ;
        RECT 253.475 -151.805 253.805 -151.475 ;
        RECT 253.475 -153.165 253.805 -152.835 ;
        RECT 253.475 -154.525 253.805 -154.195 ;
        RECT 253.475 -155.885 253.805 -155.555 ;
        RECT 253.475 -157.245 253.805 -156.915 ;
        RECT 253.475 -158.605 253.805 -158.275 ;
        RECT 253.475 -159.965 253.805 -159.635 ;
        RECT 253.475 -161.325 253.805 -160.995 ;
        RECT 253.475 -162.685 253.805 -162.355 ;
        RECT 253.475 -164.045 253.805 -163.715 ;
        RECT 253.475 -165.405 253.805 -165.075 ;
        RECT 253.475 -166.765 253.805 -166.435 ;
        RECT 253.475 -168.125 253.805 -167.795 ;
        RECT 253.475 -169.485 253.805 -169.155 ;
        RECT 253.475 -170.845 253.805 -170.515 ;
        RECT 253.475 -172.205 253.805 -171.875 ;
        RECT 253.475 -173.565 253.805 -173.235 ;
        RECT 253.475 -174.925 253.805 -174.595 ;
        RECT 253.475 -176.285 253.805 -175.955 ;
        RECT 253.475 -177.645 253.805 -177.315 ;
        RECT 253.475 -179.005 253.805 -178.675 ;
        RECT 253.475 -180.365 253.805 -180.035 ;
        RECT 253.475 -181.725 253.805 -181.395 ;
        RECT 253.475 -183.085 253.805 -182.755 ;
        RECT 253.475 -184.445 253.805 -184.115 ;
        RECT 253.475 -185.805 253.805 -185.475 ;
        RECT 253.475 -187.165 253.805 -186.835 ;
        RECT 253.475 -188.525 253.805 -188.195 ;
        RECT 253.475 -189.885 253.805 -189.555 ;
        RECT 253.475 -191.245 253.805 -190.915 ;
        RECT 253.475 -192.605 253.805 -192.275 ;
        RECT 253.475 -193.965 253.805 -193.635 ;
        RECT 253.475 -195.325 253.805 -194.995 ;
        RECT 253.475 -196.685 253.805 -196.355 ;
        RECT 253.475 -198.045 253.805 -197.715 ;
        RECT 253.475 -199.405 253.805 -199.075 ;
        RECT 253.475 -200.765 253.805 -200.435 ;
        RECT 253.475 -202.125 253.805 -201.795 ;
        RECT 253.475 -203.485 253.805 -203.155 ;
        RECT 253.475 -204.845 253.805 -204.515 ;
        RECT 253.475 -206.205 253.805 -205.875 ;
        RECT 253.475 -207.565 253.805 -207.235 ;
        RECT 253.475 -208.925 253.805 -208.595 ;
        RECT 253.475 -210.285 253.805 -209.955 ;
        RECT 253.475 -211.645 253.805 -211.315 ;
        RECT 253.475 -213.005 253.805 -212.675 ;
        RECT 253.475 -214.365 253.805 -214.035 ;
        RECT 253.475 -215.725 253.805 -215.395 ;
        RECT 253.475 -217.085 253.805 -216.755 ;
        RECT 253.475 -218.445 253.805 -218.115 ;
        RECT 253.475 -219.805 253.805 -219.475 ;
        RECT 253.475 -221.165 253.805 -220.835 ;
        RECT 253.475 -222.525 253.805 -222.195 ;
        RECT 253.475 -223.885 253.805 -223.555 ;
        RECT 253.475 -225.245 253.805 -224.915 ;
        RECT 253.475 -226.605 253.805 -226.275 ;
        RECT 253.475 -227.965 253.805 -227.635 ;
        RECT 253.475 -229.325 253.805 -228.995 ;
        RECT 253.475 -230.685 253.805 -230.355 ;
        RECT 253.475 -232.045 253.805 -231.715 ;
        RECT 253.475 -233.405 253.805 -233.075 ;
        RECT 253.475 -234.765 253.805 -234.435 ;
        RECT 253.475 -236.125 253.805 -235.795 ;
        RECT 253.475 -237.485 253.805 -237.155 ;
        RECT 253.475 -238.845 253.805 -238.515 ;
        RECT 253.475 -241.09 253.805 -239.96 ;
        RECT 253.48 -241.205 253.8 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.01 -125.535 254.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 244.04 255.165 245.17 ;
        RECT 254.835 242.595 255.165 242.925 ;
        RECT 254.835 241.235 255.165 241.565 ;
        RECT 254.835 239.875 255.165 240.205 ;
        RECT 254.835 238.515 255.165 238.845 ;
        RECT 254.835 237.155 255.165 237.485 ;
        RECT 254.84 237.155 255.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 -0.845 255.165 -0.515 ;
        RECT 254.835 -2.205 255.165 -1.875 ;
        RECT 254.835 -3.565 255.165 -3.235 ;
        RECT 254.84 -3.565 255.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 244.04 256.525 245.17 ;
        RECT 256.195 242.595 256.525 242.925 ;
        RECT 256.195 241.235 256.525 241.565 ;
        RECT 256.195 239.875 256.525 240.205 ;
        RECT 256.195 238.515 256.525 238.845 ;
        RECT 256.195 237.155 256.525 237.485 ;
        RECT 256.2 237.155 256.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 -0.845 256.525 -0.515 ;
        RECT 256.195 -2.205 256.525 -1.875 ;
        RECT 256.195 -3.565 256.525 -3.235 ;
        RECT 256.2 -3.565 256.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 244.04 257.885 245.17 ;
        RECT 257.555 242.595 257.885 242.925 ;
        RECT 257.555 241.235 257.885 241.565 ;
        RECT 257.555 239.875 257.885 240.205 ;
        RECT 257.555 238.515 257.885 238.845 ;
        RECT 257.555 237.155 257.885 237.485 ;
        RECT 257.56 237.155 257.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 -0.845 257.885 -0.515 ;
        RECT 257.555 -2.205 257.885 -1.875 ;
        RECT 257.555 -3.565 257.885 -3.235 ;
        RECT 257.56 -3.565 257.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 -123.245 257.885 -122.915 ;
        RECT 257.555 -124.605 257.885 -124.275 ;
        RECT 257.555 -125.965 257.885 -125.635 ;
        RECT 257.555 -127.325 257.885 -126.995 ;
        RECT 257.555 -128.685 257.885 -128.355 ;
        RECT 257.555 -130.045 257.885 -129.715 ;
        RECT 257.555 -131.405 257.885 -131.075 ;
        RECT 257.555 -132.765 257.885 -132.435 ;
        RECT 257.555 -134.125 257.885 -133.795 ;
        RECT 257.555 -135.485 257.885 -135.155 ;
        RECT 257.555 -136.845 257.885 -136.515 ;
        RECT 257.555 -138.205 257.885 -137.875 ;
        RECT 257.555 -139.565 257.885 -139.235 ;
        RECT 257.555 -140.925 257.885 -140.595 ;
        RECT 257.555 -142.285 257.885 -141.955 ;
        RECT 257.555 -143.645 257.885 -143.315 ;
        RECT 257.555 -145.005 257.885 -144.675 ;
        RECT 257.555 -146.365 257.885 -146.035 ;
        RECT 257.555 -147.725 257.885 -147.395 ;
        RECT 257.555 -149.085 257.885 -148.755 ;
        RECT 257.555 -150.445 257.885 -150.115 ;
        RECT 257.555 -151.805 257.885 -151.475 ;
        RECT 257.555 -153.165 257.885 -152.835 ;
        RECT 257.555 -154.525 257.885 -154.195 ;
        RECT 257.555 -155.885 257.885 -155.555 ;
        RECT 257.555 -157.245 257.885 -156.915 ;
        RECT 257.555 -158.605 257.885 -158.275 ;
        RECT 257.555 -159.965 257.885 -159.635 ;
        RECT 257.555 -161.325 257.885 -160.995 ;
        RECT 257.555 -162.685 257.885 -162.355 ;
        RECT 257.555 -164.045 257.885 -163.715 ;
        RECT 257.555 -165.405 257.885 -165.075 ;
        RECT 257.555 -166.765 257.885 -166.435 ;
        RECT 257.555 -168.125 257.885 -167.795 ;
        RECT 257.555 -169.485 257.885 -169.155 ;
        RECT 257.555 -170.845 257.885 -170.515 ;
        RECT 257.555 -172.205 257.885 -171.875 ;
        RECT 257.555 -173.565 257.885 -173.235 ;
        RECT 257.555 -174.925 257.885 -174.595 ;
        RECT 257.555 -176.285 257.885 -175.955 ;
        RECT 257.555 -177.645 257.885 -177.315 ;
        RECT 257.555 -179.005 257.885 -178.675 ;
        RECT 257.555 -180.365 257.885 -180.035 ;
        RECT 257.555 -181.725 257.885 -181.395 ;
        RECT 257.555 -183.085 257.885 -182.755 ;
        RECT 257.555 -184.445 257.885 -184.115 ;
        RECT 257.555 -185.805 257.885 -185.475 ;
        RECT 257.555 -187.165 257.885 -186.835 ;
        RECT 257.555 -188.525 257.885 -188.195 ;
        RECT 257.555 -189.885 257.885 -189.555 ;
        RECT 257.555 -191.245 257.885 -190.915 ;
        RECT 257.555 -192.605 257.885 -192.275 ;
        RECT 257.555 -193.965 257.885 -193.635 ;
        RECT 257.555 -195.325 257.885 -194.995 ;
        RECT 257.555 -196.685 257.885 -196.355 ;
        RECT 257.555 -198.045 257.885 -197.715 ;
        RECT 257.555 -199.405 257.885 -199.075 ;
        RECT 257.555 -200.765 257.885 -200.435 ;
        RECT 257.555 -202.125 257.885 -201.795 ;
        RECT 257.555 -203.485 257.885 -203.155 ;
        RECT 257.555 -204.845 257.885 -204.515 ;
        RECT 257.555 -206.205 257.885 -205.875 ;
        RECT 257.555 -207.565 257.885 -207.235 ;
        RECT 257.555 -208.925 257.885 -208.595 ;
        RECT 257.555 -210.285 257.885 -209.955 ;
        RECT 257.555 -211.645 257.885 -211.315 ;
        RECT 257.555 -213.005 257.885 -212.675 ;
        RECT 257.555 -214.365 257.885 -214.035 ;
        RECT 257.555 -215.725 257.885 -215.395 ;
        RECT 257.555 -217.085 257.885 -216.755 ;
        RECT 257.555 -218.445 257.885 -218.115 ;
        RECT 257.555 -219.805 257.885 -219.475 ;
        RECT 257.555 -221.165 257.885 -220.835 ;
        RECT 257.555 -222.525 257.885 -222.195 ;
        RECT 257.555 -223.885 257.885 -223.555 ;
        RECT 257.555 -225.245 257.885 -224.915 ;
        RECT 257.555 -226.605 257.885 -226.275 ;
        RECT 257.555 -227.965 257.885 -227.635 ;
        RECT 257.555 -229.325 257.885 -228.995 ;
        RECT 257.555 -230.685 257.885 -230.355 ;
        RECT 257.555 -232.045 257.885 -231.715 ;
        RECT 257.555 -233.405 257.885 -233.075 ;
        RECT 257.555 -234.765 257.885 -234.435 ;
        RECT 257.555 -236.125 257.885 -235.795 ;
        RECT 257.555 -237.485 257.885 -237.155 ;
        RECT 257.555 -238.845 257.885 -238.515 ;
        RECT 257.555 -241.09 257.885 -239.96 ;
        RECT 257.56 -241.205 257.88 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 244.04 259.245 245.17 ;
        RECT 258.915 242.595 259.245 242.925 ;
        RECT 258.915 241.235 259.245 241.565 ;
        RECT 258.915 239.875 259.245 240.205 ;
        RECT 258.915 238.515 259.245 238.845 ;
        RECT 258.915 237.155 259.245 237.485 ;
        RECT 258.92 237.155 259.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 -0.845 259.245 -0.515 ;
        RECT 258.915 -2.205 259.245 -1.875 ;
        RECT 258.915 -3.565 259.245 -3.235 ;
        RECT 258.92 -3.565 259.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 -123.245 259.245 -122.915 ;
        RECT 258.915 -124.605 259.245 -124.275 ;
        RECT 258.915 -125.965 259.245 -125.635 ;
        RECT 258.915 -127.325 259.245 -126.995 ;
        RECT 258.915 -128.685 259.245 -128.355 ;
        RECT 258.915 -130.045 259.245 -129.715 ;
        RECT 258.915 -131.405 259.245 -131.075 ;
        RECT 258.915 -132.765 259.245 -132.435 ;
        RECT 258.915 -134.125 259.245 -133.795 ;
        RECT 258.915 -135.485 259.245 -135.155 ;
        RECT 258.915 -136.845 259.245 -136.515 ;
        RECT 258.915 -138.205 259.245 -137.875 ;
        RECT 258.915 -139.565 259.245 -139.235 ;
        RECT 258.915 -140.925 259.245 -140.595 ;
        RECT 258.915 -142.285 259.245 -141.955 ;
        RECT 258.915 -143.645 259.245 -143.315 ;
        RECT 258.915 -145.005 259.245 -144.675 ;
        RECT 258.915 -146.365 259.245 -146.035 ;
        RECT 258.915 -147.725 259.245 -147.395 ;
        RECT 258.915 -149.085 259.245 -148.755 ;
        RECT 258.915 -150.445 259.245 -150.115 ;
        RECT 258.915 -151.805 259.245 -151.475 ;
        RECT 258.915 -153.165 259.245 -152.835 ;
        RECT 258.915 -154.525 259.245 -154.195 ;
        RECT 258.915 -155.885 259.245 -155.555 ;
        RECT 258.915 -157.245 259.245 -156.915 ;
        RECT 258.915 -158.605 259.245 -158.275 ;
        RECT 258.915 -159.965 259.245 -159.635 ;
        RECT 258.915 -161.325 259.245 -160.995 ;
        RECT 258.915 -162.685 259.245 -162.355 ;
        RECT 258.915 -164.045 259.245 -163.715 ;
        RECT 258.915 -165.405 259.245 -165.075 ;
        RECT 258.915 -166.765 259.245 -166.435 ;
        RECT 258.915 -168.125 259.245 -167.795 ;
        RECT 258.915 -169.485 259.245 -169.155 ;
        RECT 258.915 -170.845 259.245 -170.515 ;
        RECT 258.915 -172.205 259.245 -171.875 ;
        RECT 258.915 -173.565 259.245 -173.235 ;
        RECT 258.915 -174.925 259.245 -174.595 ;
        RECT 258.915 -176.285 259.245 -175.955 ;
        RECT 258.915 -177.645 259.245 -177.315 ;
        RECT 258.915 -179.005 259.245 -178.675 ;
        RECT 258.915 -180.365 259.245 -180.035 ;
        RECT 258.915 -181.725 259.245 -181.395 ;
        RECT 258.915 -183.085 259.245 -182.755 ;
        RECT 258.915 -184.445 259.245 -184.115 ;
        RECT 258.915 -185.805 259.245 -185.475 ;
        RECT 258.915 -187.165 259.245 -186.835 ;
        RECT 258.915 -188.525 259.245 -188.195 ;
        RECT 258.915 -189.885 259.245 -189.555 ;
        RECT 258.915 -191.245 259.245 -190.915 ;
        RECT 258.915 -192.605 259.245 -192.275 ;
        RECT 258.915 -193.965 259.245 -193.635 ;
        RECT 258.915 -195.325 259.245 -194.995 ;
        RECT 258.915 -196.685 259.245 -196.355 ;
        RECT 258.915 -198.045 259.245 -197.715 ;
        RECT 258.915 -199.405 259.245 -199.075 ;
        RECT 258.915 -200.765 259.245 -200.435 ;
        RECT 258.915 -202.125 259.245 -201.795 ;
        RECT 258.915 -203.485 259.245 -203.155 ;
        RECT 258.915 -204.845 259.245 -204.515 ;
        RECT 258.915 -206.205 259.245 -205.875 ;
        RECT 258.915 -207.565 259.245 -207.235 ;
        RECT 258.915 -208.925 259.245 -208.595 ;
        RECT 258.915 -210.285 259.245 -209.955 ;
        RECT 258.915 -211.645 259.245 -211.315 ;
        RECT 258.915 -213.005 259.245 -212.675 ;
        RECT 258.915 -214.365 259.245 -214.035 ;
        RECT 258.915 -215.725 259.245 -215.395 ;
        RECT 258.915 -217.085 259.245 -216.755 ;
        RECT 258.915 -218.445 259.245 -218.115 ;
        RECT 258.915 -219.805 259.245 -219.475 ;
        RECT 258.915 -221.165 259.245 -220.835 ;
        RECT 258.915 -222.525 259.245 -222.195 ;
        RECT 258.915 -223.885 259.245 -223.555 ;
        RECT 258.915 -225.245 259.245 -224.915 ;
        RECT 258.915 -226.605 259.245 -226.275 ;
        RECT 258.915 -227.965 259.245 -227.635 ;
        RECT 258.915 -229.325 259.245 -228.995 ;
        RECT 258.915 -230.685 259.245 -230.355 ;
        RECT 258.915 -232.045 259.245 -231.715 ;
        RECT 258.915 -233.405 259.245 -233.075 ;
        RECT 258.915 -234.765 259.245 -234.435 ;
        RECT 258.915 -236.125 259.245 -235.795 ;
        RECT 258.915 -237.485 259.245 -237.155 ;
        RECT 258.915 -238.845 259.245 -238.515 ;
        RECT 258.915 -241.09 259.245 -239.96 ;
        RECT 258.92 -241.205 259.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 244.04 260.605 245.17 ;
        RECT 260.275 242.595 260.605 242.925 ;
        RECT 260.275 241.235 260.605 241.565 ;
        RECT 260.275 239.875 260.605 240.205 ;
        RECT 260.275 238.515 260.605 238.845 ;
        RECT 260.275 237.155 260.605 237.485 ;
        RECT 260.28 237.155 260.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 -0.845 260.605 -0.515 ;
        RECT 260.275 -2.205 260.605 -1.875 ;
        RECT 260.275 -3.565 260.605 -3.235 ;
        RECT 260.28 -3.565 260.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 -123.245 260.605 -122.915 ;
        RECT 260.275 -124.605 260.605 -124.275 ;
        RECT 260.275 -125.965 260.605 -125.635 ;
        RECT 260.275 -127.325 260.605 -126.995 ;
        RECT 260.275 -128.685 260.605 -128.355 ;
        RECT 260.275 -130.045 260.605 -129.715 ;
        RECT 260.275 -131.405 260.605 -131.075 ;
        RECT 260.275 -132.765 260.605 -132.435 ;
        RECT 260.275 -134.125 260.605 -133.795 ;
        RECT 260.275 -135.485 260.605 -135.155 ;
        RECT 260.275 -136.845 260.605 -136.515 ;
        RECT 260.275 -138.205 260.605 -137.875 ;
        RECT 260.275 -139.565 260.605 -139.235 ;
        RECT 260.275 -140.925 260.605 -140.595 ;
        RECT 260.275 -142.285 260.605 -141.955 ;
        RECT 260.275 -143.645 260.605 -143.315 ;
        RECT 260.275 -145.005 260.605 -144.675 ;
        RECT 260.275 -146.365 260.605 -146.035 ;
        RECT 260.275 -147.725 260.605 -147.395 ;
        RECT 260.275 -149.085 260.605 -148.755 ;
        RECT 260.275 -150.445 260.605 -150.115 ;
        RECT 260.275 -151.805 260.605 -151.475 ;
        RECT 260.275 -153.165 260.605 -152.835 ;
        RECT 260.275 -154.525 260.605 -154.195 ;
        RECT 260.275 -155.885 260.605 -155.555 ;
        RECT 260.275 -157.245 260.605 -156.915 ;
        RECT 260.275 -158.605 260.605 -158.275 ;
        RECT 260.275 -159.965 260.605 -159.635 ;
        RECT 260.275 -161.325 260.605 -160.995 ;
        RECT 260.275 -162.685 260.605 -162.355 ;
        RECT 260.275 -164.045 260.605 -163.715 ;
        RECT 260.275 -165.405 260.605 -165.075 ;
        RECT 260.275 -166.765 260.605 -166.435 ;
        RECT 260.275 -168.125 260.605 -167.795 ;
        RECT 260.275 -169.485 260.605 -169.155 ;
        RECT 260.275 -170.845 260.605 -170.515 ;
        RECT 260.275 -172.205 260.605 -171.875 ;
        RECT 260.275 -173.565 260.605 -173.235 ;
        RECT 260.275 -174.925 260.605 -174.595 ;
        RECT 260.275 -176.285 260.605 -175.955 ;
        RECT 260.275 -177.645 260.605 -177.315 ;
        RECT 260.275 -179.005 260.605 -178.675 ;
        RECT 260.275 -180.365 260.605 -180.035 ;
        RECT 260.275 -181.725 260.605 -181.395 ;
        RECT 260.275 -183.085 260.605 -182.755 ;
        RECT 260.275 -184.445 260.605 -184.115 ;
        RECT 260.275 -185.805 260.605 -185.475 ;
        RECT 260.275 -187.165 260.605 -186.835 ;
        RECT 260.275 -188.525 260.605 -188.195 ;
        RECT 260.275 -189.885 260.605 -189.555 ;
        RECT 260.275 -191.245 260.605 -190.915 ;
        RECT 260.275 -192.605 260.605 -192.275 ;
        RECT 260.275 -193.965 260.605 -193.635 ;
        RECT 260.275 -195.325 260.605 -194.995 ;
        RECT 260.275 -196.685 260.605 -196.355 ;
        RECT 260.275 -198.045 260.605 -197.715 ;
        RECT 260.275 -199.405 260.605 -199.075 ;
        RECT 260.275 -200.765 260.605 -200.435 ;
        RECT 260.275 -202.125 260.605 -201.795 ;
        RECT 260.275 -203.485 260.605 -203.155 ;
        RECT 260.275 -204.845 260.605 -204.515 ;
        RECT 260.275 -206.205 260.605 -205.875 ;
        RECT 260.275 -207.565 260.605 -207.235 ;
        RECT 260.275 -208.925 260.605 -208.595 ;
        RECT 260.275 -210.285 260.605 -209.955 ;
        RECT 260.275 -211.645 260.605 -211.315 ;
        RECT 260.275 -213.005 260.605 -212.675 ;
        RECT 260.275 -214.365 260.605 -214.035 ;
        RECT 260.275 -215.725 260.605 -215.395 ;
        RECT 260.275 -217.085 260.605 -216.755 ;
        RECT 260.275 -218.445 260.605 -218.115 ;
        RECT 260.275 -219.805 260.605 -219.475 ;
        RECT 260.275 -221.165 260.605 -220.835 ;
        RECT 260.275 -222.525 260.605 -222.195 ;
        RECT 260.275 -223.885 260.605 -223.555 ;
        RECT 260.275 -225.245 260.605 -224.915 ;
        RECT 260.275 -226.605 260.605 -226.275 ;
        RECT 260.275 -227.965 260.605 -227.635 ;
        RECT 260.275 -229.325 260.605 -228.995 ;
        RECT 260.275 -230.685 260.605 -230.355 ;
        RECT 260.275 -232.045 260.605 -231.715 ;
        RECT 260.275 -233.405 260.605 -233.075 ;
        RECT 260.275 -234.765 260.605 -234.435 ;
        RECT 260.275 -236.125 260.605 -235.795 ;
        RECT 260.275 -237.485 260.605 -237.155 ;
        RECT 260.275 -238.845 260.605 -238.515 ;
        RECT 260.275 -241.09 260.605 -239.96 ;
        RECT 260.28 -241.205 260.6 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 244.04 261.965 245.17 ;
        RECT 261.635 242.595 261.965 242.925 ;
        RECT 261.635 241.235 261.965 241.565 ;
        RECT 261.635 239.875 261.965 240.205 ;
        RECT 261.635 238.515 261.965 238.845 ;
        RECT 261.635 237.155 261.965 237.485 ;
        RECT 261.64 237.155 261.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 -0.845 261.965 -0.515 ;
        RECT 261.635 -2.205 261.965 -1.875 ;
        RECT 261.635 -3.565 261.965 -3.235 ;
        RECT 261.64 -3.565 261.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 -123.245 261.965 -122.915 ;
        RECT 261.635 -124.605 261.965 -124.275 ;
        RECT 261.635 -125.965 261.965 -125.635 ;
        RECT 261.635 -127.325 261.965 -126.995 ;
        RECT 261.635 -128.685 261.965 -128.355 ;
        RECT 261.635 -130.045 261.965 -129.715 ;
        RECT 261.635 -131.405 261.965 -131.075 ;
        RECT 261.635 -132.765 261.965 -132.435 ;
        RECT 261.635 -134.125 261.965 -133.795 ;
        RECT 261.635 -135.485 261.965 -135.155 ;
        RECT 261.635 -136.845 261.965 -136.515 ;
        RECT 261.635 -138.205 261.965 -137.875 ;
        RECT 261.635 -139.565 261.965 -139.235 ;
        RECT 261.635 -140.925 261.965 -140.595 ;
        RECT 261.635 -142.285 261.965 -141.955 ;
        RECT 261.635 -143.645 261.965 -143.315 ;
        RECT 261.635 -145.005 261.965 -144.675 ;
        RECT 261.635 -146.365 261.965 -146.035 ;
        RECT 261.635 -147.725 261.965 -147.395 ;
        RECT 261.635 -149.085 261.965 -148.755 ;
        RECT 261.635 -150.445 261.965 -150.115 ;
        RECT 261.635 -151.805 261.965 -151.475 ;
        RECT 261.635 -153.165 261.965 -152.835 ;
        RECT 261.635 -154.525 261.965 -154.195 ;
        RECT 261.635 -155.885 261.965 -155.555 ;
        RECT 261.635 -157.245 261.965 -156.915 ;
        RECT 261.635 -158.605 261.965 -158.275 ;
        RECT 261.635 -159.965 261.965 -159.635 ;
        RECT 261.635 -161.325 261.965 -160.995 ;
        RECT 261.635 -162.685 261.965 -162.355 ;
        RECT 261.635 -164.045 261.965 -163.715 ;
        RECT 261.635 -165.405 261.965 -165.075 ;
        RECT 261.635 -166.765 261.965 -166.435 ;
        RECT 261.635 -168.125 261.965 -167.795 ;
        RECT 261.635 -169.485 261.965 -169.155 ;
        RECT 261.635 -170.845 261.965 -170.515 ;
        RECT 261.635 -172.205 261.965 -171.875 ;
        RECT 261.635 -173.565 261.965 -173.235 ;
        RECT 261.635 -174.925 261.965 -174.595 ;
        RECT 261.635 -176.285 261.965 -175.955 ;
        RECT 261.635 -177.645 261.965 -177.315 ;
        RECT 261.635 -179.005 261.965 -178.675 ;
        RECT 261.635 -180.365 261.965 -180.035 ;
        RECT 261.635 -181.725 261.965 -181.395 ;
        RECT 261.635 -183.085 261.965 -182.755 ;
        RECT 261.635 -184.445 261.965 -184.115 ;
        RECT 261.635 -185.805 261.965 -185.475 ;
        RECT 261.635 -187.165 261.965 -186.835 ;
        RECT 261.635 -188.525 261.965 -188.195 ;
        RECT 261.635 -189.885 261.965 -189.555 ;
        RECT 261.635 -191.245 261.965 -190.915 ;
        RECT 261.635 -192.605 261.965 -192.275 ;
        RECT 261.635 -193.965 261.965 -193.635 ;
        RECT 261.635 -195.325 261.965 -194.995 ;
        RECT 261.635 -196.685 261.965 -196.355 ;
        RECT 261.635 -198.045 261.965 -197.715 ;
        RECT 261.635 -199.405 261.965 -199.075 ;
        RECT 261.635 -200.765 261.965 -200.435 ;
        RECT 261.635 -202.125 261.965 -201.795 ;
        RECT 261.635 -203.485 261.965 -203.155 ;
        RECT 261.635 -204.845 261.965 -204.515 ;
        RECT 261.635 -206.205 261.965 -205.875 ;
        RECT 261.635 -207.565 261.965 -207.235 ;
        RECT 261.635 -208.925 261.965 -208.595 ;
        RECT 261.635 -210.285 261.965 -209.955 ;
        RECT 261.635 -211.645 261.965 -211.315 ;
        RECT 261.635 -213.005 261.965 -212.675 ;
        RECT 261.635 -214.365 261.965 -214.035 ;
        RECT 261.635 -215.725 261.965 -215.395 ;
        RECT 261.635 -217.085 261.965 -216.755 ;
        RECT 261.635 -218.445 261.965 -218.115 ;
        RECT 261.635 -219.805 261.965 -219.475 ;
        RECT 261.635 -221.165 261.965 -220.835 ;
        RECT 261.635 -222.525 261.965 -222.195 ;
        RECT 261.635 -223.885 261.965 -223.555 ;
        RECT 261.635 -225.245 261.965 -224.915 ;
        RECT 261.635 -226.605 261.965 -226.275 ;
        RECT 261.635 -227.965 261.965 -227.635 ;
        RECT 261.635 -229.325 261.965 -228.995 ;
        RECT 261.635 -230.685 261.965 -230.355 ;
        RECT 261.635 -232.045 261.965 -231.715 ;
        RECT 261.635 -233.405 261.965 -233.075 ;
        RECT 261.635 -234.765 261.965 -234.435 ;
        RECT 261.635 -236.125 261.965 -235.795 ;
        RECT 261.635 -237.485 261.965 -237.155 ;
        RECT 261.635 -238.845 261.965 -238.515 ;
        RECT 261.635 -241.09 261.965 -239.96 ;
        RECT 261.64 -241.205 261.96 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 244.04 263.325 245.17 ;
        RECT 262.995 242.595 263.325 242.925 ;
        RECT 262.995 241.235 263.325 241.565 ;
        RECT 262.995 239.875 263.325 240.205 ;
        RECT 262.995 238.515 263.325 238.845 ;
        RECT 262.995 237.155 263.325 237.485 ;
        RECT 263 237.155 263.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 -0.845 263.325 -0.515 ;
        RECT 262.995 -2.205 263.325 -1.875 ;
        RECT 262.995 -3.565 263.325 -3.235 ;
        RECT 263 -3.565 263.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 -123.245 263.325 -122.915 ;
        RECT 262.995 -124.605 263.325 -124.275 ;
        RECT 262.995 -125.965 263.325 -125.635 ;
        RECT 262.995 -127.325 263.325 -126.995 ;
        RECT 262.995 -128.685 263.325 -128.355 ;
        RECT 262.995 -130.045 263.325 -129.715 ;
        RECT 262.995 -131.405 263.325 -131.075 ;
        RECT 262.995 -132.765 263.325 -132.435 ;
        RECT 262.995 -134.125 263.325 -133.795 ;
        RECT 262.995 -135.485 263.325 -135.155 ;
        RECT 262.995 -136.845 263.325 -136.515 ;
        RECT 262.995 -138.205 263.325 -137.875 ;
        RECT 262.995 -139.565 263.325 -139.235 ;
        RECT 262.995 -140.925 263.325 -140.595 ;
        RECT 262.995 -142.285 263.325 -141.955 ;
        RECT 262.995 -143.645 263.325 -143.315 ;
        RECT 262.995 -145.005 263.325 -144.675 ;
        RECT 262.995 -146.365 263.325 -146.035 ;
        RECT 262.995 -147.725 263.325 -147.395 ;
        RECT 262.995 -149.085 263.325 -148.755 ;
        RECT 262.995 -150.445 263.325 -150.115 ;
        RECT 262.995 -151.805 263.325 -151.475 ;
        RECT 262.995 -153.165 263.325 -152.835 ;
        RECT 262.995 -154.525 263.325 -154.195 ;
        RECT 262.995 -155.885 263.325 -155.555 ;
        RECT 262.995 -157.245 263.325 -156.915 ;
        RECT 262.995 -158.605 263.325 -158.275 ;
        RECT 262.995 -159.965 263.325 -159.635 ;
        RECT 262.995 -161.325 263.325 -160.995 ;
        RECT 262.995 -162.685 263.325 -162.355 ;
        RECT 262.995 -164.045 263.325 -163.715 ;
        RECT 262.995 -165.405 263.325 -165.075 ;
        RECT 262.995 -166.765 263.325 -166.435 ;
        RECT 262.995 -168.125 263.325 -167.795 ;
        RECT 262.995 -169.485 263.325 -169.155 ;
        RECT 262.995 -170.845 263.325 -170.515 ;
        RECT 262.995 -172.205 263.325 -171.875 ;
        RECT 262.995 -173.565 263.325 -173.235 ;
        RECT 262.995 -174.925 263.325 -174.595 ;
        RECT 262.995 -176.285 263.325 -175.955 ;
        RECT 262.995 -177.645 263.325 -177.315 ;
        RECT 262.995 -179.005 263.325 -178.675 ;
        RECT 262.995 -180.365 263.325 -180.035 ;
        RECT 262.995 -181.725 263.325 -181.395 ;
        RECT 262.995 -183.085 263.325 -182.755 ;
        RECT 262.995 -184.445 263.325 -184.115 ;
        RECT 262.995 -185.805 263.325 -185.475 ;
        RECT 262.995 -187.165 263.325 -186.835 ;
        RECT 262.995 -188.525 263.325 -188.195 ;
        RECT 262.995 -189.885 263.325 -189.555 ;
        RECT 262.995 -191.245 263.325 -190.915 ;
        RECT 262.995 -192.605 263.325 -192.275 ;
        RECT 262.995 -193.965 263.325 -193.635 ;
        RECT 262.995 -195.325 263.325 -194.995 ;
        RECT 262.995 -196.685 263.325 -196.355 ;
        RECT 262.995 -198.045 263.325 -197.715 ;
        RECT 262.995 -199.405 263.325 -199.075 ;
        RECT 262.995 -200.765 263.325 -200.435 ;
        RECT 262.995 -202.125 263.325 -201.795 ;
        RECT 262.995 -203.485 263.325 -203.155 ;
        RECT 262.995 -204.845 263.325 -204.515 ;
        RECT 262.995 -206.205 263.325 -205.875 ;
        RECT 262.995 -207.565 263.325 -207.235 ;
        RECT 262.995 -208.925 263.325 -208.595 ;
        RECT 262.995 -210.285 263.325 -209.955 ;
        RECT 262.995 -211.645 263.325 -211.315 ;
        RECT 262.995 -213.005 263.325 -212.675 ;
        RECT 262.995 -214.365 263.325 -214.035 ;
        RECT 262.995 -215.725 263.325 -215.395 ;
        RECT 262.995 -217.085 263.325 -216.755 ;
        RECT 262.995 -218.445 263.325 -218.115 ;
        RECT 262.995 -219.805 263.325 -219.475 ;
        RECT 262.995 -221.165 263.325 -220.835 ;
        RECT 262.995 -222.525 263.325 -222.195 ;
        RECT 262.995 -223.885 263.325 -223.555 ;
        RECT 262.995 -225.245 263.325 -224.915 ;
        RECT 262.995 -226.605 263.325 -226.275 ;
        RECT 262.995 -227.965 263.325 -227.635 ;
        RECT 262.995 -229.325 263.325 -228.995 ;
        RECT 262.995 -230.685 263.325 -230.355 ;
        RECT 262.995 -232.045 263.325 -231.715 ;
        RECT 262.995 -233.405 263.325 -233.075 ;
        RECT 262.995 -234.765 263.325 -234.435 ;
        RECT 262.995 -236.125 263.325 -235.795 ;
        RECT 262.995 -237.485 263.325 -237.155 ;
        RECT 262.995 -238.845 263.325 -238.515 ;
        RECT 262.995 -241.09 263.325 -239.96 ;
        RECT 263 -241.205 263.32 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 244.04 264.685 245.17 ;
        RECT 264.355 242.595 264.685 242.925 ;
        RECT 264.355 241.235 264.685 241.565 ;
        RECT 264.355 239.875 264.685 240.205 ;
        RECT 264.355 238.515 264.685 238.845 ;
        RECT 264.355 237.155 264.685 237.485 ;
        RECT 264.36 237.155 264.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 -127.325 264.685 -126.995 ;
        RECT 264.355 -128.685 264.685 -128.355 ;
        RECT 264.355 -130.045 264.685 -129.715 ;
        RECT 264.355 -131.405 264.685 -131.075 ;
        RECT 264.355 -132.765 264.685 -132.435 ;
        RECT 264.355 -134.125 264.685 -133.795 ;
        RECT 264.355 -135.485 264.685 -135.155 ;
        RECT 264.355 -136.845 264.685 -136.515 ;
        RECT 264.355 -138.205 264.685 -137.875 ;
        RECT 264.355 -139.565 264.685 -139.235 ;
        RECT 264.355 -140.925 264.685 -140.595 ;
        RECT 264.355 -142.285 264.685 -141.955 ;
        RECT 264.355 -143.645 264.685 -143.315 ;
        RECT 264.355 -145.005 264.685 -144.675 ;
        RECT 264.355 -146.365 264.685 -146.035 ;
        RECT 264.355 -147.725 264.685 -147.395 ;
        RECT 264.355 -149.085 264.685 -148.755 ;
        RECT 264.355 -150.445 264.685 -150.115 ;
        RECT 264.355 -151.805 264.685 -151.475 ;
        RECT 264.355 -153.165 264.685 -152.835 ;
        RECT 264.355 -154.525 264.685 -154.195 ;
        RECT 264.355 -155.885 264.685 -155.555 ;
        RECT 264.355 -157.245 264.685 -156.915 ;
        RECT 264.355 -158.605 264.685 -158.275 ;
        RECT 264.355 -159.965 264.685 -159.635 ;
        RECT 264.355 -161.325 264.685 -160.995 ;
        RECT 264.355 -162.685 264.685 -162.355 ;
        RECT 264.355 -164.045 264.685 -163.715 ;
        RECT 264.355 -165.405 264.685 -165.075 ;
        RECT 264.355 -166.765 264.685 -166.435 ;
        RECT 264.355 -168.125 264.685 -167.795 ;
        RECT 264.355 -169.485 264.685 -169.155 ;
        RECT 264.355 -170.845 264.685 -170.515 ;
        RECT 264.355 -172.205 264.685 -171.875 ;
        RECT 264.355 -173.565 264.685 -173.235 ;
        RECT 264.355 -174.925 264.685 -174.595 ;
        RECT 264.355 -176.285 264.685 -175.955 ;
        RECT 264.355 -177.645 264.685 -177.315 ;
        RECT 264.355 -179.005 264.685 -178.675 ;
        RECT 264.355 -180.365 264.685 -180.035 ;
        RECT 264.355 -181.725 264.685 -181.395 ;
        RECT 264.355 -183.085 264.685 -182.755 ;
        RECT 264.355 -184.445 264.685 -184.115 ;
        RECT 264.355 -185.805 264.685 -185.475 ;
        RECT 264.355 -187.165 264.685 -186.835 ;
        RECT 264.355 -188.525 264.685 -188.195 ;
        RECT 264.355 -189.885 264.685 -189.555 ;
        RECT 264.355 -191.245 264.685 -190.915 ;
        RECT 264.355 -192.605 264.685 -192.275 ;
        RECT 264.355 -193.965 264.685 -193.635 ;
        RECT 264.355 -195.325 264.685 -194.995 ;
        RECT 264.355 -196.685 264.685 -196.355 ;
        RECT 264.355 -198.045 264.685 -197.715 ;
        RECT 264.355 -199.405 264.685 -199.075 ;
        RECT 264.355 -200.765 264.685 -200.435 ;
        RECT 264.355 -202.125 264.685 -201.795 ;
        RECT 264.355 -203.485 264.685 -203.155 ;
        RECT 264.355 -204.845 264.685 -204.515 ;
        RECT 264.355 -206.205 264.685 -205.875 ;
        RECT 264.355 -207.565 264.685 -207.235 ;
        RECT 264.355 -208.925 264.685 -208.595 ;
        RECT 264.355 -210.285 264.685 -209.955 ;
        RECT 264.355 -211.645 264.685 -211.315 ;
        RECT 264.355 -213.005 264.685 -212.675 ;
        RECT 264.355 -214.365 264.685 -214.035 ;
        RECT 264.355 -215.725 264.685 -215.395 ;
        RECT 264.355 -217.085 264.685 -216.755 ;
        RECT 264.355 -218.445 264.685 -218.115 ;
        RECT 264.355 -219.805 264.685 -219.475 ;
        RECT 264.355 -221.165 264.685 -220.835 ;
        RECT 264.355 -222.525 264.685 -222.195 ;
        RECT 264.355 -223.885 264.685 -223.555 ;
        RECT 264.355 -225.245 264.685 -224.915 ;
        RECT 264.355 -226.605 264.685 -226.275 ;
        RECT 264.355 -227.965 264.685 -227.635 ;
        RECT 264.355 -229.325 264.685 -228.995 ;
        RECT 264.355 -230.685 264.685 -230.355 ;
        RECT 264.355 -232.045 264.685 -231.715 ;
        RECT 264.355 -233.405 264.685 -233.075 ;
        RECT 264.355 -234.765 264.685 -234.435 ;
        RECT 264.355 -236.125 264.685 -235.795 ;
        RECT 264.355 -237.485 264.685 -237.155 ;
        RECT 264.355 -238.845 264.685 -238.515 ;
        RECT 264.355 -241.09 264.685 -239.96 ;
        RECT 264.36 -241.205 264.68 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.91 -125.535 265.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.715 244.04 266.045 245.17 ;
        RECT 265.715 242.595 266.045 242.925 ;
        RECT 265.715 241.235 266.045 241.565 ;
        RECT 265.715 239.875 266.045 240.205 ;
        RECT 265.715 238.515 266.045 238.845 ;
        RECT 265.715 237.155 266.045 237.485 ;
        RECT 265.72 237.155 266.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.715 -0.845 266.045 -0.515 ;
        RECT 265.715 -2.205 266.045 -1.875 ;
        RECT 265.715 -3.565 266.045 -3.235 ;
        RECT 265.72 -3.565 266.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 244.04 267.405 245.17 ;
        RECT 267.075 242.595 267.405 242.925 ;
        RECT 267.075 241.235 267.405 241.565 ;
        RECT 267.075 239.875 267.405 240.205 ;
        RECT 267.075 238.515 267.405 238.845 ;
        RECT 267.075 237.155 267.405 237.485 ;
        RECT 267.08 237.155 267.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 -0.845 267.405 -0.515 ;
        RECT 267.075 -2.205 267.405 -1.875 ;
        RECT 267.075 -3.565 267.405 -3.235 ;
        RECT 267.08 -3.565 267.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 244.04 268.765 245.17 ;
        RECT 268.435 242.595 268.765 242.925 ;
        RECT 268.435 241.235 268.765 241.565 ;
        RECT 268.435 239.875 268.765 240.205 ;
        RECT 268.435 238.515 268.765 238.845 ;
        RECT 268.435 237.155 268.765 237.485 ;
        RECT 268.44 237.155 268.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 -0.845 268.765 -0.515 ;
        RECT 268.435 -2.205 268.765 -1.875 ;
        RECT 268.435 -3.565 268.765 -3.235 ;
        RECT 268.44 -3.565 268.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 -123.245 268.765 -122.915 ;
        RECT 268.435 -124.605 268.765 -124.275 ;
        RECT 268.435 -125.965 268.765 -125.635 ;
        RECT 268.435 -127.325 268.765 -126.995 ;
        RECT 268.435 -128.685 268.765 -128.355 ;
        RECT 268.435 -130.045 268.765 -129.715 ;
        RECT 268.435 -131.405 268.765 -131.075 ;
        RECT 268.435 -132.765 268.765 -132.435 ;
        RECT 268.435 -134.125 268.765 -133.795 ;
        RECT 268.435 -135.485 268.765 -135.155 ;
        RECT 268.435 -136.845 268.765 -136.515 ;
        RECT 268.435 -138.205 268.765 -137.875 ;
        RECT 268.435 -139.565 268.765 -139.235 ;
        RECT 268.435 -140.925 268.765 -140.595 ;
        RECT 268.435 -142.285 268.765 -141.955 ;
        RECT 268.435 -143.645 268.765 -143.315 ;
        RECT 268.435 -145.005 268.765 -144.675 ;
        RECT 268.435 -146.365 268.765 -146.035 ;
        RECT 268.435 -147.725 268.765 -147.395 ;
        RECT 268.435 -149.085 268.765 -148.755 ;
        RECT 268.435 -150.445 268.765 -150.115 ;
        RECT 268.435 -151.805 268.765 -151.475 ;
        RECT 268.435 -153.165 268.765 -152.835 ;
        RECT 268.435 -154.525 268.765 -154.195 ;
        RECT 268.435 -155.885 268.765 -155.555 ;
        RECT 268.435 -157.245 268.765 -156.915 ;
        RECT 268.435 -158.605 268.765 -158.275 ;
        RECT 268.435 -159.965 268.765 -159.635 ;
        RECT 268.435 -161.325 268.765 -160.995 ;
        RECT 268.435 -162.685 268.765 -162.355 ;
        RECT 268.435 -164.045 268.765 -163.715 ;
        RECT 268.435 -165.405 268.765 -165.075 ;
        RECT 268.435 -166.765 268.765 -166.435 ;
        RECT 268.435 -168.125 268.765 -167.795 ;
        RECT 268.435 -169.485 268.765 -169.155 ;
        RECT 268.435 -170.845 268.765 -170.515 ;
        RECT 268.435 -172.205 268.765 -171.875 ;
        RECT 268.435 -173.565 268.765 -173.235 ;
        RECT 268.435 -174.925 268.765 -174.595 ;
        RECT 268.435 -176.285 268.765 -175.955 ;
        RECT 268.435 -177.645 268.765 -177.315 ;
        RECT 268.435 -179.005 268.765 -178.675 ;
        RECT 268.435 -180.365 268.765 -180.035 ;
        RECT 268.435 -181.725 268.765 -181.395 ;
        RECT 268.435 -183.085 268.765 -182.755 ;
        RECT 268.435 -184.445 268.765 -184.115 ;
        RECT 268.435 -185.805 268.765 -185.475 ;
        RECT 268.435 -187.165 268.765 -186.835 ;
        RECT 268.435 -188.525 268.765 -188.195 ;
        RECT 268.435 -189.885 268.765 -189.555 ;
        RECT 268.435 -191.245 268.765 -190.915 ;
        RECT 268.435 -192.605 268.765 -192.275 ;
        RECT 268.435 -193.965 268.765 -193.635 ;
        RECT 268.435 -195.325 268.765 -194.995 ;
        RECT 268.435 -196.685 268.765 -196.355 ;
        RECT 268.435 -198.045 268.765 -197.715 ;
        RECT 268.435 -199.405 268.765 -199.075 ;
        RECT 268.435 -200.765 268.765 -200.435 ;
        RECT 268.435 -202.125 268.765 -201.795 ;
        RECT 268.435 -203.485 268.765 -203.155 ;
        RECT 268.435 -204.845 268.765 -204.515 ;
        RECT 268.435 -206.205 268.765 -205.875 ;
        RECT 268.435 -207.565 268.765 -207.235 ;
        RECT 268.435 -208.925 268.765 -208.595 ;
        RECT 268.435 -210.285 268.765 -209.955 ;
        RECT 268.435 -211.645 268.765 -211.315 ;
        RECT 268.435 -213.005 268.765 -212.675 ;
        RECT 268.435 -214.365 268.765 -214.035 ;
        RECT 268.435 -215.725 268.765 -215.395 ;
        RECT 268.435 -217.085 268.765 -216.755 ;
        RECT 268.435 -218.445 268.765 -218.115 ;
        RECT 268.435 -219.805 268.765 -219.475 ;
        RECT 268.435 -221.165 268.765 -220.835 ;
        RECT 268.435 -222.525 268.765 -222.195 ;
        RECT 268.435 -223.885 268.765 -223.555 ;
        RECT 268.435 -225.245 268.765 -224.915 ;
        RECT 268.435 -226.605 268.765 -226.275 ;
        RECT 268.435 -227.965 268.765 -227.635 ;
        RECT 268.435 -229.325 268.765 -228.995 ;
        RECT 268.435 -230.685 268.765 -230.355 ;
        RECT 268.435 -232.045 268.765 -231.715 ;
        RECT 268.435 -233.405 268.765 -233.075 ;
        RECT 268.435 -234.765 268.765 -234.435 ;
        RECT 268.435 -236.125 268.765 -235.795 ;
        RECT 268.435 -237.485 268.765 -237.155 ;
        RECT 268.435 -238.845 268.765 -238.515 ;
        RECT 268.435 -241.09 268.765 -239.96 ;
        RECT 268.44 -241.205 268.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 244.04 270.125 245.17 ;
        RECT 269.795 242.595 270.125 242.925 ;
        RECT 269.795 241.235 270.125 241.565 ;
        RECT 269.795 239.875 270.125 240.205 ;
        RECT 269.795 238.515 270.125 238.845 ;
        RECT 269.795 237.155 270.125 237.485 ;
        RECT 269.8 237.155 270.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 -0.845 270.125 -0.515 ;
        RECT 269.795 -2.205 270.125 -1.875 ;
        RECT 269.795 -3.565 270.125 -3.235 ;
        RECT 269.8 -3.565 270.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 -123.245 270.125 -122.915 ;
        RECT 269.795 -124.605 270.125 -124.275 ;
        RECT 269.795 -125.965 270.125 -125.635 ;
        RECT 269.795 -127.325 270.125 -126.995 ;
        RECT 269.795 -128.685 270.125 -128.355 ;
        RECT 269.795 -130.045 270.125 -129.715 ;
        RECT 269.795 -131.405 270.125 -131.075 ;
        RECT 269.795 -132.765 270.125 -132.435 ;
        RECT 269.795 -134.125 270.125 -133.795 ;
        RECT 269.795 -135.485 270.125 -135.155 ;
        RECT 269.795 -136.845 270.125 -136.515 ;
        RECT 269.795 -138.205 270.125 -137.875 ;
        RECT 269.795 -139.565 270.125 -139.235 ;
        RECT 269.795 -140.925 270.125 -140.595 ;
        RECT 269.795 -142.285 270.125 -141.955 ;
        RECT 269.795 -143.645 270.125 -143.315 ;
        RECT 269.795 -145.005 270.125 -144.675 ;
        RECT 269.795 -146.365 270.125 -146.035 ;
        RECT 269.795 -147.725 270.125 -147.395 ;
        RECT 269.795 -149.085 270.125 -148.755 ;
        RECT 269.795 -150.445 270.125 -150.115 ;
        RECT 269.795 -151.805 270.125 -151.475 ;
        RECT 269.795 -153.165 270.125 -152.835 ;
        RECT 269.795 -154.525 270.125 -154.195 ;
        RECT 269.795 -155.885 270.125 -155.555 ;
        RECT 269.795 -157.245 270.125 -156.915 ;
        RECT 269.795 -158.605 270.125 -158.275 ;
        RECT 269.795 -159.965 270.125 -159.635 ;
        RECT 269.795 -161.325 270.125 -160.995 ;
        RECT 269.795 -162.685 270.125 -162.355 ;
        RECT 269.795 -164.045 270.125 -163.715 ;
        RECT 269.795 -165.405 270.125 -165.075 ;
        RECT 269.795 -166.765 270.125 -166.435 ;
        RECT 269.795 -168.125 270.125 -167.795 ;
        RECT 269.795 -169.485 270.125 -169.155 ;
        RECT 269.795 -170.845 270.125 -170.515 ;
        RECT 269.795 -172.205 270.125 -171.875 ;
        RECT 269.795 -173.565 270.125 -173.235 ;
        RECT 269.795 -174.925 270.125 -174.595 ;
        RECT 269.795 -176.285 270.125 -175.955 ;
        RECT 269.795 -177.645 270.125 -177.315 ;
        RECT 269.795 -179.005 270.125 -178.675 ;
        RECT 269.795 -180.365 270.125 -180.035 ;
        RECT 269.795 -181.725 270.125 -181.395 ;
        RECT 269.795 -183.085 270.125 -182.755 ;
        RECT 269.795 -184.445 270.125 -184.115 ;
        RECT 269.795 -185.805 270.125 -185.475 ;
        RECT 269.795 -187.165 270.125 -186.835 ;
        RECT 269.795 -188.525 270.125 -188.195 ;
        RECT 269.795 -189.885 270.125 -189.555 ;
        RECT 269.795 -191.245 270.125 -190.915 ;
        RECT 269.795 -192.605 270.125 -192.275 ;
        RECT 269.795 -193.965 270.125 -193.635 ;
        RECT 269.795 -195.325 270.125 -194.995 ;
        RECT 269.795 -196.685 270.125 -196.355 ;
        RECT 269.795 -198.045 270.125 -197.715 ;
        RECT 269.795 -199.405 270.125 -199.075 ;
        RECT 269.795 -200.765 270.125 -200.435 ;
        RECT 269.795 -202.125 270.125 -201.795 ;
        RECT 269.795 -203.485 270.125 -203.155 ;
        RECT 269.795 -204.845 270.125 -204.515 ;
        RECT 269.795 -206.205 270.125 -205.875 ;
        RECT 269.795 -207.565 270.125 -207.235 ;
        RECT 269.795 -208.925 270.125 -208.595 ;
        RECT 269.795 -210.285 270.125 -209.955 ;
        RECT 269.795 -211.645 270.125 -211.315 ;
        RECT 269.795 -213.005 270.125 -212.675 ;
        RECT 269.795 -214.365 270.125 -214.035 ;
        RECT 269.795 -215.725 270.125 -215.395 ;
        RECT 269.795 -217.085 270.125 -216.755 ;
        RECT 269.795 -218.445 270.125 -218.115 ;
        RECT 269.795 -219.805 270.125 -219.475 ;
        RECT 269.795 -221.165 270.125 -220.835 ;
        RECT 269.795 -222.525 270.125 -222.195 ;
        RECT 269.795 -223.885 270.125 -223.555 ;
        RECT 269.795 -225.245 270.125 -224.915 ;
        RECT 269.795 -226.605 270.125 -226.275 ;
        RECT 269.795 -227.965 270.125 -227.635 ;
        RECT 269.795 -229.325 270.125 -228.995 ;
        RECT 269.795 -230.685 270.125 -230.355 ;
        RECT 269.795 -232.045 270.125 -231.715 ;
        RECT 269.795 -233.405 270.125 -233.075 ;
        RECT 269.795 -234.765 270.125 -234.435 ;
        RECT 269.795 -236.125 270.125 -235.795 ;
        RECT 269.795 -237.485 270.125 -237.155 ;
        RECT 269.795 -238.845 270.125 -238.515 ;
        RECT 269.795 -241.09 270.125 -239.96 ;
        RECT 269.8 -241.205 270.12 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 244.04 271.485 245.17 ;
        RECT 271.155 242.595 271.485 242.925 ;
        RECT 271.155 241.235 271.485 241.565 ;
        RECT 271.155 239.875 271.485 240.205 ;
        RECT 271.155 238.515 271.485 238.845 ;
        RECT 271.155 237.155 271.485 237.485 ;
        RECT 271.16 237.155 271.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 -0.845 271.485 -0.515 ;
        RECT 271.155 -2.205 271.485 -1.875 ;
        RECT 271.155 -3.565 271.485 -3.235 ;
        RECT 271.16 -3.565 271.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 -150.445 271.485 -150.115 ;
        RECT 271.155 -151.805 271.485 -151.475 ;
        RECT 271.155 -153.165 271.485 -152.835 ;
        RECT 271.155 -154.525 271.485 -154.195 ;
        RECT 271.155 -155.885 271.485 -155.555 ;
        RECT 271.155 -157.245 271.485 -156.915 ;
        RECT 271.155 -158.605 271.485 -158.275 ;
        RECT 271.155 -159.965 271.485 -159.635 ;
        RECT 271.155 -161.325 271.485 -160.995 ;
        RECT 271.155 -162.685 271.485 -162.355 ;
        RECT 271.155 -164.045 271.485 -163.715 ;
        RECT 271.155 -165.405 271.485 -165.075 ;
        RECT 271.155 -166.765 271.485 -166.435 ;
        RECT 271.155 -168.125 271.485 -167.795 ;
        RECT 271.155 -169.485 271.485 -169.155 ;
        RECT 271.155 -170.845 271.485 -170.515 ;
        RECT 271.155 -172.205 271.485 -171.875 ;
        RECT 271.155 -173.565 271.485 -173.235 ;
        RECT 271.155 -174.925 271.485 -174.595 ;
        RECT 271.155 -176.285 271.485 -175.955 ;
        RECT 271.155 -177.645 271.485 -177.315 ;
        RECT 271.155 -179.005 271.485 -178.675 ;
        RECT 271.155 -180.365 271.485 -180.035 ;
        RECT 271.155 -181.725 271.485 -181.395 ;
        RECT 271.155 -183.085 271.485 -182.755 ;
        RECT 271.155 -184.445 271.485 -184.115 ;
        RECT 271.155 -185.805 271.485 -185.475 ;
        RECT 271.155 -187.165 271.485 -186.835 ;
        RECT 271.155 -188.525 271.485 -188.195 ;
        RECT 271.155 -189.885 271.485 -189.555 ;
        RECT 271.155 -191.245 271.485 -190.915 ;
        RECT 271.155 -192.605 271.485 -192.275 ;
        RECT 271.155 -193.965 271.485 -193.635 ;
        RECT 271.155 -195.325 271.485 -194.995 ;
        RECT 271.155 -196.685 271.485 -196.355 ;
        RECT 271.155 -198.045 271.485 -197.715 ;
        RECT 271.155 -199.405 271.485 -199.075 ;
        RECT 271.155 -200.765 271.485 -200.435 ;
        RECT 271.155 -202.125 271.485 -201.795 ;
        RECT 271.155 -203.485 271.485 -203.155 ;
        RECT 271.155 -204.845 271.485 -204.515 ;
        RECT 271.155 -206.205 271.485 -205.875 ;
        RECT 271.155 -207.565 271.485 -207.235 ;
        RECT 271.155 -208.925 271.485 -208.595 ;
        RECT 271.155 -210.285 271.485 -209.955 ;
        RECT 271.155 -211.645 271.485 -211.315 ;
        RECT 271.155 -213.005 271.485 -212.675 ;
        RECT 271.155 -214.365 271.485 -214.035 ;
        RECT 271.155 -215.725 271.485 -215.395 ;
        RECT 271.155 -217.085 271.485 -216.755 ;
        RECT 271.155 -218.445 271.485 -218.115 ;
        RECT 271.155 -219.805 271.485 -219.475 ;
        RECT 271.155 -221.165 271.485 -220.835 ;
        RECT 271.155 -222.525 271.485 -222.195 ;
        RECT 271.155 -223.885 271.485 -223.555 ;
        RECT 271.155 -225.245 271.485 -224.915 ;
        RECT 271.155 -226.605 271.485 -226.275 ;
        RECT 271.155 -227.965 271.485 -227.635 ;
        RECT 271.155 -229.325 271.485 -228.995 ;
        RECT 271.155 -230.685 271.485 -230.355 ;
        RECT 271.155 -232.045 271.485 -231.715 ;
        RECT 271.155 -233.405 271.485 -233.075 ;
        RECT 271.155 -234.765 271.485 -234.435 ;
        RECT 271.155 -236.125 271.485 -235.795 ;
        RECT 271.155 -237.485 271.485 -237.155 ;
        RECT 271.155 -238.845 271.485 -238.515 ;
        RECT 271.155 -241.09 271.485 -239.96 ;
        RECT 271.16 -241.205 271.48 -122.24 ;
        RECT 271.155 -123.245 271.485 -122.915 ;
        RECT 271.155 -124.605 271.485 -124.275 ;
        RECT 271.155 -125.965 271.485 -125.635 ;
        RECT 271.155 -127.325 271.485 -126.995 ;
        RECT 271.155 -128.685 271.485 -128.355 ;
        RECT 271.155 -130.045 271.485 -129.715 ;
        RECT 271.155 -131.405 271.485 -131.075 ;
        RECT 271.155 -132.765 271.485 -132.435 ;
        RECT 271.155 -134.125 271.485 -133.795 ;
        RECT 271.155 -135.485 271.485 -135.155 ;
        RECT 271.155 -136.845 271.485 -136.515 ;
        RECT 271.155 -138.205 271.485 -137.875 ;
        RECT 271.155 -139.565 271.485 -139.235 ;
        RECT 271.155 -140.925 271.485 -140.595 ;
        RECT 271.155 -142.285 271.485 -141.955 ;
        RECT 271.155 -143.645 271.485 -143.315 ;
        RECT 271.155 -145.005 271.485 -144.675 ;
        RECT 271.155 -146.365 271.485 -146.035 ;
        RECT 271.155 -147.725 271.485 -147.395 ;
        RECT 271.155 -149.085 271.485 -148.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 -123.245 237.485 -122.915 ;
        RECT 237.155 -124.605 237.485 -124.275 ;
        RECT 237.155 -125.965 237.485 -125.635 ;
        RECT 237.155 -127.325 237.485 -126.995 ;
        RECT 237.155 -128.685 237.485 -128.355 ;
        RECT 237.155 -130.045 237.485 -129.715 ;
        RECT 237.155 -131.405 237.485 -131.075 ;
        RECT 237.155 -132.765 237.485 -132.435 ;
        RECT 237.155 -134.125 237.485 -133.795 ;
        RECT 237.155 -135.485 237.485 -135.155 ;
        RECT 237.155 -136.845 237.485 -136.515 ;
        RECT 237.155 -138.205 237.485 -137.875 ;
        RECT 237.155 -139.565 237.485 -139.235 ;
        RECT 237.155 -140.925 237.485 -140.595 ;
        RECT 237.155 -142.285 237.485 -141.955 ;
        RECT 237.155 -143.645 237.485 -143.315 ;
        RECT 237.155 -145.005 237.485 -144.675 ;
        RECT 237.155 -146.365 237.485 -146.035 ;
        RECT 237.155 -147.725 237.485 -147.395 ;
        RECT 237.155 -149.085 237.485 -148.755 ;
        RECT 237.155 -150.445 237.485 -150.115 ;
        RECT 237.155 -151.805 237.485 -151.475 ;
        RECT 237.155 -153.165 237.485 -152.835 ;
        RECT 237.155 -154.525 237.485 -154.195 ;
        RECT 237.155 -155.885 237.485 -155.555 ;
        RECT 237.155 -157.245 237.485 -156.915 ;
        RECT 237.155 -158.605 237.485 -158.275 ;
        RECT 237.155 -159.965 237.485 -159.635 ;
        RECT 237.155 -161.325 237.485 -160.995 ;
        RECT 237.155 -162.685 237.485 -162.355 ;
        RECT 237.155 -164.045 237.485 -163.715 ;
        RECT 237.155 -165.405 237.485 -165.075 ;
        RECT 237.155 -166.765 237.485 -166.435 ;
        RECT 237.155 -168.125 237.485 -167.795 ;
        RECT 237.155 -169.485 237.485 -169.155 ;
        RECT 237.155 -170.845 237.485 -170.515 ;
        RECT 237.155 -172.205 237.485 -171.875 ;
        RECT 237.155 -173.565 237.485 -173.235 ;
        RECT 237.155 -174.925 237.485 -174.595 ;
        RECT 237.155 -176.285 237.485 -175.955 ;
        RECT 237.155 -177.645 237.485 -177.315 ;
        RECT 237.155 -179.005 237.485 -178.675 ;
        RECT 237.155 -180.365 237.485 -180.035 ;
        RECT 237.155 -181.725 237.485 -181.395 ;
        RECT 237.155 -183.085 237.485 -182.755 ;
        RECT 237.155 -184.445 237.485 -184.115 ;
        RECT 237.155 -185.805 237.485 -185.475 ;
        RECT 237.155 -187.165 237.485 -186.835 ;
        RECT 237.155 -188.525 237.485 -188.195 ;
        RECT 237.155 -189.885 237.485 -189.555 ;
        RECT 237.155 -191.245 237.485 -190.915 ;
        RECT 237.155 -192.605 237.485 -192.275 ;
        RECT 237.155 -193.965 237.485 -193.635 ;
        RECT 237.155 -195.325 237.485 -194.995 ;
        RECT 237.155 -196.685 237.485 -196.355 ;
        RECT 237.155 -198.045 237.485 -197.715 ;
        RECT 237.155 -199.405 237.485 -199.075 ;
        RECT 237.155 -200.765 237.485 -200.435 ;
        RECT 237.155 -202.125 237.485 -201.795 ;
        RECT 237.155 -203.485 237.485 -203.155 ;
        RECT 237.155 -204.845 237.485 -204.515 ;
        RECT 237.155 -206.205 237.485 -205.875 ;
        RECT 237.155 -207.565 237.485 -207.235 ;
        RECT 237.155 -208.925 237.485 -208.595 ;
        RECT 237.155 -210.285 237.485 -209.955 ;
        RECT 237.155 -211.645 237.485 -211.315 ;
        RECT 237.155 -213.005 237.485 -212.675 ;
        RECT 237.155 -214.365 237.485 -214.035 ;
        RECT 237.155 -215.725 237.485 -215.395 ;
        RECT 237.155 -217.085 237.485 -216.755 ;
        RECT 237.155 -218.445 237.485 -218.115 ;
        RECT 237.155 -219.805 237.485 -219.475 ;
        RECT 237.155 -221.165 237.485 -220.835 ;
        RECT 237.155 -222.525 237.485 -222.195 ;
        RECT 237.155 -223.885 237.485 -223.555 ;
        RECT 237.155 -225.245 237.485 -224.915 ;
        RECT 237.155 -226.605 237.485 -226.275 ;
        RECT 237.155 -227.965 237.485 -227.635 ;
        RECT 237.155 -229.325 237.485 -228.995 ;
        RECT 237.155 -230.685 237.485 -230.355 ;
        RECT 237.155 -232.045 237.485 -231.715 ;
        RECT 237.155 -233.405 237.485 -233.075 ;
        RECT 237.155 -234.765 237.485 -234.435 ;
        RECT 237.155 -236.125 237.485 -235.795 ;
        RECT 237.155 -237.485 237.485 -237.155 ;
        RECT 237.155 -238.845 237.485 -238.515 ;
        RECT 237.155 -241.09 237.485 -239.96 ;
        RECT 237.16 -241.205 237.48 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 244.04 238.845 245.17 ;
        RECT 238.515 242.595 238.845 242.925 ;
        RECT 238.515 241.235 238.845 241.565 ;
        RECT 238.515 239.875 238.845 240.205 ;
        RECT 238.515 238.515 238.845 238.845 ;
        RECT 238.515 237.155 238.845 237.485 ;
        RECT 238.52 237.155 238.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 -0.845 238.845 -0.515 ;
        RECT 238.515 -2.205 238.845 -1.875 ;
        RECT 238.515 -3.565 238.845 -3.235 ;
        RECT 238.52 -3.565 238.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 -123.245 238.845 -122.915 ;
        RECT 238.515 -124.605 238.845 -124.275 ;
        RECT 238.515 -125.965 238.845 -125.635 ;
        RECT 238.515 -127.325 238.845 -126.995 ;
        RECT 238.515 -128.685 238.845 -128.355 ;
        RECT 238.515 -130.045 238.845 -129.715 ;
        RECT 238.515 -131.405 238.845 -131.075 ;
        RECT 238.515 -132.765 238.845 -132.435 ;
        RECT 238.515 -134.125 238.845 -133.795 ;
        RECT 238.515 -135.485 238.845 -135.155 ;
        RECT 238.515 -136.845 238.845 -136.515 ;
        RECT 238.515 -138.205 238.845 -137.875 ;
        RECT 238.515 -139.565 238.845 -139.235 ;
        RECT 238.515 -140.925 238.845 -140.595 ;
        RECT 238.515 -142.285 238.845 -141.955 ;
        RECT 238.515 -143.645 238.845 -143.315 ;
        RECT 238.515 -145.005 238.845 -144.675 ;
        RECT 238.515 -146.365 238.845 -146.035 ;
        RECT 238.515 -147.725 238.845 -147.395 ;
        RECT 238.515 -149.085 238.845 -148.755 ;
        RECT 238.515 -150.445 238.845 -150.115 ;
        RECT 238.515 -151.805 238.845 -151.475 ;
        RECT 238.515 -153.165 238.845 -152.835 ;
        RECT 238.515 -154.525 238.845 -154.195 ;
        RECT 238.515 -155.885 238.845 -155.555 ;
        RECT 238.515 -157.245 238.845 -156.915 ;
        RECT 238.515 -158.605 238.845 -158.275 ;
        RECT 238.515 -159.965 238.845 -159.635 ;
        RECT 238.515 -161.325 238.845 -160.995 ;
        RECT 238.515 -162.685 238.845 -162.355 ;
        RECT 238.515 -164.045 238.845 -163.715 ;
        RECT 238.515 -165.405 238.845 -165.075 ;
        RECT 238.515 -166.765 238.845 -166.435 ;
        RECT 238.515 -168.125 238.845 -167.795 ;
        RECT 238.515 -169.485 238.845 -169.155 ;
        RECT 238.515 -170.845 238.845 -170.515 ;
        RECT 238.515 -172.205 238.845 -171.875 ;
        RECT 238.515 -173.565 238.845 -173.235 ;
        RECT 238.515 -174.925 238.845 -174.595 ;
        RECT 238.515 -176.285 238.845 -175.955 ;
        RECT 238.515 -177.645 238.845 -177.315 ;
        RECT 238.515 -179.005 238.845 -178.675 ;
        RECT 238.515 -180.365 238.845 -180.035 ;
        RECT 238.515 -181.725 238.845 -181.395 ;
        RECT 238.515 -183.085 238.845 -182.755 ;
        RECT 238.515 -184.445 238.845 -184.115 ;
        RECT 238.515 -185.805 238.845 -185.475 ;
        RECT 238.515 -187.165 238.845 -186.835 ;
        RECT 238.515 -188.525 238.845 -188.195 ;
        RECT 238.515 -189.885 238.845 -189.555 ;
        RECT 238.515 -191.245 238.845 -190.915 ;
        RECT 238.515 -192.605 238.845 -192.275 ;
        RECT 238.515 -193.965 238.845 -193.635 ;
        RECT 238.515 -195.325 238.845 -194.995 ;
        RECT 238.515 -196.685 238.845 -196.355 ;
        RECT 238.515 -198.045 238.845 -197.715 ;
        RECT 238.515 -199.405 238.845 -199.075 ;
        RECT 238.515 -200.765 238.845 -200.435 ;
        RECT 238.515 -202.125 238.845 -201.795 ;
        RECT 238.515 -203.485 238.845 -203.155 ;
        RECT 238.515 -204.845 238.845 -204.515 ;
        RECT 238.515 -206.205 238.845 -205.875 ;
        RECT 238.515 -207.565 238.845 -207.235 ;
        RECT 238.515 -208.925 238.845 -208.595 ;
        RECT 238.515 -210.285 238.845 -209.955 ;
        RECT 238.515 -211.645 238.845 -211.315 ;
        RECT 238.515 -213.005 238.845 -212.675 ;
        RECT 238.515 -214.365 238.845 -214.035 ;
        RECT 238.515 -215.725 238.845 -215.395 ;
        RECT 238.515 -217.085 238.845 -216.755 ;
        RECT 238.515 -218.445 238.845 -218.115 ;
        RECT 238.515 -219.805 238.845 -219.475 ;
        RECT 238.515 -221.165 238.845 -220.835 ;
        RECT 238.515 -222.525 238.845 -222.195 ;
        RECT 238.515 -223.885 238.845 -223.555 ;
        RECT 238.515 -225.245 238.845 -224.915 ;
        RECT 238.515 -226.605 238.845 -226.275 ;
        RECT 238.515 -227.965 238.845 -227.635 ;
        RECT 238.515 -229.325 238.845 -228.995 ;
        RECT 238.515 -230.685 238.845 -230.355 ;
        RECT 238.515 -232.045 238.845 -231.715 ;
        RECT 238.515 -233.405 238.845 -233.075 ;
        RECT 238.515 -234.765 238.845 -234.435 ;
        RECT 238.515 -236.125 238.845 -235.795 ;
        RECT 238.515 -237.485 238.845 -237.155 ;
        RECT 238.515 -238.845 238.845 -238.515 ;
        RECT 238.515 -241.09 238.845 -239.96 ;
        RECT 238.52 -241.205 238.84 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 244.04 240.205 245.17 ;
        RECT 239.875 242.595 240.205 242.925 ;
        RECT 239.875 241.235 240.205 241.565 ;
        RECT 239.875 239.875 240.205 240.205 ;
        RECT 239.875 238.515 240.205 238.845 ;
        RECT 239.875 237.155 240.205 237.485 ;
        RECT 239.88 237.155 240.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 -0.845 240.205 -0.515 ;
        RECT 239.875 -2.205 240.205 -1.875 ;
        RECT 239.875 -3.565 240.205 -3.235 ;
        RECT 239.88 -3.565 240.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 -123.245 240.205 -122.915 ;
        RECT 239.875 -124.605 240.205 -124.275 ;
        RECT 239.875 -125.965 240.205 -125.635 ;
        RECT 239.875 -127.325 240.205 -126.995 ;
        RECT 239.875 -128.685 240.205 -128.355 ;
        RECT 239.875 -130.045 240.205 -129.715 ;
        RECT 239.875 -131.405 240.205 -131.075 ;
        RECT 239.875 -132.765 240.205 -132.435 ;
        RECT 239.875 -134.125 240.205 -133.795 ;
        RECT 239.875 -135.485 240.205 -135.155 ;
        RECT 239.875 -136.845 240.205 -136.515 ;
        RECT 239.875 -138.205 240.205 -137.875 ;
        RECT 239.875 -139.565 240.205 -139.235 ;
        RECT 239.875 -140.925 240.205 -140.595 ;
        RECT 239.875 -142.285 240.205 -141.955 ;
        RECT 239.875 -143.645 240.205 -143.315 ;
        RECT 239.875 -145.005 240.205 -144.675 ;
        RECT 239.875 -146.365 240.205 -146.035 ;
        RECT 239.875 -147.725 240.205 -147.395 ;
        RECT 239.875 -149.085 240.205 -148.755 ;
        RECT 239.875 -150.445 240.205 -150.115 ;
        RECT 239.875 -151.805 240.205 -151.475 ;
        RECT 239.875 -153.165 240.205 -152.835 ;
        RECT 239.875 -154.525 240.205 -154.195 ;
        RECT 239.875 -155.885 240.205 -155.555 ;
        RECT 239.875 -157.245 240.205 -156.915 ;
        RECT 239.875 -158.605 240.205 -158.275 ;
        RECT 239.875 -159.965 240.205 -159.635 ;
        RECT 239.875 -161.325 240.205 -160.995 ;
        RECT 239.875 -162.685 240.205 -162.355 ;
        RECT 239.875 -164.045 240.205 -163.715 ;
        RECT 239.875 -165.405 240.205 -165.075 ;
        RECT 239.875 -166.765 240.205 -166.435 ;
        RECT 239.875 -168.125 240.205 -167.795 ;
        RECT 239.875 -169.485 240.205 -169.155 ;
        RECT 239.875 -170.845 240.205 -170.515 ;
        RECT 239.875 -172.205 240.205 -171.875 ;
        RECT 239.875 -173.565 240.205 -173.235 ;
        RECT 239.875 -174.925 240.205 -174.595 ;
        RECT 239.875 -176.285 240.205 -175.955 ;
        RECT 239.875 -177.645 240.205 -177.315 ;
        RECT 239.875 -179.005 240.205 -178.675 ;
        RECT 239.875 -180.365 240.205 -180.035 ;
        RECT 239.875 -181.725 240.205 -181.395 ;
        RECT 239.875 -183.085 240.205 -182.755 ;
        RECT 239.875 -184.445 240.205 -184.115 ;
        RECT 239.875 -185.805 240.205 -185.475 ;
        RECT 239.875 -187.165 240.205 -186.835 ;
        RECT 239.875 -188.525 240.205 -188.195 ;
        RECT 239.875 -189.885 240.205 -189.555 ;
        RECT 239.875 -191.245 240.205 -190.915 ;
        RECT 239.875 -192.605 240.205 -192.275 ;
        RECT 239.875 -193.965 240.205 -193.635 ;
        RECT 239.875 -195.325 240.205 -194.995 ;
        RECT 239.875 -196.685 240.205 -196.355 ;
        RECT 239.875 -198.045 240.205 -197.715 ;
        RECT 239.875 -199.405 240.205 -199.075 ;
        RECT 239.875 -200.765 240.205 -200.435 ;
        RECT 239.875 -202.125 240.205 -201.795 ;
        RECT 239.875 -203.485 240.205 -203.155 ;
        RECT 239.875 -204.845 240.205 -204.515 ;
        RECT 239.875 -206.205 240.205 -205.875 ;
        RECT 239.875 -207.565 240.205 -207.235 ;
        RECT 239.875 -208.925 240.205 -208.595 ;
        RECT 239.875 -210.285 240.205 -209.955 ;
        RECT 239.875 -211.645 240.205 -211.315 ;
        RECT 239.875 -213.005 240.205 -212.675 ;
        RECT 239.875 -214.365 240.205 -214.035 ;
        RECT 239.875 -215.725 240.205 -215.395 ;
        RECT 239.875 -217.085 240.205 -216.755 ;
        RECT 239.875 -218.445 240.205 -218.115 ;
        RECT 239.875 -219.805 240.205 -219.475 ;
        RECT 239.875 -221.165 240.205 -220.835 ;
        RECT 239.875 -222.525 240.205 -222.195 ;
        RECT 239.875 -223.885 240.205 -223.555 ;
        RECT 239.875 -225.245 240.205 -224.915 ;
        RECT 239.875 -226.605 240.205 -226.275 ;
        RECT 239.875 -227.965 240.205 -227.635 ;
        RECT 239.875 -229.325 240.205 -228.995 ;
        RECT 239.875 -230.685 240.205 -230.355 ;
        RECT 239.875 -232.045 240.205 -231.715 ;
        RECT 239.875 -233.405 240.205 -233.075 ;
        RECT 239.875 -234.765 240.205 -234.435 ;
        RECT 239.875 -236.125 240.205 -235.795 ;
        RECT 239.875 -237.485 240.205 -237.155 ;
        RECT 239.875 -238.845 240.205 -238.515 ;
        RECT 239.875 -241.09 240.205 -239.96 ;
        RECT 239.88 -241.205 240.2 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 244.04 241.565 245.17 ;
        RECT 241.235 242.595 241.565 242.925 ;
        RECT 241.235 241.235 241.565 241.565 ;
        RECT 241.235 239.875 241.565 240.205 ;
        RECT 241.235 238.515 241.565 238.845 ;
        RECT 241.235 237.155 241.565 237.485 ;
        RECT 241.24 237.155 241.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 -0.845 241.565 -0.515 ;
        RECT 241.235 -2.205 241.565 -1.875 ;
        RECT 241.235 -3.565 241.565 -3.235 ;
        RECT 241.24 -3.565 241.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 -123.245 241.565 -122.915 ;
        RECT 241.235 -124.605 241.565 -124.275 ;
        RECT 241.235 -125.965 241.565 -125.635 ;
        RECT 241.235 -127.325 241.565 -126.995 ;
        RECT 241.235 -128.685 241.565 -128.355 ;
        RECT 241.235 -130.045 241.565 -129.715 ;
        RECT 241.235 -131.405 241.565 -131.075 ;
        RECT 241.235 -132.765 241.565 -132.435 ;
        RECT 241.235 -134.125 241.565 -133.795 ;
        RECT 241.235 -135.485 241.565 -135.155 ;
        RECT 241.235 -136.845 241.565 -136.515 ;
        RECT 241.235 -138.205 241.565 -137.875 ;
        RECT 241.235 -139.565 241.565 -139.235 ;
        RECT 241.235 -140.925 241.565 -140.595 ;
        RECT 241.235 -142.285 241.565 -141.955 ;
        RECT 241.235 -143.645 241.565 -143.315 ;
        RECT 241.235 -145.005 241.565 -144.675 ;
        RECT 241.235 -146.365 241.565 -146.035 ;
        RECT 241.235 -147.725 241.565 -147.395 ;
        RECT 241.235 -149.085 241.565 -148.755 ;
        RECT 241.235 -150.445 241.565 -150.115 ;
        RECT 241.235 -151.805 241.565 -151.475 ;
        RECT 241.235 -153.165 241.565 -152.835 ;
        RECT 241.235 -154.525 241.565 -154.195 ;
        RECT 241.235 -155.885 241.565 -155.555 ;
        RECT 241.235 -157.245 241.565 -156.915 ;
        RECT 241.235 -158.605 241.565 -158.275 ;
        RECT 241.235 -159.965 241.565 -159.635 ;
        RECT 241.235 -161.325 241.565 -160.995 ;
        RECT 241.235 -162.685 241.565 -162.355 ;
        RECT 241.235 -164.045 241.565 -163.715 ;
        RECT 241.235 -165.405 241.565 -165.075 ;
        RECT 241.235 -166.765 241.565 -166.435 ;
        RECT 241.235 -168.125 241.565 -167.795 ;
        RECT 241.235 -169.485 241.565 -169.155 ;
        RECT 241.235 -170.845 241.565 -170.515 ;
        RECT 241.235 -172.205 241.565 -171.875 ;
        RECT 241.235 -173.565 241.565 -173.235 ;
        RECT 241.235 -174.925 241.565 -174.595 ;
        RECT 241.235 -176.285 241.565 -175.955 ;
        RECT 241.235 -177.645 241.565 -177.315 ;
        RECT 241.235 -179.005 241.565 -178.675 ;
        RECT 241.235 -180.365 241.565 -180.035 ;
        RECT 241.235 -181.725 241.565 -181.395 ;
        RECT 241.235 -183.085 241.565 -182.755 ;
        RECT 241.235 -184.445 241.565 -184.115 ;
        RECT 241.235 -185.805 241.565 -185.475 ;
        RECT 241.235 -187.165 241.565 -186.835 ;
        RECT 241.235 -188.525 241.565 -188.195 ;
        RECT 241.235 -189.885 241.565 -189.555 ;
        RECT 241.235 -191.245 241.565 -190.915 ;
        RECT 241.235 -192.605 241.565 -192.275 ;
        RECT 241.235 -193.965 241.565 -193.635 ;
        RECT 241.235 -195.325 241.565 -194.995 ;
        RECT 241.235 -196.685 241.565 -196.355 ;
        RECT 241.235 -198.045 241.565 -197.715 ;
        RECT 241.235 -199.405 241.565 -199.075 ;
        RECT 241.235 -200.765 241.565 -200.435 ;
        RECT 241.235 -202.125 241.565 -201.795 ;
        RECT 241.235 -203.485 241.565 -203.155 ;
        RECT 241.235 -204.845 241.565 -204.515 ;
        RECT 241.235 -206.205 241.565 -205.875 ;
        RECT 241.235 -207.565 241.565 -207.235 ;
        RECT 241.235 -208.925 241.565 -208.595 ;
        RECT 241.235 -210.285 241.565 -209.955 ;
        RECT 241.235 -211.645 241.565 -211.315 ;
        RECT 241.235 -213.005 241.565 -212.675 ;
        RECT 241.235 -214.365 241.565 -214.035 ;
        RECT 241.235 -215.725 241.565 -215.395 ;
        RECT 241.235 -217.085 241.565 -216.755 ;
        RECT 241.235 -218.445 241.565 -218.115 ;
        RECT 241.235 -219.805 241.565 -219.475 ;
        RECT 241.235 -221.165 241.565 -220.835 ;
        RECT 241.235 -222.525 241.565 -222.195 ;
        RECT 241.235 -223.885 241.565 -223.555 ;
        RECT 241.235 -225.245 241.565 -224.915 ;
        RECT 241.235 -226.605 241.565 -226.275 ;
        RECT 241.235 -227.965 241.565 -227.635 ;
        RECT 241.235 -229.325 241.565 -228.995 ;
        RECT 241.235 -230.685 241.565 -230.355 ;
        RECT 241.235 -232.045 241.565 -231.715 ;
        RECT 241.235 -233.405 241.565 -233.075 ;
        RECT 241.235 -234.765 241.565 -234.435 ;
        RECT 241.235 -236.125 241.565 -235.795 ;
        RECT 241.235 -237.485 241.565 -237.155 ;
        RECT 241.235 -238.845 241.565 -238.515 ;
        RECT 241.235 -241.09 241.565 -239.96 ;
        RECT 241.24 -241.205 241.56 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 244.04 242.925 245.17 ;
        RECT 242.595 242.595 242.925 242.925 ;
        RECT 242.595 241.235 242.925 241.565 ;
        RECT 242.595 239.875 242.925 240.205 ;
        RECT 242.595 238.515 242.925 238.845 ;
        RECT 242.595 237.155 242.925 237.485 ;
        RECT 242.6 237.155 242.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 -127.325 242.925 -126.995 ;
        RECT 242.595 -128.685 242.925 -128.355 ;
        RECT 242.595 -130.045 242.925 -129.715 ;
        RECT 242.595 -131.405 242.925 -131.075 ;
        RECT 242.595 -132.765 242.925 -132.435 ;
        RECT 242.595 -134.125 242.925 -133.795 ;
        RECT 242.595 -135.485 242.925 -135.155 ;
        RECT 242.595 -136.845 242.925 -136.515 ;
        RECT 242.595 -138.205 242.925 -137.875 ;
        RECT 242.595 -139.565 242.925 -139.235 ;
        RECT 242.595 -140.925 242.925 -140.595 ;
        RECT 242.595 -142.285 242.925 -141.955 ;
        RECT 242.595 -143.645 242.925 -143.315 ;
        RECT 242.595 -145.005 242.925 -144.675 ;
        RECT 242.595 -146.365 242.925 -146.035 ;
        RECT 242.595 -147.725 242.925 -147.395 ;
        RECT 242.595 -149.085 242.925 -148.755 ;
        RECT 242.595 -150.445 242.925 -150.115 ;
        RECT 242.595 -151.805 242.925 -151.475 ;
        RECT 242.595 -153.165 242.925 -152.835 ;
        RECT 242.595 -154.525 242.925 -154.195 ;
        RECT 242.595 -155.885 242.925 -155.555 ;
        RECT 242.595 -157.245 242.925 -156.915 ;
        RECT 242.595 -158.605 242.925 -158.275 ;
        RECT 242.595 -159.965 242.925 -159.635 ;
        RECT 242.595 -161.325 242.925 -160.995 ;
        RECT 242.595 -162.685 242.925 -162.355 ;
        RECT 242.595 -164.045 242.925 -163.715 ;
        RECT 242.595 -165.405 242.925 -165.075 ;
        RECT 242.595 -166.765 242.925 -166.435 ;
        RECT 242.595 -168.125 242.925 -167.795 ;
        RECT 242.595 -169.485 242.925 -169.155 ;
        RECT 242.595 -170.845 242.925 -170.515 ;
        RECT 242.595 -172.205 242.925 -171.875 ;
        RECT 242.595 -173.565 242.925 -173.235 ;
        RECT 242.595 -174.925 242.925 -174.595 ;
        RECT 242.595 -176.285 242.925 -175.955 ;
        RECT 242.595 -177.645 242.925 -177.315 ;
        RECT 242.595 -179.005 242.925 -178.675 ;
        RECT 242.595 -180.365 242.925 -180.035 ;
        RECT 242.595 -181.725 242.925 -181.395 ;
        RECT 242.595 -183.085 242.925 -182.755 ;
        RECT 242.595 -184.445 242.925 -184.115 ;
        RECT 242.595 -185.805 242.925 -185.475 ;
        RECT 242.595 -187.165 242.925 -186.835 ;
        RECT 242.595 -188.525 242.925 -188.195 ;
        RECT 242.595 -189.885 242.925 -189.555 ;
        RECT 242.595 -191.245 242.925 -190.915 ;
        RECT 242.595 -192.605 242.925 -192.275 ;
        RECT 242.595 -193.965 242.925 -193.635 ;
        RECT 242.595 -195.325 242.925 -194.995 ;
        RECT 242.595 -196.685 242.925 -196.355 ;
        RECT 242.595 -198.045 242.925 -197.715 ;
        RECT 242.595 -199.405 242.925 -199.075 ;
        RECT 242.595 -200.765 242.925 -200.435 ;
        RECT 242.595 -202.125 242.925 -201.795 ;
        RECT 242.595 -203.485 242.925 -203.155 ;
        RECT 242.595 -204.845 242.925 -204.515 ;
        RECT 242.595 -206.205 242.925 -205.875 ;
        RECT 242.595 -207.565 242.925 -207.235 ;
        RECT 242.595 -208.925 242.925 -208.595 ;
        RECT 242.595 -210.285 242.925 -209.955 ;
        RECT 242.595 -211.645 242.925 -211.315 ;
        RECT 242.595 -213.005 242.925 -212.675 ;
        RECT 242.595 -214.365 242.925 -214.035 ;
        RECT 242.595 -215.725 242.925 -215.395 ;
        RECT 242.595 -217.085 242.925 -216.755 ;
        RECT 242.595 -218.445 242.925 -218.115 ;
        RECT 242.595 -219.805 242.925 -219.475 ;
        RECT 242.595 -221.165 242.925 -220.835 ;
        RECT 242.595 -222.525 242.925 -222.195 ;
        RECT 242.595 -223.885 242.925 -223.555 ;
        RECT 242.595 -225.245 242.925 -224.915 ;
        RECT 242.595 -226.605 242.925 -226.275 ;
        RECT 242.595 -227.965 242.925 -227.635 ;
        RECT 242.595 -229.325 242.925 -228.995 ;
        RECT 242.595 -230.685 242.925 -230.355 ;
        RECT 242.595 -232.045 242.925 -231.715 ;
        RECT 242.595 -233.405 242.925 -233.075 ;
        RECT 242.595 -234.765 242.925 -234.435 ;
        RECT 242.595 -236.125 242.925 -235.795 ;
        RECT 242.595 -237.485 242.925 -237.155 ;
        RECT 242.595 -238.845 242.925 -238.515 ;
        RECT 242.595 -241.09 242.925 -239.96 ;
        RECT 242.6 -241.205 242.92 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.11 -125.535 243.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 244.04 244.285 245.17 ;
        RECT 243.955 242.595 244.285 242.925 ;
        RECT 243.955 241.235 244.285 241.565 ;
        RECT 243.955 239.875 244.285 240.205 ;
        RECT 243.955 238.515 244.285 238.845 ;
        RECT 243.955 237.155 244.285 237.485 ;
        RECT 243.96 237.155 244.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 -0.845 244.285 -0.515 ;
        RECT 243.955 -2.205 244.285 -1.875 ;
        RECT 243.955 -3.565 244.285 -3.235 ;
        RECT 243.96 -3.565 244.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 244.04 245.645 245.17 ;
        RECT 245.315 242.595 245.645 242.925 ;
        RECT 245.315 241.235 245.645 241.565 ;
        RECT 245.315 239.875 245.645 240.205 ;
        RECT 245.315 238.515 245.645 238.845 ;
        RECT 245.315 237.155 245.645 237.485 ;
        RECT 245.32 237.155 245.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 -0.845 245.645 -0.515 ;
        RECT 245.315 -2.205 245.645 -1.875 ;
        RECT 245.315 -3.565 245.645 -3.235 ;
        RECT 245.32 -3.565 245.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 244.04 247.005 245.17 ;
        RECT 246.675 242.595 247.005 242.925 ;
        RECT 246.675 241.235 247.005 241.565 ;
        RECT 246.675 239.875 247.005 240.205 ;
        RECT 246.675 238.515 247.005 238.845 ;
        RECT 246.675 237.155 247.005 237.485 ;
        RECT 246.68 237.155 247 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 -0.845 247.005 -0.515 ;
        RECT 246.675 -2.205 247.005 -1.875 ;
        RECT 246.675 -3.565 247.005 -3.235 ;
        RECT 246.68 -3.565 247 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 -123.245 247.005 -122.915 ;
        RECT 246.675 -124.605 247.005 -124.275 ;
        RECT 246.675 -125.965 247.005 -125.635 ;
        RECT 246.675 -127.325 247.005 -126.995 ;
        RECT 246.675 -128.685 247.005 -128.355 ;
        RECT 246.675 -130.045 247.005 -129.715 ;
        RECT 246.675 -131.405 247.005 -131.075 ;
        RECT 246.675 -132.765 247.005 -132.435 ;
        RECT 246.675 -134.125 247.005 -133.795 ;
        RECT 246.675 -135.485 247.005 -135.155 ;
        RECT 246.675 -136.845 247.005 -136.515 ;
        RECT 246.675 -138.205 247.005 -137.875 ;
        RECT 246.675 -139.565 247.005 -139.235 ;
        RECT 246.675 -140.925 247.005 -140.595 ;
        RECT 246.675 -142.285 247.005 -141.955 ;
        RECT 246.675 -143.645 247.005 -143.315 ;
        RECT 246.675 -145.005 247.005 -144.675 ;
        RECT 246.675 -146.365 247.005 -146.035 ;
        RECT 246.675 -147.725 247.005 -147.395 ;
        RECT 246.675 -149.085 247.005 -148.755 ;
        RECT 246.675 -150.445 247.005 -150.115 ;
        RECT 246.675 -151.805 247.005 -151.475 ;
        RECT 246.675 -153.165 247.005 -152.835 ;
        RECT 246.675 -154.525 247.005 -154.195 ;
        RECT 246.675 -155.885 247.005 -155.555 ;
        RECT 246.675 -157.245 247.005 -156.915 ;
        RECT 246.675 -158.605 247.005 -158.275 ;
        RECT 246.675 -159.965 247.005 -159.635 ;
        RECT 246.675 -161.325 247.005 -160.995 ;
        RECT 246.675 -162.685 247.005 -162.355 ;
        RECT 246.675 -164.045 247.005 -163.715 ;
        RECT 246.675 -165.405 247.005 -165.075 ;
        RECT 246.675 -166.765 247.005 -166.435 ;
        RECT 246.675 -168.125 247.005 -167.795 ;
        RECT 246.675 -169.485 247.005 -169.155 ;
        RECT 246.675 -170.845 247.005 -170.515 ;
        RECT 246.675 -172.205 247.005 -171.875 ;
        RECT 246.675 -173.565 247.005 -173.235 ;
        RECT 246.675 -174.925 247.005 -174.595 ;
        RECT 246.675 -176.285 247.005 -175.955 ;
        RECT 246.675 -177.645 247.005 -177.315 ;
        RECT 246.675 -179.005 247.005 -178.675 ;
        RECT 246.675 -180.365 247.005 -180.035 ;
        RECT 246.675 -181.725 247.005 -181.395 ;
        RECT 246.675 -183.085 247.005 -182.755 ;
        RECT 246.675 -184.445 247.005 -184.115 ;
        RECT 246.675 -185.805 247.005 -185.475 ;
        RECT 246.675 -187.165 247.005 -186.835 ;
        RECT 246.675 -188.525 247.005 -188.195 ;
        RECT 246.675 -189.885 247.005 -189.555 ;
        RECT 246.675 -191.245 247.005 -190.915 ;
        RECT 246.675 -192.605 247.005 -192.275 ;
        RECT 246.675 -193.965 247.005 -193.635 ;
        RECT 246.675 -195.325 247.005 -194.995 ;
        RECT 246.675 -196.685 247.005 -196.355 ;
        RECT 246.675 -198.045 247.005 -197.715 ;
        RECT 246.675 -199.405 247.005 -199.075 ;
        RECT 246.675 -200.765 247.005 -200.435 ;
        RECT 246.675 -202.125 247.005 -201.795 ;
        RECT 246.675 -203.485 247.005 -203.155 ;
        RECT 246.675 -204.845 247.005 -204.515 ;
        RECT 246.675 -206.205 247.005 -205.875 ;
        RECT 246.675 -207.565 247.005 -207.235 ;
        RECT 246.675 -208.925 247.005 -208.595 ;
        RECT 246.675 -210.285 247.005 -209.955 ;
        RECT 246.675 -211.645 247.005 -211.315 ;
        RECT 246.675 -213.005 247.005 -212.675 ;
        RECT 246.675 -214.365 247.005 -214.035 ;
        RECT 246.675 -215.725 247.005 -215.395 ;
        RECT 246.675 -217.085 247.005 -216.755 ;
        RECT 246.675 -218.445 247.005 -218.115 ;
        RECT 246.675 -219.805 247.005 -219.475 ;
        RECT 246.675 -221.165 247.005 -220.835 ;
        RECT 246.675 -222.525 247.005 -222.195 ;
        RECT 246.675 -223.885 247.005 -223.555 ;
        RECT 246.675 -225.245 247.005 -224.915 ;
        RECT 246.675 -226.605 247.005 -226.275 ;
        RECT 246.675 -227.965 247.005 -227.635 ;
        RECT 246.675 -229.325 247.005 -228.995 ;
        RECT 246.675 -230.685 247.005 -230.355 ;
        RECT 246.675 -232.045 247.005 -231.715 ;
        RECT 246.675 -233.405 247.005 -233.075 ;
        RECT 246.675 -234.765 247.005 -234.435 ;
        RECT 246.675 -236.125 247.005 -235.795 ;
        RECT 246.675 -237.485 247.005 -237.155 ;
        RECT 246.675 -238.845 247.005 -238.515 ;
        RECT 246.675 -241.09 247.005 -239.96 ;
        RECT 246.68 -241.205 247 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 244.04 248.365 245.17 ;
        RECT 248.035 242.595 248.365 242.925 ;
        RECT 248.035 241.235 248.365 241.565 ;
        RECT 248.035 239.875 248.365 240.205 ;
        RECT 248.035 238.515 248.365 238.845 ;
        RECT 248.035 237.155 248.365 237.485 ;
        RECT 248.04 237.155 248.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 -0.845 248.365 -0.515 ;
        RECT 248.035 -2.205 248.365 -1.875 ;
        RECT 248.035 -3.565 248.365 -3.235 ;
        RECT 248.04 -3.565 248.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 -123.245 248.365 -122.915 ;
        RECT 248.035 -124.605 248.365 -124.275 ;
        RECT 248.035 -125.965 248.365 -125.635 ;
        RECT 248.035 -127.325 248.365 -126.995 ;
        RECT 248.035 -128.685 248.365 -128.355 ;
        RECT 248.035 -130.045 248.365 -129.715 ;
        RECT 248.035 -131.405 248.365 -131.075 ;
        RECT 248.035 -132.765 248.365 -132.435 ;
        RECT 248.035 -134.125 248.365 -133.795 ;
        RECT 248.035 -135.485 248.365 -135.155 ;
        RECT 248.035 -136.845 248.365 -136.515 ;
        RECT 248.035 -138.205 248.365 -137.875 ;
        RECT 248.035 -139.565 248.365 -139.235 ;
        RECT 248.035 -140.925 248.365 -140.595 ;
        RECT 248.035 -142.285 248.365 -141.955 ;
        RECT 248.035 -143.645 248.365 -143.315 ;
        RECT 248.035 -145.005 248.365 -144.675 ;
        RECT 248.035 -146.365 248.365 -146.035 ;
        RECT 248.035 -147.725 248.365 -147.395 ;
        RECT 248.035 -149.085 248.365 -148.755 ;
        RECT 248.035 -150.445 248.365 -150.115 ;
        RECT 248.035 -151.805 248.365 -151.475 ;
        RECT 248.035 -153.165 248.365 -152.835 ;
        RECT 248.035 -154.525 248.365 -154.195 ;
        RECT 248.035 -155.885 248.365 -155.555 ;
        RECT 248.035 -157.245 248.365 -156.915 ;
        RECT 248.035 -158.605 248.365 -158.275 ;
        RECT 248.035 -159.965 248.365 -159.635 ;
        RECT 248.035 -161.325 248.365 -160.995 ;
        RECT 248.035 -162.685 248.365 -162.355 ;
        RECT 248.035 -164.045 248.365 -163.715 ;
        RECT 248.035 -165.405 248.365 -165.075 ;
        RECT 248.035 -166.765 248.365 -166.435 ;
        RECT 248.035 -168.125 248.365 -167.795 ;
        RECT 248.035 -169.485 248.365 -169.155 ;
        RECT 248.035 -170.845 248.365 -170.515 ;
        RECT 248.035 -172.205 248.365 -171.875 ;
        RECT 248.035 -173.565 248.365 -173.235 ;
        RECT 248.035 -174.925 248.365 -174.595 ;
        RECT 248.035 -176.285 248.365 -175.955 ;
        RECT 248.035 -177.645 248.365 -177.315 ;
        RECT 248.035 -179.005 248.365 -178.675 ;
        RECT 248.035 -180.365 248.365 -180.035 ;
        RECT 248.035 -181.725 248.365 -181.395 ;
        RECT 248.035 -183.085 248.365 -182.755 ;
        RECT 248.035 -184.445 248.365 -184.115 ;
        RECT 248.035 -185.805 248.365 -185.475 ;
        RECT 248.035 -187.165 248.365 -186.835 ;
        RECT 248.035 -188.525 248.365 -188.195 ;
        RECT 248.035 -189.885 248.365 -189.555 ;
        RECT 248.035 -191.245 248.365 -190.915 ;
        RECT 248.035 -192.605 248.365 -192.275 ;
        RECT 248.035 -193.965 248.365 -193.635 ;
        RECT 248.035 -195.325 248.365 -194.995 ;
        RECT 248.035 -196.685 248.365 -196.355 ;
        RECT 248.035 -198.045 248.365 -197.715 ;
        RECT 248.035 -199.405 248.365 -199.075 ;
        RECT 248.035 -200.765 248.365 -200.435 ;
        RECT 248.035 -202.125 248.365 -201.795 ;
        RECT 248.035 -203.485 248.365 -203.155 ;
        RECT 248.035 -204.845 248.365 -204.515 ;
        RECT 248.035 -206.205 248.365 -205.875 ;
        RECT 248.035 -207.565 248.365 -207.235 ;
        RECT 248.035 -208.925 248.365 -208.595 ;
        RECT 248.035 -210.285 248.365 -209.955 ;
        RECT 248.035 -211.645 248.365 -211.315 ;
        RECT 248.035 -213.005 248.365 -212.675 ;
        RECT 248.035 -214.365 248.365 -214.035 ;
        RECT 248.035 -215.725 248.365 -215.395 ;
        RECT 248.035 -217.085 248.365 -216.755 ;
        RECT 248.035 -218.445 248.365 -218.115 ;
        RECT 248.035 -219.805 248.365 -219.475 ;
        RECT 248.035 -221.165 248.365 -220.835 ;
        RECT 248.035 -222.525 248.365 -222.195 ;
        RECT 248.035 -223.885 248.365 -223.555 ;
        RECT 248.035 -225.245 248.365 -224.915 ;
        RECT 248.035 -226.605 248.365 -226.275 ;
        RECT 248.035 -227.965 248.365 -227.635 ;
        RECT 248.035 -229.325 248.365 -228.995 ;
        RECT 248.035 -230.685 248.365 -230.355 ;
        RECT 248.035 -232.045 248.365 -231.715 ;
        RECT 248.035 -233.405 248.365 -233.075 ;
        RECT 248.035 -234.765 248.365 -234.435 ;
        RECT 248.035 -236.125 248.365 -235.795 ;
        RECT 248.035 -237.485 248.365 -237.155 ;
        RECT 248.035 -238.845 248.365 -238.515 ;
        RECT 248.035 -241.09 248.365 -239.96 ;
        RECT 248.04 -241.205 248.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 244.04 249.725 245.17 ;
        RECT 249.395 242.595 249.725 242.925 ;
        RECT 249.395 241.235 249.725 241.565 ;
        RECT 249.395 239.875 249.725 240.205 ;
        RECT 249.395 238.515 249.725 238.845 ;
        RECT 249.395 237.155 249.725 237.485 ;
        RECT 249.4 237.155 249.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 -0.845 249.725 -0.515 ;
        RECT 249.395 -2.205 249.725 -1.875 ;
        RECT 249.395 -3.565 249.725 -3.235 ;
        RECT 249.4 -3.565 249.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 -123.245 249.725 -122.915 ;
        RECT 249.395 -124.605 249.725 -124.275 ;
        RECT 249.395 -125.965 249.725 -125.635 ;
        RECT 249.395 -127.325 249.725 -126.995 ;
        RECT 249.395 -128.685 249.725 -128.355 ;
        RECT 249.395 -130.045 249.725 -129.715 ;
        RECT 249.395 -131.405 249.725 -131.075 ;
        RECT 249.395 -132.765 249.725 -132.435 ;
        RECT 249.395 -134.125 249.725 -133.795 ;
        RECT 249.395 -135.485 249.725 -135.155 ;
        RECT 249.395 -136.845 249.725 -136.515 ;
        RECT 249.395 -138.205 249.725 -137.875 ;
        RECT 249.395 -139.565 249.725 -139.235 ;
        RECT 249.395 -140.925 249.725 -140.595 ;
        RECT 249.395 -142.285 249.725 -141.955 ;
        RECT 249.395 -143.645 249.725 -143.315 ;
        RECT 249.395 -145.005 249.725 -144.675 ;
        RECT 249.395 -146.365 249.725 -146.035 ;
        RECT 249.395 -147.725 249.725 -147.395 ;
        RECT 249.395 -149.085 249.725 -148.755 ;
        RECT 249.395 -150.445 249.725 -150.115 ;
        RECT 249.395 -151.805 249.725 -151.475 ;
        RECT 249.395 -153.165 249.725 -152.835 ;
        RECT 249.395 -154.525 249.725 -154.195 ;
        RECT 249.395 -155.885 249.725 -155.555 ;
        RECT 249.395 -157.245 249.725 -156.915 ;
        RECT 249.395 -158.605 249.725 -158.275 ;
        RECT 249.395 -159.965 249.725 -159.635 ;
        RECT 249.395 -161.325 249.725 -160.995 ;
        RECT 249.395 -162.685 249.725 -162.355 ;
        RECT 249.395 -164.045 249.725 -163.715 ;
        RECT 249.395 -165.405 249.725 -165.075 ;
        RECT 249.395 -166.765 249.725 -166.435 ;
        RECT 249.395 -168.125 249.725 -167.795 ;
        RECT 249.395 -169.485 249.725 -169.155 ;
        RECT 249.395 -170.845 249.725 -170.515 ;
        RECT 249.395 -172.205 249.725 -171.875 ;
        RECT 249.395 -173.565 249.725 -173.235 ;
        RECT 249.395 -174.925 249.725 -174.595 ;
        RECT 249.395 -176.285 249.725 -175.955 ;
        RECT 249.395 -177.645 249.725 -177.315 ;
        RECT 249.395 -179.005 249.725 -178.675 ;
        RECT 249.395 -180.365 249.725 -180.035 ;
        RECT 249.395 -181.725 249.725 -181.395 ;
        RECT 249.395 -183.085 249.725 -182.755 ;
        RECT 249.395 -184.445 249.725 -184.115 ;
        RECT 249.395 -185.805 249.725 -185.475 ;
        RECT 249.395 -187.165 249.725 -186.835 ;
        RECT 249.395 -188.525 249.725 -188.195 ;
        RECT 249.395 -189.885 249.725 -189.555 ;
        RECT 249.395 -191.245 249.725 -190.915 ;
        RECT 249.395 -192.605 249.725 -192.275 ;
        RECT 249.395 -193.965 249.725 -193.635 ;
        RECT 249.395 -195.325 249.725 -194.995 ;
        RECT 249.395 -196.685 249.725 -196.355 ;
        RECT 249.395 -198.045 249.725 -197.715 ;
        RECT 249.395 -199.405 249.725 -199.075 ;
        RECT 249.395 -200.765 249.725 -200.435 ;
        RECT 249.395 -202.125 249.725 -201.795 ;
        RECT 249.395 -203.485 249.725 -203.155 ;
        RECT 249.395 -204.845 249.725 -204.515 ;
        RECT 249.395 -206.205 249.725 -205.875 ;
        RECT 249.395 -207.565 249.725 -207.235 ;
        RECT 249.395 -208.925 249.725 -208.595 ;
        RECT 249.395 -210.285 249.725 -209.955 ;
        RECT 249.395 -211.645 249.725 -211.315 ;
        RECT 249.395 -213.005 249.725 -212.675 ;
        RECT 249.395 -214.365 249.725 -214.035 ;
        RECT 249.395 -215.725 249.725 -215.395 ;
        RECT 249.395 -217.085 249.725 -216.755 ;
        RECT 249.395 -218.445 249.725 -218.115 ;
        RECT 249.395 -219.805 249.725 -219.475 ;
        RECT 249.395 -221.165 249.725 -220.835 ;
        RECT 249.395 -222.525 249.725 -222.195 ;
        RECT 249.395 -223.885 249.725 -223.555 ;
        RECT 249.395 -225.245 249.725 -224.915 ;
        RECT 249.395 -226.605 249.725 -226.275 ;
        RECT 249.395 -227.965 249.725 -227.635 ;
        RECT 249.395 -229.325 249.725 -228.995 ;
        RECT 249.395 -230.685 249.725 -230.355 ;
        RECT 249.395 -232.045 249.725 -231.715 ;
        RECT 249.395 -233.405 249.725 -233.075 ;
        RECT 249.395 -234.765 249.725 -234.435 ;
        RECT 249.395 -236.125 249.725 -235.795 ;
        RECT 249.395 -237.485 249.725 -237.155 ;
        RECT 249.395 -238.845 249.725 -238.515 ;
        RECT 249.395 -241.09 249.725 -239.96 ;
        RECT 249.4 -241.205 249.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 244.04 251.085 245.17 ;
        RECT 250.755 242.595 251.085 242.925 ;
        RECT 250.755 241.235 251.085 241.565 ;
        RECT 250.755 239.875 251.085 240.205 ;
        RECT 250.755 238.515 251.085 238.845 ;
        RECT 250.755 237.155 251.085 237.485 ;
        RECT 250.76 237.155 251.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 -0.845 251.085 -0.515 ;
        RECT 250.755 -2.205 251.085 -1.875 ;
        RECT 250.755 -3.565 251.085 -3.235 ;
        RECT 250.76 -3.565 251.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 -123.245 251.085 -122.915 ;
        RECT 250.755 -124.605 251.085 -124.275 ;
        RECT 250.755 -125.965 251.085 -125.635 ;
        RECT 250.755 -127.325 251.085 -126.995 ;
        RECT 250.755 -128.685 251.085 -128.355 ;
        RECT 250.755 -130.045 251.085 -129.715 ;
        RECT 250.755 -131.405 251.085 -131.075 ;
        RECT 250.755 -132.765 251.085 -132.435 ;
        RECT 250.755 -134.125 251.085 -133.795 ;
        RECT 250.755 -135.485 251.085 -135.155 ;
        RECT 250.755 -136.845 251.085 -136.515 ;
        RECT 250.755 -138.205 251.085 -137.875 ;
        RECT 250.755 -139.565 251.085 -139.235 ;
        RECT 250.755 -140.925 251.085 -140.595 ;
        RECT 250.755 -142.285 251.085 -141.955 ;
        RECT 250.755 -143.645 251.085 -143.315 ;
        RECT 250.755 -145.005 251.085 -144.675 ;
        RECT 250.755 -146.365 251.085 -146.035 ;
        RECT 250.755 -147.725 251.085 -147.395 ;
        RECT 250.755 -149.085 251.085 -148.755 ;
        RECT 250.755 -150.445 251.085 -150.115 ;
        RECT 250.755 -151.805 251.085 -151.475 ;
        RECT 250.755 -153.165 251.085 -152.835 ;
        RECT 250.755 -154.525 251.085 -154.195 ;
        RECT 250.755 -155.885 251.085 -155.555 ;
        RECT 250.755 -157.245 251.085 -156.915 ;
        RECT 250.755 -158.605 251.085 -158.275 ;
        RECT 250.755 -159.965 251.085 -159.635 ;
        RECT 250.755 -161.325 251.085 -160.995 ;
        RECT 250.755 -162.685 251.085 -162.355 ;
        RECT 250.755 -164.045 251.085 -163.715 ;
        RECT 250.755 -165.405 251.085 -165.075 ;
        RECT 250.755 -166.765 251.085 -166.435 ;
        RECT 250.755 -168.125 251.085 -167.795 ;
        RECT 250.755 -169.485 251.085 -169.155 ;
        RECT 250.755 -170.845 251.085 -170.515 ;
        RECT 250.755 -172.205 251.085 -171.875 ;
        RECT 250.755 -173.565 251.085 -173.235 ;
        RECT 250.755 -174.925 251.085 -174.595 ;
        RECT 250.755 -176.285 251.085 -175.955 ;
        RECT 250.755 -177.645 251.085 -177.315 ;
        RECT 250.755 -179.005 251.085 -178.675 ;
        RECT 250.755 -180.365 251.085 -180.035 ;
        RECT 250.755 -181.725 251.085 -181.395 ;
        RECT 250.755 -183.085 251.085 -182.755 ;
        RECT 250.755 -184.445 251.085 -184.115 ;
        RECT 250.755 -185.805 251.085 -185.475 ;
        RECT 250.755 -187.165 251.085 -186.835 ;
        RECT 250.755 -188.525 251.085 -188.195 ;
        RECT 250.755 -189.885 251.085 -189.555 ;
        RECT 250.755 -191.245 251.085 -190.915 ;
        RECT 250.755 -192.605 251.085 -192.275 ;
        RECT 250.755 -193.965 251.085 -193.635 ;
        RECT 250.755 -195.325 251.085 -194.995 ;
        RECT 250.755 -196.685 251.085 -196.355 ;
        RECT 250.755 -198.045 251.085 -197.715 ;
        RECT 250.755 -199.405 251.085 -199.075 ;
        RECT 250.755 -200.765 251.085 -200.435 ;
        RECT 250.755 -202.125 251.085 -201.795 ;
        RECT 250.755 -203.485 251.085 -203.155 ;
        RECT 250.755 -204.845 251.085 -204.515 ;
        RECT 250.755 -206.205 251.085 -205.875 ;
        RECT 250.755 -207.565 251.085 -207.235 ;
        RECT 250.755 -208.925 251.085 -208.595 ;
        RECT 250.755 -210.285 251.085 -209.955 ;
        RECT 250.755 -211.645 251.085 -211.315 ;
        RECT 250.755 -213.005 251.085 -212.675 ;
        RECT 250.755 -214.365 251.085 -214.035 ;
        RECT 250.755 -215.725 251.085 -215.395 ;
        RECT 250.755 -217.085 251.085 -216.755 ;
        RECT 250.755 -218.445 251.085 -218.115 ;
        RECT 250.755 -219.805 251.085 -219.475 ;
        RECT 250.755 -221.165 251.085 -220.835 ;
        RECT 250.755 -222.525 251.085 -222.195 ;
        RECT 250.755 -223.885 251.085 -223.555 ;
        RECT 250.755 -225.245 251.085 -224.915 ;
        RECT 250.755 -226.605 251.085 -226.275 ;
        RECT 250.755 -227.965 251.085 -227.635 ;
        RECT 250.755 -229.325 251.085 -228.995 ;
        RECT 250.755 -230.685 251.085 -230.355 ;
        RECT 250.755 -232.045 251.085 -231.715 ;
        RECT 250.755 -233.405 251.085 -233.075 ;
        RECT 250.755 -234.765 251.085 -234.435 ;
        RECT 250.755 -236.125 251.085 -235.795 ;
        RECT 250.755 -237.485 251.085 -237.155 ;
        RECT 250.755 -238.845 251.085 -238.515 ;
        RECT 250.755 -241.09 251.085 -239.96 ;
        RECT 250.76 -241.205 251.08 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 244.04 252.445 245.17 ;
        RECT 252.115 242.595 252.445 242.925 ;
        RECT 252.115 241.235 252.445 241.565 ;
        RECT 252.115 239.875 252.445 240.205 ;
        RECT 252.115 238.515 252.445 238.845 ;
        RECT 252.115 237.155 252.445 237.485 ;
        RECT 252.12 237.155 252.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 -0.845 252.445 -0.515 ;
        RECT 252.115 -2.205 252.445 -1.875 ;
        RECT 252.115 -3.565 252.445 -3.235 ;
        RECT 252.12 -3.565 252.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 -123.245 252.445 -122.915 ;
        RECT 252.115 -124.605 252.445 -124.275 ;
        RECT 252.115 -125.965 252.445 -125.635 ;
        RECT 252.115 -127.325 252.445 -126.995 ;
        RECT 252.115 -128.685 252.445 -128.355 ;
        RECT 252.115 -130.045 252.445 -129.715 ;
        RECT 252.115 -131.405 252.445 -131.075 ;
        RECT 252.115 -132.765 252.445 -132.435 ;
        RECT 252.115 -134.125 252.445 -133.795 ;
        RECT 252.115 -135.485 252.445 -135.155 ;
        RECT 252.115 -136.845 252.445 -136.515 ;
        RECT 252.115 -138.205 252.445 -137.875 ;
        RECT 252.115 -139.565 252.445 -139.235 ;
        RECT 252.115 -140.925 252.445 -140.595 ;
        RECT 252.115 -142.285 252.445 -141.955 ;
        RECT 252.115 -143.645 252.445 -143.315 ;
        RECT 252.115 -145.005 252.445 -144.675 ;
        RECT 252.115 -146.365 252.445 -146.035 ;
        RECT 252.115 -147.725 252.445 -147.395 ;
        RECT 252.115 -149.085 252.445 -148.755 ;
        RECT 252.115 -150.445 252.445 -150.115 ;
        RECT 252.115 -151.805 252.445 -151.475 ;
        RECT 252.115 -153.165 252.445 -152.835 ;
        RECT 252.115 -154.525 252.445 -154.195 ;
        RECT 252.115 -155.885 252.445 -155.555 ;
        RECT 252.115 -157.245 252.445 -156.915 ;
        RECT 252.115 -158.605 252.445 -158.275 ;
        RECT 252.115 -159.965 252.445 -159.635 ;
        RECT 252.115 -161.325 252.445 -160.995 ;
        RECT 252.115 -162.685 252.445 -162.355 ;
        RECT 252.115 -164.045 252.445 -163.715 ;
        RECT 252.115 -165.405 252.445 -165.075 ;
        RECT 252.115 -166.765 252.445 -166.435 ;
        RECT 252.115 -168.125 252.445 -167.795 ;
        RECT 252.115 -169.485 252.445 -169.155 ;
        RECT 252.115 -170.845 252.445 -170.515 ;
        RECT 252.115 -172.205 252.445 -171.875 ;
        RECT 252.115 -173.565 252.445 -173.235 ;
        RECT 252.115 -174.925 252.445 -174.595 ;
        RECT 252.115 -176.285 252.445 -175.955 ;
        RECT 252.115 -177.645 252.445 -177.315 ;
        RECT 252.115 -179.005 252.445 -178.675 ;
        RECT 252.115 -180.365 252.445 -180.035 ;
        RECT 252.115 -181.725 252.445 -181.395 ;
        RECT 252.115 -183.085 252.445 -182.755 ;
        RECT 252.115 -184.445 252.445 -184.115 ;
        RECT 252.115 -185.805 252.445 -185.475 ;
        RECT 252.115 -187.165 252.445 -186.835 ;
        RECT 252.115 -188.525 252.445 -188.195 ;
        RECT 252.115 -189.885 252.445 -189.555 ;
        RECT 252.115 -191.245 252.445 -190.915 ;
        RECT 252.115 -192.605 252.445 -192.275 ;
        RECT 252.115 -193.965 252.445 -193.635 ;
        RECT 252.115 -195.325 252.445 -194.995 ;
        RECT 252.115 -196.685 252.445 -196.355 ;
        RECT 252.115 -198.045 252.445 -197.715 ;
        RECT 252.115 -199.405 252.445 -199.075 ;
        RECT 252.115 -200.765 252.445 -200.435 ;
        RECT 252.115 -202.125 252.445 -201.795 ;
        RECT 252.115 -203.485 252.445 -203.155 ;
        RECT 252.115 -204.845 252.445 -204.515 ;
        RECT 252.115 -206.205 252.445 -205.875 ;
        RECT 252.115 -207.565 252.445 -207.235 ;
        RECT 252.115 -208.925 252.445 -208.595 ;
        RECT 252.115 -210.285 252.445 -209.955 ;
        RECT 252.115 -211.645 252.445 -211.315 ;
        RECT 252.115 -213.005 252.445 -212.675 ;
        RECT 252.115 -214.365 252.445 -214.035 ;
        RECT 252.115 -215.725 252.445 -215.395 ;
        RECT 252.115 -217.085 252.445 -216.755 ;
        RECT 252.115 -218.445 252.445 -218.115 ;
        RECT 252.115 -219.805 252.445 -219.475 ;
        RECT 252.115 -221.165 252.445 -220.835 ;
        RECT 252.115 -222.525 252.445 -222.195 ;
        RECT 252.115 -223.885 252.445 -223.555 ;
        RECT 252.115 -225.245 252.445 -224.915 ;
        RECT 252.115 -226.605 252.445 -226.275 ;
        RECT 252.115 -227.965 252.445 -227.635 ;
        RECT 252.115 -229.325 252.445 -228.995 ;
        RECT 252.115 -230.685 252.445 -230.355 ;
        RECT 252.115 -232.045 252.445 -231.715 ;
        RECT 252.115 -233.405 252.445 -233.075 ;
        RECT 252.115 -234.765 252.445 -234.435 ;
        RECT 252.115 -236.125 252.445 -235.795 ;
        RECT 252.115 -237.485 252.445 -237.155 ;
        RECT 252.115 -238.845 252.445 -238.515 ;
        RECT 252.115 -241.09 252.445 -239.96 ;
        RECT 252.12 -241.205 252.44 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.475 237.155 253.805 237.485 ;
        RECT 253.48 237.155 253.8 245.285 ;
        RECT 253.475 244.04 253.805 245.17 ;
        RECT 253.475 242.595 253.805 242.925 ;
        RECT 253.475 241.235 253.805 241.565 ;
        RECT 253.475 239.875 253.805 240.205 ;
        RECT 253.475 238.515 253.805 238.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 244.04 219.805 245.17 ;
        RECT 219.475 242.595 219.805 242.925 ;
        RECT 219.475 241.235 219.805 241.565 ;
        RECT 219.475 239.875 219.805 240.205 ;
        RECT 219.475 238.515 219.805 238.845 ;
        RECT 219.475 237.155 219.805 237.485 ;
        RECT 219.48 237.155 219.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 -0.845 219.805 -0.515 ;
        RECT 219.475 -2.205 219.805 -1.875 ;
        RECT 219.475 -3.565 219.805 -3.235 ;
        RECT 219.48 -3.565 219.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 -123.245 219.805 -122.915 ;
        RECT 219.475 -124.605 219.805 -124.275 ;
        RECT 219.475 -125.965 219.805 -125.635 ;
        RECT 219.475 -127.325 219.805 -126.995 ;
        RECT 219.475 -128.685 219.805 -128.355 ;
        RECT 219.475 -130.045 219.805 -129.715 ;
        RECT 219.475 -131.405 219.805 -131.075 ;
        RECT 219.475 -132.765 219.805 -132.435 ;
        RECT 219.475 -134.125 219.805 -133.795 ;
        RECT 219.475 -135.485 219.805 -135.155 ;
        RECT 219.475 -136.845 219.805 -136.515 ;
        RECT 219.475 -138.205 219.805 -137.875 ;
        RECT 219.475 -139.565 219.805 -139.235 ;
        RECT 219.475 -140.925 219.805 -140.595 ;
        RECT 219.475 -142.285 219.805 -141.955 ;
        RECT 219.475 -143.645 219.805 -143.315 ;
        RECT 219.475 -145.005 219.805 -144.675 ;
        RECT 219.475 -146.365 219.805 -146.035 ;
        RECT 219.475 -147.725 219.805 -147.395 ;
        RECT 219.475 -149.085 219.805 -148.755 ;
        RECT 219.475 -150.445 219.805 -150.115 ;
        RECT 219.475 -151.805 219.805 -151.475 ;
        RECT 219.475 -153.165 219.805 -152.835 ;
        RECT 219.475 -154.525 219.805 -154.195 ;
        RECT 219.475 -155.885 219.805 -155.555 ;
        RECT 219.475 -157.245 219.805 -156.915 ;
        RECT 219.475 -158.605 219.805 -158.275 ;
        RECT 219.475 -159.965 219.805 -159.635 ;
        RECT 219.475 -161.325 219.805 -160.995 ;
        RECT 219.475 -162.685 219.805 -162.355 ;
        RECT 219.475 -164.045 219.805 -163.715 ;
        RECT 219.475 -165.405 219.805 -165.075 ;
        RECT 219.475 -166.765 219.805 -166.435 ;
        RECT 219.475 -168.125 219.805 -167.795 ;
        RECT 219.475 -169.485 219.805 -169.155 ;
        RECT 219.475 -170.845 219.805 -170.515 ;
        RECT 219.475 -172.205 219.805 -171.875 ;
        RECT 219.475 -173.565 219.805 -173.235 ;
        RECT 219.475 -174.925 219.805 -174.595 ;
        RECT 219.475 -176.285 219.805 -175.955 ;
        RECT 219.475 -177.645 219.805 -177.315 ;
        RECT 219.475 -179.005 219.805 -178.675 ;
        RECT 219.475 -180.365 219.805 -180.035 ;
        RECT 219.475 -181.725 219.805 -181.395 ;
        RECT 219.475 -183.085 219.805 -182.755 ;
        RECT 219.475 -184.445 219.805 -184.115 ;
        RECT 219.475 -185.805 219.805 -185.475 ;
        RECT 219.475 -187.165 219.805 -186.835 ;
        RECT 219.475 -188.525 219.805 -188.195 ;
        RECT 219.475 -189.885 219.805 -189.555 ;
        RECT 219.475 -191.245 219.805 -190.915 ;
        RECT 219.475 -192.605 219.805 -192.275 ;
        RECT 219.475 -193.965 219.805 -193.635 ;
        RECT 219.475 -195.325 219.805 -194.995 ;
        RECT 219.475 -196.685 219.805 -196.355 ;
        RECT 219.475 -198.045 219.805 -197.715 ;
        RECT 219.475 -199.405 219.805 -199.075 ;
        RECT 219.475 -200.765 219.805 -200.435 ;
        RECT 219.475 -202.125 219.805 -201.795 ;
        RECT 219.475 -203.485 219.805 -203.155 ;
        RECT 219.475 -204.845 219.805 -204.515 ;
        RECT 219.475 -206.205 219.805 -205.875 ;
        RECT 219.475 -207.565 219.805 -207.235 ;
        RECT 219.475 -208.925 219.805 -208.595 ;
        RECT 219.475 -210.285 219.805 -209.955 ;
        RECT 219.475 -211.645 219.805 -211.315 ;
        RECT 219.475 -213.005 219.805 -212.675 ;
        RECT 219.475 -214.365 219.805 -214.035 ;
        RECT 219.475 -215.725 219.805 -215.395 ;
        RECT 219.475 -217.085 219.805 -216.755 ;
        RECT 219.475 -218.445 219.805 -218.115 ;
        RECT 219.475 -219.805 219.805 -219.475 ;
        RECT 219.475 -221.165 219.805 -220.835 ;
        RECT 219.475 -222.525 219.805 -222.195 ;
        RECT 219.475 -223.885 219.805 -223.555 ;
        RECT 219.475 -225.245 219.805 -224.915 ;
        RECT 219.475 -226.605 219.805 -226.275 ;
        RECT 219.475 -227.965 219.805 -227.635 ;
        RECT 219.475 -229.325 219.805 -228.995 ;
        RECT 219.475 -230.685 219.805 -230.355 ;
        RECT 219.475 -232.045 219.805 -231.715 ;
        RECT 219.475 -233.405 219.805 -233.075 ;
        RECT 219.475 -234.765 219.805 -234.435 ;
        RECT 219.475 -236.125 219.805 -235.795 ;
        RECT 219.475 -237.485 219.805 -237.155 ;
        RECT 219.475 -238.845 219.805 -238.515 ;
        RECT 219.475 -241.09 219.805 -239.96 ;
        RECT 219.48 -241.205 219.8 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 244.04 221.165 245.17 ;
        RECT 220.835 242.595 221.165 242.925 ;
        RECT 220.835 241.235 221.165 241.565 ;
        RECT 220.835 239.875 221.165 240.205 ;
        RECT 220.835 238.515 221.165 238.845 ;
        RECT 220.835 237.155 221.165 237.485 ;
        RECT 220.84 237.155 221.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 -127.325 221.165 -126.995 ;
        RECT 220.835 -128.685 221.165 -128.355 ;
        RECT 220.835 -130.045 221.165 -129.715 ;
        RECT 220.835 -131.405 221.165 -131.075 ;
        RECT 220.835 -132.765 221.165 -132.435 ;
        RECT 220.835 -134.125 221.165 -133.795 ;
        RECT 220.835 -135.485 221.165 -135.155 ;
        RECT 220.835 -136.845 221.165 -136.515 ;
        RECT 220.835 -138.205 221.165 -137.875 ;
        RECT 220.835 -139.565 221.165 -139.235 ;
        RECT 220.835 -140.925 221.165 -140.595 ;
        RECT 220.835 -142.285 221.165 -141.955 ;
        RECT 220.835 -143.645 221.165 -143.315 ;
        RECT 220.835 -145.005 221.165 -144.675 ;
        RECT 220.835 -146.365 221.165 -146.035 ;
        RECT 220.835 -147.725 221.165 -147.395 ;
        RECT 220.835 -149.085 221.165 -148.755 ;
        RECT 220.835 -150.445 221.165 -150.115 ;
        RECT 220.835 -151.805 221.165 -151.475 ;
        RECT 220.835 -153.165 221.165 -152.835 ;
        RECT 220.835 -154.525 221.165 -154.195 ;
        RECT 220.835 -155.885 221.165 -155.555 ;
        RECT 220.835 -157.245 221.165 -156.915 ;
        RECT 220.835 -158.605 221.165 -158.275 ;
        RECT 220.835 -159.965 221.165 -159.635 ;
        RECT 220.835 -161.325 221.165 -160.995 ;
        RECT 220.835 -162.685 221.165 -162.355 ;
        RECT 220.835 -164.045 221.165 -163.715 ;
        RECT 220.835 -165.405 221.165 -165.075 ;
        RECT 220.835 -166.765 221.165 -166.435 ;
        RECT 220.835 -168.125 221.165 -167.795 ;
        RECT 220.835 -169.485 221.165 -169.155 ;
        RECT 220.835 -170.845 221.165 -170.515 ;
        RECT 220.835 -172.205 221.165 -171.875 ;
        RECT 220.835 -173.565 221.165 -173.235 ;
        RECT 220.835 -174.925 221.165 -174.595 ;
        RECT 220.835 -176.285 221.165 -175.955 ;
        RECT 220.835 -177.645 221.165 -177.315 ;
        RECT 220.835 -179.005 221.165 -178.675 ;
        RECT 220.835 -180.365 221.165 -180.035 ;
        RECT 220.835 -181.725 221.165 -181.395 ;
        RECT 220.835 -183.085 221.165 -182.755 ;
        RECT 220.835 -184.445 221.165 -184.115 ;
        RECT 220.835 -185.805 221.165 -185.475 ;
        RECT 220.835 -187.165 221.165 -186.835 ;
        RECT 220.835 -188.525 221.165 -188.195 ;
        RECT 220.835 -189.885 221.165 -189.555 ;
        RECT 220.835 -191.245 221.165 -190.915 ;
        RECT 220.835 -192.605 221.165 -192.275 ;
        RECT 220.835 -193.965 221.165 -193.635 ;
        RECT 220.835 -195.325 221.165 -194.995 ;
        RECT 220.835 -196.685 221.165 -196.355 ;
        RECT 220.835 -198.045 221.165 -197.715 ;
        RECT 220.835 -199.405 221.165 -199.075 ;
        RECT 220.835 -200.765 221.165 -200.435 ;
        RECT 220.835 -202.125 221.165 -201.795 ;
        RECT 220.835 -203.485 221.165 -203.155 ;
        RECT 220.835 -204.845 221.165 -204.515 ;
        RECT 220.835 -206.205 221.165 -205.875 ;
        RECT 220.835 -207.565 221.165 -207.235 ;
        RECT 220.835 -208.925 221.165 -208.595 ;
        RECT 220.835 -210.285 221.165 -209.955 ;
        RECT 220.835 -211.645 221.165 -211.315 ;
        RECT 220.835 -213.005 221.165 -212.675 ;
        RECT 220.835 -214.365 221.165 -214.035 ;
        RECT 220.835 -215.725 221.165 -215.395 ;
        RECT 220.835 -217.085 221.165 -216.755 ;
        RECT 220.835 -218.445 221.165 -218.115 ;
        RECT 220.835 -219.805 221.165 -219.475 ;
        RECT 220.835 -221.165 221.165 -220.835 ;
        RECT 220.835 -222.525 221.165 -222.195 ;
        RECT 220.835 -223.885 221.165 -223.555 ;
        RECT 220.835 -225.245 221.165 -224.915 ;
        RECT 220.835 -226.605 221.165 -226.275 ;
        RECT 220.835 -227.965 221.165 -227.635 ;
        RECT 220.835 -229.325 221.165 -228.995 ;
        RECT 220.835 -230.685 221.165 -230.355 ;
        RECT 220.835 -232.045 221.165 -231.715 ;
        RECT 220.835 -233.405 221.165 -233.075 ;
        RECT 220.835 -234.765 221.165 -234.435 ;
        RECT 220.835 -236.125 221.165 -235.795 ;
        RECT 220.835 -237.485 221.165 -237.155 ;
        RECT 220.835 -238.845 221.165 -238.515 ;
        RECT 220.835 -241.09 221.165 -239.96 ;
        RECT 220.84 -241.205 221.16 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.31 -125.535 221.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 244.04 222.525 245.17 ;
        RECT 222.195 242.595 222.525 242.925 ;
        RECT 222.195 241.235 222.525 241.565 ;
        RECT 222.195 239.875 222.525 240.205 ;
        RECT 222.195 238.515 222.525 238.845 ;
        RECT 222.195 237.155 222.525 237.485 ;
        RECT 222.2 237.155 222.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 -0.845 222.525 -0.515 ;
        RECT 222.195 -2.205 222.525 -1.875 ;
        RECT 222.195 -3.565 222.525 -3.235 ;
        RECT 222.2 -3.565 222.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.555 244.04 223.885 245.17 ;
        RECT 223.555 242.595 223.885 242.925 ;
        RECT 223.555 241.235 223.885 241.565 ;
        RECT 223.555 239.875 223.885 240.205 ;
        RECT 223.555 238.515 223.885 238.845 ;
        RECT 223.555 237.155 223.885 237.485 ;
        RECT 223.56 237.155 223.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.555 -0.845 223.885 -0.515 ;
        RECT 223.555 -2.205 223.885 -1.875 ;
        RECT 223.555 -3.565 223.885 -3.235 ;
        RECT 223.56 -3.565 223.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 244.04 225.245 245.17 ;
        RECT 224.915 242.595 225.245 242.925 ;
        RECT 224.915 241.235 225.245 241.565 ;
        RECT 224.915 239.875 225.245 240.205 ;
        RECT 224.915 238.515 225.245 238.845 ;
        RECT 224.915 237.155 225.245 237.485 ;
        RECT 224.92 237.155 225.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 -0.845 225.245 -0.515 ;
        RECT 224.915 -2.205 225.245 -1.875 ;
        RECT 224.915 -3.565 225.245 -3.235 ;
        RECT 224.92 -3.565 225.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 -123.245 225.245 -122.915 ;
        RECT 224.915 -124.605 225.245 -124.275 ;
        RECT 224.915 -125.965 225.245 -125.635 ;
        RECT 224.915 -127.325 225.245 -126.995 ;
        RECT 224.915 -128.685 225.245 -128.355 ;
        RECT 224.915 -130.045 225.245 -129.715 ;
        RECT 224.915 -131.405 225.245 -131.075 ;
        RECT 224.915 -132.765 225.245 -132.435 ;
        RECT 224.915 -134.125 225.245 -133.795 ;
        RECT 224.915 -135.485 225.245 -135.155 ;
        RECT 224.915 -136.845 225.245 -136.515 ;
        RECT 224.915 -138.205 225.245 -137.875 ;
        RECT 224.915 -139.565 225.245 -139.235 ;
        RECT 224.915 -140.925 225.245 -140.595 ;
        RECT 224.915 -142.285 225.245 -141.955 ;
        RECT 224.915 -143.645 225.245 -143.315 ;
        RECT 224.915 -145.005 225.245 -144.675 ;
        RECT 224.915 -146.365 225.245 -146.035 ;
        RECT 224.915 -147.725 225.245 -147.395 ;
        RECT 224.915 -149.085 225.245 -148.755 ;
        RECT 224.915 -150.445 225.245 -150.115 ;
        RECT 224.915 -151.805 225.245 -151.475 ;
        RECT 224.915 -153.165 225.245 -152.835 ;
        RECT 224.915 -154.525 225.245 -154.195 ;
        RECT 224.915 -155.885 225.245 -155.555 ;
        RECT 224.915 -157.245 225.245 -156.915 ;
        RECT 224.915 -158.605 225.245 -158.275 ;
        RECT 224.915 -159.965 225.245 -159.635 ;
        RECT 224.915 -161.325 225.245 -160.995 ;
        RECT 224.915 -162.685 225.245 -162.355 ;
        RECT 224.915 -164.045 225.245 -163.715 ;
        RECT 224.915 -165.405 225.245 -165.075 ;
        RECT 224.915 -166.765 225.245 -166.435 ;
        RECT 224.915 -168.125 225.245 -167.795 ;
        RECT 224.915 -169.485 225.245 -169.155 ;
        RECT 224.915 -170.845 225.245 -170.515 ;
        RECT 224.915 -172.205 225.245 -171.875 ;
        RECT 224.915 -173.565 225.245 -173.235 ;
        RECT 224.915 -174.925 225.245 -174.595 ;
        RECT 224.915 -176.285 225.245 -175.955 ;
        RECT 224.915 -177.645 225.245 -177.315 ;
        RECT 224.915 -179.005 225.245 -178.675 ;
        RECT 224.915 -180.365 225.245 -180.035 ;
        RECT 224.915 -181.725 225.245 -181.395 ;
        RECT 224.915 -183.085 225.245 -182.755 ;
        RECT 224.915 -184.445 225.245 -184.115 ;
        RECT 224.915 -185.805 225.245 -185.475 ;
        RECT 224.915 -187.165 225.245 -186.835 ;
        RECT 224.915 -188.525 225.245 -188.195 ;
        RECT 224.915 -189.885 225.245 -189.555 ;
        RECT 224.915 -191.245 225.245 -190.915 ;
        RECT 224.915 -192.605 225.245 -192.275 ;
        RECT 224.915 -193.965 225.245 -193.635 ;
        RECT 224.915 -195.325 225.245 -194.995 ;
        RECT 224.915 -196.685 225.245 -196.355 ;
        RECT 224.915 -198.045 225.245 -197.715 ;
        RECT 224.915 -199.405 225.245 -199.075 ;
        RECT 224.915 -200.765 225.245 -200.435 ;
        RECT 224.915 -202.125 225.245 -201.795 ;
        RECT 224.915 -203.485 225.245 -203.155 ;
        RECT 224.915 -204.845 225.245 -204.515 ;
        RECT 224.915 -206.205 225.245 -205.875 ;
        RECT 224.915 -207.565 225.245 -207.235 ;
        RECT 224.915 -208.925 225.245 -208.595 ;
        RECT 224.915 -210.285 225.245 -209.955 ;
        RECT 224.915 -211.645 225.245 -211.315 ;
        RECT 224.915 -213.005 225.245 -212.675 ;
        RECT 224.915 -214.365 225.245 -214.035 ;
        RECT 224.915 -215.725 225.245 -215.395 ;
        RECT 224.915 -217.085 225.245 -216.755 ;
        RECT 224.915 -218.445 225.245 -218.115 ;
        RECT 224.915 -219.805 225.245 -219.475 ;
        RECT 224.915 -221.165 225.245 -220.835 ;
        RECT 224.915 -222.525 225.245 -222.195 ;
        RECT 224.915 -223.885 225.245 -223.555 ;
        RECT 224.915 -225.245 225.245 -224.915 ;
        RECT 224.915 -226.605 225.245 -226.275 ;
        RECT 224.915 -227.965 225.245 -227.635 ;
        RECT 224.915 -229.325 225.245 -228.995 ;
        RECT 224.915 -230.685 225.245 -230.355 ;
        RECT 224.915 -232.045 225.245 -231.715 ;
        RECT 224.915 -233.405 225.245 -233.075 ;
        RECT 224.915 -234.765 225.245 -234.435 ;
        RECT 224.915 -236.125 225.245 -235.795 ;
        RECT 224.915 -237.485 225.245 -237.155 ;
        RECT 224.915 -238.845 225.245 -238.515 ;
        RECT 224.915 -241.09 225.245 -239.96 ;
        RECT 224.92 -241.205 225.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 244.04 226.605 245.17 ;
        RECT 226.275 242.595 226.605 242.925 ;
        RECT 226.275 241.235 226.605 241.565 ;
        RECT 226.275 239.875 226.605 240.205 ;
        RECT 226.275 238.515 226.605 238.845 ;
        RECT 226.275 237.155 226.605 237.485 ;
        RECT 226.28 237.155 226.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 -0.845 226.605 -0.515 ;
        RECT 226.275 -2.205 226.605 -1.875 ;
        RECT 226.275 -3.565 226.605 -3.235 ;
        RECT 226.28 -3.565 226.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 -123.245 226.605 -122.915 ;
        RECT 226.275 -124.605 226.605 -124.275 ;
        RECT 226.275 -125.965 226.605 -125.635 ;
        RECT 226.275 -127.325 226.605 -126.995 ;
        RECT 226.275 -128.685 226.605 -128.355 ;
        RECT 226.275 -130.045 226.605 -129.715 ;
        RECT 226.275 -131.405 226.605 -131.075 ;
        RECT 226.275 -132.765 226.605 -132.435 ;
        RECT 226.275 -134.125 226.605 -133.795 ;
        RECT 226.275 -135.485 226.605 -135.155 ;
        RECT 226.275 -136.845 226.605 -136.515 ;
        RECT 226.275 -138.205 226.605 -137.875 ;
        RECT 226.275 -139.565 226.605 -139.235 ;
        RECT 226.275 -140.925 226.605 -140.595 ;
        RECT 226.275 -142.285 226.605 -141.955 ;
        RECT 226.275 -143.645 226.605 -143.315 ;
        RECT 226.275 -145.005 226.605 -144.675 ;
        RECT 226.275 -146.365 226.605 -146.035 ;
        RECT 226.275 -147.725 226.605 -147.395 ;
        RECT 226.275 -149.085 226.605 -148.755 ;
        RECT 226.275 -150.445 226.605 -150.115 ;
        RECT 226.275 -151.805 226.605 -151.475 ;
        RECT 226.275 -153.165 226.605 -152.835 ;
        RECT 226.275 -154.525 226.605 -154.195 ;
        RECT 226.275 -155.885 226.605 -155.555 ;
        RECT 226.275 -157.245 226.605 -156.915 ;
        RECT 226.275 -158.605 226.605 -158.275 ;
        RECT 226.275 -159.965 226.605 -159.635 ;
        RECT 226.275 -161.325 226.605 -160.995 ;
        RECT 226.275 -162.685 226.605 -162.355 ;
        RECT 226.275 -164.045 226.605 -163.715 ;
        RECT 226.275 -165.405 226.605 -165.075 ;
        RECT 226.275 -166.765 226.605 -166.435 ;
        RECT 226.275 -168.125 226.605 -167.795 ;
        RECT 226.275 -169.485 226.605 -169.155 ;
        RECT 226.275 -170.845 226.605 -170.515 ;
        RECT 226.275 -172.205 226.605 -171.875 ;
        RECT 226.275 -173.565 226.605 -173.235 ;
        RECT 226.275 -174.925 226.605 -174.595 ;
        RECT 226.275 -176.285 226.605 -175.955 ;
        RECT 226.275 -177.645 226.605 -177.315 ;
        RECT 226.275 -179.005 226.605 -178.675 ;
        RECT 226.275 -180.365 226.605 -180.035 ;
        RECT 226.275 -181.725 226.605 -181.395 ;
        RECT 226.275 -183.085 226.605 -182.755 ;
        RECT 226.275 -184.445 226.605 -184.115 ;
        RECT 226.275 -185.805 226.605 -185.475 ;
        RECT 226.275 -187.165 226.605 -186.835 ;
        RECT 226.275 -188.525 226.605 -188.195 ;
        RECT 226.275 -189.885 226.605 -189.555 ;
        RECT 226.275 -191.245 226.605 -190.915 ;
        RECT 226.275 -192.605 226.605 -192.275 ;
        RECT 226.275 -193.965 226.605 -193.635 ;
        RECT 226.275 -195.325 226.605 -194.995 ;
        RECT 226.275 -196.685 226.605 -196.355 ;
        RECT 226.275 -198.045 226.605 -197.715 ;
        RECT 226.275 -199.405 226.605 -199.075 ;
        RECT 226.275 -200.765 226.605 -200.435 ;
        RECT 226.275 -202.125 226.605 -201.795 ;
        RECT 226.275 -203.485 226.605 -203.155 ;
        RECT 226.275 -204.845 226.605 -204.515 ;
        RECT 226.275 -206.205 226.605 -205.875 ;
        RECT 226.275 -207.565 226.605 -207.235 ;
        RECT 226.275 -208.925 226.605 -208.595 ;
        RECT 226.275 -210.285 226.605 -209.955 ;
        RECT 226.275 -211.645 226.605 -211.315 ;
        RECT 226.275 -213.005 226.605 -212.675 ;
        RECT 226.275 -214.365 226.605 -214.035 ;
        RECT 226.275 -215.725 226.605 -215.395 ;
        RECT 226.275 -217.085 226.605 -216.755 ;
        RECT 226.275 -218.445 226.605 -218.115 ;
        RECT 226.275 -219.805 226.605 -219.475 ;
        RECT 226.275 -221.165 226.605 -220.835 ;
        RECT 226.275 -222.525 226.605 -222.195 ;
        RECT 226.275 -223.885 226.605 -223.555 ;
        RECT 226.275 -225.245 226.605 -224.915 ;
        RECT 226.275 -226.605 226.605 -226.275 ;
        RECT 226.275 -227.965 226.605 -227.635 ;
        RECT 226.275 -229.325 226.605 -228.995 ;
        RECT 226.275 -230.685 226.605 -230.355 ;
        RECT 226.275 -232.045 226.605 -231.715 ;
        RECT 226.275 -233.405 226.605 -233.075 ;
        RECT 226.275 -234.765 226.605 -234.435 ;
        RECT 226.275 -236.125 226.605 -235.795 ;
        RECT 226.275 -237.485 226.605 -237.155 ;
        RECT 226.275 -238.845 226.605 -238.515 ;
        RECT 226.275 -241.09 226.605 -239.96 ;
        RECT 226.28 -241.205 226.6 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 244.04 227.965 245.17 ;
        RECT 227.635 242.595 227.965 242.925 ;
        RECT 227.635 241.235 227.965 241.565 ;
        RECT 227.635 239.875 227.965 240.205 ;
        RECT 227.635 238.515 227.965 238.845 ;
        RECT 227.635 237.155 227.965 237.485 ;
        RECT 227.64 237.155 227.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 -0.845 227.965 -0.515 ;
        RECT 227.635 -2.205 227.965 -1.875 ;
        RECT 227.635 -3.565 227.965 -3.235 ;
        RECT 227.64 -3.565 227.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 -123.245 227.965 -122.915 ;
        RECT 227.635 -124.605 227.965 -124.275 ;
        RECT 227.635 -125.965 227.965 -125.635 ;
        RECT 227.635 -127.325 227.965 -126.995 ;
        RECT 227.635 -128.685 227.965 -128.355 ;
        RECT 227.635 -130.045 227.965 -129.715 ;
        RECT 227.635 -131.405 227.965 -131.075 ;
        RECT 227.635 -132.765 227.965 -132.435 ;
        RECT 227.635 -134.125 227.965 -133.795 ;
        RECT 227.635 -135.485 227.965 -135.155 ;
        RECT 227.635 -136.845 227.965 -136.515 ;
        RECT 227.635 -138.205 227.965 -137.875 ;
        RECT 227.635 -139.565 227.965 -139.235 ;
        RECT 227.635 -140.925 227.965 -140.595 ;
        RECT 227.635 -142.285 227.965 -141.955 ;
        RECT 227.635 -143.645 227.965 -143.315 ;
        RECT 227.635 -145.005 227.965 -144.675 ;
        RECT 227.635 -146.365 227.965 -146.035 ;
        RECT 227.635 -147.725 227.965 -147.395 ;
        RECT 227.635 -149.085 227.965 -148.755 ;
        RECT 227.635 -150.445 227.965 -150.115 ;
        RECT 227.635 -151.805 227.965 -151.475 ;
        RECT 227.635 -153.165 227.965 -152.835 ;
        RECT 227.635 -154.525 227.965 -154.195 ;
        RECT 227.635 -155.885 227.965 -155.555 ;
        RECT 227.635 -157.245 227.965 -156.915 ;
        RECT 227.635 -158.605 227.965 -158.275 ;
        RECT 227.635 -159.965 227.965 -159.635 ;
        RECT 227.635 -161.325 227.965 -160.995 ;
        RECT 227.635 -162.685 227.965 -162.355 ;
        RECT 227.635 -164.045 227.965 -163.715 ;
        RECT 227.635 -165.405 227.965 -165.075 ;
        RECT 227.635 -166.765 227.965 -166.435 ;
        RECT 227.635 -168.125 227.965 -167.795 ;
        RECT 227.635 -169.485 227.965 -169.155 ;
        RECT 227.635 -170.845 227.965 -170.515 ;
        RECT 227.635 -172.205 227.965 -171.875 ;
        RECT 227.635 -173.565 227.965 -173.235 ;
        RECT 227.635 -174.925 227.965 -174.595 ;
        RECT 227.635 -176.285 227.965 -175.955 ;
        RECT 227.635 -177.645 227.965 -177.315 ;
        RECT 227.635 -179.005 227.965 -178.675 ;
        RECT 227.635 -180.365 227.965 -180.035 ;
        RECT 227.635 -181.725 227.965 -181.395 ;
        RECT 227.635 -183.085 227.965 -182.755 ;
        RECT 227.635 -184.445 227.965 -184.115 ;
        RECT 227.635 -185.805 227.965 -185.475 ;
        RECT 227.635 -187.165 227.965 -186.835 ;
        RECT 227.635 -188.525 227.965 -188.195 ;
        RECT 227.635 -189.885 227.965 -189.555 ;
        RECT 227.635 -191.245 227.965 -190.915 ;
        RECT 227.635 -192.605 227.965 -192.275 ;
        RECT 227.635 -193.965 227.965 -193.635 ;
        RECT 227.635 -195.325 227.965 -194.995 ;
        RECT 227.635 -196.685 227.965 -196.355 ;
        RECT 227.635 -198.045 227.965 -197.715 ;
        RECT 227.635 -199.405 227.965 -199.075 ;
        RECT 227.635 -200.765 227.965 -200.435 ;
        RECT 227.635 -202.125 227.965 -201.795 ;
        RECT 227.635 -203.485 227.965 -203.155 ;
        RECT 227.635 -204.845 227.965 -204.515 ;
        RECT 227.635 -206.205 227.965 -205.875 ;
        RECT 227.635 -207.565 227.965 -207.235 ;
        RECT 227.635 -208.925 227.965 -208.595 ;
        RECT 227.635 -210.285 227.965 -209.955 ;
        RECT 227.635 -211.645 227.965 -211.315 ;
        RECT 227.635 -213.005 227.965 -212.675 ;
        RECT 227.635 -214.365 227.965 -214.035 ;
        RECT 227.635 -215.725 227.965 -215.395 ;
        RECT 227.635 -217.085 227.965 -216.755 ;
        RECT 227.635 -218.445 227.965 -218.115 ;
        RECT 227.635 -219.805 227.965 -219.475 ;
        RECT 227.635 -221.165 227.965 -220.835 ;
        RECT 227.635 -222.525 227.965 -222.195 ;
        RECT 227.635 -223.885 227.965 -223.555 ;
        RECT 227.635 -225.245 227.965 -224.915 ;
        RECT 227.635 -226.605 227.965 -226.275 ;
        RECT 227.635 -227.965 227.965 -227.635 ;
        RECT 227.635 -229.325 227.965 -228.995 ;
        RECT 227.635 -230.685 227.965 -230.355 ;
        RECT 227.635 -232.045 227.965 -231.715 ;
        RECT 227.635 -233.405 227.965 -233.075 ;
        RECT 227.635 -234.765 227.965 -234.435 ;
        RECT 227.635 -236.125 227.965 -235.795 ;
        RECT 227.635 -237.485 227.965 -237.155 ;
        RECT 227.635 -238.845 227.965 -238.515 ;
        RECT 227.635 -241.09 227.965 -239.96 ;
        RECT 227.64 -241.205 227.96 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 244.04 229.325 245.17 ;
        RECT 228.995 242.595 229.325 242.925 ;
        RECT 228.995 241.235 229.325 241.565 ;
        RECT 228.995 239.875 229.325 240.205 ;
        RECT 228.995 238.515 229.325 238.845 ;
        RECT 228.995 237.155 229.325 237.485 ;
        RECT 229 237.155 229.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 -0.845 229.325 -0.515 ;
        RECT 228.995 -2.205 229.325 -1.875 ;
        RECT 228.995 -3.565 229.325 -3.235 ;
        RECT 229 -3.565 229.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 -123.245 229.325 -122.915 ;
        RECT 228.995 -124.605 229.325 -124.275 ;
        RECT 228.995 -125.965 229.325 -125.635 ;
        RECT 228.995 -127.325 229.325 -126.995 ;
        RECT 228.995 -128.685 229.325 -128.355 ;
        RECT 228.995 -130.045 229.325 -129.715 ;
        RECT 228.995 -131.405 229.325 -131.075 ;
        RECT 228.995 -132.765 229.325 -132.435 ;
        RECT 228.995 -134.125 229.325 -133.795 ;
        RECT 228.995 -135.485 229.325 -135.155 ;
        RECT 228.995 -136.845 229.325 -136.515 ;
        RECT 228.995 -138.205 229.325 -137.875 ;
        RECT 228.995 -139.565 229.325 -139.235 ;
        RECT 228.995 -140.925 229.325 -140.595 ;
        RECT 228.995 -142.285 229.325 -141.955 ;
        RECT 228.995 -143.645 229.325 -143.315 ;
        RECT 228.995 -145.005 229.325 -144.675 ;
        RECT 228.995 -146.365 229.325 -146.035 ;
        RECT 228.995 -147.725 229.325 -147.395 ;
        RECT 228.995 -149.085 229.325 -148.755 ;
        RECT 228.995 -150.445 229.325 -150.115 ;
        RECT 228.995 -151.805 229.325 -151.475 ;
        RECT 228.995 -153.165 229.325 -152.835 ;
        RECT 228.995 -154.525 229.325 -154.195 ;
        RECT 228.995 -155.885 229.325 -155.555 ;
        RECT 228.995 -157.245 229.325 -156.915 ;
        RECT 228.995 -158.605 229.325 -158.275 ;
        RECT 228.995 -159.965 229.325 -159.635 ;
        RECT 228.995 -161.325 229.325 -160.995 ;
        RECT 228.995 -162.685 229.325 -162.355 ;
        RECT 228.995 -164.045 229.325 -163.715 ;
        RECT 228.995 -165.405 229.325 -165.075 ;
        RECT 228.995 -166.765 229.325 -166.435 ;
        RECT 228.995 -168.125 229.325 -167.795 ;
        RECT 228.995 -169.485 229.325 -169.155 ;
        RECT 228.995 -170.845 229.325 -170.515 ;
        RECT 228.995 -172.205 229.325 -171.875 ;
        RECT 228.995 -173.565 229.325 -173.235 ;
        RECT 228.995 -174.925 229.325 -174.595 ;
        RECT 228.995 -176.285 229.325 -175.955 ;
        RECT 228.995 -177.645 229.325 -177.315 ;
        RECT 228.995 -179.005 229.325 -178.675 ;
        RECT 228.995 -180.365 229.325 -180.035 ;
        RECT 228.995 -181.725 229.325 -181.395 ;
        RECT 228.995 -183.085 229.325 -182.755 ;
        RECT 228.995 -184.445 229.325 -184.115 ;
        RECT 228.995 -185.805 229.325 -185.475 ;
        RECT 228.995 -187.165 229.325 -186.835 ;
        RECT 228.995 -188.525 229.325 -188.195 ;
        RECT 228.995 -189.885 229.325 -189.555 ;
        RECT 228.995 -191.245 229.325 -190.915 ;
        RECT 228.995 -192.605 229.325 -192.275 ;
        RECT 228.995 -193.965 229.325 -193.635 ;
        RECT 228.995 -195.325 229.325 -194.995 ;
        RECT 228.995 -196.685 229.325 -196.355 ;
        RECT 228.995 -198.045 229.325 -197.715 ;
        RECT 228.995 -199.405 229.325 -199.075 ;
        RECT 228.995 -200.765 229.325 -200.435 ;
        RECT 228.995 -202.125 229.325 -201.795 ;
        RECT 228.995 -203.485 229.325 -203.155 ;
        RECT 228.995 -204.845 229.325 -204.515 ;
        RECT 228.995 -206.205 229.325 -205.875 ;
        RECT 228.995 -207.565 229.325 -207.235 ;
        RECT 228.995 -208.925 229.325 -208.595 ;
        RECT 228.995 -210.285 229.325 -209.955 ;
        RECT 228.995 -211.645 229.325 -211.315 ;
        RECT 228.995 -213.005 229.325 -212.675 ;
        RECT 228.995 -214.365 229.325 -214.035 ;
        RECT 228.995 -215.725 229.325 -215.395 ;
        RECT 228.995 -217.085 229.325 -216.755 ;
        RECT 228.995 -218.445 229.325 -218.115 ;
        RECT 228.995 -219.805 229.325 -219.475 ;
        RECT 228.995 -221.165 229.325 -220.835 ;
        RECT 228.995 -222.525 229.325 -222.195 ;
        RECT 228.995 -223.885 229.325 -223.555 ;
        RECT 228.995 -225.245 229.325 -224.915 ;
        RECT 228.995 -226.605 229.325 -226.275 ;
        RECT 228.995 -227.965 229.325 -227.635 ;
        RECT 228.995 -229.325 229.325 -228.995 ;
        RECT 228.995 -230.685 229.325 -230.355 ;
        RECT 228.995 -232.045 229.325 -231.715 ;
        RECT 228.995 -233.405 229.325 -233.075 ;
        RECT 228.995 -234.765 229.325 -234.435 ;
        RECT 228.995 -236.125 229.325 -235.795 ;
        RECT 228.995 -237.485 229.325 -237.155 ;
        RECT 228.995 -238.845 229.325 -238.515 ;
        RECT 228.995 -241.09 229.325 -239.96 ;
        RECT 229 -241.205 229.32 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 244.04 230.685 245.17 ;
        RECT 230.355 242.595 230.685 242.925 ;
        RECT 230.355 241.235 230.685 241.565 ;
        RECT 230.355 239.875 230.685 240.205 ;
        RECT 230.355 238.515 230.685 238.845 ;
        RECT 230.355 237.155 230.685 237.485 ;
        RECT 230.36 237.155 230.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 -0.845 230.685 -0.515 ;
        RECT 230.355 -2.205 230.685 -1.875 ;
        RECT 230.355 -3.565 230.685 -3.235 ;
        RECT 230.36 -3.565 230.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 -123.245 230.685 -122.915 ;
        RECT 230.355 -124.605 230.685 -124.275 ;
        RECT 230.355 -125.965 230.685 -125.635 ;
        RECT 230.355 -127.325 230.685 -126.995 ;
        RECT 230.355 -128.685 230.685 -128.355 ;
        RECT 230.355 -130.045 230.685 -129.715 ;
        RECT 230.355 -131.405 230.685 -131.075 ;
        RECT 230.355 -132.765 230.685 -132.435 ;
        RECT 230.355 -134.125 230.685 -133.795 ;
        RECT 230.355 -135.485 230.685 -135.155 ;
        RECT 230.355 -136.845 230.685 -136.515 ;
        RECT 230.355 -138.205 230.685 -137.875 ;
        RECT 230.355 -139.565 230.685 -139.235 ;
        RECT 230.355 -140.925 230.685 -140.595 ;
        RECT 230.355 -142.285 230.685 -141.955 ;
        RECT 230.355 -143.645 230.685 -143.315 ;
        RECT 230.355 -145.005 230.685 -144.675 ;
        RECT 230.355 -146.365 230.685 -146.035 ;
        RECT 230.355 -147.725 230.685 -147.395 ;
        RECT 230.355 -149.085 230.685 -148.755 ;
        RECT 230.355 -150.445 230.685 -150.115 ;
        RECT 230.355 -151.805 230.685 -151.475 ;
        RECT 230.355 -153.165 230.685 -152.835 ;
        RECT 230.355 -154.525 230.685 -154.195 ;
        RECT 230.355 -155.885 230.685 -155.555 ;
        RECT 230.355 -157.245 230.685 -156.915 ;
        RECT 230.355 -158.605 230.685 -158.275 ;
        RECT 230.355 -159.965 230.685 -159.635 ;
        RECT 230.355 -161.325 230.685 -160.995 ;
        RECT 230.355 -162.685 230.685 -162.355 ;
        RECT 230.355 -164.045 230.685 -163.715 ;
        RECT 230.355 -165.405 230.685 -165.075 ;
        RECT 230.355 -166.765 230.685 -166.435 ;
        RECT 230.355 -168.125 230.685 -167.795 ;
        RECT 230.355 -169.485 230.685 -169.155 ;
        RECT 230.355 -170.845 230.685 -170.515 ;
        RECT 230.355 -172.205 230.685 -171.875 ;
        RECT 230.355 -173.565 230.685 -173.235 ;
        RECT 230.355 -174.925 230.685 -174.595 ;
        RECT 230.355 -176.285 230.685 -175.955 ;
        RECT 230.355 -177.645 230.685 -177.315 ;
        RECT 230.355 -179.005 230.685 -178.675 ;
        RECT 230.355 -180.365 230.685 -180.035 ;
        RECT 230.355 -181.725 230.685 -181.395 ;
        RECT 230.355 -183.085 230.685 -182.755 ;
        RECT 230.355 -184.445 230.685 -184.115 ;
        RECT 230.355 -185.805 230.685 -185.475 ;
        RECT 230.355 -187.165 230.685 -186.835 ;
        RECT 230.355 -188.525 230.685 -188.195 ;
        RECT 230.355 -189.885 230.685 -189.555 ;
        RECT 230.355 -191.245 230.685 -190.915 ;
        RECT 230.355 -192.605 230.685 -192.275 ;
        RECT 230.355 -193.965 230.685 -193.635 ;
        RECT 230.355 -195.325 230.685 -194.995 ;
        RECT 230.355 -196.685 230.685 -196.355 ;
        RECT 230.355 -198.045 230.685 -197.715 ;
        RECT 230.355 -199.405 230.685 -199.075 ;
        RECT 230.355 -200.765 230.685 -200.435 ;
        RECT 230.355 -202.125 230.685 -201.795 ;
        RECT 230.355 -203.485 230.685 -203.155 ;
        RECT 230.355 -204.845 230.685 -204.515 ;
        RECT 230.355 -206.205 230.685 -205.875 ;
        RECT 230.355 -207.565 230.685 -207.235 ;
        RECT 230.355 -208.925 230.685 -208.595 ;
        RECT 230.355 -210.285 230.685 -209.955 ;
        RECT 230.355 -211.645 230.685 -211.315 ;
        RECT 230.355 -213.005 230.685 -212.675 ;
        RECT 230.355 -214.365 230.685 -214.035 ;
        RECT 230.355 -215.725 230.685 -215.395 ;
        RECT 230.355 -217.085 230.685 -216.755 ;
        RECT 230.355 -218.445 230.685 -218.115 ;
        RECT 230.355 -219.805 230.685 -219.475 ;
        RECT 230.355 -221.165 230.685 -220.835 ;
        RECT 230.355 -222.525 230.685 -222.195 ;
        RECT 230.355 -223.885 230.685 -223.555 ;
        RECT 230.355 -225.245 230.685 -224.915 ;
        RECT 230.355 -226.605 230.685 -226.275 ;
        RECT 230.355 -227.965 230.685 -227.635 ;
        RECT 230.355 -229.325 230.685 -228.995 ;
        RECT 230.355 -230.685 230.685 -230.355 ;
        RECT 230.355 -232.045 230.685 -231.715 ;
        RECT 230.355 -233.405 230.685 -233.075 ;
        RECT 230.355 -234.765 230.685 -234.435 ;
        RECT 230.355 -236.125 230.685 -235.795 ;
        RECT 230.355 -237.485 230.685 -237.155 ;
        RECT 230.355 -238.845 230.685 -238.515 ;
        RECT 230.355 -241.09 230.685 -239.96 ;
        RECT 230.36 -241.205 230.68 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 244.04 232.045 245.17 ;
        RECT 231.715 242.595 232.045 242.925 ;
        RECT 231.715 241.235 232.045 241.565 ;
        RECT 231.715 239.875 232.045 240.205 ;
        RECT 231.715 238.515 232.045 238.845 ;
        RECT 231.715 237.155 232.045 237.485 ;
        RECT 231.72 237.155 232.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 -127.325 232.045 -126.995 ;
        RECT 231.715 -128.685 232.045 -128.355 ;
        RECT 231.715 -130.045 232.045 -129.715 ;
        RECT 231.715 -131.405 232.045 -131.075 ;
        RECT 231.715 -132.765 232.045 -132.435 ;
        RECT 231.715 -134.125 232.045 -133.795 ;
        RECT 231.715 -135.485 232.045 -135.155 ;
        RECT 231.715 -136.845 232.045 -136.515 ;
        RECT 231.715 -138.205 232.045 -137.875 ;
        RECT 231.715 -139.565 232.045 -139.235 ;
        RECT 231.715 -140.925 232.045 -140.595 ;
        RECT 231.715 -142.285 232.045 -141.955 ;
        RECT 231.715 -143.645 232.045 -143.315 ;
        RECT 231.715 -145.005 232.045 -144.675 ;
        RECT 231.715 -146.365 232.045 -146.035 ;
        RECT 231.715 -147.725 232.045 -147.395 ;
        RECT 231.715 -149.085 232.045 -148.755 ;
        RECT 231.715 -150.445 232.045 -150.115 ;
        RECT 231.715 -151.805 232.045 -151.475 ;
        RECT 231.715 -153.165 232.045 -152.835 ;
        RECT 231.715 -154.525 232.045 -154.195 ;
        RECT 231.715 -155.885 232.045 -155.555 ;
        RECT 231.715 -157.245 232.045 -156.915 ;
        RECT 231.715 -158.605 232.045 -158.275 ;
        RECT 231.715 -159.965 232.045 -159.635 ;
        RECT 231.715 -161.325 232.045 -160.995 ;
        RECT 231.715 -162.685 232.045 -162.355 ;
        RECT 231.715 -164.045 232.045 -163.715 ;
        RECT 231.715 -165.405 232.045 -165.075 ;
        RECT 231.715 -166.765 232.045 -166.435 ;
        RECT 231.715 -168.125 232.045 -167.795 ;
        RECT 231.715 -169.485 232.045 -169.155 ;
        RECT 231.715 -170.845 232.045 -170.515 ;
        RECT 231.715 -172.205 232.045 -171.875 ;
        RECT 231.715 -173.565 232.045 -173.235 ;
        RECT 231.715 -174.925 232.045 -174.595 ;
        RECT 231.715 -176.285 232.045 -175.955 ;
        RECT 231.715 -177.645 232.045 -177.315 ;
        RECT 231.715 -179.005 232.045 -178.675 ;
        RECT 231.715 -180.365 232.045 -180.035 ;
        RECT 231.715 -181.725 232.045 -181.395 ;
        RECT 231.715 -183.085 232.045 -182.755 ;
        RECT 231.715 -184.445 232.045 -184.115 ;
        RECT 231.715 -185.805 232.045 -185.475 ;
        RECT 231.715 -187.165 232.045 -186.835 ;
        RECT 231.715 -188.525 232.045 -188.195 ;
        RECT 231.715 -189.885 232.045 -189.555 ;
        RECT 231.715 -191.245 232.045 -190.915 ;
        RECT 231.715 -192.605 232.045 -192.275 ;
        RECT 231.715 -193.965 232.045 -193.635 ;
        RECT 231.715 -195.325 232.045 -194.995 ;
        RECT 231.715 -196.685 232.045 -196.355 ;
        RECT 231.715 -198.045 232.045 -197.715 ;
        RECT 231.715 -199.405 232.045 -199.075 ;
        RECT 231.715 -200.765 232.045 -200.435 ;
        RECT 231.715 -202.125 232.045 -201.795 ;
        RECT 231.715 -203.485 232.045 -203.155 ;
        RECT 231.715 -204.845 232.045 -204.515 ;
        RECT 231.715 -206.205 232.045 -205.875 ;
        RECT 231.715 -207.565 232.045 -207.235 ;
        RECT 231.715 -208.925 232.045 -208.595 ;
        RECT 231.715 -210.285 232.045 -209.955 ;
        RECT 231.715 -211.645 232.045 -211.315 ;
        RECT 231.715 -213.005 232.045 -212.675 ;
        RECT 231.715 -214.365 232.045 -214.035 ;
        RECT 231.715 -215.725 232.045 -215.395 ;
        RECT 231.715 -217.085 232.045 -216.755 ;
        RECT 231.715 -218.445 232.045 -218.115 ;
        RECT 231.715 -219.805 232.045 -219.475 ;
        RECT 231.715 -221.165 232.045 -220.835 ;
        RECT 231.715 -222.525 232.045 -222.195 ;
        RECT 231.715 -223.885 232.045 -223.555 ;
        RECT 231.715 -225.245 232.045 -224.915 ;
        RECT 231.715 -226.605 232.045 -226.275 ;
        RECT 231.715 -227.965 232.045 -227.635 ;
        RECT 231.715 -229.325 232.045 -228.995 ;
        RECT 231.715 -230.685 232.045 -230.355 ;
        RECT 231.715 -232.045 232.045 -231.715 ;
        RECT 231.715 -233.405 232.045 -233.075 ;
        RECT 231.715 -234.765 232.045 -234.435 ;
        RECT 231.715 -236.125 232.045 -235.795 ;
        RECT 231.715 -237.485 232.045 -237.155 ;
        RECT 231.715 -238.845 232.045 -238.515 ;
        RECT 231.715 -241.09 232.045 -239.96 ;
        RECT 231.72 -241.205 232.04 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.21 -125.535 232.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 244.04 233.405 245.17 ;
        RECT 233.075 242.595 233.405 242.925 ;
        RECT 233.075 241.235 233.405 241.565 ;
        RECT 233.075 239.875 233.405 240.205 ;
        RECT 233.075 238.515 233.405 238.845 ;
        RECT 233.075 237.155 233.405 237.485 ;
        RECT 233.08 237.155 233.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 -0.845 233.405 -0.515 ;
        RECT 233.075 -2.205 233.405 -1.875 ;
        RECT 233.075 -3.565 233.405 -3.235 ;
        RECT 233.08 -3.565 233.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 244.04 234.765 245.17 ;
        RECT 234.435 242.595 234.765 242.925 ;
        RECT 234.435 241.235 234.765 241.565 ;
        RECT 234.435 239.875 234.765 240.205 ;
        RECT 234.435 238.515 234.765 238.845 ;
        RECT 234.435 237.155 234.765 237.485 ;
        RECT 234.44 237.155 234.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 -0.845 234.765 -0.515 ;
        RECT 234.435 -2.205 234.765 -1.875 ;
        RECT 234.435 -3.565 234.765 -3.235 ;
        RECT 234.44 -3.565 234.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 244.04 236.125 245.17 ;
        RECT 235.795 242.595 236.125 242.925 ;
        RECT 235.795 241.235 236.125 241.565 ;
        RECT 235.795 239.875 236.125 240.205 ;
        RECT 235.795 238.515 236.125 238.845 ;
        RECT 235.795 237.155 236.125 237.485 ;
        RECT 235.8 237.155 236.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 -0.845 236.125 -0.515 ;
        RECT 235.795 -2.205 236.125 -1.875 ;
        RECT 235.795 -3.565 236.125 -3.235 ;
        RECT 235.8 -3.565 236.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 -123.245 236.125 -122.915 ;
        RECT 235.795 -124.605 236.125 -124.275 ;
        RECT 235.795 -125.965 236.125 -125.635 ;
        RECT 235.795 -127.325 236.125 -126.995 ;
        RECT 235.795 -128.685 236.125 -128.355 ;
        RECT 235.795 -130.045 236.125 -129.715 ;
        RECT 235.795 -131.405 236.125 -131.075 ;
        RECT 235.795 -132.765 236.125 -132.435 ;
        RECT 235.795 -134.125 236.125 -133.795 ;
        RECT 235.795 -135.485 236.125 -135.155 ;
        RECT 235.795 -136.845 236.125 -136.515 ;
        RECT 235.795 -138.205 236.125 -137.875 ;
        RECT 235.795 -139.565 236.125 -139.235 ;
        RECT 235.795 -140.925 236.125 -140.595 ;
        RECT 235.795 -142.285 236.125 -141.955 ;
        RECT 235.795 -143.645 236.125 -143.315 ;
        RECT 235.795 -145.005 236.125 -144.675 ;
        RECT 235.795 -146.365 236.125 -146.035 ;
        RECT 235.795 -147.725 236.125 -147.395 ;
        RECT 235.795 -149.085 236.125 -148.755 ;
        RECT 235.795 -150.445 236.125 -150.115 ;
        RECT 235.795 -151.805 236.125 -151.475 ;
        RECT 235.795 -153.165 236.125 -152.835 ;
        RECT 235.795 -154.525 236.125 -154.195 ;
        RECT 235.795 -155.885 236.125 -155.555 ;
        RECT 235.795 -157.245 236.125 -156.915 ;
        RECT 235.795 -158.605 236.125 -158.275 ;
        RECT 235.795 -159.965 236.125 -159.635 ;
        RECT 235.795 -161.325 236.125 -160.995 ;
        RECT 235.795 -162.685 236.125 -162.355 ;
        RECT 235.795 -164.045 236.125 -163.715 ;
        RECT 235.795 -165.405 236.125 -165.075 ;
        RECT 235.795 -166.765 236.125 -166.435 ;
        RECT 235.795 -168.125 236.125 -167.795 ;
        RECT 235.795 -169.485 236.125 -169.155 ;
        RECT 235.795 -170.845 236.125 -170.515 ;
        RECT 235.795 -172.205 236.125 -171.875 ;
        RECT 235.795 -173.565 236.125 -173.235 ;
        RECT 235.795 -174.925 236.125 -174.595 ;
        RECT 235.795 -176.285 236.125 -175.955 ;
        RECT 235.795 -177.645 236.125 -177.315 ;
        RECT 235.795 -179.005 236.125 -178.675 ;
        RECT 235.795 -180.365 236.125 -180.035 ;
        RECT 235.795 -181.725 236.125 -181.395 ;
        RECT 235.795 -183.085 236.125 -182.755 ;
        RECT 235.795 -184.445 236.125 -184.115 ;
        RECT 235.795 -185.805 236.125 -185.475 ;
        RECT 235.795 -187.165 236.125 -186.835 ;
        RECT 235.795 -188.525 236.125 -188.195 ;
        RECT 235.795 -189.885 236.125 -189.555 ;
        RECT 235.795 -191.245 236.125 -190.915 ;
        RECT 235.795 -192.605 236.125 -192.275 ;
        RECT 235.795 -193.965 236.125 -193.635 ;
        RECT 235.795 -195.325 236.125 -194.995 ;
        RECT 235.795 -196.685 236.125 -196.355 ;
        RECT 235.795 -198.045 236.125 -197.715 ;
        RECT 235.795 -199.405 236.125 -199.075 ;
        RECT 235.795 -200.765 236.125 -200.435 ;
        RECT 235.795 -202.125 236.125 -201.795 ;
        RECT 235.795 -203.485 236.125 -203.155 ;
        RECT 235.795 -204.845 236.125 -204.515 ;
        RECT 235.795 -206.205 236.125 -205.875 ;
        RECT 235.795 -207.565 236.125 -207.235 ;
        RECT 235.795 -208.925 236.125 -208.595 ;
        RECT 235.795 -210.285 236.125 -209.955 ;
        RECT 235.795 -211.645 236.125 -211.315 ;
        RECT 235.795 -213.005 236.125 -212.675 ;
        RECT 235.795 -214.365 236.125 -214.035 ;
        RECT 235.795 -215.725 236.125 -215.395 ;
        RECT 235.795 -217.085 236.125 -216.755 ;
        RECT 235.795 -218.445 236.125 -218.115 ;
        RECT 235.795 -219.805 236.125 -219.475 ;
        RECT 235.795 -221.165 236.125 -220.835 ;
        RECT 235.795 -222.525 236.125 -222.195 ;
        RECT 235.795 -223.885 236.125 -223.555 ;
        RECT 235.795 -225.245 236.125 -224.915 ;
        RECT 235.795 -226.605 236.125 -226.275 ;
        RECT 235.795 -227.965 236.125 -227.635 ;
        RECT 235.795 -229.325 236.125 -228.995 ;
        RECT 235.795 -230.685 236.125 -230.355 ;
        RECT 235.795 -232.045 236.125 -231.715 ;
        RECT 235.795 -233.405 236.125 -233.075 ;
        RECT 235.795 -234.765 236.125 -234.435 ;
        RECT 235.795 -236.125 236.125 -235.795 ;
        RECT 235.795 -237.485 236.125 -237.155 ;
        RECT 235.795 -238.845 236.125 -238.515 ;
        RECT 235.795 -241.09 236.125 -239.96 ;
        RECT 235.8 -241.205 236.12 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 244.04 237.485 245.17 ;
        RECT 237.155 242.595 237.485 242.925 ;
        RECT 237.155 241.235 237.485 241.565 ;
        RECT 237.155 239.875 237.485 240.205 ;
        RECT 237.155 238.515 237.485 238.845 ;
        RECT 237.155 237.155 237.485 237.485 ;
        RECT 237.16 237.155 237.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.16 -3.565 237.48 -0.515 ;
        RECT 237.155 -0.845 237.485 -0.515 ;
        RECT 237.155 -2.205 237.485 -1.875 ;
        RECT 237.155 -3.565 237.485 -3.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.51 -125.535 199.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 244.04 200.765 245.17 ;
        RECT 200.435 242.595 200.765 242.925 ;
        RECT 200.435 241.235 200.765 241.565 ;
        RECT 200.435 239.875 200.765 240.205 ;
        RECT 200.435 238.515 200.765 238.845 ;
        RECT 200.435 237.155 200.765 237.485 ;
        RECT 200.44 237.155 200.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 -0.845 200.765 -0.515 ;
        RECT 200.435 -2.205 200.765 -1.875 ;
        RECT 200.435 -3.565 200.765 -3.235 ;
        RECT 200.44 -3.565 200.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 244.04 202.125 245.17 ;
        RECT 201.795 242.595 202.125 242.925 ;
        RECT 201.795 241.235 202.125 241.565 ;
        RECT 201.795 239.875 202.125 240.205 ;
        RECT 201.795 238.515 202.125 238.845 ;
        RECT 201.795 237.155 202.125 237.485 ;
        RECT 201.8 237.155 202.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 -0.845 202.125 -0.515 ;
        RECT 201.795 -2.205 202.125 -1.875 ;
        RECT 201.795 -3.565 202.125 -3.235 ;
        RECT 201.8 -3.565 202.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 244.04 203.485 245.17 ;
        RECT 203.155 242.595 203.485 242.925 ;
        RECT 203.155 241.235 203.485 241.565 ;
        RECT 203.155 239.875 203.485 240.205 ;
        RECT 203.155 238.515 203.485 238.845 ;
        RECT 203.155 237.155 203.485 237.485 ;
        RECT 203.16 237.155 203.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 -0.845 203.485 -0.515 ;
        RECT 203.155 -2.205 203.485 -1.875 ;
        RECT 203.155 -3.565 203.485 -3.235 ;
        RECT 203.16 -3.565 203.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 -123.245 203.485 -122.915 ;
        RECT 203.155 -124.605 203.485 -124.275 ;
        RECT 203.155 -125.965 203.485 -125.635 ;
        RECT 203.155 -127.325 203.485 -126.995 ;
        RECT 203.155 -128.685 203.485 -128.355 ;
        RECT 203.155 -130.045 203.485 -129.715 ;
        RECT 203.155 -131.405 203.485 -131.075 ;
        RECT 203.155 -132.765 203.485 -132.435 ;
        RECT 203.155 -134.125 203.485 -133.795 ;
        RECT 203.155 -135.485 203.485 -135.155 ;
        RECT 203.155 -136.845 203.485 -136.515 ;
        RECT 203.155 -138.205 203.485 -137.875 ;
        RECT 203.155 -139.565 203.485 -139.235 ;
        RECT 203.155 -140.925 203.485 -140.595 ;
        RECT 203.155 -142.285 203.485 -141.955 ;
        RECT 203.155 -143.645 203.485 -143.315 ;
        RECT 203.155 -145.005 203.485 -144.675 ;
        RECT 203.155 -146.365 203.485 -146.035 ;
        RECT 203.155 -147.725 203.485 -147.395 ;
        RECT 203.155 -149.085 203.485 -148.755 ;
        RECT 203.155 -150.445 203.485 -150.115 ;
        RECT 203.155 -151.805 203.485 -151.475 ;
        RECT 203.155 -153.165 203.485 -152.835 ;
        RECT 203.155 -154.525 203.485 -154.195 ;
        RECT 203.155 -155.885 203.485 -155.555 ;
        RECT 203.155 -157.245 203.485 -156.915 ;
        RECT 203.155 -158.605 203.485 -158.275 ;
        RECT 203.155 -159.965 203.485 -159.635 ;
        RECT 203.155 -161.325 203.485 -160.995 ;
        RECT 203.155 -162.685 203.485 -162.355 ;
        RECT 203.155 -164.045 203.485 -163.715 ;
        RECT 203.155 -165.405 203.485 -165.075 ;
        RECT 203.155 -166.765 203.485 -166.435 ;
        RECT 203.155 -168.125 203.485 -167.795 ;
        RECT 203.155 -169.485 203.485 -169.155 ;
        RECT 203.155 -170.845 203.485 -170.515 ;
        RECT 203.155 -172.205 203.485 -171.875 ;
        RECT 203.155 -173.565 203.485 -173.235 ;
        RECT 203.155 -174.925 203.485 -174.595 ;
        RECT 203.155 -176.285 203.485 -175.955 ;
        RECT 203.155 -177.645 203.485 -177.315 ;
        RECT 203.155 -179.005 203.485 -178.675 ;
        RECT 203.155 -180.365 203.485 -180.035 ;
        RECT 203.155 -181.725 203.485 -181.395 ;
        RECT 203.155 -183.085 203.485 -182.755 ;
        RECT 203.155 -184.445 203.485 -184.115 ;
        RECT 203.155 -185.805 203.485 -185.475 ;
        RECT 203.155 -187.165 203.485 -186.835 ;
        RECT 203.155 -188.525 203.485 -188.195 ;
        RECT 203.155 -189.885 203.485 -189.555 ;
        RECT 203.155 -191.245 203.485 -190.915 ;
        RECT 203.155 -192.605 203.485 -192.275 ;
        RECT 203.155 -193.965 203.485 -193.635 ;
        RECT 203.155 -195.325 203.485 -194.995 ;
        RECT 203.155 -196.685 203.485 -196.355 ;
        RECT 203.155 -198.045 203.485 -197.715 ;
        RECT 203.155 -199.405 203.485 -199.075 ;
        RECT 203.155 -200.765 203.485 -200.435 ;
        RECT 203.155 -202.125 203.485 -201.795 ;
        RECT 203.155 -203.485 203.485 -203.155 ;
        RECT 203.155 -204.845 203.485 -204.515 ;
        RECT 203.155 -206.205 203.485 -205.875 ;
        RECT 203.155 -207.565 203.485 -207.235 ;
        RECT 203.155 -208.925 203.485 -208.595 ;
        RECT 203.155 -210.285 203.485 -209.955 ;
        RECT 203.155 -211.645 203.485 -211.315 ;
        RECT 203.155 -213.005 203.485 -212.675 ;
        RECT 203.155 -214.365 203.485 -214.035 ;
        RECT 203.155 -215.725 203.485 -215.395 ;
        RECT 203.155 -217.085 203.485 -216.755 ;
        RECT 203.155 -218.445 203.485 -218.115 ;
        RECT 203.155 -219.805 203.485 -219.475 ;
        RECT 203.155 -221.165 203.485 -220.835 ;
        RECT 203.155 -222.525 203.485 -222.195 ;
        RECT 203.155 -223.885 203.485 -223.555 ;
        RECT 203.155 -225.245 203.485 -224.915 ;
        RECT 203.155 -226.605 203.485 -226.275 ;
        RECT 203.155 -227.965 203.485 -227.635 ;
        RECT 203.155 -229.325 203.485 -228.995 ;
        RECT 203.155 -230.685 203.485 -230.355 ;
        RECT 203.155 -232.045 203.485 -231.715 ;
        RECT 203.155 -233.405 203.485 -233.075 ;
        RECT 203.155 -234.765 203.485 -234.435 ;
        RECT 203.155 -236.125 203.485 -235.795 ;
        RECT 203.155 -237.485 203.485 -237.155 ;
        RECT 203.155 -238.845 203.485 -238.515 ;
        RECT 203.155 -241.09 203.485 -239.96 ;
        RECT 203.16 -241.205 203.48 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 244.04 204.845 245.17 ;
        RECT 204.515 242.595 204.845 242.925 ;
        RECT 204.515 241.235 204.845 241.565 ;
        RECT 204.515 239.875 204.845 240.205 ;
        RECT 204.515 238.515 204.845 238.845 ;
        RECT 204.515 237.155 204.845 237.485 ;
        RECT 204.52 237.155 204.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 -0.845 204.845 -0.515 ;
        RECT 204.515 -2.205 204.845 -1.875 ;
        RECT 204.515 -3.565 204.845 -3.235 ;
        RECT 204.52 -3.565 204.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 -123.245 204.845 -122.915 ;
        RECT 204.515 -124.605 204.845 -124.275 ;
        RECT 204.515 -125.965 204.845 -125.635 ;
        RECT 204.515 -127.325 204.845 -126.995 ;
        RECT 204.515 -128.685 204.845 -128.355 ;
        RECT 204.515 -130.045 204.845 -129.715 ;
        RECT 204.515 -131.405 204.845 -131.075 ;
        RECT 204.515 -132.765 204.845 -132.435 ;
        RECT 204.515 -134.125 204.845 -133.795 ;
        RECT 204.515 -135.485 204.845 -135.155 ;
        RECT 204.515 -136.845 204.845 -136.515 ;
        RECT 204.515 -138.205 204.845 -137.875 ;
        RECT 204.515 -139.565 204.845 -139.235 ;
        RECT 204.515 -140.925 204.845 -140.595 ;
        RECT 204.515 -142.285 204.845 -141.955 ;
        RECT 204.515 -143.645 204.845 -143.315 ;
        RECT 204.515 -145.005 204.845 -144.675 ;
        RECT 204.515 -146.365 204.845 -146.035 ;
        RECT 204.515 -147.725 204.845 -147.395 ;
        RECT 204.515 -149.085 204.845 -148.755 ;
        RECT 204.515 -150.445 204.845 -150.115 ;
        RECT 204.515 -151.805 204.845 -151.475 ;
        RECT 204.515 -153.165 204.845 -152.835 ;
        RECT 204.515 -154.525 204.845 -154.195 ;
        RECT 204.515 -155.885 204.845 -155.555 ;
        RECT 204.515 -157.245 204.845 -156.915 ;
        RECT 204.515 -158.605 204.845 -158.275 ;
        RECT 204.515 -159.965 204.845 -159.635 ;
        RECT 204.515 -161.325 204.845 -160.995 ;
        RECT 204.515 -162.685 204.845 -162.355 ;
        RECT 204.515 -164.045 204.845 -163.715 ;
        RECT 204.515 -165.405 204.845 -165.075 ;
        RECT 204.515 -166.765 204.845 -166.435 ;
        RECT 204.515 -168.125 204.845 -167.795 ;
        RECT 204.515 -169.485 204.845 -169.155 ;
        RECT 204.515 -170.845 204.845 -170.515 ;
        RECT 204.515 -172.205 204.845 -171.875 ;
        RECT 204.515 -173.565 204.845 -173.235 ;
        RECT 204.515 -174.925 204.845 -174.595 ;
        RECT 204.515 -176.285 204.845 -175.955 ;
        RECT 204.515 -177.645 204.845 -177.315 ;
        RECT 204.515 -179.005 204.845 -178.675 ;
        RECT 204.515 -180.365 204.845 -180.035 ;
        RECT 204.515 -181.725 204.845 -181.395 ;
        RECT 204.515 -183.085 204.845 -182.755 ;
        RECT 204.515 -184.445 204.845 -184.115 ;
        RECT 204.515 -185.805 204.845 -185.475 ;
        RECT 204.515 -187.165 204.845 -186.835 ;
        RECT 204.515 -188.525 204.845 -188.195 ;
        RECT 204.515 -189.885 204.845 -189.555 ;
        RECT 204.515 -191.245 204.845 -190.915 ;
        RECT 204.515 -192.605 204.845 -192.275 ;
        RECT 204.515 -193.965 204.845 -193.635 ;
        RECT 204.515 -195.325 204.845 -194.995 ;
        RECT 204.515 -196.685 204.845 -196.355 ;
        RECT 204.515 -198.045 204.845 -197.715 ;
        RECT 204.515 -199.405 204.845 -199.075 ;
        RECT 204.515 -200.765 204.845 -200.435 ;
        RECT 204.515 -202.125 204.845 -201.795 ;
        RECT 204.515 -203.485 204.845 -203.155 ;
        RECT 204.515 -204.845 204.845 -204.515 ;
        RECT 204.515 -206.205 204.845 -205.875 ;
        RECT 204.515 -207.565 204.845 -207.235 ;
        RECT 204.515 -208.925 204.845 -208.595 ;
        RECT 204.515 -210.285 204.845 -209.955 ;
        RECT 204.515 -211.645 204.845 -211.315 ;
        RECT 204.515 -213.005 204.845 -212.675 ;
        RECT 204.515 -214.365 204.845 -214.035 ;
        RECT 204.515 -215.725 204.845 -215.395 ;
        RECT 204.515 -217.085 204.845 -216.755 ;
        RECT 204.515 -218.445 204.845 -218.115 ;
        RECT 204.515 -219.805 204.845 -219.475 ;
        RECT 204.515 -221.165 204.845 -220.835 ;
        RECT 204.515 -222.525 204.845 -222.195 ;
        RECT 204.515 -223.885 204.845 -223.555 ;
        RECT 204.515 -225.245 204.845 -224.915 ;
        RECT 204.515 -226.605 204.845 -226.275 ;
        RECT 204.515 -227.965 204.845 -227.635 ;
        RECT 204.515 -229.325 204.845 -228.995 ;
        RECT 204.515 -230.685 204.845 -230.355 ;
        RECT 204.515 -232.045 204.845 -231.715 ;
        RECT 204.515 -233.405 204.845 -233.075 ;
        RECT 204.515 -234.765 204.845 -234.435 ;
        RECT 204.515 -236.125 204.845 -235.795 ;
        RECT 204.515 -237.485 204.845 -237.155 ;
        RECT 204.515 -238.845 204.845 -238.515 ;
        RECT 204.515 -241.09 204.845 -239.96 ;
        RECT 204.52 -241.205 204.84 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 244.04 206.205 245.17 ;
        RECT 205.875 242.595 206.205 242.925 ;
        RECT 205.875 241.235 206.205 241.565 ;
        RECT 205.875 239.875 206.205 240.205 ;
        RECT 205.875 238.515 206.205 238.845 ;
        RECT 205.875 237.155 206.205 237.485 ;
        RECT 205.88 237.155 206.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 -0.845 206.205 -0.515 ;
        RECT 205.875 -2.205 206.205 -1.875 ;
        RECT 205.875 -3.565 206.205 -3.235 ;
        RECT 205.88 -3.565 206.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 -123.245 206.205 -122.915 ;
        RECT 205.875 -124.605 206.205 -124.275 ;
        RECT 205.875 -125.965 206.205 -125.635 ;
        RECT 205.875 -127.325 206.205 -126.995 ;
        RECT 205.875 -128.685 206.205 -128.355 ;
        RECT 205.875 -130.045 206.205 -129.715 ;
        RECT 205.875 -131.405 206.205 -131.075 ;
        RECT 205.875 -132.765 206.205 -132.435 ;
        RECT 205.875 -134.125 206.205 -133.795 ;
        RECT 205.875 -135.485 206.205 -135.155 ;
        RECT 205.875 -136.845 206.205 -136.515 ;
        RECT 205.875 -138.205 206.205 -137.875 ;
        RECT 205.875 -139.565 206.205 -139.235 ;
        RECT 205.875 -140.925 206.205 -140.595 ;
        RECT 205.875 -142.285 206.205 -141.955 ;
        RECT 205.875 -143.645 206.205 -143.315 ;
        RECT 205.875 -145.005 206.205 -144.675 ;
        RECT 205.875 -146.365 206.205 -146.035 ;
        RECT 205.875 -147.725 206.205 -147.395 ;
        RECT 205.875 -149.085 206.205 -148.755 ;
        RECT 205.875 -150.445 206.205 -150.115 ;
        RECT 205.875 -151.805 206.205 -151.475 ;
        RECT 205.875 -153.165 206.205 -152.835 ;
        RECT 205.875 -154.525 206.205 -154.195 ;
        RECT 205.875 -155.885 206.205 -155.555 ;
        RECT 205.875 -157.245 206.205 -156.915 ;
        RECT 205.875 -158.605 206.205 -158.275 ;
        RECT 205.875 -159.965 206.205 -159.635 ;
        RECT 205.875 -161.325 206.205 -160.995 ;
        RECT 205.875 -162.685 206.205 -162.355 ;
        RECT 205.875 -164.045 206.205 -163.715 ;
        RECT 205.875 -165.405 206.205 -165.075 ;
        RECT 205.875 -166.765 206.205 -166.435 ;
        RECT 205.875 -168.125 206.205 -167.795 ;
        RECT 205.875 -169.485 206.205 -169.155 ;
        RECT 205.875 -170.845 206.205 -170.515 ;
        RECT 205.875 -172.205 206.205 -171.875 ;
        RECT 205.875 -173.565 206.205 -173.235 ;
        RECT 205.875 -174.925 206.205 -174.595 ;
        RECT 205.875 -176.285 206.205 -175.955 ;
        RECT 205.875 -177.645 206.205 -177.315 ;
        RECT 205.875 -179.005 206.205 -178.675 ;
        RECT 205.875 -180.365 206.205 -180.035 ;
        RECT 205.875 -181.725 206.205 -181.395 ;
        RECT 205.875 -183.085 206.205 -182.755 ;
        RECT 205.875 -184.445 206.205 -184.115 ;
        RECT 205.875 -185.805 206.205 -185.475 ;
        RECT 205.875 -187.165 206.205 -186.835 ;
        RECT 205.875 -188.525 206.205 -188.195 ;
        RECT 205.875 -189.885 206.205 -189.555 ;
        RECT 205.875 -191.245 206.205 -190.915 ;
        RECT 205.875 -192.605 206.205 -192.275 ;
        RECT 205.875 -193.965 206.205 -193.635 ;
        RECT 205.875 -195.325 206.205 -194.995 ;
        RECT 205.875 -196.685 206.205 -196.355 ;
        RECT 205.875 -198.045 206.205 -197.715 ;
        RECT 205.875 -199.405 206.205 -199.075 ;
        RECT 205.875 -200.765 206.205 -200.435 ;
        RECT 205.875 -202.125 206.205 -201.795 ;
        RECT 205.875 -203.485 206.205 -203.155 ;
        RECT 205.875 -204.845 206.205 -204.515 ;
        RECT 205.875 -206.205 206.205 -205.875 ;
        RECT 205.875 -207.565 206.205 -207.235 ;
        RECT 205.875 -208.925 206.205 -208.595 ;
        RECT 205.875 -210.285 206.205 -209.955 ;
        RECT 205.875 -211.645 206.205 -211.315 ;
        RECT 205.875 -213.005 206.205 -212.675 ;
        RECT 205.875 -214.365 206.205 -214.035 ;
        RECT 205.875 -215.725 206.205 -215.395 ;
        RECT 205.875 -217.085 206.205 -216.755 ;
        RECT 205.875 -218.445 206.205 -218.115 ;
        RECT 205.875 -219.805 206.205 -219.475 ;
        RECT 205.875 -221.165 206.205 -220.835 ;
        RECT 205.875 -222.525 206.205 -222.195 ;
        RECT 205.875 -223.885 206.205 -223.555 ;
        RECT 205.875 -225.245 206.205 -224.915 ;
        RECT 205.875 -226.605 206.205 -226.275 ;
        RECT 205.875 -227.965 206.205 -227.635 ;
        RECT 205.875 -229.325 206.205 -228.995 ;
        RECT 205.875 -230.685 206.205 -230.355 ;
        RECT 205.875 -232.045 206.205 -231.715 ;
        RECT 205.875 -233.405 206.205 -233.075 ;
        RECT 205.875 -234.765 206.205 -234.435 ;
        RECT 205.875 -236.125 206.205 -235.795 ;
        RECT 205.875 -237.485 206.205 -237.155 ;
        RECT 205.875 -238.845 206.205 -238.515 ;
        RECT 205.875 -241.09 206.205 -239.96 ;
        RECT 205.88 -241.205 206.2 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 244.04 207.565 245.17 ;
        RECT 207.235 242.595 207.565 242.925 ;
        RECT 207.235 241.235 207.565 241.565 ;
        RECT 207.235 239.875 207.565 240.205 ;
        RECT 207.235 238.515 207.565 238.845 ;
        RECT 207.235 237.155 207.565 237.485 ;
        RECT 207.24 237.155 207.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 -0.845 207.565 -0.515 ;
        RECT 207.235 -2.205 207.565 -1.875 ;
        RECT 207.235 -3.565 207.565 -3.235 ;
        RECT 207.24 -3.565 207.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 -123.245 207.565 -122.915 ;
        RECT 207.235 -124.605 207.565 -124.275 ;
        RECT 207.235 -125.965 207.565 -125.635 ;
        RECT 207.235 -127.325 207.565 -126.995 ;
        RECT 207.235 -128.685 207.565 -128.355 ;
        RECT 207.235 -130.045 207.565 -129.715 ;
        RECT 207.235 -131.405 207.565 -131.075 ;
        RECT 207.235 -132.765 207.565 -132.435 ;
        RECT 207.235 -134.125 207.565 -133.795 ;
        RECT 207.235 -135.485 207.565 -135.155 ;
        RECT 207.235 -136.845 207.565 -136.515 ;
        RECT 207.235 -138.205 207.565 -137.875 ;
        RECT 207.235 -139.565 207.565 -139.235 ;
        RECT 207.235 -140.925 207.565 -140.595 ;
        RECT 207.235 -142.285 207.565 -141.955 ;
        RECT 207.235 -143.645 207.565 -143.315 ;
        RECT 207.235 -145.005 207.565 -144.675 ;
        RECT 207.235 -146.365 207.565 -146.035 ;
        RECT 207.235 -147.725 207.565 -147.395 ;
        RECT 207.235 -149.085 207.565 -148.755 ;
        RECT 207.235 -150.445 207.565 -150.115 ;
        RECT 207.235 -151.805 207.565 -151.475 ;
        RECT 207.235 -153.165 207.565 -152.835 ;
        RECT 207.235 -154.525 207.565 -154.195 ;
        RECT 207.235 -155.885 207.565 -155.555 ;
        RECT 207.235 -157.245 207.565 -156.915 ;
        RECT 207.235 -158.605 207.565 -158.275 ;
        RECT 207.235 -159.965 207.565 -159.635 ;
        RECT 207.235 -161.325 207.565 -160.995 ;
        RECT 207.235 -162.685 207.565 -162.355 ;
        RECT 207.235 -164.045 207.565 -163.715 ;
        RECT 207.235 -165.405 207.565 -165.075 ;
        RECT 207.235 -166.765 207.565 -166.435 ;
        RECT 207.235 -168.125 207.565 -167.795 ;
        RECT 207.235 -169.485 207.565 -169.155 ;
        RECT 207.235 -170.845 207.565 -170.515 ;
        RECT 207.235 -172.205 207.565 -171.875 ;
        RECT 207.235 -173.565 207.565 -173.235 ;
        RECT 207.235 -174.925 207.565 -174.595 ;
        RECT 207.235 -176.285 207.565 -175.955 ;
        RECT 207.235 -177.645 207.565 -177.315 ;
        RECT 207.235 -179.005 207.565 -178.675 ;
        RECT 207.235 -180.365 207.565 -180.035 ;
        RECT 207.235 -181.725 207.565 -181.395 ;
        RECT 207.235 -183.085 207.565 -182.755 ;
        RECT 207.235 -184.445 207.565 -184.115 ;
        RECT 207.235 -185.805 207.565 -185.475 ;
        RECT 207.235 -187.165 207.565 -186.835 ;
        RECT 207.235 -188.525 207.565 -188.195 ;
        RECT 207.235 -189.885 207.565 -189.555 ;
        RECT 207.235 -191.245 207.565 -190.915 ;
        RECT 207.235 -192.605 207.565 -192.275 ;
        RECT 207.235 -193.965 207.565 -193.635 ;
        RECT 207.235 -195.325 207.565 -194.995 ;
        RECT 207.235 -196.685 207.565 -196.355 ;
        RECT 207.235 -198.045 207.565 -197.715 ;
        RECT 207.235 -199.405 207.565 -199.075 ;
        RECT 207.235 -200.765 207.565 -200.435 ;
        RECT 207.235 -202.125 207.565 -201.795 ;
        RECT 207.235 -203.485 207.565 -203.155 ;
        RECT 207.235 -204.845 207.565 -204.515 ;
        RECT 207.235 -206.205 207.565 -205.875 ;
        RECT 207.235 -207.565 207.565 -207.235 ;
        RECT 207.235 -208.925 207.565 -208.595 ;
        RECT 207.235 -210.285 207.565 -209.955 ;
        RECT 207.235 -211.645 207.565 -211.315 ;
        RECT 207.235 -213.005 207.565 -212.675 ;
        RECT 207.235 -214.365 207.565 -214.035 ;
        RECT 207.235 -215.725 207.565 -215.395 ;
        RECT 207.235 -217.085 207.565 -216.755 ;
        RECT 207.235 -218.445 207.565 -218.115 ;
        RECT 207.235 -219.805 207.565 -219.475 ;
        RECT 207.235 -221.165 207.565 -220.835 ;
        RECT 207.235 -222.525 207.565 -222.195 ;
        RECT 207.235 -223.885 207.565 -223.555 ;
        RECT 207.235 -225.245 207.565 -224.915 ;
        RECT 207.235 -226.605 207.565 -226.275 ;
        RECT 207.235 -227.965 207.565 -227.635 ;
        RECT 207.235 -229.325 207.565 -228.995 ;
        RECT 207.235 -230.685 207.565 -230.355 ;
        RECT 207.235 -232.045 207.565 -231.715 ;
        RECT 207.235 -233.405 207.565 -233.075 ;
        RECT 207.235 -234.765 207.565 -234.435 ;
        RECT 207.235 -236.125 207.565 -235.795 ;
        RECT 207.235 -237.485 207.565 -237.155 ;
        RECT 207.235 -238.845 207.565 -238.515 ;
        RECT 207.235 -241.09 207.565 -239.96 ;
        RECT 207.24 -241.205 207.56 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 244.04 208.925 245.17 ;
        RECT 208.595 242.595 208.925 242.925 ;
        RECT 208.595 241.235 208.925 241.565 ;
        RECT 208.595 239.875 208.925 240.205 ;
        RECT 208.595 238.515 208.925 238.845 ;
        RECT 208.595 237.155 208.925 237.485 ;
        RECT 208.6 237.155 208.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 -0.845 208.925 -0.515 ;
        RECT 208.595 -2.205 208.925 -1.875 ;
        RECT 208.595 -3.565 208.925 -3.235 ;
        RECT 208.6 -3.565 208.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 -123.245 208.925 -122.915 ;
        RECT 208.595 -124.605 208.925 -124.275 ;
        RECT 208.595 -125.965 208.925 -125.635 ;
        RECT 208.595 -127.325 208.925 -126.995 ;
        RECT 208.595 -128.685 208.925 -128.355 ;
        RECT 208.595 -130.045 208.925 -129.715 ;
        RECT 208.595 -131.405 208.925 -131.075 ;
        RECT 208.595 -132.765 208.925 -132.435 ;
        RECT 208.595 -134.125 208.925 -133.795 ;
        RECT 208.595 -135.485 208.925 -135.155 ;
        RECT 208.595 -136.845 208.925 -136.515 ;
        RECT 208.595 -138.205 208.925 -137.875 ;
        RECT 208.595 -139.565 208.925 -139.235 ;
        RECT 208.595 -140.925 208.925 -140.595 ;
        RECT 208.595 -142.285 208.925 -141.955 ;
        RECT 208.595 -143.645 208.925 -143.315 ;
        RECT 208.595 -145.005 208.925 -144.675 ;
        RECT 208.595 -146.365 208.925 -146.035 ;
        RECT 208.595 -147.725 208.925 -147.395 ;
        RECT 208.595 -149.085 208.925 -148.755 ;
        RECT 208.595 -150.445 208.925 -150.115 ;
        RECT 208.595 -151.805 208.925 -151.475 ;
        RECT 208.595 -153.165 208.925 -152.835 ;
        RECT 208.595 -154.525 208.925 -154.195 ;
        RECT 208.595 -155.885 208.925 -155.555 ;
        RECT 208.595 -157.245 208.925 -156.915 ;
        RECT 208.595 -158.605 208.925 -158.275 ;
        RECT 208.595 -159.965 208.925 -159.635 ;
        RECT 208.595 -161.325 208.925 -160.995 ;
        RECT 208.595 -162.685 208.925 -162.355 ;
        RECT 208.595 -164.045 208.925 -163.715 ;
        RECT 208.595 -165.405 208.925 -165.075 ;
        RECT 208.595 -166.765 208.925 -166.435 ;
        RECT 208.595 -168.125 208.925 -167.795 ;
        RECT 208.595 -169.485 208.925 -169.155 ;
        RECT 208.595 -170.845 208.925 -170.515 ;
        RECT 208.595 -172.205 208.925 -171.875 ;
        RECT 208.595 -173.565 208.925 -173.235 ;
        RECT 208.595 -174.925 208.925 -174.595 ;
        RECT 208.595 -176.285 208.925 -175.955 ;
        RECT 208.595 -177.645 208.925 -177.315 ;
        RECT 208.595 -179.005 208.925 -178.675 ;
        RECT 208.595 -180.365 208.925 -180.035 ;
        RECT 208.595 -181.725 208.925 -181.395 ;
        RECT 208.595 -183.085 208.925 -182.755 ;
        RECT 208.595 -184.445 208.925 -184.115 ;
        RECT 208.595 -185.805 208.925 -185.475 ;
        RECT 208.595 -187.165 208.925 -186.835 ;
        RECT 208.595 -188.525 208.925 -188.195 ;
        RECT 208.595 -189.885 208.925 -189.555 ;
        RECT 208.595 -191.245 208.925 -190.915 ;
        RECT 208.595 -192.605 208.925 -192.275 ;
        RECT 208.595 -193.965 208.925 -193.635 ;
        RECT 208.595 -195.325 208.925 -194.995 ;
        RECT 208.595 -196.685 208.925 -196.355 ;
        RECT 208.595 -198.045 208.925 -197.715 ;
        RECT 208.595 -199.405 208.925 -199.075 ;
        RECT 208.595 -200.765 208.925 -200.435 ;
        RECT 208.595 -202.125 208.925 -201.795 ;
        RECT 208.595 -203.485 208.925 -203.155 ;
        RECT 208.595 -204.845 208.925 -204.515 ;
        RECT 208.595 -206.205 208.925 -205.875 ;
        RECT 208.595 -207.565 208.925 -207.235 ;
        RECT 208.595 -208.925 208.925 -208.595 ;
        RECT 208.595 -210.285 208.925 -209.955 ;
        RECT 208.595 -211.645 208.925 -211.315 ;
        RECT 208.595 -213.005 208.925 -212.675 ;
        RECT 208.595 -214.365 208.925 -214.035 ;
        RECT 208.595 -215.725 208.925 -215.395 ;
        RECT 208.595 -217.085 208.925 -216.755 ;
        RECT 208.595 -218.445 208.925 -218.115 ;
        RECT 208.595 -219.805 208.925 -219.475 ;
        RECT 208.595 -221.165 208.925 -220.835 ;
        RECT 208.595 -222.525 208.925 -222.195 ;
        RECT 208.595 -223.885 208.925 -223.555 ;
        RECT 208.595 -225.245 208.925 -224.915 ;
        RECT 208.595 -226.605 208.925 -226.275 ;
        RECT 208.595 -227.965 208.925 -227.635 ;
        RECT 208.595 -229.325 208.925 -228.995 ;
        RECT 208.595 -230.685 208.925 -230.355 ;
        RECT 208.595 -232.045 208.925 -231.715 ;
        RECT 208.595 -233.405 208.925 -233.075 ;
        RECT 208.595 -234.765 208.925 -234.435 ;
        RECT 208.595 -236.125 208.925 -235.795 ;
        RECT 208.595 -237.485 208.925 -237.155 ;
        RECT 208.595 -238.845 208.925 -238.515 ;
        RECT 208.595 -241.09 208.925 -239.96 ;
        RECT 208.6 -241.205 208.92 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 244.04 210.285 245.17 ;
        RECT 209.955 242.595 210.285 242.925 ;
        RECT 209.955 241.235 210.285 241.565 ;
        RECT 209.955 239.875 210.285 240.205 ;
        RECT 209.955 238.515 210.285 238.845 ;
        RECT 209.955 237.155 210.285 237.485 ;
        RECT 209.96 237.155 210.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 -127.325 210.285 -126.995 ;
        RECT 209.955 -128.685 210.285 -128.355 ;
        RECT 209.955 -130.045 210.285 -129.715 ;
        RECT 209.955 -131.405 210.285 -131.075 ;
        RECT 209.955 -132.765 210.285 -132.435 ;
        RECT 209.955 -134.125 210.285 -133.795 ;
        RECT 209.955 -135.485 210.285 -135.155 ;
        RECT 209.955 -136.845 210.285 -136.515 ;
        RECT 209.955 -138.205 210.285 -137.875 ;
        RECT 209.955 -139.565 210.285 -139.235 ;
        RECT 209.955 -140.925 210.285 -140.595 ;
        RECT 209.955 -142.285 210.285 -141.955 ;
        RECT 209.955 -143.645 210.285 -143.315 ;
        RECT 209.955 -145.005 210.285 -144.675 ;
        RECT 209.955 -146.365 210.285 -146.035 ;
        RECT 209.955 -147.725 210.285 -147.395 ;
        RECT 209.955 -149.085 210.285 -148.755 ;
        RECT 209.955 -150.445 210.285 -150.115 ;
        RECT 209.955 -151.805 210.285 -151.475 ;
        RECT 209.955 -153.165 210.285 -152.835 ;
        RECT 209.955 -154.525 210.285 -154.195 ;
        RECT 209.955 -155.885 210.285 -155.555 ;
        RECT 209.955 -157.245 210.285 -156.915 ;
        RECT 209.955 -158.605 210.285 -158.275 ;
        RECT 209.955 -159.965 210.285 -159.635 ;
        RECT 209.955 -161.325 210.285 -160.995 ;
        RECT 209.955 -162.685 210.285 -162.355 ;
        RECT 209.955 -164.045 210.285 -163.715 ;
        RECT 209.955 -165.405 210.285 -165.075 ;
        RECT 209.955 -166.765 210.285 -166.435 ;
        RECT 209.955 -168.125 210.285 -167.795 ;
        RECT 209.955 -169.485 210.285 -169.155 ;
        RECT 209.955 -170.845 210.285 -170.515 ;
        RECT 209.955 -172.205 210.285 -171.875 ;
        RECT 209.955 -173.565 210.285 -173.235 ;
        RECT 209.955 -174.925 210.285 -174.595 ;
        RECT 209.955 -176.285 210.285 -175.955 ;
        RECT 209.955 -177.645 210.285 -177.315 ;
        RECT 209.955 -179.005 210.285 -178.675 ;
        RECT 209.955 -180.365 210.285 -180.035 ;
        RECT 209.955 -181.725 210.285 -181.395 ;
        RECT 209.955 -183.085 210.285 -182.755 ;
        RECT 209.955 -184.445 210.285 -184.115 ;
        RECT 209.955 -185.805 210.285 -185.475 ;
        RECT 209.955 -187.165 210.285 -186.835 ;
        RECT 209.955 -188.525 210.285 -188.195 ;
        RECT 209.955 -189.885 210.285 -189.555 ;
        RECT 209.955 -191.245 210.285 -190.915 ;
        RECT 209.955 -192.605 210.285 -192.275 ;
        RECT 209.955 -193.965 210.285 -193.635 ;
        RECT 209.955 -195.325 210.285 -194.995 ;
        RECT 209.955 -196.685 210.285 -196.355 ;
        RECT 209.955 -198.045 210.285 -197.715 ;
        RECT 209.955 -199.405 210.285 -199.075 ;
        RECT 209.955 -200.765 210.285 -200.435 ;
        RECT 209.955 -202.125 210.285 -201.795 ;
        RECT 209.955 -203.485 210.285 -203.155 ;
        RECT 209.955 -204.845 210.285 -204.515 ;
        RECT 209.955 -206.205 210.285 -205.875 ;
        RECT 209.955 -207.565 210.285 -207.235 ;
        RECT 209.955 -208.925 210.285 -208.595 ;
        RECT 209.955 -210.285 210.285 -209.955 ;
        RECT 209.955 -211.645 210.285 -211.315 ;
        RECT 209.955 -213.005 210.285 -212.675 ;
        RECT 209.955 -214.365 210.285 -214.035 ;
        RECT 209.955 -215.725 210.285 -215.395 ;
        RECT 209.955 -217.085 210.285 -216.755 ;
        RECT 209.955 -218.445 210.285 -218.115 ;
        RECT 209.955 -219.805 210.285 -219.475 ;
        RECT 209.955 -221.165 210.285 -220.835 ;
        RECT 209.955 -222.525 210.285 -222.195 ;
        RECT 209.955 -223.885 210.285 -223.555 ;
        RECT 209.955 -225.245 210.285 -224.915 ;
        RECT 209.955 -226.605 210.285 -226.275 ;
        RECT 209.955 -227.965 210.285 -227.635 ;
        RECT 209.955 -229.325 210.285 -228.995 ;
        RECT 209.955 -230.685 210.285 -230.355 ;
        RECT 209.955 -232.045 210.285 -231.715 ;
        RECT 209.955 -233.405 210.285 -233.075 ;
        RECT 209.955 -234.765 210.285 -234.435 ;
        RECT 209.955 -236.125 210.285 -235.795 ;
        RECT 209.955 -237.485 210.285 -237.155 ;
        RECT 209.955 -238.845 210.285 -238.515 ;
        RECT 209.955 -241.09 210.285 -239.96 ;
        RECT 209.96 -241.205 210.28 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.41 -125.535 210.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 244.04 211.645 245.17 ;
        RECT 211.315 242.595 211.645 242.925 ;
        RECT 211.315 241.235 211.645 241.565 ;
        RECT 211.315 239.875 211.645 240.205 ;
        RECT 211.315 238.515 211.645 238.845 ;
        RECT 211.315 237.155 211.645 237.485 ;
        RECT 211.32 237.155 211.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 -0.845 211.645 -0.515 ;
        RECT 211.315 -2.205 211.645 -1.875 ;
        RECT 211.315 -3.565 211.645 -3.235 ;
        RECT 211.32 -3.565 211.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 244.04 213.005 245.17 ;
        RECT 212.675 242.595 213.005 242.925 ;
        RECT 212.675 241.235 213.005 241.565 ;
        RECT 212.675 239.875 213.005 240.205 ;
        RECT 212.675 238.515 213.005 238.845 ;
        RECT 212.675 237.155 213.005 237.485 ;
        RECT 212.68 237.155 213 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 -0.845 213.005 -0.515 ;
        RECT 212.675 -2.205 213.005 -1.875 ;
        RECT 212.675 -3.565 213.005 -3.235 ;
        RECT 212.68 -3.565 213 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 244.04 214.365 245.17 ;
        RECT 214.035 242.595 214.365 242.925 ;
        RECT 214.035 241.235 214.365 241.565 ;
        RECT 214.035 239.875 214.365 240.205 ;
        RECT 214.035 238.515 214.365 238.845 ;
        RECT 214.035 237.155 214.365 237.485 ;
        RECT 214.04 237.155 214.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 -0.845 214.365 -0.515 ;
        RECT 214.035 -2.205 214.365 -1.875 ;
        RECT 214.035 -3.565 214.365 -3.235 ;
        RECT 214.04 -3.565 214.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 -123.245 214.365 -122.915 ;
        RECT 214.035 -124.605 214.365 -124.275 ;
        RECT 214.035 -125.965 214.365 -125.635 ;
        RECT 214.035 -127.325 214.365 -126.995 ;
        RECT 214.035 -128.685 214.365 -128.355 ;
        RECT 214.035 -130.045 214.365 -129.715 ;
        RECT 214.035 -131.405 214.365 -131.075 ;
        RECT 214.035 -132.765 214.365 -132.435 ;
        RECT 214.035 -134.125 214.365 -133.795 ;
        RECT 214.035 -135.485 214.365 -135.155 ;
        RECT 214.035 -136.845 214.365 -136.515 ;
        RECT 214.035 -138.205 214.365 -137.875 ;
        RECT 214.035 -139.565 214.365 -139.235 ;
        RECT 214.035 -140.925 214.365 -140.595 ;
        RECT 214.035 -142.285 214.365 -141.955 ;
        RECT 214.035 -143.645 214.365 -143.315 ;
        RECT 214.035 -145.005 214.365 -144.675 ;
        RECT 214.035 -146.365 214.365 -146.035 ;
        RECT 214.035 -147.725 214.365 -147.395 ;
        RECT 214.035 -149.085 214.365 -148.755 ;
        RECT 214.035 -150.445 214.365 -150.115 ;
        RECT 214.035 -151.805 214.365 -151.475 ;
        RECT 214.035 -153.165 214.365 -152.835 ;
        RECT 214.035 -154.525 214.365 -154.195 ;
        RECT 214.035 -155.885 214.365 -155.555 ;
        RECT 214.035 -157.245 214.365 -156.915 ;
        RECT 214.035 -158.605 214.365 -158.275 ;
        RECT 214.035 -159.965 214.365 -159.635 ;
        RECT 214.035 -161.325 214.365 -160.995 ;
        RECT 214.035 -162.685 214.365 -162.355 ;
        RECT 214.035 -164.045 214.365 -163.715 ;
        RECT 214.035 -165.405 214.365 -165.075 ;
        RECT 214.035 -166.765 214.365 -166.435 ;
        RECT 214.035 -168.125 214.365 -167.795 ;
        RECT 214.035 -169.485 214.365 -169.155 ;
        RECT 214.035 -170.845 214.365 -170.515 ;
        RECT 214.035 -172.205 214.365 -171.875 ;
        RECT 214.035 -173.565 214.365 -173.235 ;
        RECT 214.035 -174.925 214.365 -174.595 ;
        RECT 214.035 -176.285 214.365 -175.955 ;
        RECT 214.035 -177.645 214.365 -177.315 ;
        RECT 214.035 -179.005 214.365 -178.675 ;
        RECT 214.035 -180.365 214.365 -180.035 ;
        RECT 214.035 -181.725 214.365 -181.395 ;
        RECT 214.035 -183.085 214.365 -182.755 ;
        RECT 214.035 -184.445 214.365 -184.115 ;
        RECT 214.035 -185.805 214.365 -185.475 ;
        RECT 214.035 -187.165 214.365 -186.835 ;
        RECT 214.035 -188.525 214.365 -188.195 ;
        RECT 214.035 -189.885 214.365 -189.555 ;
        RECT 214.035 -191.245 214.365 -190.915 ;
        RECT 214.035 -192.605 214.365 -192.275 ;
        RECT 214.035 -193.965 214.365 -193.635 ;
        RECT 214.035 -195.325 214.365 -194.995 ;
        RECT 214.035 -196.685 214.365 -196.355 ;
        RECT 214.035 -198.045 214.365 -197.715 ;
        RECT 214.035 -199.405 214.365 -199.075 ;
        RECT 214.035 -200.765 214.365 -200.435 ;
        RECT 214.035 -202.125 214.365 -201.795 ;
        RECT 214.035 -203.485 214.365 -203.155 ;
        RECT 214.035 -204.845 214.365 -204.515 ;
        RECT 214.035 -206.205 214.365 -205.875 ;
        RECT 214.035 -207.565 214.365 -207.235 ;
        RECT 214.035 -208.925 214.365 -208.595 ;
        RECT 214.035 -210.285 214.365 -209.955 ;
        RECT 214.035 -211.645 214.365 -211.315 ;
        RECT 214.035 -213.005 214.365 -212.675 ;
        RECT 214.035 -214.365 214.365 -214.035 ;
        RECT 214.035 -215.725 214.365 -215.395 ;
        RECT 214.035 -217.085 214.365 -216.755 ;
        RECT 214.035 -218.445 214.365 -218.115 ;
        RECT 214.035 -219.805 214.365 -219.475 ;
        RECT 214.035 -221.165 214.365 -220.835 ;
        RECT 214.035 -222.525 214.365 -222.195 ;
        RECT 214.035 -223.885 214.365 -223.555 ;
        RECT 214.035 -225.245 214.365 -224.915 ;
        RECT 214.035 -226.605 214.365 -226.275 ;
        RECT 214.035 -227.965 214.365 -227.635 ;
        RECT 214.035 -229.325 214.365 -228.995 ;
        RECT 214.035 -230.685 214.365 -230.355 ;
        RECT 214.035 -232.045 214.365 -231.715 ;
        RECT 214.035 -233.405 214.365 -233.075 ;
        RECT 214.035 -234.765 214.365 -234.435 ;
        RECT 214.035 -236.125 214.365 -235.795 ;
        RECT 214.035 -237.485 214.365 -237.155 ;
        RECT 214.035 -238.845 214.365 -238.515 ;
        RECT 214.035 -241.09 214.365 -239.96 ;
        RECT 214.04 -241.205 214.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 244.04 215.725 245.17 ;
        RECT 215.395 242.595 215.725 242.925 ;
        RECT 215.395 241.235 215.725 241.565 ;
        RECT 215.395 239.875 215.725 240.205 ;
        RECT 215.395 238.515 215.725 238.845 ;
        RECT 215.395 237.155 215.725 237.485 ;
        RECT 215.4 237.155 215.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 -0.845 215.725 -0.515 ;
        RECT 215.395 -2.205 215.725 -1.875 ;
        RECT 215.395 -3.565 215.725 -3.235 ;
        RECT 215.4 -3.565 215.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 -123.245 215.725 -122.915 ;
        RECT 215.395 -124.605 215.725 -124.275 ;
        RECT 215.395 -125.965 215.725 -125.635 ;
        RECT 215.395 -127.325 215.725 -126.995 ;
        RECT 215.395 -128.685 215.725 -128.355 ;
        RECT 215.395 -130.045 215.725 -129.715 ;
        RECT 215.395 -131.405 215.725 -131.075 ;
        RECT 215.395 -132.765 215.725 -132.435 ;
        RECT 215.395 -134.125 215.725 -133.795 ;
        RECT 215.395 -135.485 215.725 -135.155 ;
        RECT 215.395 -136.845 215.725 -136.515 ;
        RECT 215.395 -138.205 215.725 -137.875 ;
        RECT 215.395 -139.565 215.725 -139.235 ;
        RECT 215.395 -140.925 215.725 -140.595 ;
        RECT 215.395 -142.285 215.725 -141.955 ;
        RECT 215.395 -143.645 215.725 -143.315 ;
        RECT 215.395 -145.005 215.725 -144.675 ;
        RECT 215.395 -146.365 215.725 -146.035 ;
        RECT 215.395 -147.725 215.725 -147.395 ;
        RECT 215.395 -149.085 215.725 -148.755 ;
        RECT 215.395 -150.445 215.725 -150.115 ;
        RECT 215.395 -151.805 215.725 -151.475 ;
        RECT 215.395 -153.165 215.725 -152.835 ;
        RECT 215.395 -154.525 215.725 -154.195 ;
        RECT 215.395 -155.885 215.725 -155.555 ;
        RECT 215.395 -157.245 215.725 -156.915 ;
        RECT 215.395 -158.605 215.725 -158.275 ;
        RECT 215.395 -159.965 215.725 -159.635 ;
        RECT 215.395 -161.325 215.725 -160.995 ;
        RECT 215.395 -162.685 215.725 -162.355 ;
        RECT 215.395 -164.045 215.725 -163.715 ;
        RECT 215.395 -165.405 215.725 -165.075 ;
        RECT 215.395 -166.765 215.725 -166.435 ;
        RECT 215.395 -168.125 215.725 -167.795 ;
        RECT 215.395 -169.485 215.725 -169.155 ;
        RECT 215.395 -170.845 215.725 -170.515 ;
        RECT 215.395 -172.205 215.725 -171.875 ;
        RECT 215.395 -173.565 215.725 -173.235 ;
        RECT 215.395 -174.925 215.725 -174.595 ;
        RECT 215.395 -176.285 215.725 -175.955 ;
        RECT 215.395 -177.645 215.725 -177.315 ;
        RECT 215.395 -179.005 215.725 -178.675 ;
        RECT 215.395 -180.365 215.725 -180.035 ;
        RECT 215.395 -181.725 215.725 -181.395 ;
        RECT 215.395 -183.085 215.725 -182.755 ;
        RECT 215.395 -184.445 215.725 -184.115 ;
        RECT 215.395 -185.805 215.725 -185.475 ;
        RECT 215.395 -187.165 215.725 -186.835 ;
        RECT 215.395 -188.525 215.725 -188.195 ;
        RECT 215.395 -189.885 215.725 -189.555 ;
        RECT 215.395 -191.245 215.725 -190.915 ;
        RECT 215.395 -192.605 215.725 -192.275 ;
        RECT 215.395 -193.965 215.725 -193.635 ;
        RECT 215.395 -195.325 215.725 -194.995 ;
        RECT 215.395 -196.685 215.725 -196.355 ;
        RECT 215.395 -198.045 215.725 -197.715 ;
        RECT 215.395 -199.405 215.725 -199.075 ;
        RECT 215.395 -200.765 215.725 -200.435 ;
        RECT 215.395 -202.125 215.725 -201.795 ;
        RECT 215.395 -203.485 215.725 -203.155 ;
        RECT 215.395 -204.845 215.725 -204.515 ;
        RECT 215.395 -206.205 215.725 -205.875 ;
        RECT 215.395 -207.565 215.725 -207.235 ;
        RECT 215.395 -208.925 215.725 -208.595 ;
        RECT 215.395 -210.285 215.725 -209.955 ;
        RECT 215.395 -211.645 215.725 -211.315 ;
        RECT 215.395 -213.005 215.725 -212.675 ;
        RECT 215.395 -214.365 215.725 -214.035 ;
        RECT 215.395 -215.725 215.725 -215.395 ;
        RECT 215.395 -217.085 215.725 -216.755 ;
        RECT 215.395 -218.445 215.725 -218.115 ;
        RECT 215.395 -219.805 215.725 -219.475 ;
        RECT 215.395 -221.165 215.725 -220.835 ;
        RECT 215.395 -222.525 215.725 -222.195 ;
        RECT 215.395 -223.885 215.725 -223.555 ;
        RECT 215.395 -225.245 215.725 -224.915 ;
        RECT 215.395 -226.605 215.725 -226.275 ;
        RECT 215.395 -227.965 215.725 -227.635 ;
        RECT 215.395 -229.325 215.725 -228.995 ;
        RECT 215.395 -230.685 215.725 -230.355 ;
        RECT 215.395 -232.045 215.725 -231.715 ;
        RECT 215.395 -233.405 215.725 -233.075 ;
        RECT 215.395 -234.765 215.725 -234.435 ;
        RECT 215.395 -236.125 215.725 -235.795 ;
        RECT 215.395 -237.485 215.725 -237.155 ;
        RECT 215.395 -238.845 215.725 -238.515 ;
        RECT 215.395 -241.09 215.725 -239.96 ;
        RECT 215.4 -241.205 215.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 244.04 217.085 245.17 ;
        RECT 216.755 242.595 217.085 242.925 ;
        RECT 216.755 241.235 217.085 241.565 ;
        RECT 216.755 239.875 217.085 240.205 ;
        RECT 216.755 238.515 217.085 238.845 ;
        RECT 216.755 237.155 217.085 237.485 ;
        RECT 216.76 237.155 217.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 -0.845 217.085 -0.515 ;
        RECT 216.755 -2.205 217.085 -1.875 ;
        RECT 216.755 -3.565 217.085 -3.235 ;
        RECT 216.76 -3.565 217.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 -123.245 217.085 -122.915 ;
        RECT 216.755 -124.605 217.085 -124.275 ;
        RECT 216.755 -125.965 217.085 -125.635 ;
        RECT 216.755 -127.325 217.085 -126.995 ;
        RECT 216.755 -128.685 217.085 -128.355 ;
        RECT 216.755 -130.045 217.085 -129.715 ;
        RECT 216.755 -131.405 217.085 -131.075 ;
        RECT 216.755 -132.765 217.085 -132.435 ;
        RECT 216.755 -134.125 217.085 -133.795 ;
        RECT 216.755 -135.485 217.085 -135.155 ;
        RECT 216.755 -136.845 217.085 -136.515 ;
        RECT 216.755 -138.205 217.085 -137.875 ;
        RECT 216.755 -139.565 217.085 -139.235 ;
        RECT 216.755 -140.925 217.085 -140.595 ;
        RECT 216.755 -142.285 217.085 -141.955 ;
        RECT 216.755 -143.645 217.085 -143.315 ;
        RECT 216.755 -145.005 217.085 -144.675 ;
        RECT 216.755 -146.365 217.085 -146.035 ;
        RECT 216.755 -147.725 217.085 -147.395 ;
        RECT 216.755 -149.085 217.085 -148.755 ;
        RECT 216.755 -150.445 217.085 -150.115 ;
        RECT 216.755 -151.805 217.085 -151.475 ;
        RECT 216.755 -153.165 217.085 -152.835 ;
        RECT 216.755 -154.525 217.085 -154.195 ;
        RECT 216.755 -155.885 217.085 -155.555 ;
        RECT 216.755 -157.245 217.085 -156.915 ;
        RECT 216.755 -158.605 217.085 -158.275 ;
        RECT 216.755 -159.965 217.085 -159.635 ;
        RECT 216.755 -161.325 217.085 -160.995 ;
        RECT 216.755 -162.685 217.085 -162.355 ;
        RECT 216.755 -164.045 217.085 -163.715 ;
        RECT 216.755 -165.405 217.085 -165.075 ;
        RECT 216.755 -166.765 217.085 -166.435 ;
        RECT 216.755 -168.125 217.085 -167.795 ;
        RECT 216.755 -169.485 217.085 -169.155 ;
        RECT 216.755 -170.845 217.085 -170.515 ;
        RECT 216.755 -172.205 217.085 -171.875 ;
        RECT 216.755 -173.565 217.085 -173.235 ;
        RECT 216.755 -174.925 217.085 -174.595 ;
        RECT 216.755 -176.285 217.085 -175.955 ;
        RECT 216.755 -177.645 217.085 -177.315 ;
        RECT 216.755 -179.005 217.085 -178.675 ;
        RECT 216.755 -180.365 217.085 -180.035 ;
        RECT 216.755 -181.725 217.085 -181.395 ;
        RECT 216.755 -183.085 217.085 -182.755 ;
        RECT 216.755 -184.445 217.085 -184.115 ;
        RECT 216.755 -185.805 217.085 -185.475 ;
        RECT 216.755 -187.165 217.085 -186.835 ;
        RECT 216.755 -188.525 217.085 -188.195 ;
        RECT 216.755 -189.885 217.085 -189.555 ;
        RECT 216.755 -191.245 217.085 -190.915 ;
        RECT 216.755 -192.605 217.085 -192.275 ;
        RECT 216.755 -193.965 217.085 -193.635 ;
        RECT 216.755 -195.325 217.085 -194.995 ;
        RECT 216.755 -196.685 217.085 -196.355 ;
        RECT 216.755 -198.045 217.085 -197.715 ;
        RECT 216.755 -199.405 217.085 -199.075 ;
        RECT 216.755 -200.765 217.085 -200.435 ;
        RECT 216.755 -202.125 217.085 -201.795 ;
        RECT 216.755 -203.485 217.085 -203.155 ;
        RECT 216.755 -204.845 217.085 -204.515 ;
        RECT 216.755 -206.205 217.085 -205.875 ;
        RECT 216.755 -207.565 217.085 -207.235 ;
        RECT 216.755 -208.925 217.085 -208.595 ;
        RECT 216.755 -210.285 217.085 -209.955 ;
        RECT 216.755 -211.645 217.085 -211.315 ;
        RECT 216.755 -213.005 217.085 -212.675 ;
        RECT 216.755 -214.365 217.085 -214.035 ;
        RECT 216.755 -215.725 217.085 -215.395 ;
        RECT 216.755 -217.085 217.085 -216.755 ;
        RECT 216.755 -218.445 217.085 -218.115 ;
        RECT 216.755 -219.805 217.085 -219.475 ;
        RECT 216.755 -221.165 217.085 -220.835 ;
        RECT 216.755 -222.525 217.085 -222.195 ;
        RECT 216.755 -223.885 217.085 -223.555 ;
        RECT 216.755 -225.245 217.085 -224.915 ;
        RECT 216.755 -226.605 217.085 -226.275 ;
        RECT 216.755 -227.965 217.085 -227.635 ;
        RECT 216.755 -229.325 217.085 -228.995 ;
        RECT 216.755 -230.685 217.085 -230.355 ;
        RECT 216.755 -232.045 217.085 -231.715 ;
        RECT 216.755 -233.405 217.085 -233.075 ;
        RECT 216.755 -234.765 217.085 -234.435 ;
        RECT 216.755 -236.125 217.085 -235.795 ;
        RECT 216.755 -237.485 217.085 -237.155 ;
        RECT 216.755 -238.845 217.085 -238.515 ;
        RECT 216.755 -241.09 217.085 -239.96 ;
        RECT 216.76 -241.205 217.08 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 244.04 218.445 245.17 ;
        RECT 218.115 242.595 218.445 242.925 ;
        RECT 218.115 241.235 218.445 241.565 ;
        RECT 218.115 239.875 218.445 240.205 ;
        RECT 218.115 238.515 218.445 238.845 ;
        RECT 218.115 237.155 218.445 237.485 ;
        RECT 218.12 237.155 218.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 -0.845 218.445 -0.515 ;
        RECT 218.115 -2.205 218.445 -1.875 ;
        RECT 218.115 -3.565 218.445 -3.235 ;
        RECT 218.12 -3.565 218.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 -217.085 218.445 -216.755 ;
        RECT 218.115 -218.445 218.445 -218.115 ;
        RECT 218.115 -219.805 218.445 -219.475 ;
        RECT 218.115 -221.165 218.445 -220.835 ;
        RECT 218.115 -222.525 218.445 -222.195 ;
        RECT 218.115 -223.885 218.445 -223.555 ;
        RECT 218.115 -225.245 218.445 -224.915 ;
        RECT 218.115 -226.605 218.445 -226.275 ;
        RECT 218.115 -227.965 218.445 -227.635 ;
        RECT 218.115 -229.325 218.445 -228.995 ;
        RECT 218.115 -230.685 218.445 -230.355 ;
        RECT 218.115 -232.045 218.445 -231.715 ;
        RECT 218.115 -233.405 218.445 -233.075 ;
        RECT 218.115 -234.765 218.445 -234.435 ;
        RECT 218.115 -236.125 218.445 -235.795 ;
        RECT 218.115 -237.485 218.445 -237.155 ;
        RECT 218.115 -238.845 218.445 -238.515 ;
        RECT 218.115 -241.09 218.445 -239.96 ;
        RECT 218.12 -241.205 218.44 -122.24 ;
        RECT 218.115 -123.245 218.445 -122.915 ;
        RECT 218.115 -124.605 218.445 -124.275 ;
        RECT 218.115 -125.965 218.445 -125.635 ;
        RECT 218.115 -127.325 218.445 -126.995 ;
        RECT 218.115 -128.685 218.445 -128.355 ;
        RECT 218.115 -130.045 218.445 -129.715 ;
        RECT 218.115 -131.405 218.445 -131.075 ;
        RECT 218.115 -132.765 218.445 -132.435 ;
        RECT 218.115 -134.125 218.445 -133.795 ;
        RECT 218.115 -135.485 218.445 -135.155 ;
        RECT 218.115 -136.845 218.445 -136.515 ;
        RECT 218.115 -138.205 218.445 -137.875 ;
        RECT 218.115 -139.565 218.445 -139.235 ;
        RECT 218.115 -140.925 218.445 -140.595 ;
        RECT 218.115 -142.285 218.445 -141.955 ;
        RECT 218.115 -143.645 218.445 -143.315 ;
        RECT 218.115 -145.005 218.445 -144.675 ;
        RECT 218.115 -146.365 218.445 -146.035 ;
        RECT 218.115 -147.725 218.445 -147.395 ;
        RECT 218.115 -149.085 218.445 -148.755 ;
        RECT 218.115 -150.445 218.445 -150.115 ;
        RECT 218.115 -151.805 218.445 -151.475 ;
        RECT 218.115 -153.165 218.445 -152.835 ;
        RECT 218.115 -154.525 218.445 -154.195 ;
        RECT 218.115 -155.885 218.445 -155.555 ;
        RECT 218.115 -157.245 218.445 -156.915 ;
        RECT 218.115 -158.605 218.445 -158.275 ;
        RECT 218.115 -159.965 218.445 -159.635 ;
        RECT 218.115 -161.325 218.445 -160.995 ;
        RECT 218.115 -162.685 218.445 -162.355 ;
        RECT 218.115 -164.045 218.445 -163.715 ;
        RECT 218.115 -165.405 218.445 -165.075 ;
        RECT 218.115 -166.765 218.445 -166.435 ;
        RECT 218.115 -168.125 218.445 -167.795 ;
        RECT 218.115 -169.485 218.445 -169.155 ;
        RECT 218.115 -170.845 218.445 -170.515 ;
        RECT 218.115 -172.205 218.445 -171.875 ;
        RECT 218.115 -173.565 218.445 -173.235 ;
        RECT 218.115 -174.925 218.445 -174.595 ;
        RECT 218.115 -176.285 218.445 -175.955 ;
        RECT 218.115 -177.645 218.445 -177.315 ;
        RECT 218.115 -179.005 218.445 -178.675 ;
        RECT 218.115 -180.365 218.445 -180.035 ;
        RECT 218.115 -181.725 218.445 -181.395 ;
        RECT 218.115 -183.085 218.445 -182.755 ;
        RECT 218.115 -184.445 218.445 -184.115 ;
        RECT 218.115 -185.805 218.445 -185.475 ;
        RECT 218.115 -187.165 218.445 -186.835 ;
        RECT 218.115 -188.525 218.445 -188.195 ;
        RECT 218.115 -189.885 218.445 -189.555 ;
        RECT 218.115 -191.245 218.445 -190.915 ;
        RECT 218.115 -192.605 218.445 -192.275 ;
        RECT 218.115 -193.965 218.445 -193.635 ;
        RECT 218.115 -195.325 218.445 -194.995 ;
        RECT 218.115 -196.685 218.445 -196.355 ;
        RECT 218.115 -198.045 218.445 -197.715 ;
        RECT 218.115 -199.405 218.445 -199.075 ;
        RECT 218.115 -200.765 218.445 -200.435 ;
        RECT 218.115 -202.125 218.445 -201.795 ;
        RECT 218.115 -203.485 218.445 -203.155 ;
        RECT 218.115 -204.845 218.445 -204.515 ;
        RECT 218.115 -206.205 218.445 -205.875 ;
        RECT 218.115 -207.565 218.445 -207.235 ;
        RECT 218.115 -208.925 218.445 -208.595 ;
        RECT 218.115 -210.285 218.445 -209.955 ;
        RECT 218.115 -211.645 218.445 -211.315 ;
        RECT 218.115 -213.005 218.445 -212.675 ;
        RECT 218.115 -214.365 218.445 -214.035 ;
        RECT 218.115 -215.725 218.445 -215.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 244.04 184.445 245.17 ;
        RECT 184.115 242.595 184.445 242.925 ;
        RECT 184.115 241.235 184.445 241.565 ;
        RECT 184.115 239.875 184.445 240.205 ;
        RECT 184.115 238.515 184.445 238.845 ;
        RECT 184.115 237.155 184.445 237.485 ;
        RECT 184.12 237.155 184.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -0.845 184.445 -0.515 ;
        RECT 184.115 -2.205 184.445 -1.875 ;
        RECT 184.115 -3.565 184.445 -3.235 ;
        RECT 184.12 -3.565 184.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -123.245 184.445 -122.915 ;
        RECT 184.115 -124.605 184.445 -124.275 ;
        RECT 184.115 -125.965 184.445 -125.635 ;
        RECT 184.115 -127.325 184.445 -126.995 ;
        RECT 184.115 -128.685 184.445 -128.355 ;
        RECT 184.115 -130.045 184.445 -129.715 ;
        RECT 184.115 -131.405 184.445 -131.075 ;
        RECT 184.115 -132.765 184.445 -132.435 ;
        RECT 184.115 -134.125 184.445 -133.795 ;
        RECT 184.115 -135.485 184.445 -135.155 ;
        RECT 184.115 -136.845 184.445 -136.515 ;
        RECT 184.115 -138.205 184.445 -137.875 ;
        RECT 184.115 -139.565 184.445 -139.235 ;
        RECT 184.115 -140.925 184.445 -140.595 ;
        RECT 184.115 -142.285 184.445 -141.955 ;
        RECT 184.115 -143.645 184.445 -143.315 ;
        RECT 184.115 -145.005 184.445 -144.675 ;
        RECT 184.115 -146.365 184.445 -146.035 ;
        RECT 184.115 -147.725 184.445 -147.395 ;
        RECT 184.115 -149.085 184.445 -148.755 ;
        RECT 184.115 -150.445 184.445 -150.115 ;
        RECT 184.115 -151.805 184.445 -151.475 ;
        RECT 184.115 -153.165 184.445 -152.835 ;
        RECT 184.115 -154.525 184.445 -154.195 ;
        RECT 184.115 -155.885 184.445 -155.555 ;
        RECT 184.115 -157.245 184.445 -156.915 ;
        RECT 184.115 -158.605 184.445 -158.275 ;
        RECT 184.115 -159.965 184.445 -159.635 ;
        RECT 184.115 -161.325 184.445 -160.995 ;
        RECT 184.115 -162.685 184.445 -162.355 ;
        RECT 184.115 -164.045 184.445 -163.715 ;
        RECT 184.115 -165.405 184.445 -165.075 ;
        RECT 184.115 -166.765 184.445 -166.435 ;
        RECT 184.115 -168.125 184.445 -167.795 ;
        RECT 184.115 -169.485 184.445 -169.155 ;
        RECT 184.115 -170.845 184.445 -170.515 ;
        RECT 184.115 -172.205 184.445 -171.875 ;
        RECT 184.115 -173.565 184.445 -173.235 ;
        RECT 184.115 -174.925 184.445 -174.595 ;
        RECT 184.115 -176.285 184.445 -175.955 ;
        RECT 184.115 -177.645 184.445 -177.315 ;
        RECT 184.115 -179.005 184.445 -178.675 ;
        RECT 184.115 -180.365 184.445 -180.035 ;
        RECT 184.115 -181.725 184.445 -181.395 ;
        RECT 184.115 -183.085 184.445 -182.755 ;
        RECT 184.115 -184.445 184.445 -184.115 ;
        RECT 184.115 -185.805 184.445 -185.475 ;
        RECT 184.115 -187.165 184.445 -186.835 ;
        RECT 184.115 -188.525 184.445 -188.195 ;
        RECT 184.115 -189.885 184.445 -189.555 ;
        RECT 184.115 -191.245 184.445 -190.915 ;
        RECT 184.115 -192.605 184.445 -192.275 ;
        RECT 184.115 -193.965 184.445 -193.635 ;
        RECT 184.115 -195.325 184.445 -194.995 ;
        RECT 184.115 -196.685 184.445 -196.355 ;
        RECT 184.115 -198.045 184.445 -197.715 ;
        RECT 184.115 -199.405 184.445 -199.075 ;
        RECT 184.115 -200.765 184.445 -200.435 ;
        RECT 184.115 -202.125 184.445 -201.795 ;
        RECT 184.115 -203.485 184.445 -203.155 ;
        RECT 184.115 -204.845 184.445 -204.515 ;
        RECT 184.115 -206.205 184.445 -205.875 ;
        RECT 184.115 -207.565 184.445 -207.235 ;
        RECT 184.115 -208.925 184.445 -208.595 ;
        RECT 184.115 -210.285 184.445 -209.955 ;
        RECT 184.115 -211.645 184.445 -211.315 ;
        RECT 184.115 -213.005 184.445 -212.675 ;
        RECT 184.115 -214.365 184.445 -214.035 ;
        RECT 184.115 -215.725 184.445 -215.395 ;
        RECT 184.115 -217.085 184.445 -216.755 ;
        RECT 184.115 -218.445 184.445 -218.115 ;
        RECT 184.115 -219.805 184.445 -219.475 ;
        RECT 184.115 -221.165 184.445 -220.835 ;
        RECT 184.115 -222.525 184.445 -222.195 ;
        RECT 184.115 -223.885 184.445 -223.555 ;
        RECT 184.115 -225.245 184.445 -224.915 ;
        RECT 184.115 -226.605 184.445 -226.275 ;
        RECT 184.115 -227.965 184.445 -227.635 ;
        RECT 184.115 -229.325 184.445 -228.995 ;
        RECT 184.115 -230.685 184.445 -230.355 ;
        RECT 184.115 -232.045 184.445 -231.715 ;
        RECT 184.115 -233.405 184.445 -233.075 ;
        RECT 184.115 -234.765 184.445 -234.435 ;
        RECT 184.115 -236.125 184.445 -235.795 ;
        RECT 184.115 -237.485 184.445 -237.155 ;
        RECT 184.115 -238.845 184.445 -238.515 ;
        RECT 184.115 -241.09 184.445 -239.96 ;
        RECT 184.12 -241.205 184.44 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 244.04 185.805 245.17 ;
        RECT 185.475 242.595 185.805 242.925 ;
        RECT 185.475 241.235 185.805 241.565 ;
        RECT 185.475 239.875 185.805 240.205 ;
        RECT 185.475 238.515 185.805 238.845 ;
        RECT 185.475 237.155 185.805 237.485 ;
        RECT 185.48 237.155 185.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 -0.845 185.805 -0.515 ;
        RECT 185.475 -2.205 185.805 -1.875 ;
        RECT 185.475 -3.565 185.805 -3.235 ;
        RECT 185.48 -3.565 185.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 -123.245 185.805 -122.915 ;
        RECT 185.475 -124.605 185.805 -124.275 ;
        RECT 185.475 -125.965 185.805 -125.635 ;
        RECT 185.475 -127.325 185.805 -126.995 ;
        RECT 185.475 -128.685 185.805 -128.355 ;
        RECT 185.475 -130.045 185.805 -129.715 ;
        RECT 185.475 -131.405 185.805 -131.075 ;
        RECT 185.475 -132.765 185.805 -132.435 ;
        RECT 185.475 -134.125 185.805 -133.795 ;
        RECT 185.475 -135.485 185.805 -135.155 ;
        RECT 185.475 -136.845 185.805 -136.515 ;
        RECT 185.475 -138.205 185.805 -137.875 ;
        RECT 185.475 -139.565 185.805 -139.235 ;
        RECT 185.475 -140.925 185.805 -140.595 ;
        RECT 185.475 -142.285 185.805 -141.955 ;
        RECT 185.475 -143.645 185.805 -143.315 ;
        RECT 185.475 -145.005 185.805 -144.675 ;
        RECT 185.475 -146.365 185.805 -146.035 ;
        RECT 185.475 -147.725 185.805 -147.395 ;
        RECT 185.475 -149.085 185.805 -148.755 ;
        RECT 185.475 -150.445 185.805 -150.115 ;
        RECT 185.475 -151.805 185.805 -151.475 ;
        RECT 185.475 -153.165 185.805 -152.835 ;
        RECT 185.475 -154.525 185.805 -154.195 ;
        RECT 185.475 -155.885 185.805 -155.555 ;
        RECT 185.475 -157.245 185.805 -156.915 ;
        RECT 185.475 -158.605 185.805 -158.275 ;
        RECT 185.475 -159.965 185.805 -159.635 ;
        RECT 185.475 -161.325 185.805 -160.995 ;
        RECT 185.475 -162.685 185.805 -162.355 ;
        RECT 185.475 -164.045 185.805 -163.715 ;
        RECT 185.475 -165.405 185.805 -165.075 ;
        RECT 185.475 -166.765 185.805 -166.435 ;
        RECT 185.475 -168.125 185.805 -167.795 ;
        RECT 185.475 -169.485 185.805 -169.155 ;
        RECT 185.475 -170.845 185.805 -170.515 ;
        RECT 185.475 -172.205 185.805 -171.875 ;
        RECT 185.475 -173.565 185.805 -173.235 ;
        RECT 185.475 -174.925 185.805 -174.595 ;
        RECT 185.475 -176.285 185.805 -175.955 ;
        RECT 185.475 -177.645 185.805 -177.315 ;
        RECT 185.475 -179.005 185.805 -178.675 ;
        RECT 185.475 -180.365 185.805 -180.035 ;
        RECT 185.475 -181.725 185.805 -181.395 ;
        RECT 185.475 -183.085 185.805 -182.755 ;
        RECT 185.475 -184.445 185.805 -184.115 ;
        RECT 185.475 -185.805 185.805 -185.475 ;
        RECT 185.475 -187.165 185.805 -186.835 ;
        RECT 185.475 -188.525 185.805 -188.195 ;
        RECT 185.475 -189.885 185.805 -189.555 ;
        RECT 185.475 -191.245 185.805 -190.915 ;
        RECT 185.475 -192.605 185.805 -192.275 ;
        RECT 185.475 -193.965 185.805 -193.635 ;
        RECT 185.475 -195.325 185.805 -194.995 ;
        RECT 185.475 -196.685 185.805 -196.355 ;
        RECT 185.475 -198.045 185.805 -197.715 ;
        RECT 185.475 -199.405 185.805 -199.075 ;
        RECT 185.475 -200.765 185.805 -200.435 ;
        RECT 185.475 -202.125 185.805 -201.795 ;
        RECT 185.475 -203.485 185.805 -203.155 ;
        RECT 185.475 -204.845 185.805 -204.515 ;
        RECT 185.475 -206.205 185.805 -205.875 ;
        RECT 185.475 -207.565 185.805 -207.235 ;
        RECT 185.475 -208.925 185.805 -208.595 ;
        RECT 185.475 -210.285 185.805 -209.955 ;
        RECT 185.475 -211.645 185.805 -211.315 ;
        RECT 185.475 -213.005 185.805 -212.675 ;
        RECT 185.475 -214.365 185.805 -214.035 ;
        RECT 185.475 -215.725 185.805 -215.395 ;
        RECT 185.475 -217.085 185.805 -216.755 ;
        RECT 185.475 -218.445 185.805 -218.115 ;
        RECT 185.475 -219.805 185.805 -219.475 ;
        RECT 185.475 -221.165 185.805 -220.835 ;
        RECT 185.475 -222.525 185.805 -222.195 ;
        RECT 185.475 -223.885 185.805 -223.555 ;
        RECT 185.475 -225.245 185.805 -224.915 ;
        RECT 185.475 -226.605 185.805 -226.275 ;
        RECT 185.475 -227.965 185.805 -227.635 ;
        RECT 185.475 -229.325 185.805 -228.995 ;
        RECT 185.475 -230.685 185.805 -230.355 ;
        RECT 185.475 -232.045 185.805 -231.715 ;
        RECT 185.475 -233.405 185.805 -233.075 ;
        RECT 185.475 -234.765 185.805 -234.435 ;
        RECT 185.475 -236.125 185.805 -235.795 ;
        RECT 185.475 -237.485 185.805 -237.155 ;
        RECT 185.475 -238.845 185.805 -238.515 ;
        RECT 185.475 -241.09 185.805 -239.96 ;
        RECT 185.48 -241.205 185.8 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 244.04 187.165 245.17 ;
        RECT 186.835 242.595 187.165 242.925 ;
        RECT 186.835 241.235 187.165 241.565 ;
        RECT 186.835 239.875 187.165 240.205 ;
        RECT 186.835 238.515 187.165 238.845 ;
        RECT 186.835 237.155 187.165 237.485 ;
        RECT 186.84 237.155 187.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 -0.845 187.165 -0.515 ;
        RECT 186.835 -2.205 187.165 -1.875 ;
        RECT 186.835 -3.565 187.165 -3.235 ;
        RECT 186.84 -3.565 187.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 -123.245 187.165 -122.915 ;
        RECT 186.835 -124.605 187.165 -124.275 ;
        RECT 186.835 -125.965 187.165 -125.635 ;
        RECT 186.835 -127.325 187.165 -126.995 ;
        RECT 186.835 -128.685 187.165 -128.355 ;
        RECT 186.835 -130.045 187.165 -129.715 ;
        RECT 186.835 -131.405 187.165 -131.075 ;
        RECT 186.835 -132.765 187.165 -132.435 ;
        RECT 186.835 -134.125 187.165 -133.795 ;
        RECT 186.835 -135.485 187.165 -135.155 ;
        RECT 186.835 -136.845 187.165 -136.515 ;
        RECT 186.835 -138.205 187.165 -137.875 ;
        RECT 186.835 -139.565 187.165 -139.235 ;
        RECT 186.835 -140.925 187.165 -140.595 ;
        RECT 186.835 -142.285 187.165 -141.955 ;
        RECT 186.835 -143.645 187.165 -143.315 ;
        RECT 186.835 -145.005 187.165 -144.675 ;
        RECT 186.835 -146.365 187.165 -146.035 ;
        RECT 186.835 -147.725 187.165 -147.395 ;
        RECT 186.835 -149.085 187.165 -148.755 ;
        RECT 186.835 -150.445 187.165 -150.115 ;
        RECT 186.835 -151.805 187.165 -151.475 ;
        RECT 186.835 -153.165 187.165 -152.835 ;
        RECT 186.835 -154.525 187.165 -154.195 ;
        RECT 186.835 -155.885 187.165 -155.555 ;
        RECT 186.835 -157.245 187.165 -156.915 ;
        RECT 186.835 -158.605 187.165 -158.275 ;
        RECT 186.835 -159.965 187.165 -159.635 ;
        RECT 186.835 -161.325 187.165 -160.995 ;
        RECT 186.835 -162.685 187.165 -162.355 ;
        RECT 186.835 -164.045 187.165 -163.715 ;
        RECT 186.835 -165.405 187.165 -165.075 ;
        RECT 186.835 -166.765 187.165 -166.435 ;
        RECT 186.835 -168.125 187.165 -167.795 ;
        RECT 186.835 -169.485 187.165 -169.155 ;
        RECT 186.835 -170.845 187.165 -170.515 ;
        RECT 186.835 -172.205 187.165 -171.875 ;
        RECT 186.835 -173.565 187.165 -173.235 ;
        RECT 186.835 -174.925 187.165 -174.595 ;
        RECT 186.835 -176.285 187.165 -175.955 ;
        RECT 186.835 -177.645 187.165 -177.315 ;
        RECT 186.835 -179.005 187.165 -178.675 ;
        RECT 186.835 -180.365 187.165 -180.035 ;
        RECT 186.835 -181.725 187.165 -181.395 ;
        RECT 186.835 -183.085 187.165 -182.755 ;
        RECT 186.835 -184.445 187.165 -184.115 ;
        RECT 186.835 -185.805 187.165 -185.475 ;
        RECT 186.835 -187.165 187.165 -186.835 ;
        RECT 186.835 -188.525 187.165 -188.195 ;
        RECT 186.835 -189.885 187.165 -189.555 ;
        RECT 186.835 -191.245 187.165 -190.915 ;
        RECT 186.835 -192.605 187.165 -192.275 ;
        RECT 186.835 -193.965 187.165 -193.635 ;
        RECT 186.835 -195.325 187.165 -194.995 ;
        RECT 186.835 -196.685 187.165 -196.355 ;
        RECT 186.835 -198.045 187.165 -197.715 ;
        RECT 186.835 -199.405 187.165 -199.075 ;
        RECT 186.835 -200.765 187.165 -200.435 ;
        RECT 186.835 -202.125 187.165 -201.795 ;
        RECT 186.835 -203.485 187.165 -203.155 ;
        RECT 186.835 -204.845 187.165 -204.515 ;
        RECT 186.835 -206.205 187.165 -205.875 ;
        RECT 186.835 -207.565 187.165 -207.235 ;
        RECT 186.835 -208.925 187.165 -208.595 ;
        RECT 186.835 -210.285 187.165 -209.955 ;
        RECT 186.835 -211.645 187.165 -211.315 ;
        RECT 186.835 -213.005 187.165 -212.675 ;
        RECT 186.835 -214.365 187.165 -214.035 ;
        RECT 186.835 -215.725 187.165 -215.395 ;
        RECT 186.835 -217.085 187.165 -216.755 ;
        RECT 186.835 -218.445 187.165 -218.115 ;
        RECT 186.835 -219.805 187.165 -219.475 ;
        RECT 186.835 -221.165 187.165 -220.835 ;
        RECT 186.835 -222.525 187.165 -222.195 ;
        RECT 186.835 -223.885 187.165 -223.555 ;
        RECT 186.835 -225.245 187.165 -224.915 ;
        RECT 186.835 -226.605 187.165 -226.275 ;
        RECT 186.835 -227.965 187.165 -227.635 ;
        RECT 186.835 -229.325 187.165 -228.995 ;
        RECT 186.835 -230.685 187.165 -230.355 ;
        RECT 186.835 -232.045 187.165 -231.715 ;
        RECT 186.835 -233.405 187.165 -233.075 ;
        RECT 186.835 -234.765 187.165 -234.435 ;
        RECT 186.835 -236.125 187.165 -235.795 ;
        RECT 186.835 -237.485 187.165 -237.155 ;
        RECT 186.835 -238.845 187.165 -238.515 ;
        RECT 186.835 -241.09 187.165 -239.96 ;
        RECT 186.84 -241.205 187.16 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 244.04 188.525 245.17 ;
        RECT 188.195 242.595 188.525 242.925 ;
        RECT 188.195 241.235 188.525 241.565 ;
        RECT 188.195 239.875 188.525 240.205 ;
        RECT 188.195 238.515 188.525 238.845 ;
        RECT 188.195 237.155 188.525 237.485 ;
        RECT 188.2 237.155 188.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 -127.325 188.525 -126.995 ;
        RECT 188.195 -128.685 188.525 -128.355 ;
        RECT 188.195 -130.045 188.525 -129.715 ;
        RECT 188.195 -131.405 188.525 -131.075 ;
        RECT 188.195 -132.765 188.525 -132.435 ;
        RECT 188.195 -134.125 188.525 -133.795 ;
        RECT 188.195 -135.485 188.525 -135.155 ;
        RECT 188.195 -136.845 188.525 -136.515 ;
        RECT 188.195 -138.205 188.525 -137.875 ;
        RECT 188.195 -139.565 188.525 -139.235 ;
        RECT 188.195 -140.925 188.525 -140.595 ;
        RECT 188.195 -142.285 188.525 -141.955 ;
        RECT 188.195 -143.645 188.525 -143.315 ;
        RECT 188.195 -145.005 188.525 -144.675 ;
        RECT 188.195 -146.365 188.525 -146.035 ;
        RECT 188.195 -147.725 188.525 -147.395 ;
        RECT 188.195 -149.085 188.525 -148.755 ;
        RECT 188.195 -150.445 188.525 -150.115 ;
        RECT 188.195 -151.805 188.525 -151.475 ;
        RECT 188.195 -153.165 188.525 -152.835 ;
        RECT 188.195 -154.525 188.525 -154.195 ;
        RECT 188.195 -155.885 188.525 -155.555 ;
        RECT 188.195 -157.245 188.525 -156.915 ;
        RECT 188.195 -158.605 188.525 -158.275 ;
        RECT 188.195 -159.965 188.525 -159.635 ;
        RECT 188.195 -161.325 188.525 -160.995 ;
        RECT 188.195 -162.685 188.525 -162.355 ;
        RECT 188.195 -164.045 188.525 -163.715 ;
        RECT 188.195 -165.405 188.525 -165.075 ;
        RECT 188.195 -166.765 188.525 -166.435 ;
        RECT 188.195 -168.125 188.525 -167.795 ;
        RECT 188.195 -169.485 188.525 -169.155 ;
        RECT 188.195 -170.845 188.525 -170.515 ;
        RECT 188.195 -172.205 188.525 -171.875 ;
        RECT 188.195 -173.565 188.525 -173.235 ;
        RECT 188.195 -174.925 188.525 -174.595 ;
        RECT 188.195 -176.285 188.525 -175.955 ;
        RECT 188.195 -177.645 188.525 -177.315 ;
        RECT 188.195 -179.005 188.525 -178.675 ;
        RECT 188.195 -180.365 188.525 -180.035 ;
        RECT 188.195 -181.725 188.525 -181.395 ;
        RECT 188.195 -183.085 188.525 -182.755 ;
        RECT 188.195 -184.445 188.525 -184.115 ;
        RECT 188.195 -185.805 188.525 -185.475 ;
        RECT 188.195 -187.165 188.525 -186.835 ;
        RECT 188.195 -188.525 188.525 -188.195 ;
        RECT 188.195 -189.885 188.525 -189.555 ;
        RECT 188.195 -191.245 188.525 -190.915 ;
        RECT 188.195 -192.605 188.525 -192.275 ;
        RECT 188.195 -193.965 188.525 -193.635 ;
        RECT 188.195 -195.325 188.525 -194.995 ;
        RECT 188.195 -196.685 188.525 -196.355 ;
        RECT 188.195 -198.045 188.525 -197.715 ;
        RECT 188.195 -199.405 188.525 -199.075 ;
        RECT 188.195 -200.765 188.525 -200.435 ;
        RECT 188.195 -202.125 188.525 -201.795 ;
        RECT 188.195 -203.485 188.525 -203.155 ;
        RECT 188.195 -204.845 188.525 -204.515 ;
        RECT 188.195 -206.205 188.525 -205.875 ;
        RECT 188.195 -207.565 188.525 -207.235 ;
        RECT 188.195 -208.925 188.525 -208.595 ;
        RECT 188.195 -210.285 188.525 -209.955 ;
        RECT 188.195 -211.645 188.525 -211.315 ;
        RECT 188.195 -213.005 188.525 -212.675 ;
        RECT 188.195 -214.365 188.525 -214.035 ;
        RECT 188.195 -215.725 188.525 -215.395 ;
        RECT 188.195 -217.085 188.525 -216.755 ;
        RECT 188.195 -218.445 188.525 -218.115 ;
        RECT 188.195 -219.805 188.525 -219.475 ;
        RECT 188.195 -221.165 188.525 -220.835 ;
        RECT 188.195 -222.525 188.525 -222.195 ;
        RECT 188.195 -223.885 188.525 -223.555 ;
        RECT 188.195 -225.245 188.525 -224.915 ;
        RECT 188.195 -226.605 188.525 -226.275 ;
        RECT 188.195 -227.965 188.525 -227.635 ;
        RECT 188.195 -229.325 188.525 -228.995 ;
        RECT 188.195 -230.685 188.525 -230.355 ;
        RECT 188.195 -232.045 188.525 -231.715 ;
        RECT 188.195 -233.405 188.525 -233.075 ;
        RECT 188.195 -234.765 188.525 -234.435 ;
        RECT 188.195 -236.125 188.525 -235.795 ;
        RECT 188.195 -237.485 188.525 -237.155 ;
        RECT 188.195 -238.845 188.525 -238.515 ;
        RECT 188.195 -241.09 188.525 -239.96 ;
        RECT 188.2 -241.205 188.52 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.61 -125.535 188.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 244.04 189.885 245.17 ;
        RECT 189.555 242.595 189.885 242.925 ;
        RECT 189.555 241.235 189.885 241.565 ;
        RECT 189.555 239.875 189.885 240.205 ;
        RECT 189.555 238.515 189.885 238.845 ;
        RECT 189.555 237.155 189.885 237.485 ;
        RECT 189.56 237.155 189.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 -0.845 189.885 -0.515 ;
        RECT 189.555 -2.205 189.885 -1.875 ;
        RECT 189.555 -3.565 189.885 -3.235 ;
        RECT 189.56 -3.565 189.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 244.04 191.245 245.17 ;
        RECT 190.915 242.595 191.245 242.925 ;
        RECT 190.915 241.235 191.245 241.565 ;
        RECT 190.915 239.875 191.245 240.205 ;
        RECT 190.915 238.515 191.245 238.845 ;
        RECT 190.915 237.155 191.245 237.485 ;
        RECT 190.92 237.155 191.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 -0.845 191.245 -0.515 ;
        RECT 190.915 -2.205 191.245 -1.875 ;
        RECT 190.915 -3.565 191.245 -3.235 ;
        RECT 190.92 -3.565 191.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 244.04 192.605 245.17 ;
        RECT 192.275 242.595 192.605 242.925 ;
        RECT 192.275 241.235 192.605 241.565 ;
        RECT 192.275 239.875 192.605 240.205 ;
        RECT 192.275 238.515 192.605 238.845 ;
        RECT 192.275 237.155 192.605 237.485 ;
        RECT 192.28 237.155 192.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 -0.845 192.605 -0.515 ;
        RECT 192.275 -2.205 192.605 -1.875 ;
        RECT 192.275 -3.565 192.605 -3.235 ;
        RECT 192.28 -3.565 192.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 -123.245 192.605 -122.915 ;
        RECT 192.275 -124.605 192.605 -124.275 ;
        RECT 192.275 -125.965 192.605 -125.635 ;
        RECT 192.275 -127.325 192.605 -126.995 ;
        RECT 192.275 -128.685 192.605 -128.355 ;
        RECT 192.275 -130.045 192.605 -129.715 ;
        RECT 192.275 -131.405 192.605 -131.075 ;
        RECT 192.275 -132.765 192.605 -132.435 ;
        RECT 192.275 -134.125 192.605 -133.795 ;
        RECT 192.275 -135.485 192.605 -135.155 ;
        RECT 192.275 -136.845 192.605 -136.515 ;
        RECT 192.275 -138.205 192.605 -137.875 ;
        RECT 192.275 -139.565 192.605 -139.235 ;
        RECT 192.275 -140.925 192.605 -140.595 ;
        RECT 192.275 -142.285 192.605 -141.955 ;
        RECT 192.275 -143.645 192.605 -143.315 ;
        RECT 192.275 -145.005 192.605 -144.675 ;
        RECT 192.275 -146.365 192.605 -146.035 ;
        RECT 192.275 -147.725 192.605 -147.395 ;
        RECT 192.275 -149.085 192.605 -148.755 ;
        RECT 192.275 -150.445 192.605 -150.115 ;
        RECT 192.275 -151.805 192.605 -151.475 ;
        RECT 192.275 -153.165 192.605 -152.835 ;
        RECT 192.275 -154.525 192.605 -154.195 ;
        RECT 192.275 -155.885 192.605 -155.555 ;
        RECT 192.275 -157.245 192.605 -156.915 ;
        RECT 192.275 -158.605 192.605 -158.275 ;
        RECT 192.275 -159.965 192.605 -159.635 ;
        RECT 192.275 -161.325 192.605 -160.995 ;
        RECT 192.275 -162.685 192.605 -162.355 ;
        RECT 192.275 -164.045 192.605 -163.715 ;
        RECT 192.275 -165.405 192.605 -165.075 ;
        RECT 192.275 -166.765 192.605 -166.435 ;
        RECT 192.275 -168.125 192.605 -167.795 ;
        RECT 192.275 -169.485 192.605 -169.155 ;
        RECT 192.275 -170.845 192.605 -170.515 ;
        RECT 192.275 -172.205 192.605 -171.875 ;
        RECT 192.275 -173.565 192.605 -173.235 ;
        RECT 192.275 -174.925 192.605 -174.595 ;
        RECT 192.275 -176.285 192.605 -175.955 ;
        RECT 192.275 -177.645 192.605 -177.315 ;
        RECT 192.275 -179.005 192.605 -178.675 ;
        RECT 192.275 -180.365 192.605 -180.035 ;
        RECT 192.275 -181.725 192.605 -181.395 ;
        RECT 192.275 -183.085 192.605 -182.755 ;
        RECT 192.275 -184.445 192.605 -184.115 ;
        RECT 192.275 -185.805 192.605 -185.475 ;
        RECT 192.275 -187.165 192.605 -186.835 ;
        RECT 192.275 -188.525 192.605 -188.195 ;
        RECT 192.275 -189.885 192.605 -189.555 ;
        RECT 192.275 -191.245 192.605 -190.915 ;
        RECT 192.275 -192.605 192.605 -192.275 ;
        RECT 192.275 -193.965 192.605 -193.635 ;
        RECT 192.275 -195.325 192.605 -194.995 ;
        RECT 192.275 -196.685 192.605 -196.355 ;
        RECT 192.275 -198.045 192.605 -197.715 ;
        RECT 192.275 -199.405 192.605 -199.075 ;
        RECT 192.275 -200.765 192.605 -200.435 ;
        RECT 192.275 -202.125 192.605 -201.795 ;
        RECT 192.275 -203.485 192.605 -203.155 ;
        RECT 192.275 -204.845 192.605 -204.515 ;
        RECT 192.275 -206.205 192.605 -205.875 ;
        RECT 192.275 -207.565 192.605 -207.235 ;
        RECT 192.275 -208.925 192.605 -208.595 ;
        RECT 192.275 -210.285 192.605 -209.955 ;
        RECT 192.275 -211.645 192.605 -211.315 ;
        RECT 192.275 -213.005 192.605 -212.675 ;
        RECT 192.275 -214.365 192.605 -214.035 ;
        RECT 192.275 -215.725 192.605 -215.395 ;
        RECT 192.275 -217.085 192.605 -216.755 ;
        RECT 192.275 -218.445 192.605 -218.115 ;
        RECT 192.275 -219.805 192.605 -219.475 ;
        RECT 192.275 -221.165 192.605 -220.835 ;
        RECT 192.275 -222.525 192.605 -222.195 ;
        RECT 192.275 -223.885 192.605 -223.555 ;
        RECT 192.275 -225.245 192.605 -224.915 ;
        RECT 192.275 -226.605 192.605 -226.275 ;
        RECT 192.275 -227.965 192.605 -227.635 ;
        RECT 192.275 -229.325 192.605 -228.995 ;
        RECT 192.275 -230.685 192.605 -230.355 ;
        RECT 192.275 -232.045 192.605 -231.715 ;
        RECT 192.275 -233.405 192.605 -233.075 ;
        RECT 192.275 -234.765 192.605 -234.435 ;
        RECT 192.275 -236.125 192.605 -235.795 ;
        RECT 192.275 -237.485 192.605 -237.155 ;
        RECT 192.275 -238.845 192.605 -238.515 ;
        RECT 192.275 -241.09 192.605 -239.96 ;
        RECT 192.28 -241.205 192.6 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 244.04 193.965 245.17 ;
        RECT 193.635 242.595 193.965 242.925 ;
        RECT 193.635 241.235 193.965 241.565 ;
        RECT 193.635 239.875 193.965 240.205 ;
        RECT 193.635 238.515 193.965 238.845 ;
        RECT 193.635 237.155 193.965 237.485 ;
        RECT 193.64 237.155 193.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 -0.845 193.965 -0.515 ;
        RECT 193.635 -2.205 193.965 -1.875 ;
        RECT 193.635 -3.565 193.965 -3.235 ;
        RECT 193.64 -3.565 193.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 -123.245 193.965 -122.915 ;
        RECT 193.635 -124.605 193.965 -124.275 ;
        RECT 193.635 -125.965 193.965 -125.635 ;
        RECT 193.635 -127.325 193.965 -126.995 ;
        RECT 193.635 -128.685 193.965 -128.355 ;
        RECT 193.635 -130.045 193.965 -129.715 ;
        RECT 193.635 -131.405 193.965 -131.075 ;
        RECT 193.635 -132.765 193.965 -132.435 ;
        RECT 193.635 -134.125 193.965 -133.795 ;
        RECT 193.635 -135.485 193.965 -135.155 ;
        RECT 193.635 -136.845 193.965 -136.515 ;
        RECT 193.635 -138.205 193.965 -137.875 ;
        RECT 193.635 -139.565 193.965 -139.235 ;
        RECT 193.635 -140.925 193.965 -140.595 ;
        RECT 193.635 -142.285 193.965 -141.955 ;
        RECT 193.635 -143.645 193.965 -143.315 ;
        RECT 193.635 -145.005 193.965 -144.675 ;
        RECT 193.635 -146.365 193.965 -146.035 ;
        RECT 193.635 -147.725 193.965 -147.395 ;
        RECT 193.635 -149.085 193.965 -148.755 ;
        RECT 193.635 -150.445 193.965 -150.115 ;
        RECT 193.635 -151.805 193.965 -151.475 ;
        RECT 193.635 -153.165 193.965 -152.835 ;
        RECT 193.635 -154.525 193.965 -154.195 ;
        RECT 193.635 -155.885 193.965 -155.555 ;
        RECT 193.635 -157.245 193.965 -156.915 ;
        RECT 193.635 -158.605 193.965 -158.275 ;
        RECT 193.635 -159.965 193.965 -159.635 ;
        RECT 193.635 -161.325 193.965 -160.995 ;
        RECT 193.635 -162.685 193.965 -162.355 ;
        RECT 193.635 -164.045 193.965 -163.715 ;
        RECT 193.635 -165.405 193.965 -165.075 ;
        RECT 193.635 -166.765 193.965 -166.435 ;
        RECT 193.635 -168.125 193.965 -167.795 ;
        RECT 193.635 -169.485 193.965 -169.155 ;
        RECT 193.635 -170.845 193.965 -170.515 ;
        RECT 193.635 -172.205 193.965 -171.875 ;
        RECT 193.635 -173.565 193.965 -173.235 ;
        RECT 193.635 -174.925 193.965 -174.595 ;
        RECT 193.635 -176.285 193.965 -175.955 ;
        RECT 193.635 -177.645 193.965 -177.315 ;
        RECT 193.635 -179.005 193.965 -178.675 ;
        RECT 193.635 -180.365 193.965 -180.035 ;
        RECT 193.635 -181.725 193.965 -181.395 ;
        RECT 193.635 -183.085 193.965 -182.755 ;
        RECT 193.635 -184.445 193.965 -184.115 ;
        RECT 193.635 -185.805 193.965 -185.475 ;
        RECT 193.635 -187.165 193.965 -186.835 ;
        RECT 193.635 -188.525 193.965 -188.195 ;
        RECT 193.635 -189.885 193.965 -189.555 ;
        RECT 193.635 -191.245 193.965 -190.915 ;
        RECT 193.635 -192.605 193.965 -192.275 ;
        RECT 193.635 -193.965 193.965 -193.635 ;
        RECT 193.635 -195.325 193.965 -194.995 ;
        RECT 193.635 -196.685 193.965 -196.355 ;
        RECT 193.635 -198.045 193.965 -197.715 ;
        RECT 193.635 -199.405 193.965 -199.075 ;
        RECT 193.635 -200.765 193.965 -200.435 ;
        RECT 193.635 -202.125 193.965 -201.795 ;
        RECT 193.635 -203.485 193.965 -203.155 ;
        RECT 193.635 -204.845 193.965 -204.515 ;
        RECT 193.635 -206.205 193.965 -205.875 ;
        RECT 193.635 -207.565 193.965 -207.235 ;
        RECT 193.635 -208.925 193.965 -208.595 ;
        RECT 193.635 -210.285 193.965 -209.955 ;
        RECT 193.635 -211.645 193.965 -211.315 ;
        RECT 193.635 -213.005 193.965 -212.675 ;
        RECT 193.635 -214.365 193.965 -214.035 ;
        RECT 193.635 -215.725 193.965 -215.395 ;
        RECT 193.635 -217.085 193.965 -216.755 ;
        RECT 193.635 -218.445 193.965 -218.115 ;
        RECT 193.635 -219.805 193.965 -219.475 ;
        RECT 193.635 -221.165 193.965 -220.835 ;
        RECT 193.635 -222.525 193.965 -222.195 ;
        RECT 193.635 -223.885 193.965 -223.555 ;
        RECT 193.635 -225.245 193.965 -224.915 ;
        RECT 193.635 -226.605 193.965 -226.275 ;
        RECT 193.635 -227.965 193.965 -227.635 ;
        RECT 193.635 -229.325 193.965 -228.995 ;
        RECT 193.635 -230.685 193.965 -230.355 ;
        RECT 193.635 -232.045 193.965 -231.715 ;
        RECT 193.635 -233.405 193.965 -233.075 ;
        RECT 193.635 -234.765 193.965 -234.435 ;
        RECT 193.635 -236.125 193.965 -235.795 ;
        RECT 193.635 -237.485 193.965 -237.155 ;
        RECT 193.635 -238.845 193.965 -238.515 ;
        RECT 193.635 -241.09 193.965 -239.96 ;
        RECT 193.64 -241.205 193.96 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 244.04 195.325 245.17 ;
        RECT 194.995 242.595 195.325 242.925 ;
        RECT 194.995 241.235 195.325 241.565 ;
        RECT 194.995 239.875 195.325 240.205 ;
        RECT 194.995 238.515 195.325 238.845 ;
        RECT 194.995 237.155 195.325 237.485 ;
        RECT 195 237.155 195.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 -0.845 195.325 -0.515 ;
        RECT 194.995 -2.205 195.325 -1.875 ;
        RECT 194.995 -3.565 195.325 -3.235 ;
        RECT 195 -3.565 195.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 -123.245 195.325 -122.915 ;
        RECT 194.995 -124.605 195.325 -124.275 ;
        RECT 194.995 -125.965 195.325 -125.635 ;
        RECT 194.995 -127.325 195.325 -126.995 ;
        RECT 194.995 -128.685 195.325 -128.355 ;
        RECT 194.995 -130.045 195.325 -129.715 ;
        RECT 194.995 -131.405 195.325 -131.075 ;
        RECT 194.995 -132.765 195.325 -132.435 ;
        RECT 194.995 -134.125 195.325 -133.795 ;
        RECT 194.995 -135.485 195.325 -135.155 ;
        RECT 194.995 -136.845 195.325 -136.515 ;
        RECT 194.995 -138.205 195.325 -137.875 ;
        RECT 194.995 -139.565 195.325 -139.235 ;
        RECT 194.995 -140.925 195.325 -140.595 ;
        RECT 194.995 -142.285 195.325 -141.955 ;
        RECT 194.995 -143.645 195.325 -143.315 ;
        RECT 194.995 -145.005 195.325 -144.675 ;
        RECT 194.995 -146.365 195.325 -146.035 ;
        RECT 194.995 -147.725 195.325 -147.395 ;
        RECT 194.995 -149.085 195.325 -148.755 ;
        RECT 194.995 -150.445 195.325 -150.115 ;
        RECT 194.995 -151.805 195.325 -151.475 ;
        RECT 194.995 -153.165 195.325 -152.835 ;
        RECT 194.995 -154.525 195.325 -154.195 ;
        RECT 194.995 -155.885 195.325 -155.555 ;
        RECT 194.995 -157.245 195.325 -156.915 ;
        RECT 194.995 -158.605 195.325 -158.275 ;
        RECT 194.995 -159.965 195.325 -159.635 ;
        RECT 194.995 -161.325 195.325 -160.995 ;
        RECT 194.995 -162.685 195.325 -162.355 ;
        RECT 194.995 -164.045 195.325 -163.715 ;
        RECT 194.995 -165.405 195.325 -165.075 ;
        RECT 194.995 -166.765 195.325 -166.435 ;
        RECT 194.995 -168.125 195.325 -167.795 ;
        RECT 194.995 -169.485 195.325 -169.155 ;
        RECT 194.995 -170.845 195.325 -170.515 ;
        RECT 194.995 -172.205 195.325 -171.875 ;
        RECT 194.995 -173.565 195.325 -173.235 ;
        RECT 194.995 -174.925 195.325 -174.595 ;
        RECT 194.995 -176.285 195.325 -175.955 ;
        RECT 194.995 -177.645 195.325 -177.315 ;
        RECT 194.995 -179.005 195.325 -178.675 ;
        RECT 194.995 -180.365 195.325 -180.035 ;
        RECT 194.995 -181.725 195.325 -181.395 ;
        RECT 194.995 -183.085 195.325 -182.755 ;
        RECT 194.995 -184.445 195.325 -184.115 ;
        RECT 194.995 -185.805 195.325 -185.475 ;
        RECT 194.995 -187.165 195.325 -186.835 ;
        RECT 194.995 -188.525 195.325 -188.195 ;
        RECT 194.995 -189.885 195.325 -189.555 ;
        RECT 194.995 -191.245 195.325 -190.915 ;
        RECT 194.995 -192.605 195.325 -192.275 ;
        RECT 194.995 -193.965 195.325 -193.635 ;
        RECT 194.995 -195.325 195.325 -194.995 ;
        RECT 194.995 -196.685 195.325 -196.355 ;
        RECT 194.995 -198.045 195.325 -197.715 ;
        RECT 194.995 -199.405 195.325 -199.075 ;
        RECT 194.995 -200.765 195.325 -200.435 ;
        RECT 194.995 -202.125 195.325 -201.795 ;
        RECT 194.995 -203.485 195.325 -203.155 ;
        RECT 194.995 -204.845 195.325 -204.515 ;
        RECT 194.995 -206.205 195.325 -205.875 ;
        RECT 194.995 -207.565 195.325 -207.235 ;
        RECT 194.995 -208.925 195.325 -208.595 ;
        RECT 194.995 -210.285 195.325 -209.955 ;
        RECT 194.995 -211.645 195.325 -211.315 ;
        RECT 194.995 -213.005 195.325 -212.675 ;
        RECT 194.995 -214.365 195.325 -214.035 ;
        RECT 194.995 -215.725 195.325 -215.395 ;
        RECT 194.995 -217.085 195.325 -216.755 ;
        RECT 194.995 -218.445 195.325 -218.115 ;
        RECT 194.995 -219.805 195.325 -219.475 ;
        RECT 194.995 -221.165 195.325 -220.835 ;
        RECT 194.995 -222.525 195.325 -222.195 ;
        RECT 194.995 -223.885 195.325 -223.555 ;
        RECT 194.995 -225.245 195.325 -224.915 ;
        RECT 194.995 -226.605 195.325 -226.275 ;
        RECT 194.995 -227.965 195.325 -227.635 ;
        RECT 194.995 -229.325 195.325 -228.995 ;
        RECT 194.995 -230.685 195.325 -230.355 ;
        RECT 194.995 -232.045 195.325 -231.715 ;
        RECT 194.995 -233.405 195.325 -233.075 ;
        RECT 194.995 -234.765 195.325 -234.435 ;
        RECT 194.995 -236.125 195.325 -235.795 ;
        RECT 194.995 -237.485 195.325 -237.155 ;
        RECT 194.995 -238.845 195.325 -238.515 ;
        RECT 194.995 -241.09 195.325 -239.96 ;
        RECT 195 -241.205 195.32 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 244.04 196.685 245.17 ;
        RECT 196.355 242.595 196.685 242.925 ;
        RECT 196.355 241.235 196.685 241.565 ;
        RECT 196.355 239.875 196.685 240.205 ;
        RECT 196.355 238.515 196.685 238.845 ;
        RECT 196.355 237.155 196.685 237.485 ;
        RECT 196.36 237.155 196.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -0.845 196.685 -0.515 ;
        RECT 196.355 -2.205 196.685 -1.875 ;
        RECT 196.355 -3.565 196.685 -3.235 ;
        RECT 196.36 -3.565 196.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -123.245 196.685 -122.915 ;
        RECT 196.355 -124.605 196.685 -124.275 ;
        RECT 196.355 -125.965 196.685 -125.635 ;
        RECT 196.355 -127.325 196.685 -126.995 ;
        RECT 196.355 -128.685 196.685 -128.355 ;
        RECT 196.355 -130.045 196.685 -129.715 ;
        RECT 196.355 -131.405 196.685 -131.075 ;
        RECT 196.355 -132.765 196.685 -132.435 ;
        RECT 196.355 -134.125 196.685 -133.795 ;
        RECT 196.355 -135.485 196.685 -135.155 ;
        RECT 196.355 -136.845 196.685 -136.515 ;
        RECT 196.355 -138.205 196.685 -137.875 ;
        RECT 196.355 -139.565 196.685 -139.235 ;
        RECT 196.355 -140.925 196.685 -140.595 ;
        RECT 196.355 -142.285 196.685 -141.955 ;
        RECT 196.355 -143.645 196.685 -143.315 ;
        RECT 196.355 -145.005 196.685 -144.675 ;
        RECT 196.355 -146.365 196.685 -146.035 ;
        RECT 196.355 -147.725 196.685 -147.395 ;
        RECT 196.355 -149.085 196.685 -148.755 ;
        RECT 196.355 -150.445 196.685 -150.115 ;
        RECT 196.355 -151.805 196.685 -151.475 ;
        RECT 196.355 -153.165 196.685 -152.835 ;
        RECT 196.355 -154.525 196.685 -154.195 ;
        RECT 196.355 -155.885 196.685 -155.555 ;
        RECT 196.355 -157.245 196.685 -156.915 ;
        RECT 196.355 -158.605 196.685 -158.275 ;
        RECT 196.355 -159.965 196.685 -159.635 ;
        RECT 196.355 -161.325 196.685 -160.995 ;
        RECT 196.355 -162.685 196.685 -162.355 ;
        RECT 196.355 -164.045 196.685 -163.715 ;
        RECT 196.355 -165.405 196.685 -165.075 ;
        RECT 196.355 -166.765 196.685 -166.435 ;
        RECT 196.355 -168.125 196.685 -167.795 ;
        RECT 196.355 -169.485 196.685 -169.155 ;
        RECT 196.355 -170.845 196.685 -170.515 ;
        RECT 196.355 -172.205 196.685 -171.875 ;
        RECT 196.355 -173.565 196.685 -173.235 ;
        RECT 196.355 -174.925 196.685 -174.595 ;
        RECT 196.355 -176.285 196.685 -175.955 ;
        RECT 196.355 -177.645 196.685 -177.315 ;
        RECT 196.355 -179.005 196.685 -178.675 ;
        RECT 196.355 -180.365 196.685 -180.035 ;
        RECT 196.355 -181.725 196.685 -181.395 ;
        RECT 196.355 -183.085 196.685 -182.755 ;
        RECT 196.355 -184.445 196.685 -184.115 ;
        RECT 196.355 -185.805 196.685 -185.475 ;
        RECT 196.355 -187.165 196.685 -186.835 ;
        RECT 196.355 -188.525 196.685 -188.195 ;
        RECT 196.355 -189.885 196.685 -189.555 ;
        RECT 196.355 -191.245 196.685 -190.915 ;
        RECT 196.355 -192.605 196.685 -192.275 ;
        RECT 196.355 -193.965 196.685 -193.635 ;
        RECT 196.355 -195.325 196.685 -194.995 ;
        RECT 196.355 -196.685 196.685 -196.355 ;
        RECT 196.355 -198.045 196.685 -197.715 ;
        RECT 196.355 -199.405 196.685 -199.075 ;
        RECT 196.355 -200.765 196.685 -200.435 ;
        RECT 196.355 -202.125 196.685 -201.795 ;
        RECT 196.355 -203.485 196.685 -203.155 ;
        RECT 196.355 -204.845 196.685 -204.515 ;
        RECT 196.355 -206.205 196.685 -205.875 ;
        RECT 196.355 -207.565 196.685 -207.235 ;
        RECT 196.355 -208.925 196.685 -208.595 ;
        RECT 196.355 -210.285 196.685 -209.955 ;
        RECT 196.355 -211.645 196.685 -211.315 ;
        RECT 196.355 -213.005 196.685 -212.675 ;
        RECT 196.355 -214.365 196.685 -214.035 ;
        RECT 196.355 -215.725 196.685 -215.395 ;
        RECT 196.355 -217.085 196.685 -216.755 ;
        RECT 196.355 -218.445 196.685 -218.115 ;
        RECT 196.355 -219.805 196.685 -219.475 ;
        RECT 196.355 -221.165 196.685 -220.835 ;
        RECT 196.355 -222.525 196.685 -222.195 ;
        RECT 196.355 -223.885 196.685 -223.555 ;
        RECT 196.355 -225.245 196.685 -224.915 ;
        RECT 196.355 -226.605 196.685 -226.275 ;
        RECT 196.355 -227.965 196.685 -227.635 ;
        RECT 196.355 -229.325 196.685 -228.995 ;
        RECT 196.355 -230.685 196.685 -230.355 ;
        RECT 196.355 -232.045 196.685 -231.715 ;
        RECT 196.355 -233.405 196.685 -233.075 ;
        RECT 196.355 -234.765 196.685 -234.435 ;
        RECT 196.355 -236.125 196.685 -235.795 ;
        RECT 196.355 -237.485 196.685 -237.155 ;
        RECT 196.355 -238.845 196.685 -238.515 ;
        RECT 196.355 -241.09 196.685 -239.96 ;
        RECT 196.36 -241.205 196.68 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 244.04 198.045 245.17 ;
        RECT 197.715 242.595 198.045 242.925 ;
        RECT 197.715 241.235 198.045 241.565 ;
        RECT 197.715 239.875 198.045 240.205 ;
        RECT 197.715 238.515 198.045 238.845 ;
        RECT 197.715 237.155 198.045 237.485 ;
        RECT 197.72 237.155 198.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 -0.845 198.045 -0.515 ;
        RECT 197.715 -2.205 198.045 -1.875 ;
        RECT 197.715 -3.565 198.045 -3.235 ;
        RECT 197.72 -3.565 198.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 -123.245 198.045 -122.915 ;
        RECT 197.715 -124.605 198.045 -124.275 ;
        RECT 197.715 -125.965 198.045 -125.635 ;
        RECT 197.715 -127.325 198.045 -126.995 ;
        RECT 197.715 -128.685 198.045 -128.355 ;
        RECT 197.715 -130.045 198.045 -129.715 ;
        RECT 197.715 -131.405 198.045 -131.075 ;
        RECT 197.715 -132.765 198.045 -132.435 ;
        RECT 197.715 -134.125 198.045 -133.795 ;
        RECT 197.715 -135.485 198.045 -135.155 ;
        RECT 197.715 -136.845 198.045 -136.515 ;
        RECT 197.715 -138.205 198.045 -137.875 ;
        RECT 197.715 -139.565 198.045 -139.235 ;
        RECT 197.715 -140.925 198.045 -140.595 ;
        RECT 197.715 -142.285 198.045 -141.955 ;
        RECT 197.715 -143.645 198.045 -143.315 ;
        RECT 197.715 -145.005 198.045 -144.675 ;
        RECT 197.715 -146.365 198.045 -146.035 ;
        RECT 197.715 -147.725 198.045 -147.395 ;
        RECT 197.715 -149.085 198.045 -148.755 ;
        RECT 197.715 -150.445 198.045 -150.115 ;
        RECT 197.715 -151.805 198.045 -151.475 ;
        RECT 197.715 -153.165 198.045 -152.835 ;
        RECT 197.715 -154.525 198.045 -154.195 ;
        RECT 197.715 -155.885 198.045 -155.555 ;
        RECT 197.715 -157.245 198.045 -156.915 ;
        RECT 197.715 -158.605 198.045 -158.275 ;
        RECT 197.715 -159.965 198.045 -159.635 ;
        RECT 197.715 -161.325 198.045 -160.995 ;
        RECT 197.715 -162.685 198.045 -162.355 ;
        RECT 197.715 -164.045 198.045 -163.715 ;
        RECT 197.715 -165.405 198.045 -165.075 ;
        RECT 197.715 -166.765 198.045 -166.435 ;
        RECT 197.715 -168.125 198.045 -167.795 ;
        RECT 197.715 -169.485 198.045 -169.155 ;
        RECT 197.715 -170.845 198.045 -170.515 ;
        RECT 197.715 -172.205 198.045 -171.875 ;
        RECT 197.715 -173.565 198.045 -173.235 ;
        RECT 197.715 -174.925 198.045 -174.595 ;
        RECT 197.715 -176.285 198.045 -175.955 ;
        RECT 197.715 -177.645 198.045 -177.315 ;
        RECT 197.715 -179.005 198.045 -178.675 ;
        RECT 197.715 -180.365 198.045 -180.035 ;
        RECT 197.715 -181.725 198.045 -181.395 ;
        RECT 197.715 -183.085 198.045 -182.755 ;
        RECT 197.715 -184.445 198.045 -184.115 ;
        RECT 197.715 -185.805 198.045 -185.475 ;
        RECT 197.715 -187.165 198.045 -186.835 ;
        RECT 197.715 -188.525 198.045 -188.195 ;
        RECT 197.715 -189.885 198.045 -189.555 ;
        RECT 197.715 -191.245 198.045 -190.915 ;
        RECT 197.715 -192.605 198.045 -192.275 ;
        RECT 197.715 -193.965 198.045 -193.635 ;
        RECT 197.715 -195.325 198.045 -194.995 ;
        RECT 197.715 -196.685 198.045 -196.355 ;
        RECT 197.715 -198.045 198.045 -197.715 ;
        RECT 197.715 -199.405 198.045 -199.075 ;
        RECT 197.715 -200.765 198.045 -200.435 ;
        RECT 197.715 -202.125 198.045 -201.795 ;
        RECT 197.715 -203.485 198.045 -203.155 ;
        RECT 197.715 -204.845 198.045 -204.515 ;
        RECT 197.715 -206.205 198.045 -205.875 ;
        RECT 197.715 -207.565 198.045 -207.235 ;
        RECT 197.715 -208.925 198.045 -208.595 ;
        RECT 197.715 -210.285 198.045 -209.955 ;
        RECT 197.715 -211.645 198.045 -211.315 ;
        RECT 197.715 -213.005 198.045 -212.675 ;
        RECT 197.715 -214.365 198.045 -214.035 ;
        RECT 197.715 -215.725 198.045 -215.395 ;
        RECT 197.715 -217.085 198.045 -216.755 ;
        RECT 197.715 -218.445 198.045 -218.115 ;
        RECT 197.715 -219.805 198.045 -219.475 ;
        RECT 197.715 -221.165 198.045 -220.835 ;
        RECT 197.715 -222.525 198.045 -222.195 ;
        RECT 197.715 -223.885 198.045 -223.555 ;
        RECT 197.715 -225.245 198.045 -224.915 ;
        RECT 197.715 -226.605 198.045 -226.275 ;
        RECT 197.715 -227.965 198.045 -227.635 ;
        RECT 197.715 -229.325 198.045 -228.995 ;
        RECT 197.715 -230.685 198.045 -230.355 ;
        RECT 197.715 -232.045 198.045 -231.715 ;
        RECT 197.715 -233.405 198.045 -233.075 ;
        RECT 197.715 -234.765 198.045 -234.435 ;
        RECT 197.715 -236.125 198.045 -235.795 ;
        RECT 197.715 -237.485 198.045 -237.155 ;
        RECT 197.715 -238.845 198.045 -238.515 ;
        RECT 197.715 -241.09 198.045 -239.96 ;
        RECT 197.72 -241.205 198.04 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 244.04 199.405 245.17 ;
        RECT 199.075 242.595 199.405 242.925 ;
        RECT 199.075 241.235 199.405 241.565 ;
        RECT 199.075 239.875 199.405 240.205 ;
        RECT 199.075 238.515 199.405 238.845 ;
        RECT 199.075 237.155 199.405 237.485 ;
        RECT 199.08 237.155 199.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 -181.725 199.405 -181.395 ;
        RECT 199.075 -183.085 199.405 -182.755 ;
        RECT 199.075 -184.445 199.405 -184.115 ;
        RECT 199.075 -185.805 199.405 -185.475 ;
        RECT 199.075 -187.165 199.405 -186.835 ;
        RECT 199.075 -188.525 199.405 -188.195 ;
        RECT 199.075 -189.885 199.405 -189.555 ;
        RECT 199.075 -191.245 199.405 -190.915 ;
        RECT 199.075 -192.605 199.405 -192.275 ;
        RECT 199.075 -193.965 199.405 -193.635 ;
        RECT 199.075 -195.325 199.405 -194.995 ;
        RECT 199.075 -196.685 199.405 -196.355 ;
        RECT 199.075 -198.045 199.405 -197.715 ;
        RECT 199.075 -199.405 199.405 -199.075 ;
        RECT 199.075 -200.765 199.405 -200.435 ;
        RECT 199.075 -202.125 199.405 -201.795 ;
        RECT 199.075 -203.485 199.405 -203.155 ;
        RECT 199.075 -204.845 199.405 -204.515 ;
        RECT 199.075 -206.205 199.405 -205.875 ;
        RECT 199.075 -207.565 199.405 -207.235 ;
        RECT 199.075 -208.925 199.405 -208.595 ;
        RECT 199.075 -210.285 199.405 -209.955 ;
        RECT 199.075 -211.645 199.405 -211.315 ;
        RECT 199.075 -213.005 199.405 -212.675 ;
        RECT 199.075 -214.365 199.405 -214.035 ;
        RECT 199.075 -215.725 199.405 -215.395 ;
        RECT 199.075 -217.085 199.405 -216.755 ;
        RECT 199.075 -218.445 199.405 -218.115 ;
        RECT 199.075 -219.805 199.405 -219.475 ;
        RECT 199.075 -221.165 199.405 -220.835 ;
        RECT 199.075 -222.525 199.405 -222.195 ;
        RECT 199.075 -223.885 199.405 -223.555 ;
        RECT 199.075 -225.245 199.405 -224.915 ;
        RECT 199.075 -226.605 199.405 -226.275 ;
        RECT 199.075 -227.965 199.405 -227.635 ;
        RECT 199.075 -229.325 199.405 -228.995 ;
        RECT 199.075 -230.685 199.405 -230.355 ;
        RECT 199.075 -232.045 199.405 -231.715 ;
        RECT 199.075 -233.405 199.405 -233.075 ;
        RECT 199.075 -234.765 199.405 -234.435 ;
        RECT 199.075 -236.125 199.405 -235.795 ;
        RECT 199.075 -237.485 199.405 -237.155 ;
        RECT 199.075 -238.845 199.405 -238.515 ;
        RECT 199.075 -241.09 199.405 -239.96 ;
        RECT 199.08 -241.205 199.4 -126.32 ;
        RECT 199.075 -127.325 199.405 -126.995 ;
        RECT 199.075 -128.685 199.405 -128.355 ;
        RECT 199.075 -130.045 199.405 -129.715 ;
        RECT 199.075 -131.405 199.405 -131.075 ;
        RECT 199.075 -132.765 199.405 -132.435 ;
        RECT 199.075 -134.125 199.405 -133.795 ;
        RECT 199.075 -135.485 199.405 -135.155 ;
        RECT 199.075 -136.845 199.405 -136.515 ;
        RECT 199.075 -138.205 199.405 -137.875 ;
        RECT 199.075 -139.565 199.405 -139.235 ;
        RECT 199.075 -140.925 199.405 -140.595 ;
        RECT 199.075 -142.285 199.405 -141.955 ;
        RECT 199.075 -143.645 199.405 -143.315 ;
        RECT 199.075 -145.005 199.405 -144.675 ;
        RECT 199.075 -146.365 199.405 -146.035 ;
        RECT 199.075 -147.725 199.405 -147.395 ;
        RECT 199.075 -149.085 199.405 -148.755 ;
        RECT 199.075 -150.445 199.405 -150.115 ;
        RECT 199.075 -151.805 199.405 -151.475 ;
        RECT 199.075 -153.165 199.405 -152.835 ;
        RECT 199.075 -154.525 199.405 -154.195 ;
        RECT 199.075 -155.885 199.405 -155.555 ;
        RECT 199.075 -157.245 199.405 -156.915 ;
        RECT 199.075 -158.605 199.405 -158.275 ;
        RECT 199.075 -159.965 199.405 -159.635 ;
        RECT 199.075 -161.325 199.405 -160.995 ;
        RECT 199.075 -162.685 199.405 -162.355 ;
        RECT 199.075 -164.045 199.405 -163.715 ;
        RECT 199.075 -165.405 199.405 -165.075 ;
        RECT 199.075 -166.765 199.405 -166.435 ;
        RECT 199.075 -168.125 199.405 -167.795 ;
        RECT 199.075 -169.485 199.405 -169.155 ;
        RECT 199.075 -170.845 199.405 -170.515 ;
        RECT 199.075 -172.205 199.405 -171.875 ;
        RECT 199.075 -173.565 199.405 -173.235 ;
        RECT 199.075 -174.925 199.405 -174.595 ;
        RECT 199.075 -176.285 199.405 -175.955 ;
        RECT 199.075 -177.645 199.405 -177.315 ;
        RECT 199.075 -179.005 199.405 -178.675 ;
        RECT 199.075 -180.365 199.405 -180.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 244.04 165.405 245.17 ;
        RECT 165.075 242.595 165.405 242.925 ;
        RECT 165.075 241.235 165.405 241.565 ;
        RECT 165.075 239.875 165.405 240.205 ;
        RECT 165.075 238.515 165.405 238.845 ;
        RECT 165.075 237.155 165.405 237.485 ;
        RECT 165.08 237.155 165.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -0.845 165.405 -0.515 ;
        RECT 165.075 -2.205 165.405 -1.875 ;
        RECT 165.075 -3.565 165.405 -3.235 ;
        RECT 165.08 -3.565 165.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -123.245 165.405 -122.915 ;
        RECT 165.075 -124.605 165.405 -124.275 ;
        RECT 165.075 -125.965 165.405 -125.635 ;
        RECT 165.075 -127.325 165.405 -126.995 ;
        RECT 165.075 -128.685 165.405 -128.355 ;
        RECT 165.075 -130.045 165.405 -129.715 ;
        RECT 165.075 -131.405 165.405 -131.075 ;
        RECT 165.075 -132.765 165.405 -132.435 ;
        RECT 165.075 -134.125 165.405 -133.795 ;
        RECT 165.075 -135.485 165.405 -135.155 ;
        RECT 165.075 -136.845 165.405 -136.515 ;
        RECT 165.075 -138.205 165.405 -137.875 ;
        RECT 165.075 -139.565 165.405 -139.235 ;
        RECT 165.075 -140.925 165.405 -140.595 ;
        RECT 165.075 -142.285 165.405 -141.955 ;
        RECT 165.075 -143.645 165.405 -143.315 ;
        RECT 165.075 -145.005 165.405 -144.675 ;
        RECT 165.075 -146.365 165.405 -146.035 ;
        RECT 165.075 -147.725 165.405 -147.395 ;
        RECT 165.075 -149.085 165.405 -148.755 ;
        RECT 165.075 -150.445 165.405 -150.115 ;
        RECT 165.075 -151.805 165.405 -151.475 ;
        RECT 165.075 -153.165 165.405 -152.835 ;
        RECT 165.075 -154.525 165.405 -154.195 ;
        RECT 165.075 -155.885 165.405 -155.555 ;
        RECT 165.075 -157.245 165.405 -156.915 ;
        RECT 165.075 -158.605 165.405 -158.275 ;
        RECT 165.075 -159.965 165.405 -159.635 ;
        RECT 165.075 -161.325 165.405 -160.995 ;
        RECT 165.075 -162.685 165.405 -162.355 ;
        RECT 165.075 -164.045 165.405 -163.715 ;
        RECT 165.075 -165.405 165.405 -165.075 ;
        RECT 165.075 -166.765 165.405 -166.435 ;
        RECT 165.075 -168.125 165.405 -167.795 ;
        RECT 165.075 -169.485 165.405 -169.155 ;
        RECT 165.075 -170.845 165.405 -170.515 ;
        RECT 165.075 -172.205 165.405 -171.875 ;
        RECT 165.075 -173.565 165.405 -173.235 ;
        RECT 165.075 -174.925 165.405 -174.595 ;
        RECT 165.075 -176.285 165.405 -175.955 ;
        RECT 165.075 -177.645 165.405 -177.315 ;
        RECT 165.075 -179.005 165.405 -178.675 ;
        RECT 165.075 -180.365 165.405 -180.035 ;
        RECT 165.075 -181.725 165.405 -181.395 ;
        RECT 165.075 -183.085 165.405 -182.755 ;
        RECT 165.075 -184.445 165.405 -184.115 ;
        RECT 165.075 -185.805 165.405 -185.475 ;
        RECT 165.075 -187.165 165.405 -186.835 ;
        RECT 165.075 -188.525 165.405 -188.195 ;
        RECT 165.075 -189.885 165.405 -189.555 ;
        RECT 165.075 -191.245 165.405 -190.915 ;
        RECT 165.075 -192.605 165.405 -192.275 ;
        RECT 165.075 -193.965 165.405 -193.635 ;
        RECT 165.075 -195.325 165.405 -194.995 ;
        RECT 165.075 -196.685 165.405 -196.355 ;
        RECT 165.075 -198.045 165.405 -197.715 ;
        RECT 165.075 -199.405 165.405 -199.075 ;
        RECT 165.075 -200.765 165.405 -200.435 ;
        RECT 165.075 -202.125 165.405 -201.795 ;
        RECT 165.075 -203.485 165.405 -203.155 ;
        RECT 165.075 -204.845 165.405 -204.515 ;
        RECT 165.075 -206.205 165.405 -205.875 ;
        RECT 165.075 -207.565 165.405 -207.235 ;
        RECT 165.075 -208.925 165.405 -208.595 ;
        RECT 165.075 -210.285 165.405 -209.955 ;
        RECT 165.075 -211.645 165.405 -211.315 ;
        RECT 165.075 -213.005 165.405 -212.675 ;
        RECT 165.075 -214.365 165.405 -214.035 ;
        RECT 165.075 -215.725 165.405 -215.395 ;
        RECT 165.075 -217.085 165.405 -216.755 ;
        RECT 165.075 -218.445 165.405 -218.115 ;
        RECT 165.075 -219.805 165.405 -219.475 ;
        RECT 165.075 -221.165 165.405 -220.835 ;
        RECT 165.075 -222.525 165.405 -222.195 ;
        RECT 165.075 -223.885 165.405 -223.555 ;
        RECT 165.075 -225.245 165.405 -224.915 ;
        RECT 165.075 -226.605 165.405 -226.275 ;
        RECT 165.075 -227.965 165.405 -227.635 ;
        RECT 165.075 -229.325 165.405 -228.995 ;
        RECT 165.075 -230.685 165.405 -230.355 ;
        RECT 165.075 -232.045 165.405 -231.715 ;
        RECT 165.075 -233.405 165.405 -233.075 ;
        RECT 165.075 -234.765 165.405 -234.435 ;
        RECT 165.075 -236.125 165.405 -235.795 ;
        RECT 165.075 -237.485 165.405 -237.155 ;
        RECT 165.075 -238.845 165.405 -238.515 ;
        RECT 165.075 -241.09 165.405 -239.96 ;
        RECT 165.08 -241.205 165.4 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 244.04 166.765 245.17 ;
        RECT 166.435 242.595 166.765 242.925 ;
        RECT 166.435 241.235 166.765 241.565 ;
        RECT 166.435 239.875 166.765 240.205 ;
        RECT 166.435 238.515 166.765 238.845 ;
        RECT 166.435 237.155 166.765 237.485 ;
        RECT 166.44 237.155 166.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -127.325 166.765 -126.995 ;
        RECT 166.435 -128.685 166.765 -128.355 ;
        RECT 166.435 -130.045 166.765 -129.715 ;
        RECT 166.435 -131.405 166.765 -131.075 ;
        RECT 166.435 -132.765 166.765 -132.435 ;
        RECT 166.435 -134.125 166.765 -133.795 ;
        RECT 166.435 -135.485 166.765 -135.155 ;
        RECT 166.435 -136.845 166.765 -136.515 ;
        RECT 166.435 -138.205 166.765 -137.875 ;
        RECT 166.435 -139.565 166.765 -139.235 ;
        RECT 166.435 -140.925 166.765 -140.595 ;
        RECT 166.435 -142.285 166.765 -141.955 ;
        RECT 166.435 -143.645 166.765 -143.315 ;
        RECT 166.435 -145.005 166.765 -144.675 ;
        RECT 166.435 -146.365 166.765 -146.035 ;
        RECT 166.435 -147.725 166.765 -147.395 ;
        RECT 166.435 -149.085 166.765 -148.755 ;
        RECT 166.435 -150.445 166.765 -150.115 ;
        RECT 166.435 -151.805 166.765 -151.475 ;
        RECT 166.435 -153.165 166.765 -152.835 ;
        RECT 166.435 -154.525 166.765 -154.195 ;
        RECT 166.435 -155.885 166.765 -155.555 ;
        RECT 166.435 -157.245 166.765 -156.915 ;
        RECT 166.435 -158.605 166.765 -158.275 ;
        RECT 166.435 -159.965 166.765 -159.635 ;
        RECT 166.435 -161.325 166.765 -160.995 ;
        RECT 166.435 -162.685 166.765 -162.355 ;
        RECT 166.435 -164.045 166.765 -163.715 ;
        RECT 166.435 -165.405 166.765 -165.075 ;
        RECT 166.435 -166.765 166.765 -166.435 ;
        RECT 166.435 -168.125 166.765 -167.795 ;
        RECT 166.435 -169.485 166.765 -169.155 ;
        RECT 166.435 -170.845 166.765 -170.515 ;
        RECT 166.435 -172.205 166.765 -171.875 ;
        RECT 166.435 -173.565 166.765 -173.235 ;
        RECT 166.435 -174.925 166.765 -174.595 ;
        RECT 166.435 -176.285 166.765 -175.955 ;
        RECT 166.435 -177.645 166.765 -177.315 ;
        RECT 166.435 -179.005 166.765 -178.675 ;
        RECT 166.435 -180.365 166.765 -180.035 ;
        RECT 166.435 -181.725 166.765 -181.395 ;
        RECT 166.435 -183.085 166.765 -182.755 ;
        RECT 166.435 -184.445 166.765 -184.115 ;
        RECT 166.435 -185.805 166.765 -185.475 ;
        RECT 166.435 -187.165 166.765 -186.835 ;
        RECT 166.435 -188.525 166.765 -188.195 ;
        RECT 166.435 -189.885 166.765 -189.555 ;
        RECT 166.435 -191.245 166.765 -190.915 ;
        RECT 166.435 -192.605 166.765 -192.275 ;
        RECT 166.435 -193.965 166.765 -193.635 ;
        RECT 166.435 -195.325 166.765 -194.995 ;
        RECT 166.435 -196.685 166.765 -196.355 ;
        RECT 166.435 -198.045 166.765 -197.715 ;
        RECT 166.435 -199.405 166.765 -199.075 ;
        RECT 166.435 -200.765 166.765 -200.435 ;
        RECT 166.435 -202.125 166.765 -201.795 ;
        RECT 166.435 -203.485 166.765 -203.155 ;
        RECT 166.435 -204.845 166.765 -204.515 ;
        RECT 166.435 -206.205 166.765 -205.875 ;
        RECT 166.435 -207.565 166.765 -207.235 ;
        RECT 166.435 -208.925 166.765 -208.595 ;
        RECT 166.435 -210.285 166.765 -209.955 ;
        RECT 166.435 -211.645 166.765 -211.315 ;
        RECT 166.435 -213.005 166.765 -212.675 ;
        RECT 166.435 -214.365 166.765 -214.035 ;
        RECT 166.435 -215.725 166.765 -215.395 ;
        RECT 166.435 -217.085 166.765 -216.755 ;
        RECT 166.435 -218.445 166.765 -218.115 ;
        RECT 166.435 -219.805 166.765 -219.475 ;
        RECT 166.435 -221.165 166.765 -220.835 ;
        RECT 166.435 -222.525 166.765 -222.195 ;
        RECT 166.435 -223.885 166.765 -223.555 ;
        RECT 166.435 -225.245 166.765 -224.915 ;
        RECT 166.435 -226.605 166.765 -226.275 ;
        RECT 166.435 -227.965 166.765 -227.635 ;
        RECT 166.435 -229.325 166.765 -228.995 ;
        RECT 166.435 -230.685 166.765 -230.355 ;
        RECT 166.435 -232.045 166.765 -231.715 ;
        RECT 166.435 -233.405 166.765 -233.075 ;
        RECT 166.435 -234.765 166.765 -234.435 ;
        RECT 166.435 -236.125 166.765 -235.795 ;
        RECT 166.435 -237.485 166.765 -237.155 ;
        RECT 166.435 -238.845 166.765 -238.515 ;
        RECT 166.435 -241.09 166.765 -239.96 ;
        RECT 166.44 -241.205 166.76 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.81 -125.535 167.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 244.04 168.125 245.17 ;
        RECT 167.795 242.595 168.125 242.925 ;
        RECT 167.795 241.235 168.125 241.565 ;
        RECT 167.795 239.875 168.125 240.205 ;
        RECT 167.795 238.515 168.125 238.845 ;
        RECT 167.795 237.155 168.125 237.485 ;
        RECT 167.8 237.155 168.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 -0.845 168.125 -0.515 ;
        RECT 167.795 -2.205 168.125 -1.875 ;
        RECT 167.795 -3.565 168.125 -3.235 ;
        RECT 167.8 -3.565 168.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 244.04 169.485 245.17 ;
        RECT 169.155 242.595 169.485 242.925 ;
        RECT 169.155 241.235 169.485 241.565 ;
        RECT 169.155 239.875 169.485 240.205 ;
        RECT 169.155 238.515 169.485 238.845 ;
        RECT 169.155 237.155 169.485 237.485 ;
        RECT 169.16 237.155 169.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 -0.845 169.485 -0.515 ;
        RECT 169.155 -2.205 169.485 -1.875 ;
        RECT 169.155 -3.565 169.485 -3.235 ;
        RECT 169.16 -3.565 169.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 244.04 170.845 245.17 ;
        RECT 170.515 242.595 170.845 242.925 ;
        RECT 170.515 241.235 170.845 241.565 ;
        RECT 170.515 239.875 170.845 240.205 ;
        RECT 170.515 238.515 170.845 238.845 ;
        RECT 170.515 237.155 170.845 237.485 ;
        RECT 170.52 237.155 170.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 -0.845 170.845 -0.515 ;
        RECT 170.515 -2.205 170.845 -1.875 ;
        RECT 170.515 -3.565 170.845 -3.235 ;
        RECT 170.52 -3.565 170.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 -123.245 170.845 -122.915 ;
        RECT 170.515 -124.605 170.845 -124.275 ;
        RECT 170.515 -125.965 170.845 -125.635 ;
        RECT 170.515 -127.325 170.845 -126.995 ;
        RECT 170.515 -128.685 170.845 -128.355 ;
        RECT 170.515 -130.045 170.845 -129.715 ;
        RECT 170.515 -131.405 170.845 -131.075 ;
        RECT 170.515 -132.765 170.845 -132.435 ;
        RECT 170.515 -134.125 170.845 -133.795 ;
        RECT 170.515 -135.485 170.845 -135.155 ;
        RECT 170.515 -136.845 170.845 -136.515 ;
        RECT 170.515 -138.205 170.845 -137.875 ;
        RECT 170.515 -139.565 170.845 -139.235 ;
        RECT 170.515 -140.925 170.845 -140.595 ;
        RECT 170.515 -142.285 170.845 -141.955 ;
        RECT 170.515 -143.645 170.845 -143.315 ;
        RECT 170.515 -145.005 170.845 -144.675 ;
        RECT 170.515 -146.365 170.845 -146.035 ;
        RECT 170.515 -147.725 170.845 -147.395 ;
        RECT 170.515 -149.085 170.845 -148.755 ;
        RECT 170.515 -150.445 170.845 -150.115 ;
        RECT 170.515 -151.805 170.845 -151.475 ;
        RECT 170.515 -153.165 170.845 -152.835 ;
        RECT 170.515 -154.525 170.845 -154.195 ;
        RECT 170.515 -155.885 170.845 -155.555 ;
        RECT 170.515 -157.245 170.845 -156.915 ;
        RECT 170.515 -158.605 170.845 -158.275 ;
        RECT 170.515 -159.965 170.845 -159.635 ;
        RECT 170.515 -161.325 170.845 -160.995 ;
        RECT 170.515 -162.685 170.845 -162.355 ;
        RECT 170.515 -164.045 170.845 -163.715 ;
        RECT 170.515 -165.405 170.845 -165.075 ;
        RECT 170.515 -166.765 170.845 -166.435 ;
        RECT 170.515 -168.125 170.845 -167.795 ;
        RECT 170.515 -169.485 170.845 -169.155 ;
        RECT 170.515 -170.845 170.845 -170.515 ;
        RECT 170.515 -172.205 170.845 -171.875 ;
        RECT 170.515 -173.565 170.845 -173.235 ;
        RECT 170.515 -174.925 170.845 -174.595 ;
        RECT 170.515 -176.285 170.845 -175.955 ;
        RECT 170.515 -177.645 170.845 -177.315 ;
        RECT 170.515 -179.005 170.845 -178.675 ;
        RECT 170.515 -180.365 170.845 -180.035 ;
        RECT 170.515 -181.725 170.845 -181.395 ;
        RECT 170.515 -183.085 170.845 -182.755 ;
        RECT 170.515 -184.445 170.845 -184.115 ;
        RECT 170.515 -185.805 170.845 -185.475 ;
        RECT 170.515 -187.165 170.845 -186.835 ;
        RECT 170.515 -188.525 170.845 -188.195 ;
        RECT 170.515 -189.885 170.845 -189.555 ;
        RECT 170.515 -191.245 170.845 -190.915 ;
        RECT 170.515 -192.605 170.845 -192.275 ;
        RECT 170.515 -193.965 170.845 -193.635 ;
        RECT 170.515 -195.325 170.845 -194.995 ;
        RECT 170.515 -196.685 170.845 -196.355 ;
        RECT 170.515 -198.045 170.845 -197.715 ;
        RECT 170.515 -199.405 170.845 -199.075 ;
        RECT 170.515 -200.765 170.845 -200.435 ;
        RECT 170.515 -202.125 170.845 -201.795 ;
        RECT 170.515 -203.485 170.845 -203.155 ;
        RECT 170.515 -204.845 170.845 -204.515 ;
        RECT 170.515 -206.205 170.845 -205.875 ;
        RECT 170.515 -207.565 170.845 -207.235 ;
        RECT 170.515 -208.925 170.845 -208.595 ;
        RECT 170.515 -210.285 170.845 -209.955 ;
        RECT 170.515 -211.645 170.845 -211.315 ;
        RECT 170.515 -213.005 170.845 -212.675 ;
        RECT 170.515 -214.365 170.845 -214.035 ;
        RECT 170.515 -215.725 170.845 -215.395 ;
        RECT 170.515 -217.085 170.845 -216.755 ;
        RECT 170.515 -218.445 170.845 -218.115 ;
        RECT 170.515 -219.805 170.845 -219.475 ;
        RECT 170.515 -221.165 170.845 -220.835 ;
        RECT 170.515 -222.525 170.845 -222.195 ;
        RECT 170.515 -223.885 170.845 -223.555 ;
        RECT 170.515 -225.245 170.845 -224.915 ;
        RECT 170.515 -226.605 170.845 -226.275 ;
        RECT 170.515 -227.965 170.845 -227.635 ;
        RECT 170.515 -229.325 170.845 -228.995 ;
        RECT 170.515 -230.685 170.845 -230.355 ;
        RECT 170.515 -232.045 170.845 -231.715 ;
        RECT 170.515 -233.405 170.845 -233.075 ;
        RECT 170.515 -234.765 170.845 -234.435 ;
        RECT 170.515 -236.125 170.845 -235.795 ;
        RECT 170.515 -237.485 170.845 -237.155 ;
        RECT 170.515 -238.845 170.845 -238.515 ;
        RECT 170.515 -241.09 170.845 -239.96 ;
        RECT 170.52 -241.205 170.84 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 244.04 172.205 245.17 ;
        RECT 171.875 242.595 172.205 242.925 ;
        RECT 171.875 241.235 172.205 241.565 ;
        RECT 171.875 239.875 172.205 240.205 ;
        RECT 171.875 238.515 172.205 238.845 ;
        RECT 171.875 237.155 172.205 237.485 ;
        RECT 171.88 237.155 172.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -0.845 172.205 -0.515 ;
        RECT 171.875 -2.205 172.205 -1.875 ;
        RECT 171.875 -3.565 172.205 -3.235 ;
        RECT 171.88 -3.565 172.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -123.245 172.205 -122.915 ;
        RECT 171.875 -124.605 172.205 -124.275 ;
        RECT 171.875 -125.965 172.205 -125.635 ;
        RECT 171.875 -127.325 172.205 -126.995 ;
        RECT 171.875 -128.685 172.205 -128.355 ;
        RECT 171.875 -130.045 172.205 -129.715 ;
        RECT 171.875 -131.405 172.205 -131.075 ;
        RECT 171.875 -132.765 172.205 -132.435 ;
        RECT 171.875 -134.125 172.205 -133.795 ;
        RECT 171.875 -135.485 172.205 -135.155 ;
        RECT 171.875 -136.845 172.205 -136.515 ;
        RECT 171.875 -138.205 172.205 -137.875 ;
        RECT 171.875 -139.565 172.205 -139.235 ;
        RECT 171.875 -140.925 172.205 -140.595 ;
        RECT 171.875 -142.285 172.205 -141.955 ;
        RECT 171.875 -143.645 172.205 -143.315 ;
        RECT 171.875 -145.005 172.205 -144.675 ;
        RECT 171.875 -146.365 172.205 -146.035 ;
        RECT 171.875 -147.725 172.205 -147.395 ;
        RECT 171.875 -149.085 172.205 -148.755 ;
        RECT 171.875 -150.445 172.205 -150.115 ;
        RECT 171.875 -151.805 172.205 -151.475 ;
        RECT 171.875 -153.165 172.205 -152.835 ;
        RECT 171.875 -154.525 172.205 -154.195 ;
        RECT 171.875 -155.885 172.205 -155.555 ;
        RECT 171.875 -157.245 172.205 -156.915 ;
        RECT 171.875 -158.605 172.205 -158.275 ;
        RECT 171.875 -159.965 172.205 -159.635 ;
        RECT 171.875 -161.325 172.205 -160.995 ;
        RECT 171.875 -162.685 172.205 -162.355 ;
        RECT 171.875 -164.045 172.205 -163.715 ;
        RECT 171.875 -165.405 172.205 -165.075 ;
        RECT 171.875 -166.765 172.205 -166.435 ;
        RECT 171.875 -168.125 172.205 -167.795 ;
        RECT 171.875 -169.485 172.205 -169.155 ;
        RECT 171.875 -170.845 172.205 -170.515 ;
        RECT 171.875 -172.205 172.205 -171.875 ;
        RECT 171.875 -173.565 172.205 -173.235 ;
        RECT 171.875 -174.925 172.205 -174.595 ;
        RECT 171.875 -176.285 172.205 -175.955 ;
        RECT 171.875 -177.645 172.205 -177.315 ;
        RECT 171.875 -179.005 172.205 -178.675 ;
        RECT 171.875 -180.365 172.205 -180.035 ;
        RECT 171.875 -181.725 172.205 -181.395 ;
        RECT 171.875 -183.085 172.205 -182.755 ;
        RECT 171.875 -184.445 172.205 -184.115 ;
        RECT 171.875 -185.805 172.205 -185.475 ;
        RECT 171.875 -187.165 172.205 -186.835 ;
        RECT 171.875 -188.525 172.205 -188.195 ;
        RECT 171.875 -189.885 172.205 -189.555 ;
        RECT 171.875 -191.245 172.205 -190.915 ;
        RECT 171.875 -192.605 172.205 -192.275 ;
        RECT 171.875 -193.965 172.205 -193.635 ;
        RECT 171.875 -195.325 172.205 -194.995 ;
        RECT 171.875 -196.685 172.205 -196.355 ;
        RECT 171.875 -198.045 172.205 -197.715 ;
        RECT 171.875 -199.405 172.205 -199.075 ;
        RECT 171.875 -200.765 172.205 -200.435 ;
        RECT 171.875 -202.125 172.205 -201.795 ;
        RECT 171.875 -203.485 172.205 -203.155 ;
        RECT 171.875 -204.845 172.205 -204.515 ;
        RECT 171.875 -206.205 172.205 -205.875 ;
        RECT 171.875 -207.565 172.205 -207.235 ;
        RECT 171.875 -208.925 172.205 -208.595 ;
        RECT 171.875 -210.285 172.205 -209.955 ;
        RECT 171.875 -211.645 172.205 -211.315 ;
        RECT 171.875 -213.005 172.205 -212.675 ;
        RECT 171.875 -214.365 172.205 -214.035 ;
        RECT 171.875 -215.725 172.205 -215.395 ;
        RECT 171.875 -217.085 172.205 -216.755 ;
        RECT 171.875 -218.445 172.205 -218.115 ;
        RECT 171.875 -219.805 172.205 -219.475 ;
        RECT 171.875 -221.165 172.205 -220.835 ;
        RECT 171.875 -222.525 172.205 -222.195 ;
        RECT 171.875 -223.885 172.205 -223.555 ;
        RECT 171.875 -225.245 172.205 -224.915 ;
        RECT 171.875 -226.605 172.205 -226.275 ;
        RECT 171.875 -227.965 172.205 -227.635 ;
        RECT 171.875 -229.325 172.205 -228.995 ;
        RECT 171.875 -230.685 172.205 -230.355 ;
        RECT 171.875 -232.045 172.205 -231.715 ;
        RECT 171.875 -233.405 172.205 -233.075 ;
        RECT 171.875 -234.765 172.205 -234.435 ;
        RECT 171.875 -236.125 172.205 -235.795 ;
        RECT 171.875 -237.485 172.205 -237.155 ;
        RECT 171.875 -238.845 172.205 -238.515 ;
        RECT 171.875 -241.09 172.205 -239.96 ;
        RECT 171.88 -241.205 172.2 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 244.04 173.565 245.17 ;
        RECT 173.235 242.595 173.565 242.925 ;
        RECT 173.235 241.235 173.565 241.565 ;
        RECT 173.235 239.875 173.565 240.205 ;
        RECT 173.235 238.515 173.565 238.845 ;
        RECT 173.235 237.155 173.565 237.485 ;
        RECT 173.24 237.155 173.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 -0.845 173.565 -0.515 ;
        RECT 173.235 -2.205 173.565 -1.875 ;
        RECT 173.235 -3.565 173.565 -3.235 ;
        RECT 173.24 -3.565 173.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 -123.245 173.565 -122.915 ;
        RECT 173.235 -124.605 173.565 -124.275 ;
        RECT 173.235 -125.965 173.565 -125.635 ;
        RECT 173.235 -127.325 173.565 -126.995 ;
        RECT 173.235 -128.685 173.565 -128.355 ;
        RECT 173.235 -130.045 173.565 -129.715 ;
        RECT 173.235 -131.405 173.565 -131.075 ;
        RECT 173.235 -132.765 173.565 -132.435 ;
        RECT 173.235 -134.125 173.565 -133.795 ;
        RECT 173.235 -135.485 173.565 -135.155 ;
        RECT 173.235 -136.845 173.565 -136.515 ;
        RECT 173.235 -138.205 173.565 -137.875 ;
        RECT 173.235 -139.565 173.565 -139.235 ;
        RECT 173.235 -140.925 173.565 -140.595 ;
        RECT 173.235 -142.285 173.565 -141.955 ;
        RECT 173.235 -143.645 173.565 -143.315 ;
        RECT 173.235 -145.005 173.565 -144.675 ;
        RECT 173.235 -146.365 173.565 -146.035 ;
        RECT 173.235 -147.725 173.565 -147.395 ;
        RECT 173.235 -149.085 173.565 -148.755 ;
        RECT 173.235 -150.445 173.565 -150.115 ;
        RECT 173.235 -151.805 173.565 -151.475 ;
        RECT 173.235 -153.165 173.565 -152.835 ;
        RECT 173.235 -154.525 173.565 -154.195 ;
        RECT 173.235 -155.885 173.565 -155.555 ;
        RECT 173.235 -157.245 173.565 -156.915 ;
        RECT 173.235 -158.605 173.565 -158.275 ;
        RECT 173.235 -159.965 173.565 -159.635 ;
        RECT 173.235 -161.325 173.565 -160.995 ;
        RECT 173.235 -162.685 173.565 -162.355 ;
        RECT 173.235 -164.045 173.565 -163.715 ;
        RECT 173.235 -165.405 173.565 -165.075 ;
        RECT 173.235 -166.765 173.565 -166.435 ;
        RECT 173.235 -168.125 173.565 -167.795 ;
        RECT 173.235 -169.485 173.565 -169.155 ;
        RECT 173.235 -170.845 173.565 -170.515 ;
        RECT 173.235 -172.205 173.565 -171.875 ;
        RECT 173.235 -173.565 173.565 -173.235 ;
        RECT 173.235 -174.925 173.565 -174.595 ;
        RECT 173.235 -176.285 173.565 -175.955 ;
        RECT 173.235 -177.645 173.565 -177.315 ;
        RECT 173.235 -179.005 173.565 -178.675 ;
        RECT 173.235 -180.365 173.565 -180.035 ;
        RECT 173.235 -181.725 173.565 -181.395 ;
        RECT 173.235 -183.085 173.565 -182.755 ;
        RECT 173.235 -184.445 173.565 -184.115 ;
        RECT 173.235 -185.805 173.565 -185.475 ;
        RECT 173.235 -187.165 173.565 -186.835 ;
        RECT 173.235 -188.525 173.565 -188.195 ;
        RECT 173.235 -189.885 173.565 -189.555 ;
        RECT 173.235 -191.245 173.565 -190.915 ;
        RECT 173.235 -192.605 173.565 -192.275 ;
        RECT 173.235 -193.965 173.565 -193.635 ;
        RECT 173.235 -195.325 173.565 -194.995 ;
        RECT 173.235 -196.685 173.565 -196.355 ;
        RECT 173.235 -198.045 173.565 -197.715 ;
        RECT 173.235 -199.405 173.565 -199.075 ;
        RECT 173.235 -200.765 173.565 -200.435 ;
        RECT 173.235 -202.125 173.565 -201.795 ;
        RECT 173.235 -203.485 173.565 -203.155 ;
        RECT 173.235 -204.845 173.565 -204.515 ;
        RECT 173.235 -206.205 173.565 -205.875 ;
        RECT 173.235 -207.565 173.565 -207.235 ;
        RECT 173.235 -208.925 173.565 -208.595 ;
        RECT 173.235 -210.285 173.565 -209.955 ;
        RECT 173.235 -211.645 173.565 -211.315 ;
        RECT 173.235 -213.005 173.565 -212.675 ;
        RECT 173.235 -214.365 173.565 -214.035 ;
        RECT 173.235 -215.725 173.565 -215.395 ;
        RECT 173.235 -217.085 173.565 -216.755 ;
        RECT 173.235 -218.445 173.565 -218.115 ;
        RECT 173.235 -219.805 173.565 -219.475 ;
        RECT 173.235 -221.165 173.565 -220.835 ;
        RECT 173.235 -222.525 173.565 -222.195 ;
        RECT 173.235 -223.885 173.565 -223.555 ;
        RECT 173.235 -225.245 173.565 -224.915 ;
        RECT 173.235 -226.605 173.565 -226.275 ;
        RECT 173.235 -227.965 173.565 -227.635 ;
        RECT 173.235 -229.325 173.565 -228.995 ;
        RECT 173.235 -230.685 173.565 -230.355 ;
        RECT 173.235 -232.045 173.565 -231.715 ;
        RECT 173.235 -233.405 173.565 -233.075 ;
        RECT 173.235 -234.765 173.565 -234.435 ;
        RECT 173.235 -236.125 173.565 -235.795 ;
        RECT 173.235 -237.485 173.565 -237.155 ;
        RECT 173.235 -238.845 173.565 -238.515 ;
        RECT 173.235 -241.09 173.565 -239.96 ;
        RECT 173.24 -241.205 173.56 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 244.04 174.925 245.17 ;
        RECT 174.595 242.595 174.925 242.925 ;
        RECT 174.595 241.235 174.925 241.565 ;
        RECT 174.595 239.875 174.925 240.205 ;
        RECT 174.595 238.515 174.925 238.845 ;
        RECT 174.595 237.155 174.925 237.485 ;
        RECT 174.6 237.155 174.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 -0.845 174.925 -0.515 ;
        RECT 174.595 -2.205 174.925 -1.875 ;
        RECT 174.595 -3.565 174.925 -3.235 ;
        RECT 174.6 -3.565 174.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 -123.245 174.925 -122.915 ;
        RECT 174.595 -124.605 174.925 -124.275 ;
        RECT 174.595 -125.965 174.925 -125.635 ;
        RECT 174.595 -127.325 174.925 -126.995 ;
        RECT 174.595 -128.685 174.925 -128.355 ;
        RECT 174.595 -130.045 174.925 -129.715 ;
        RECT 174.595 -131.405 174.925 -131.075 ;
        RECT 174.595 -132.765 174.925 -132.435 ;
        RECT 174.595 -134.125 174.925 -133.795 ;
        RECT 174.595 -135.485 174.925 -135.155 ;
        RECT 174.595 -136.845 174.925 -136.515 ;
        RECT 174.595 -138.205 174.925 -137.875 ;
        RECT 174.595 -139.565 174.925 -139.235 ;
        RECT 174.595 -140.925 174.925 -140.595 ;
        RECT 174.595 -142.285 174.925 -141.955 ;
        RECT 174.595 -143.645 174.925 -143.315 ;
        RECT 174.595 -145.005 174.925 -144.675 ;
        RECT 174.595 -146.365 174.925 -146.035 ;
        RECT 174.595 -147.725 174.925 -147.395 ;
        RECT 174.595 -149.085 174.925 -148.755 ;
        RECT 174.595 -150.445 174.925 -150.115 ;
        RECT 174.595 -151.805 174.925 -151.475 ;
        RECT 174.595 -153.165 174.925 -152.835 ;
        RECT 174.595 -154.525 174.925 -154.195 ;
        RECT 174.595 -155.885 174.925 -155.555 ;
        RECT 174.595 -157.245 174.925 -156.915 ;
        RECT 174.595 -158.605 174.925 -158.275 ;
        RECT 174.595 -159.965 174.925 -159.635 ;
        RECT 174.595 -161.325 174.925 -160.995 ;
        RECT 174.595 -162.685 174.925 -162.355 ;
        RECT 174.595 -164.045 174.925 -163.715 ;
        RECT 174.595 -165.405 174.925 -165.075 ;
        RECT 174.595 -166.765 174.925 -166.435 ;
        RECT 174.595 -168.125 174.925 -167.795 ;
        RECT 174.595 -169.485 174.925 -169.155 ;
        RECT 174.595 -170.845 174.925 -170.515 ;
        RECT 174.595 -172.205 174.925 -171.875 ;
        RECT 174.595 -173.565 174.925 -173.235 ;
        RECT 174.595 -174.925 174.925 -174.595 ;
        RECT 174.595 -176.285 174.925 -175.955 ;
        RECT 174.595 -177.645 174.925 -177.315 ;
        RECT 174.595 -179.005 174.925 -178.675 ;
        RECT 174.595 -180.365 174.925 -180.035 ;
        RECT 174.595 -181.725 174.925 -181.395 ;
        RECT 174.595 -183.085 174.925 -182.755 ;
        RECT 174.595 -184.445 174.925 -184.115 ;
        RECT 174.595 -185.805 174.925 -185.475 ;
        RECT 174.595 -187.165 174.925 -186.835 ;
        RECT 174.595 -188.525 174.925 -188.195 ;
        RECT 174.595 -189.885 174.925 -189.555 ;
        RECT 174.595 -191.245 174.925 -190.915 ;
        RECT 174.595 -192.605 174.925 -192.275 ;
        RECT 174.595 -193.965 174.925 -193.635 ;
        RECT 174.595 -195.325 174.925 -194.995 ;
        RECT 174.595 -196.685 174.925 -196.355 ;
        RECT 174.595 -198.045 174.925 -197.715 ;
        RECT 174.595 -199.405 174.925 -199.075 ;
        RECT 174.595 -200.765 174.925 -200.435 ;
        RECT 174.595 -202.125 174.925 -201.795 ;
        RECT 174.595 -203.485 174.925 -203.155 ;
        RECT 174.595 -204.845 174.925 -204.515 ;
        RECT 174.595 -206.205 174.925 -205.875 ;
        RECT 174.595 -207.565 174.925 -207.235 ;
        RECT 174.595 -208.925 174.925 -208.595 ;
        RECT 174.595 -210.285 174.925 -209.955 ;
        RECT 174.595 -211.645 174.925 -211.315 ;
        RECT 174.595 -213.005 174.925 -212.675 ;
        RECT 174.595 -214.365 174.925 -214.035 ;
        RECT 174.595 -215.725 174.925 -215.395 ;
        RECT 174.595 -217.085 174.925 -216.755 ;
        RECT 174.595 -218.445 174.925 -218.115 ;
        RECT 174.595 -219.805 174.925 -219.475 ;
        RECT 174.595 -221.165 174.925 -220.835 ;
        RECT 174.595 -222.525 174.925 -222.195 ;
        RECT 174.595 -223.885 174.925 -223.555 ;
        RECT 174.595 -225.245 174.925 -224.915 ;
        RECT 174.595 -226.605 174.925 -226.275 ;
        RECT 174.595 -227.965 174.925 -227.635 ;
        RECT 174.595 -229.325 174.925 -228.995 ;
        RECT 174.595 -230.685 174.925 -230.355 ;
        RECT 174.595 -232.045 174.925 -231.715 ;
        RECT 174.595 -233.405 174.925 -233.075 ;
        RECT 174.595 -234.765 174.925 -234.435 ;
        RECT 174.595 -236.125 174.925 -235.795 ;
        RECT 174.595 -237.485 174.925 -237.155 ;
        RECT 174.595 -238.845 174.925 -238.515 ;
        RECT 174.595 -241.09 174.925 -239.96 ;
        RECT 174.6 -241.205 174.92 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 244.04 176.285 245.17 ;
        RECT 175.955 242.595 176.285 242.925 ;
        RECT 175.955 241.235 176.285 241.565 ;
        RECT 175.955 239.875 176.285 240.205 ;
        RECT 175.955 238.515 176.285 238.845 ;
        RECT 175.955 237.155 176.285 237.485 ;
        RECT 175.96 237.155 176.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 -0.845 176.285 -0.515 ;
        RECT 175.955 -2.205 176.285 -1.875 ;
        RECT 175.955 -3.565 176.285 -3.235 ;
        RECT 175.96 -3.565 176.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 -123.245 176.285 -122.915 ;
        RECT 175.955 -124.605 176.285 -124.275 ;
        RECT 175.955 -125.965 176.285 -125.635 ;
        RECT 175.955 -127.325 176.285 -126.995 ;
        RECT 175.955 -128.685 176.285 -128.355 ;
        RECT 175.955 -130.045 176.285 -129.715 ;
        RECT 175.955 -131.405 176.285 -131.075 ;
        RECT 175.955 -132.765 176.285 -132.435 ;
        RECT 175.955 -134.125 176.285 -133.795 ;
        RECT 175.955 -135.485 176.285 -135.155 ;
        RECT 175.955 -136.845 176.285 -136.515 ;
        RECT 175.955 -138.205 176.285 -137.875 ;
        RECT 175.955 -139.565 176.285 -139.235 ;
        RECT 175.955 -140.925 176.285 -140.595 ;
        RECT 175.955 -142.285 176.285 -141.955 ;
        RECT 175.955 -143.645 176.285 -143.315 ;
        RECT 175.955 -145.005 176.285 -144.675 ;
        RECT 175.955 -146.365 176.285 -146.035 ;
        RECT 175.955 -147.725 176.285 -147.395 ;
        RECT 175.955 -149.085 176.285 -148.755 ;
        RECT 175.955 -150.445 176.285 -150.115 ;
        RECT 175.955 -151.805 176.285 -151.475 ;
        RECT 175.955 -153.165 176.285 -152.835 ;
        RECT 175.955 -154.525 176.285 -154.195 ;
        RECT 175.955 -155.885 176.285 -155.555 ;
        RECT 175.955 -157.245 176.285 -156.915 ;
        RECT 175.955 -158.605 176.285 -158.275 ;
        RECT 175.955 -159.965 176.285 -159.635 ;
        RECT 175.955 -161.325 176.285 -160.995 ;
        RECT 175.955 -162.685 176.285 -162.355 ;
        RECT 175.955 -164.045 176.285 -163.715 ;
        RECT 175.955 -165.405 176.285 -165.075 ;
        RECT 175.955 -166.765 176.285 -166.435 ;
        RECT 175.955 -168.125 176.285 -167.795 ;
        RECT 175.955 -169.485 176.285 -169.155 ;
        RECT 175.955 -170.845 176.285 -170.515 ;
        RECT 175.955 -172.205 176.285 -171.875 ;
        RECT 175.955 -173.565 176.285 -173.235 ;
        RECT 175.955 -174.925 176.285 -174.595 ;
        RECT 175.955 -176.285 176.285 -175.955 ;
        RECT 175.955 -177.645 176.285 -177.315 ;
        RECT 175.955 -179.005 176.285 -178.675 ;
        RECT 175.955 -180.365 176.285 -180.035 ;
        RECT 175.955 -181.725 176.285 -181.395 ;
        RECT 175.955 -183.085 176.285 -182.755 ;
        RECT 175.955 -184.445 176.285 -184.115 ;
        RECT 175.955 -185.805 176.285 -185.475 ;
        RECT 175.955 -187.165 176.285 -186.835 ;
        RECT 175.955 -188.525 176.285 -188.195 ;
        RECT 175.955 -189.885 176.285 -189.555 ;
        RECT 175.955 -191.245 176.285 -190.915 ;
        RECT 175.955 -192.605 176.285 -192.275 ;
        RECT 175.955 -193.965 176.285 -193.635 ;
        RECT 175.955 -195.325 176.285 -194.995 ;
        RECT 175.955 -196.685 176.285 -196.355 ;
        RECT 175.955 -198.045 176.285 -197.715 ;
        RECT 175.955 -199.405 176.285 -199.075 ;
        RECT 175.955 -200.765 176.285 -200.435 ;
        RECT 175.955 -202.125 176.285 -201.795 ;
        RECT 175.955 -203.485 176.285 -203.155 ;
        RECT 175.955 -204.845 176.285 -204.515 ;
        RECT 175.955 -206.205 176.285 -205.875 ;
        RECT 175.955 -207.565 176.285 -207.235 ;
        RECT 175.955 -208.925 176.285 -208.595 ;
        RECT 175.955 -210.285 176.285 -209.955 ;
        RECT 175.955 -211.645 176.285 -211.315 ;
        RECT 175.955 -213.005 176.285 -212.675 ;
        RECT 175.955 -214.365 176.285 -214.035 ;
        RECT 175.955 -215.725 176.285 -215.395 ;
        RECT 175.955 -217.085 176.285 -216.755 ;
        RECT 175.955 -218.445 176.285 -218.115 ;
        RECT 175.955 -219.805 176.285 -219.475 ;
        RECT 175.955 -221.165 176.285 -220.835 ;
        RECT 175.955 -222.525 176.285 -222.195 ;
        RECT 175.955 -223.885 176.285 -223.555 ;
        RECT 175.955 -225.245 176.285 -224.915 ;
        RECT 175.955 -226.605 176.285 -226.275 ;
        RECT 175.955 -227.965 176.285 -227.635 ;
        RECT 175.955 -229.325 176.285 -228.995 ;
        RECT 175.955 -230.685 176.285 -230.355 ;
        RECT 175.955 -232.045 176.285 -231.715 ;
        RECT 175.955 -233.405 176.285 -233.075 ;
        RECT 175.955 -234.765 176.285 -234.435 ;
        RECT 175.955 -236.125 176.285 -235.795 ;
        RECT 175.955 -237.485 176.285 -237.155 ;
        RECT 175.955 -238.845 176.285 -238.515 ;
        RECT 175.955 -241.09 176.285 -239.96 ;
        RECT 175.96 -241.205 176.28 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 244.04 177.645 245.17 ;
        RECT 177.315 242.595 177.645 242.925 ;
        RECT 177.315 241.235 177.645 241.565 ;
        RECT 177.315 239.875 177.645 240.205 ;
        RECT 177.315 238.515 177.645 238.845 ;
        RECT 177.315 237.155 177.645 237.485 ;
        RECT 177.32 237.155 177.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 -127.325 177.645 -126.995 ;
        RECT 177.315 -128.685 177.645 -128.355 ;
        RECT 177.315 -130.045 177.645 -129.715 ;
        RECT 177.315 -131.405 177.645 -131.075 ;
        RECT 177.315 -132.765 177.645 -132.435 ;
        RECT 177.315 -134.125 177.645 -133.795 ;
        RECT 177.315 -135.485 177.645 -135.155 ;
        RECT 177.315 -136.845 177.645 -136.515 ;
        RECT 177.315 -138.205 177.645 -137.875 ;
        RECT 177.315 -139.565 177.645 -139.235 ;
        RECT 177.315 -140.925 177.645 -140.595 ;
        RECT 177.315 -142.285 177.645 -141.955 ;
        RECT 177.315 -143.645 177.645 -143.315 ;
        RECT 177.315 -145.005 177.645 -144.675 ;
        RECT 177.315 -146.365 177.645 -146.035 ;
        RECT 177.315 -147.725 177.645 -147.395 ;
        RECT 177.315 -149.085 177.645 -148.755 ;
        RECT 177.315 -150.445 177.645 -150.115 ;
        RECT 177.315 -151.805 177.645 -151.475 ;
        RECT 177.315 -153.165 177.645 -152.835 ;
        RECT 177.315 -154.525 177.645 -154.195 ;
        RECT 177.315 -155.885 177.645 -155.555 ;
        RECT 177.315 -157.245 177.645 -156.915 ;
        RECT 177.315 -158.605 177.645 -158.275 ;
        RECT 177.315 -159.965 177.645 -159.635 ;
        RECT 177.315 -161.325 177.645 -160.995 ;
        RECT 177.315 -162.685 177.645 -162.355 ;
        RECT 177.315 -164.045 177.645 -163.715 ;
        RECT 177.315 -165.405 177.645 -165.075 ;
        RECT 177.315 -166.765 177.645 -166.435 ;
        RECT 177.315 -168.125 177.645 -167.795 ;
        RECT 177.315 -169.485 177.645 -169.155 ;
        RECT 177.315 -170.845 177.645 -170.515 ;
        RECT 177.315 -172.205 177.645 -171.875 ;
        RECT 177.315 -173.565 177.645 -173.235 ;
        RECT 177.315 -174.925 177.645 -174.595 ;
        RECT 177.315 -176.285 177.645 -175.955 ;
        RECT 177.315 -177.645 177.645 -177.315 ;
        RECT 177.315 -179.005 177.645 -178.675 ;
        RECT 177.315 -180.365 177.645 -180.035 ;
        RECT 177.315 -181.725 177.645 -181.395 ;
        RECT 177.315 -183.085 177.645 -182.755 ;
        RECT 177.315 -184.445 177.645 -184.115 ;
        RECT 177.315 -185.805 177.645 -185.475 ;
        RECT 177.315 -187.165 177.645 -186.835 ;
        RECT 177.315 -188.525 177.645 -188.195 ;
        RECT 177.315 -189.885 177.645 -189.555 ;
        RECT 177.315 -191.245 177.645 -190.915 ;
        RECT 177.315 -192.605 177.645 -192.275 ;
        RECT 177.315 -193.965 177.645 -193.635 ;
        RECT 177.315 -195.325 177.645 -194.995 ;
        RECT 177.315 -196.685 177.645 -196.355 ;
        RECT 177.315 -198.045 177.645 -197.715 ;
        RECT 177.315 -199.405 177.645 -199.075 ;
        RECT 177.315 -200.765 177.645 -200.435 ;
        RECT 177.315 -202.125 177.645 -201.795 ;
        RECT 177.315 -203.485 177.645 -203.155 ;
        RECT 177.315 -204.845 177.645 -204.515 ;
        RECT 177.315 -206.205 177.645 -205.875 ;
        RECT 177.315 -207.565 177.645 -207.235 ;
        RECT 177.315 -208.925 177.645 -208.595 ;
        RECT 177.315 -210.285 177.645 -209.955 ;
        RECT 177.315 -211.645 177.645 -211.315 ;
        RECT 177.315 -213.005 177.645 -212.675 ;
        RECT 177.315 -214.365 177.645 -214.035 ;
        RECT 177.315 -215.725 177.645 -215.395 ;
        RECT 177.315 -217.085 177.645 -216.755 ;
        RECT 177.315 -218.445 177.645 -218.115 ;
        RECT 177.315 -219.805 177.645 -219.475 ;
        RECT 177.315 -221.165 177.645 -220.835 ;
        RECT 177.315 -222.525 177.645 -222.195 ;
        RECT 177.315 -223.885 177.645 -223.555 ;
        RECT 177.315 -225.245 177.645 -224.915 ;
        RECT 177.315 -226.605 177.645 -226.275 ;
        RECT 177.315 -227.965 177.645 -227.635 ;
        RECT 177.315 -229.325 177.645 -228.995 ;
        RECT 177.315 -230.685 177.645 -230.355 ;
        RECT 177.315 -232.045 177.645 -231.715 ;
        RECT 177.315 -233.405 177.645 -233.075 ;
        RECT 177.315 -234.765 177.645 -234.435 ;
        RECT 177.315 -236.125 177.645 -235.795 ;
        RECT 177.315 -237.485 177.645 -237.155 ;
        RECT 177.315 -238.845 177.645 -238.515 ;
        RECT 177.315 -241.09 177.645 -239.96 ;
        RECT 177.32 -241.205 177.64 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.71 -125.535 178.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 244.04 179.005 245.17 ;
        RECT 178.675 242.595 179.005 242.925 ;
        RECT 178.675 241.235 179.005 241.565 ;
        RECT 178.675 239.875 179.005 240.205 ;
        RECT 178.675 238.515 179.005 238.845 ;
        RECT 178.675 237.155 179.005 237.485 ;
        RECT 178.68 237.155 179 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 -0.845 179.005 -0.515 ;
        RECT 178.675 -2.205 179.005 -1.875 ;
        RECT 178.675 -3.565 179.005 -3.235 ;
        RECT 178.68 -3.565 179 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 244.04 180.365 245.17 ;
        RECT 180.035 242.595 180.365 242.925 ;
        RECT 180.035 241.235 180.365 241.565 ;
        RECT 180.035 239.875 180.365 240.205 ;
        RECT 180.035 238.515 180.365 238.845 ;
        RECT 180.035 237.155 180.365 237.485 ;
        RECT 180.04 237.155 180.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 -0.845 180.365 -0.515 ;
        RECT 180.035 -2.205 180.365 -1.875 ;
        RECT 180.035 -3.565 180.365 -3.235 ;
        RECT 180.04 -3.565 180.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 244.04 181.725 245.17 ;
        RECT 181.395 242.595 181.725 242.925 ;
        RECT 181.395 241.235 181.725 241.565 ;
        RECT 181.395 239.875 181.725 240.205 ;
        RECT 181.395 238.515 181.725 238.845 ;
        RECT 181.395 237.155 181.725 237.485 ;
        RECT 181.4 237.155 181.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 -0.845 181.725 -0.515 ;
        RECT 181.395 -2.205 181.725 -1.875 ;
        RECT 181.395 -3.565 181.725 -3.235 ;
        RECT 181.4 -3.565 181.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 -123.245 181.725 -122.915 ;
        RECT 181.395 -124.605 181.725 -124.275 ;
        RECT 181.395 -125.965 181.725 -125.635 ;
        RECT 181.395 -127.325 181.725 -126.995 ;
        RECT 181.395 -128.685 181.725 -128.355 ;
        RECT 181.395 -130.045 181.725 -129.715 ;
        RECT 181.395 -131.405 181.725 -131.075 ;
        RECT 181.395 -132.765 181.725 -132.435 ;
        RECT 181.395 -134.125 181.725 -133.795 ;
        RECT 181.395 -135.485 181.725 -135.155 ;
        RECT 181.395 -136.845 181.725 -136.515 ;
        RECT 181.395 -138.205 181.725 -137.875 ;
        RECT 181.395 -139.565 181.725 -139.235 ;
        RECT 181.395 -140.925 181.725 -140.595 ;
        RECT 181.395 -142.285 181.725 -141.955 ;
        RECT 181.395 -143.645 181.725 -143.315 ;
        RECT 181.395 -145.005 181.725 -144.675 ;
        RECT 181.395 -146.365 181.725 -146.035 ;
        RECT 181.395 -147.725 181.725 -147.395 ;
        RECT 181.395 -149.085 181.725 -148.755 ;
        RECT 181.395 -150.445 181.725 -150.115 ;
        RECT 181.395 -151.805 181.725 -151.475 ;
        RECT 181.395 -153.165 181.725 -152.835 ;
        RECT 181.395 -154.525 181.725 -154.195 ;
        RECT 181.395 -155.885 181.725 -155.555 ;
        RECT 181.395 -157.245 181.725 -156.915 ;
        RECT 181.395 -158.605 181.725 -158.275 ;
        RECT 181.395 -159.965 181.725 -159.635 ;
        RECT 181.395 -161.325 181.725 -160.995 ;
        RECT 181.395 -162.685 181.725 -162.355 ;
        RECT 181.395 -164.045 181.725 -163.715 ;
        RECT 181.395 -165.405 181.725 -165.075 ;
        RECT 181.395 -166.765 181.725 -166.435 ;
        RECT 181.395 -168.125 181.725 -167.795 ;
        RECT 181.395 -169.485 181.725 -169.155 ;
        RECT 181.395 -170.845 181.725 -170.515 ;
        RECT 181.395 -172.205 181.725 -171.875 ;
        RECT 181.395 -173.565 181.725 -173.235 ;
        RECT 181.395 -174.925 181.725 -174.595 ;
        RECT 181.395 -176.285 181.725 -175.955 ;
        RECT 181.395 -177.645 181.725 -177.315 ;
        RECT 181.395 -179.005 181.725 -178.675 ;
        RECT 181.395 -180.365 181.725 -180.035 ;
        RECT 181.395 -181.725 181.725 -181.395 ;
        RECT 181.395 -183.085 181.725 -182.755 ;
        RECT 181.395 -184.445 181.725 -184.115 ;
        RECT 181.395 -185.805 181.725 -185.475 ;
        RECT 181.395 -187.165 181.725 -186.835 ;
        RECT 181.395 -188.525 181.725 -188.195 ;
        RECT 181.395 -189.885 181.725 -189.555 ;
        RECT 181.395 -191.245 181.725 -190.915 ;
        RECT 181.395 -192.605 181.725 -192.275 ;
        RECT 181.395 -193.965 181.725 -193.635 ;
        RECT 181.395 -195.325 181.725 -194.995 ;
        RECT 181.395 -196.685 181.725 -196.355 ;
        RECT 181.395 -198.045 181.725 -197.715 ;
        RECT 181.395 -199.405 181.725 -199.075 ;
        RECT 181.395 -200.765 181.725 -200.435 ;
        RECT 181.395 -202.125 181.725 -201.795 ;
        RECT 181.395 -203.485 181.725 -203.155 ;
        RECT 181.395 -204.845 181.725 -204.515 ;
        RECT 181.395 -206.205 181.725 -205.875 ;
        RECT 181.395 -207.565 181.725 -207.235 ;
        RECT 181.395 -208.925 181.725 -208.595 ;
        RECT 181.395 -210.285 181.725 -209.955 ;
        RECT 181.395 -211.645 181.725 -211.315 ;
        RECT 181.395 -213.005 181.725 -212.675 ;
        RECT 181.395 -214.365 181.725 -214.035 ;
        RECT 181.395 -215.725 181.725 -215.395 ;
        RECT 181.395 -217.085 181.725 -216.755 ;
        RECT 181.395 -218.445 181.725 -218.115 ;
        RECT 181.395 -219.805 181.725 -219.475 ;
        RECT 181.395 -221.165 181.725 -220.835 ;
        RECT 181.395 -222.525 181.725 -222.195 ;
        RECT 181.395 -223.885 181.725 -223.555 ;
        RECT 181.395 -225.245 181.725 -224.915 ;
        RECT 181.395 -226.605 181.725 -226.275 ;
        RECT 181.395 -227.965 181.725 -227.635 ;
        RECT 181.395 -229.325 181.725 -228.995 ;
        RECT 181.395 -230.685 181.725 -230.355 ;
        RECT 181.395 -232.045 181.725 -231.715 ;
        RECT 181.395 -233.405 181.725 -233.075 ;
        RECT 181.395 -234.765 181.725 -234.435 ;
        RECT 181.395 -236.125 181.725 -235.795 ;
        RECT 181.395 -237.485 181.725 -237.155 ;
        RECT 181.395 -238.845 181.725 -238.515 ;
        RECT 181.395 -241.09 181.725 -239.96 ;
        RECT 181.4 -241.205 181.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 244.04 183.085 245.17 ;
        RECT 182.755 242.595 183.085 242.925 ;
        RECT 182.755 241.235 183.085 241.565 ;
        RECT 182.755 239.875 183.085 240.205 ;
        RECT 182.755 238.515 183.085 238.845 ;
        RECT 182.755 237.155 183.085 237.485 ;
        RECT 182.76 237.155 183.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 -0.845 183.085 -0.515 ;
        RECT 182.755 -2.205 183.085 -1.875 ;
        RECT 182.755 -3.565 183.085 -3.235 ;
        RECT 182.76 -3.565 183.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 -179.005 183.085 -178.675 ;
        RECT 182.755 -180.365 183.085 -180.035 ;
        RECT 182.755 -181.725 183.085 -181.395 ;
        RECT 182.755 -183.085 183.085 -182.755 ;
        RECT 182.755 -184.445 183.085 -184.115 ;
        RECT 182.755 -185.805 183.085 -185.475 ;
        RECT 182.755 -187.165 183.085 -186.835 ;
        RECT 182.755 -188.525 183.085 -188.195 ;
        RECT 182.755 -189.885 183.085 -189.555 ;
        RECT 182.755 -191.245 183.085 -190.915 ;
        RECT 182.755 -192.605 183.085 -192.275 ;
        RECT 182.755 -193.965 183.085 -193.635 ;
        RECT 182.755 -195.325 183.085 -194.995 ;
        RECT 182.755 -196.685 183.085 -196.355 ;
        RECT 182.755 -198.045 183.085 -197.715 ;
        RECT 182.755 -199.405 183.085 -199.075 ;
        RECT 182.755 -200.765 183.085 -200.435 ;
        RECT 182.755 -202.125 183.085 -201.795 ;
        RECT 182.755 -203.485 183.085 -203.155 ;
        RECT 182.755 -204.845 183.085 -204.515 ;
        RECT 182.755 -206.205 183.085 -205.875 ;
        RECT 182.755 -207.565 183.085 -207.235 ;
        RECT 182.755 -208.925 183.085 -208.595 ;
        RECT 182.755 -210.285 183.085 -209.955 ;
        RECT 182.755 -211.645 183.085 -211.315 ;
        RECT 182.755 -213.005 183.085 -212.675 ;
        RECT 182.755 -214.365 183.085 -214.035 ;
        RECT 182.755 -215.725 183.085 -215.395 ;
        RECT 182.755 -217.085 183.085 -216.755 ;
        RECT 182.755 -218.445 183.085 -218.115 ;
        RECT 182.755 -219.805 183.085 -219.475 ;
        RECT 182.755 -221.165 183.085 -220.835 ;
        RECT 182.755 -222.525 183.085 -222.195 ;
        RECT 182.755 -223.885 183.085 -223.555 ;
        RECT 182.755 -225.245 183.085 -224.915 ;
        RECT 182.755 -226.605 183.085 -226.275 ;
        RECT 182.755 -227.965 183.085 -227.635 ;
        RECT 182.755 -229.325 183.085 -228.995 ;
        RECT 182.755 -230.685 183.085 -230.355 ;
        RECT 182.755 -232.045 183.085 -231.715 ;
        RECT 182.755 -233.405 183.085 -233.075 ;
        RECT 182.755 -234.765 183.085 -234.435 ;
        RECT 182.755 -236.125 183.085 -235.795 ;
        RECT 182.755 -237.485 183.085 -237.155 ;
        RECT 182.755 -238.845 183.085 -238.515 ;
        RECT 182.755 -241.09 183.085 -239.96 ;
        RECT 182.76 -241.205 183.08 -122.24 ;
        RECT 182.755 -123.245 183.085 -122.915 ;
        RECT 182.755 -124.605 183.085 -124.275 ;
        RECT 182.755 -125.965 183.085 -125.635 ;
        RECT 182.755 -127.325 183.085 -126.995 ;
        RECT 182.755 -128.685 183.085 -128.355 ;
        RECT 182.755 -130.045 183.085 -129.715 ;
        RECT 182.755 -131.405 183.085 -131.075 ;
        RECT 182.755 -132.765 183.085 -132.435 ;
        RECT 182.755 -134.125 183.085 -133.795 ;
        RECT 182.755 -135.485 183.085 -135.155 ;
        RECT 182.755 -136.845 183.085 -136.515 ;
        RECT 182.755 -138.205 183.085 -137.875 ;
        RECT 182.755 -139.565 183.085 -139.235 ;
        RECT 182.755 -140.925 183.085 -140.595 ;
        RECT 182.755 -142.285 183.085 -141.955 ;
        RECT 182.755 -143.645 183.085 -143.315 ;
        RECT 182.755 -145.005 183.085 -144.675 ;
        RECT 182.755 -146.365 183.085 -146.035 ;
        RECT 182.755 -147.725 183.085 -147.395 ;
        RECT 182.755 -149.085 183.085 -148.755 ;
        RECT 182.755 -150.445 183.085 -150.115 ;
        RECT 182.755 -151.805 183.085 -151.475 ;
        RECT 182.755 -153.165 183.085 -152.835 ;
        RECT 182.755 -154.525 183.085 -154.195 ;
        RECT 182.755 -155.885 183.085 -155.555 ;
        RECT 182.755 -157.245 183.085 -156.915 ;
        RECT 182.755 -158.605 183.085 -158.275 ;
        RECT 182.755 -159.965 183.085 -159.635 ;
        RECT 182.755 -161.325 183.085 -160.995 ;
        RECT 182.755 -162.685 183.085 -162.355 ;
        RECT 182.755 -164.045 183.085 -163.715 ;
        RECT 182.755 -165.405 183.085 -165.075 ;
        RECT 182.755 -166.765 183.085 -166.435 ;
        RECT 182.755 -168.125 183.085 -167.795 ;
        RECT 182.755 -169.485 183.085 -169.155 ;
        RECT 182.755 -170.845 183.085 -170.515 ;
        RECT 182.755 -172.205 183.085 -171.875 ;
        RECT 182.755 -173.565 183.085 -173.235 ;
        RECT 182.755 -174.925 183.085 -174.595 ;
        RECT 182.755 -176.285 183.085 -175.955 ;
        RECT 182.755 -177.645 183.085 -177.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 244.04 147.725 245.17 ;
        RECT 147.395 242.595 147.725 242.925 ;
        RECT 147.395 241.235 147.725 241.565 ;
        RECT 147.395 239.875 147.725 240.205 ;
        RECT 147.395 238.515 147.725 238.845 ;
        RECT 147.395 237.155 147.725 237.485 ;
        RECT 147.4 237.155 147.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 -0.845 147.725 -0.515 ;
        RECT 147.395 -2.205 147.725 -1.875 ;
        RECT 147.395 -3.565 147.725 -3.235 ;
        RECT 147.4 -3.565 147.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 244.04 149.085 245.17 ;
        RECT 148.755 242.595 149.085 242.925 ;
        RECT 148.755 241.235 149.085 241.565 ;
        RECT 148.755 239.875 149.085 240.205 ;
        RECT 148.755 238.515 149.085 238.845 ;
        RECT 148.755 237.155 149.085 237.485 ;
        RECT 148.76 237.155 149.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 -0.845 149.085 -0.515 ;
        RECT 148.755 -2.205 149.085 -1.875 ;
        RECT 148.755 -3.565 149.085 -3.235 ;
        RECT 148.76 -3.565 149.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 -123.245 149.085 -122.915 ;
        RECT 148.755 -124.605 149.085 -124.275 ;
        RECT 148.755 -125.965 149.085 -125.635 ;
        RECT 148.755 -127.325 149.085 -126.995 ;
        RECT 148.755 -128.685 149.085 -128.355 ;
        RECT 148.755 -130.045 149.085 -129.715 ;
        RECT 148.755 -131.405 149.085 -131.075 ;
        RECT 148.755 -132.765 149.085 -132.435 ;
        RECT 148.755 -134.125 149.085 -133.795 ;
        RECT 148.755 -135.485 149.085 -135.155 ;
        RECT 148.755 -136.845 149.085 -136.515 ;
        RECT 148.755 -138.205 149.085 -137.875 ;
        RECT 148.755 -139.565 149.085 -139.235 ;
        RECT 148.755 -140.925 149.085 -140.595 ;
        RECT 148.755 -142.285 149.085 -141.955 ;
        RECT 148.755 -143.645 149.085 -143.315 ;
        RECT 148.755 -145.005 149.085 -144.675 ;
        RECT 148.755 -146.365 149.085 -146.035 ;
        RECT 148.755 -147.725 149.085 -147.395 ;
        RECT 148.755 -149.085 149.085 -148.755 ;
        RECT 148.755 -150.445 149.085 -150.115 ;
        RECT 148.755 -151.805 149.085 -151.475 ;
        RECT 148.755 -153.165 149.085 -152.835 ;
        RECT 148.755 -154.525 149.085 -154.195 ;
        RECT 148.755 -155.885 149.085 -155.555 ;
        RECT 148.755 -157.245 149.085 -156.915 ;
        RECT 148.755 -158.605 149.085 -158.275 ;
        RECT 148.755 -159.965 149.085 -159.635 ;
        RECT 148.755 -161.325 149.085 -160.995 ;
        RECT 148.755 -162.685 149.085 -162.355 ;
        RECT 148.755 -164.045 149.085 -163.715 ;
        RECT 148.755 -165.405 149.085 -165.075 ;
        RECT 148.755 -166.765 149.085 -166.435 ;
        RECT 148.755 -168.125 149.085 -167.795 ;
        RECT 148.755 -169.485 149.085 -169.155 ;
        RECT 148.755 -170.845 149.085 -170.515 ;
        RECT 148.755 -172.205 149.085 -171.875 ;
        RECT 148.755 -173.565 149.085 -173.235 ;
        RECT 148.755 -174.925 149.085 -174.595 ;
        RECT 148.755 -176.285 149.085 -175.955 ;
        RECT 148.755 -177.645 149.085 -177.315 ;
        RECT 148.755 -179.005 149.085 -178.675 ;
        RECT 148.755 -180.365 149.085 -180.035 ;
        RECT 148.755 -181.725 149.085 -181.395 ;
        RECT 148.755 -183.085 149.085 -182.755 ;
        RECT 148.755 -184.445 149.085 -184.115 ;
        RECT 148.755 -185.805 149.085 -185.475 ;
        RECT 148.755 -187.165 149.085 -186.835 ;
        RECT 148.755 -188.525 149.085 -188.195 ;
        RECT 148.755 -189.885 149.085 -189.555 ;
        RECT 148.755 -191.245 149.085 -190.915 ;
        RECT 148.755 -192.605 149.085 -192.275 ;
        RECT 148.755 -193.965 149.085 -193.635 ;
        RECT 148.755 -195.325 149.085 -194.995 ;
        RECT 148.755 -196.685 149.085 -196.355 ;
        RECT 148.755 -198.045 149.085 -197.715 ;
        RECT 148.755 -199.405 149.085 -199.075 ;
        RECT 148.755 -200.765 149.085 -200.435 ;
        RECT 148.755 -202.125 149.085 -201.795 ;
        RECT 148.755 -203.485 149.085 -203.155 ;
        RECT 148.755 -204.845 149.085 -204.515 ;
        RECT 148.755 -206.205 149.085 -205.875 ;
        RECT 148.755 -207.565 149.085 -207.235 ;
        RECT 148.755 -208.925 149.085 -208.595 ;
        RECT 148.755 -210.285 149.085 -209.955 ;
        RECT 148.755 -211.645 149.085 -211.315 ;
        RECT 148.755 -213.005 149.085 -212.675 ;
        RECT 148.755 -214.365 149.085 -214.035 ;
        RECT 148.755 -215.725 149.085 -215.395 ;
        RECT 148.755 -217.085 149.085 -216.755 ;
        RECT 148.755 -218.445 149.085 -218.115 ;
        RECT 148.755 -219.805 149.085 -219.475 ;
        RECT 148.755 -221.165 149.085 -220.835 ;
        RECT 148.755 -222.525 149.085 -222.195 ;
        RECT 148.755 -223.885 149.085 -223.555 ;
        RECT 148.755 -225.245 149.085 -224.915 ;
        RECT 148.755 -226.605 149.085 -226.275 ;
        RECT 148.755 -227.965 149.085 -227.635 ;
        RECT 148.755 -229.325 149.085 -228.995 ;
        RECT 148.755 -230.685 149.085 -230.355 ;
        RECT 148.755 -232.045 149.085 -231.715 ;
        RECT 148.755 -233.405 149.085 -233.075 ;
        RECT 148.755 -234.765 149.085 -234.435 ;
        RECT 148.755 -236.125 149.085 -235.795 ;
        RECT 148.755 -237.485 149.085 -237.155 ;
        RECT 148.755 -238.845 149.085 -238.515 ;
        RECT 148.755 -241.09 149.085 -239.96 ;
        RECT 148.76 -241.205 149.08 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 244.04 150.445 245.17 ;
        RECT 150.115 242.595 150.445 242.925 ;
        RECT 150.115 241.235 150.445 241.565 ;
        RECT 150.115 239.875 150.445 240.205 ;
        RECT 150.115 238.515 150.445 238.845 ;
        RECT 150.115 237.155 150.445 237.485 ;
        RECT 150.12 237.155 150.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 -0.845 150.445 -0.515 ;
        RECT 150.115 -2.205 150.445 -1.875 ;
        RECT 150.115 -3.565 150.445 -3.235 ;
        RECT 150.12 -3.565 150.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 -123.245 150.445 -122.915 ;
        RECT 150.115 -124.605 150.445 -124.275 ;
        RECT 150.115 -125.965 150.445 -125.635 ;
        RECT 150.115 -127.325 150.445 -126.995 ;
        RECT 150.115 -128.685 150.445 -128.355 ;
        RECT 150.115 -130.045 150.445 -129.715 ;
        RECT 150.115 -131.405 150.445 -131.075 ;
        RECT 150.115 -132.765 150.445 -132.435 ;
        RECT 150.115 -134.125 150.445 -133.795 ;
        RECT 150.115 -135.485 150.445 -135.155 ;
        RECT 150.115 -136.845 150.445 -136.515 ;
        RECT 150.115 -138.205 150.445 -137.875 ;
        RECT 150.115 -139.565 150.445 -139.235 ;
        RECT 150.115 -140.925 150.445 -140.595 ;
        RECT 150.115 -142.285 150.445 -141.955 ;
        RECT 150.115 -143.645 150.445 -143.315 ;
        RECT 150.115 -145.005 150.445 -144.675 ;
        RECT 150.115 -146.365 150.445 -146.035 ;
        RECT 150.115 -147.725 150.445 -147.395 ;
        RECT 150.115 -149.085 150.445 -148.755 ;
        RECT 150.115 -150.445 150.445 -150.115 ;
        RECT 150.115 -151.805 150.445 -151.475 ;
        RECT 150.115 -153.165 150.445 -152.835 ;
        RECT 150.115 -154.525 150.445 -154.195 ;
        RECT 150.115 -155.885 150.445 -155.555 ;
        RECT 150.115 -157.245 150.445 -156.915 ;
        RECT 150.115 -158.605 150.445 -158.275 ;
        RECT 150.115 -159.965 150.445 -159.635 ;
        RECT 150.115 -161.325 150.445 -160.995 ;
        RECT 150.115 -162.685 150.445 -162.355 ;
        RECT 150.115 -164.045 150.445 -163.715 ;
        RECT 150.115 -165.405 150.445 -165.075 ;
        RECT 150.115 -166.765 150.445 -166.435 ;
        RECT 150.115 -168.125 150.445 -167.795 ;
        RECT 150.115 -169.485 150.445 -169.155 ;
        RECT 150.115 -170.845 150.445 -170.515 ;
        RECT 150.115 -172.205 150.445 -171.875 ;
        RECT 150.115 -173.565 150.445 -173.235 ;
        RECT 150.115 -174.925 150.445 -174.595 ;
        RECT 150.115 -176.285 150.445 -175.955 ;
        RECT 150.115 -177.645 150.445 -177.315 ;
        RECT 150.115 -179.005 150.445 -178.675 ;
        RECT 150.115 -180.365 150.445 -180.035 ;
        RECT 150.115 -181.725 150.445 -181.395 ;
        RECT 150.115 -183.085 150.445 -182.755 ;
        RECT 150.115 -184.445 150.445 -184.115 ;
        RECT 150.115 -185.805 150.445 -185.475 ;
        RECT 150.115 -187.165 150.445 -186.835 ;
        RECT 150.115 -188.525 150.445 -188.195 ;
        RECT 150.115 -189.885 150.445 -189.555 ;
        RECT 150.115 -191.245 150.445 -190.915 ;
        RECT 150.115 -192.605 150.445 -192.275 ;
        RECT 150.115 -193.965 150.445 -193.635 ;
        RECT 150.115 -195.325 150.445 -194.995 ;
        RECT 150.115 -196.685 150.445 -196.355 ;
        RECT 150.115 -198.045 150.445 -197.715 ;
        RECT 150.115 -199.405 150.445 -199.075 ;
        RECT 150.115 -200.765 150.445 -200.435 ;
        RECT 150.115 -202.125 150.445 -201.795 ;
        RECT 150.115 -203.485 150.445 -203.155 ;
        RECT 150.115 -204.845 150.445 -204.515 ;
        RECT 150.115 -206.205 150.445 -205.875 ;
        RECT 150.115 -207.565 150.445 -207.235 ;
        RECT 150.115 -208.925 150.445 -208.595 ;
        RECT 150.115 -210.285 150.445 -209.955 ;
        RECT 150.115 -211.645 150.445 -211.315 ;
        RECT 150.115 -213.005 150.445 -212.675 ;
        RECT 150.115 -214.365 150.445 -214.035 ;
        RECT 150.115 -215.725 150.445 -215.395 ;
        RECT 150.115 -217.085 150.445 -216.755 ;
        RECT 150.115 -218.445 150.445 -218.115 ;
        RECT 150.115 -219.805 150.445 -219.475 ;
        RECT 150.115 -221.165 150.445 -220.835 ;
        RECT 150.115 -222.525 150.445 -222.195 ;
        RECT 150.115 -223.885 150.445 -223.555 ;
        RECT 150.115 -225.245 150.445 -224.915 ;
        RECT 150.115 -226.605 150.445 -226.275 ;
        RECT 150.115 -227.965 150.445 -227.635 ;
        RECT 150.115 -229.325 150.445 -228.995 ;
        RECT 150.115 -230.685 150.445 -230.355 ;
        RECT 150.115 -232.045 150.445 -231.715 ;
        RECT 150.115 -233.405 150.445 -233.075 ;
        RECT 150.115 -234.765 150.445 -234.435 ;
        RECT 150.115 -236.125 150.445 -235.795 ;
        RECT 150.115 -237.485 150.445 -237.155 ;
        RECT 150.115 -238.845 150.445 -238.515 ;
        RECT 150.115 -241.09 150.445 -239.96 ;
        RECT 150.12 -241.205 150.44 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 244.04 151.805 245.17 ;
        RECT 151.475 242.595 151.805 242.925 ;
        RECT 151.475 241.235 151.805 241.565 ;
        RECT 151.475 239.875 151.805 240.205 ;
        RECT 151.475 238.515 151.805 238.845 ;
        RECT 151.475 237.155 151.805 237.485 ;
        RECT 151.48 237.155 151.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 -0.845 151.805 -0.515 ;
        RECT 151.475 -2.205 151.805 -1.875 ;
        RECT 151.475 -3.565 151.805 -3.235 ;
        RECT 151.48 -3.565 151.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 -123.245 151.805 -122.915 ;
        RECT 151.475 -124.605 151.805 -124.275 ;
        RECT 151.475 -125.965 151.805 -125.635 ;
        RECT 151.475 -127.325 151.805 -126.995 ;
        RECT 151.475 -128.685 151.805 -128.355 ;
        RECT 151.475 -130.045 151.805 -129.715 ;
        RECT 151.475 -131.405 151.805 -131.075 ;
        RECT 151.475 -132.765 151.805 -132.435 ;
        RECT 151.475 -134.125 151.805 -133.795 ;
        RECT 151.475 -135.485 151.805 -135.155 ;
        RECT 151.475 -136.845 151.805 -136.515 ;
        RECT 151.475 -138.205 151.805 -137.875 ;
        RECT 151.475 -139.565 151.805 -139.235 ;
        RECT 151.475 -140.925 151.805 -140.595 ;
        RECT 151.475 -142.285 151.805 -141.955 ;
        RECT 151.475 -143.645 151.805 -143.315 ;
        RECT 151.475 -145.005 151.805 -144.675 ;
        RECT 151.475 -146.365 151.805 -146.035 ;
        RECT 151.475 -147.725 151.805 -147.395 ;
        RECT 151.475 -149.085 151.805 -148.755 ;
        RECT 151.475 -150.445 151.805 -150.115 ;
        RECT 151.475 -151.805 151.805 -151.475 ;
        RECT 151.475 -153.165 151.805 -152.835 ;
        RECT 151.475 -154.525 151.805 -154.195 ;
        RECT 151.475 -155.885 151.805 -155.555 ;
        RECT 151.475 -157.245 151.805 -156.915 ;
        RECT 151.475 -158.605 151.805 -158.275 ;
        RECT 151.475 -159.965 151.805 -159.635 ;
        RECT 151.475 -161.325 151.805 -160.995 ;
        RECT 151.475 -162.685 151.805 -162.355 ;
        RECT 151.475 -164.045 151.805 -163.715 ;
        RECT 151.475 -165.405 151.805 -165.075 ;
        RECT 151.475 -166.765 151.805 -166.435 ;
        RECT 151.475 -168.125 151.805 -167.795 ;
        RECT 151.475 -169.485 151.805 -169.155 ;
        RECT 151.475 -170.845 151.805 -170.515 ;
        RECT 151.475 -172.205 151.805 -171.875 ;
        RECT 151.475 -173.565 151.805 -173.235 ;
        RECT 151.475 -174.925 151.805 -174.595 ;
        RECT 151.475 -176.285 151.805 -175.955 ;
        RECT 151.475 -177.645 151.805 -177.315 ;
        RECT 151.475 -179.005 151.805 -178.675 ;
        RECT 151.475 -180.365 151.805 -180.035 ;
        RECT 151.475 -181.725 151.805 -181.395 ;
        RECT 151.475 -183.085 151.805 -182.755 ;
        RECT 151.475 -184.445 151.805 -184.115 ;
        RECT 151.475 -185.805 151.805 -185.475 ;
        RECT 151.475 -187.165 151.805 -186.835 ;
        RECT 151.475 -188.525 151.805 -188.195 ;
        RECT 151.475 -189.885 151.805 -189.555 ;
        RECT 151.475 -191.245 151.805 -190.915 ;
        RECT 151.475 -192.605 151.805 -192.275 ;
        RECT 151.475 -193.965 151.805 -193.635 ;
        RECT 151.475 -195.325 151.805 -194.995 ;
        RECT 151.475 -196.685 151.805 -196.355 ;
        RECT 151.475 -198.045 151.805 -197.715 ;
        RECT 151.475 -199.405 151.805 -199.075 ;
        RECT 151.475 -200.765 151.805 -200.435 ;
        RECT 151.475 -202.125 151.805 -201.795 ;
        RECT 151.475 -203.485 151.805 -203.155 ;
        RECT 151.475 -204.845 151.805 -204.515 ;
        RECT 151.475 -206.205 151.805 -205.875 ;
        RECT 151.475 -207.565 151.805 -207.235 ;
        RECT 151.475 -208.925 151.805 -208.595 ;
        RECT 151.475 -210.285 151.805 -209.955 ;
        RECT 151.475 -211.645 151.805 -211.315 ;
        RECT 151.475 -213.005 151.805 -212.675 ;
        RECT 151.475 -214.365 151.805 -214.035 ;
        RECT 151.475 -215.725 151.805 -215.395 ;
        RECT 151.475 -217.085 151.805 -216.755 ;
        RECT 151.475 -218.445 151.805 -218.115 ;
        RECT 151.475 -219.805 151.805 -219.475 ;
        RECT 151.475 -221.165 151.805 -220.835 ;
        RECT 151.475 -222.525 151.805 -222.195 ;
        RECT 151.475 -223.885 151.805 -223.555 ;
        RECT 151.475 -225.245 151.805 -224.915 ;
        RECT 151.475 -226.605 151.805 -226.275 ;
        RECT 151.475 -227.965 151.805 -227.635 ;
        RECT 151.475 -229.325 151.805 -228.995 ;
        RECT 151.475 -230.685 151.805 -230.355 ;
        RECT 151.475 -232.045 151.805 -231.715 ;
        RECT 151.475 -233.405 151.805 -233.075 ;
        RECT 151.475 -234.765 151.805 -234.435 ;
        RECT 151.475 -236.125 151.805 -235.795 ;
        RECT 151.475 -237.485 151.805 -237.155 ;
        RECT 151.475 -238.845 151.805 -238.515 ;
        RECT 151.475 -241.09 151.805 -239.96 ;
        RECT 151.48 -241.205 151.8 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 244.04 153.165 245.17 ;
        RECT 152.835 242.595 153.165 242.925 ;
        RECT 152.835 241.235 153.165 241.565 ;
        RECT 152.835 239.875 153.165 240.205 ;
        RECT 152.835 238.515 153.165 238.845 ;
        RECT 152.835 237.155 153.165 237.485 ;
        RECT 152.84 237.155 153.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 -0.845 153.165 -0.515 ;
        RECT 152.835 -2.205 153.165 -1.875 ;
        RECT 152.835 -3.565 153.165 -3.235 ;
        RECT 152.84 -3.565 153.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 -123.245 153.165 -122.915 ;
        RECT 152.835 -124.605 153.165 -124.275 ;
        RECT 152.835 -125.965 153.165 -125.635 ;
        RECT 152.835 -127.325 153.165 -126.995 ;
        RECT 152.835 -128.685 153.165 -128.355 ;
        RECT 152.835 -130.045 153.165 -129.715 ;
        RECT 152.835 -131.405 153.165 -131.075 ;
        RECT 152.835 -132.765 153.165 -132.435 ;
        RECT 152.835 -134.125 153.165 -133.795 ;
        RECT 152.835 -135.485 153.165 -135.155 ;
        RECT 152.835 -136.845 153.165 -136.515 ;
        RECT 152.835 -138.205 153.165 -137.875 ;
        RECT 152.835 -139.565 153.165 -139.235 ;
        RECT 152.835 -140.925 153.165 -140.595 ;
        RECT 152.835 -142.285 153.165 -141.955 ;
        RECT 152.835 -143.645 153.165 -143.315 ;
        RECT 152.835 -145.005 153.165 -144.675 ;
        RECT 152.835 -146.365 153.165 -146.035 ;
        RECT 152.835 -147.725 153.165 -147.395 ;
        RECT 152.835 -149.085 153.165 -148.755 ;
        RECT 152.835 -150.445 153.165 -150.115 ;
        RECT 152.835 -151.805 153.165 -151.475 ;
        RECT 152.835 -153.165 153.165 -152.835 ;
        RECT 152.835 -154.525 153.165 -154.195 ;
        RECT 152.835 -155.885 153.165 -155.555 ;
        RECT 152.835 -157.245 153.165 -156.915 ;
        RECT 152.835 -158.605 153.165 -158.275 ;
        RECT 152.835 -159.965 153.165 -159.635 ;
        RECT 152.835 -161.325 153.165 -160.995 ;
        RECT 152.835 -162.685 153.165 -162.355 ;
        RECT 152.835 -164.045 153.165 -163.715 ;
        RECT 152.835 -165.405 153.165 -165.075 ;
        RECT 152.835 -166.765 153.165 -166.435 ;
        RECT 152.835 -168.125 153.165 -167.795 ;
        RECT 152.835 -169.485 153.165 -169.155 ;
        RECT 152.835 -170.845 153.165 -170.515 ;
        RECT 152.835 -172.205 153.165 -171.875 ;
        RECT 152.835 -173.565 153.165 -173.235 ;
        RECT 152.835 -174.925 153.165 -174.595 ;
        RECT 152.835 -176.285 153.165 -175.955 ;
        RECT 152.835 -177.645 153.165 -177.315 ;
        RECT 152.835 -179.005 153.165 -178.675 ;
        RECT 152.835 -180.365 153.165 -180.035 ;
        RECT 152.835 -181.725 153.165 -181.395 ;
        RECT 152.835 -183.085 153.165 -182.755 ;
        RECT 152.835 -184.445 153.165 -184.115 ;
        RECT 152.835 -185.805 153.165 -185.475 ;
        RECT 152.835 -187.165 153.165 -186.835 ;
        RECT 152.835 -188.525 153.165 -188.195 ;
        RECT 152.835 -189.885 153.165 -189.555 ;
        RECT 152.835 -191.245 153.165 -190.915 ;
        RECT 152.835 -192.605 153.165 -192.275 ;
        RECT 152.835 -193.965 153.165 -193.635 ;
        RECT 152.835 -195.325 153.165 -194.995 ;
        RECT 152.835 -196.685 153.165 -196.355 ;
        RECT 152.835 -198.045 153.165 -197.715 ;
        RECT 152.835 -199.405 153.165 -199.075 ;
        RECT 152.835 -200.765 153.165 -200.435 ;
        RECT 152.835 -202.125 153.165 -201.795 ;
        RECT 152.835 -203.485 153.165 -203.155 ;
        RECT 152.835 -204.845 153.165 -204.515 ;
        RECT 152.835 -206.205 153.165 -205.875 ;
        RECT 152.835 -207.565 153.165 -207.235 ;
        RECT 152.835 -208.925 153.165 -208.595 ;
        RECT 152.835 -210.285 153.165 -209.955 ;
        RECT 152.835 -211.645 153.165 -211.315 ;
        RECT 152.835 -213.005 153.165 -212.675 ;
        RECT 152.835 -214.365 153.165 -214.035 ;
        RECT 152.835 -215.725 153.165 -215.395 ;
        RECT 152.835 -217.085 153.165 -216.755 ;
        RECT 152.835 -218.445 153.165 -218.115 ;
        RECT 152.835 -219.805 153.165 -219.475 ;
        RECT 152.835 -221.165 153.165 -220.835 ;
        RECT 152.835 -222.525 153.165 -222.195 ;
        RECT 152.835 -223.885 153.165 -223.555 ;
        RECT 152.835 -225.245 153.165 -224.915 ;
        RECT 152.835 -226.605 153.165 -226.275 ;
        RECT 152.835 -227.965 153.165 -227.635 ;
        RECT 152.835 -229.325 153.165 -228.995 ;
        RECT 152.835 -230.685 153.165 -230.355 ;
        RECT 152.835 -232.045 153.165 -231.715 ;
        RECT 152.835 -233.405 153.165 -233.075 ;
        RECT 152.835 -234.765 153.165 -234.435 ;
        RECT 152.835 -236.125 153.165 -235.795 ;
        RECT 152.835 -237.485 153.165 -237.155 ;
        RECT 152.835 -238.845 153.165 -238.515 ;
        RECT 152.835 -241.09 153.165 -239.96 ;
        RECT 152.84 -241.205 153.16 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 244.04 154.525 245.17 ;
        RECT 154.195 242.595 154.525 242.925 ;
        RECT 154.195 241.235 154.525 241.565 ;
        RECT 154.195 239.875 154.525 240.205 ;
        RECT 154.195 238.515 154.525 238.845 ;
        RECT 154.195 237.155 154.525 237.485 ;
        RECT 154.2 237.155 154.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -0.845 154.525 -0.515 ;
        RECT 154.195 -2.205 154.525 -1.875 ;
        RECT 154.195 -3.565 154.525 -3.235 ;
        RECT 154.2 -3.565 154.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -123.245 154.525 -122.915 ;
        RECT 154.195 -124.605 154.525 -124.275 ;
        RECT 154.195 -125.965 154.525 -125.635 ;
        RECT 154.195 -127.325 154.525 -126.995 ;
        RECT 154.195 -128.685 154.525 -128.355 ;
        RECT 154.195 -130.045 154.525 -129.715 ;
        RECT 154.195 -131.405 154.525 -131.075 ;
        RECT 154.195 -132.765 154.525 -132.435 ;
        RECT 154.195 -134.125 154.525 -133.795 ;
        RECT 154.195 -135.485 154.525 -135.155 ;
        RECT 154.195 -136.845 154.525 -136.515 ;
        RECT 154.195 -138.205 154.525 -137.875 ;
        RECT 154.195 -139.565 154.525 -139.235 ;
        RECT 154.195 -140.925 154.525 -140.595 ;
        RECT 154.195 -142.285 154.525 -141.955 ;
        RECT 154.195 -143.645 154.525 -143.315 ;
        RECT 154.195 -145.005 154.525 -144.675 ;
        RECT 154.195 -146.365 154.525 -146.035 ;
        RECT 154.195 -147.725 154.525 -147.395 ;
        RECT 154.195 -149.085 154.525 -148.755 ;
        RECT 154.195 -150.445 154.525 -150.115 ;
        RECT 154.195 -151.805 154.525 -151.475 ;
        RECT 154.195 -153.165 154.525 -152.835 ;
        RECT 154.195 -154.525 154.525 -154.195 ;
        RECT 154.195 -155.885 154.525 -155.555 ;
        RECT 154.195 -157.245 154.525 -156.915 ;
        RECT 154.195 -158.605 154.525 -158.275 ;
        RECT 154.195 -159.965 154.525 -159.635 ;
        RECT 154.195 -161.325 154.525 -160.995 ;
        RECT 154.195 -162.685 154.525 -162.355 ;
        RECT 154.195 -164.045 154.525 -163.715 ;
        RECT 154.195 -165.405 154.525 -165.075 ;
        RECT 154.195 -166.765 154.525 -166.435 ;
        RECT 154.195 -168.125 154.525 -167.795 ;
        RECT 154.195 -169.485 154.525 -169.155 ;
        RECT 154.195 -170.845 154.525 -170.515 ;
        RECT 154.195 -172.205 154.525 -171.875 ;
        RECT 154.195 -173.565 154.525 -173.235 ;
        RECT 154.195 -174.925 154.525 -174.595 ;
        RECT 154.195 -176.285 154.525 -175.955 ;
        RECT 154.195 -177.645 154.525 -177.315 ;
        RECT 154.195 -179.005 154.525 -178.675 ;
        RECT 154.195 -180.365 154.525 -180.035 ;
        RECT 154.195 -181.725 154.525 -181.395 ;
        RECT 154.195 -183.085 154.525 -182.755 ;
        RECT 154.195 -184.445 154.525 -184.115 ;
        RECT 154.195 -185.805 154.525 -185.475 ;
        RECT 154.195 -187.165 154.525 -186.835 ;
        RECT 154.195 -188.525 154.525 -188.195 ;
        RECT 154.195 -189.885 154.525 -189.555 ;
        RECT 154.195 -191.245 154.525 -190.915 ;
        RECT 154.195 -192.605 154.525 -192.275 ;
        RECT 154.195 -193.965 154.525 -193.635 ;
        RECT 154.195 -195.325 154.525 -194.995 ;
        RECT 154.195 -196.685 154.525 -196.355 ;
        RECT 154.195 -198.045 154.525 -197.715 ;
        RECT 154.195 -199.405 154.525 -199.075 ;
        RECT 154.195 -200.765 154.525 -200.435 ;
        RECT 154.195 -202.125 154.525 -201.795 ;
        RECT 154.195 -203.485 154.525 -203.155 ;
        RECT 154.195 -204.845 154.525 -204.515 ;
        RECT 154.195 -206.205 154.525 -205.875 ;
        RECT 154.195 -207.565 154.525 -207.235 ;
        RECT 154.195 -208.925 154.525 -208.595 ;
        RECT 154.195 -210.285 154.525 -209.955 ;
        RECT 154.195 -211.645 154.525 -211.315 ;
        RECT 154.195 -213.005 154.525 -212.675 ;
        RECT 154.195 -214.365 154.525 -214.035 ;
        RECT 154.195 -215.725 154.525 -215.395 ;
        RECT 154.195 -217.085 154.525 -216.755 ;
        RECT 154.195 -218.445 154.525 -218.115 ;
        RECT 154.195 -219.805 154.525 -219.475 ;
        RECT 154.195 -221.165 154.525 -220.835 ;
        RECT 154.195 -222.525 154.525 -222.195 ;
        RECT 154.195 -223.885 154.525 -223.555 ;
        RECT 154.195 -225.245 154.525 -224.915 ;
        RECT 154.195 -226.605 154.525 -226.275 ;
        RECT 154.195 -227.965 154.525 -227.635 ;
        RECT 154.195 -229.325 154.525 -228.995 ;
        RECT 154.195 -230.685 154.525 -230.355 ;
        RECT 154.195 -232.045 154.525 -231.715 ;
        RECT 154.195 -233.405 154.525 -233.075 ;
        RECT 154.195 -234.765 154.525 -234.435 ;
        RECT 154.195 -236.125 154.525 -235.795 ;
        RECT 154.195 -237.485 154.525 -237.155 ;
        RECT 154.195 -238.845 154.525 -238.515 ;
        RECT 154.195 -241.09 154.525 -239.96 ;
        RECT 154.2 -241.205 154.52 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 244.04 155.885 245.17 ;
        RECT 155.555 242.595 155.885 242.925 ;
        RECT 155.555 241.235 155.885 241.565 ;
        RECT 155.555 239.875 155.885 240.205 ;
        RECT 155.555 238.515 155.885 238.845 ;
        RECT 155.555 237.155 155.885 237.485 ;
        RECT 155.56 237.155 155.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 -127.325 155.885 -126.995 ;
        RECT 155.555 -128.685 155.885 -128.355 ;
        RECT 155.555 -130.045 155.885 -129.715 ;
        RECT 155.555 -131.405 155.885 -131.075 ;
        RECT 155.555 -132.765 155.885 -132.435 ;
        RECT 155.555 -134.125 155.885 -133.795 ;
        RECT 155.555 -135.485 155.885 -135.155 ;
        RECT 155.555 -136.845 155.885 -136.515 ;
        RECT 155.555 -138.205 155.885 -137.875 ;
        RECT 155.555 -139.565 155.885 -139.235 ;
        RECT 155.555 -140.925 155.885 -140.595 ;
        RECT 155.555 -142.285 155.885 -141.955 ;
        RECT 155.555 -143.645 155.885 -143.315 ;
        RECT 155.555 -145.005 155.885 -144.675 ;
        RECT 155.555 -146.365 155.885 -146.035 ;
        RECT 155.555 -147.725 155.885 -147.395 ;
        RECT 155.555 -149.085 155.885 -148.755 ;
        RECT 155.555 -150.445 155.885 -150.115 ;
        RECT 155.555 -151.805 155.885 -151.475 ;
        RECT 155.555 -153.165 155.885 -152.835 ;
        RECT 155.555 -154.525 155.885 -154.195 ;
        RECT 155.555 -155.885 155.885 -155.555 ;
        RECT 155.555 -157.245 155.885 -156.915 ;
        RECT 155.555 -158.605 155.885 -158.275 ;
        RECT 155.555 -159.965 155.885 -159.635 ;
        RECT 155.555 -161.325 155.885 -160.995 ;
        RECT 155.555 -162.685 155.885 -162.355 ;
        RECT 155.555 -164.045 155.885 -163.715 ;
        RECT 155.555 -165.405 155.885 -165.075 ;
        RECT 155.555 -166.765 155.885 -166.435 ;
        RECT 155.555 -168.125 155.885 -167.795 ;
        RECT 155.555 -169.485 155.885 -169.155 ;
        RECT 155.555 -170.845 155.885 -170.515 ;
        RECT 155.555 -172.205 155.885 -171.875 ;
        RECT 155.555 -173.565 155.885 -173.235 ;
        RECT 155.555 -174.925 155.885 -174.595 ;
        RECT 155.555 -176.285 155.885 -175.955 ;
        RECT 155.555 -177.645 155.885 -177.315 ;
        RECT 155.555 -179.005 155.885 -178.675 ;
        RECT 155.555 -180.365 155.885 -180.035 ;
        RECT 155.555 -181.725 155.885 -181.395 ;
        RECT 155.555 -183.085 155.885 -182.755 ;
        RECT 155.555 -184.445 155.885 -184.115 ;
        RECT 155.555 -185.805 155.885 -185.475 ;
        RECT 155.555 -187.165 155.885 -186.835 ;
        RECT 155.555 -188.525 155.885 -188.195 ;
        RECT 155.555 -189.885 155.885 -189.555 ;
        RECT 155.555 -191.245 155.885 -190.915 ;
        RECT 155.555 -192.605 155.885 -192.275 ;
        RECT 155.555 -193.965 155.885 -193.635 ;
        RECT 155.555 -195.325 155.885 -194.995 ;
        RECT 155.555 -196.685 155.885 -196.355 ;
        RECT 155.555 -198.045 155.885 -197.715 ;
        RECT 155.555 -199.405 155.885 -199.075 ;
        RECT 155.555 -200.765 155.885 -200.435 ;
        RECT 155.555 -202.125 155.885 -201.795 ;
        RECT 155.555 -203.485 155.885 -203.155 ;
        RECT 155.555 -204.845 155.885 -204.515 ;
        RECT 155.555 -206.205 155.885 -205.875 ;
        RECT 155.555 -207.565 155.885 -207.235 ;
        RECT 155.555 -208.925 155.885 -208.595 ;
        RECT 155.555 -210.285 155.885 -209.955 ;
        RECT 155.555 -211.645 155.885 -211.315 ;
        RECT 155.555 -213.005 155.885 -212.675 ;
        RECT 155.555 -214.365 155.885 -214.035 ;
        RECT 155.555 -215.725 155.885 -215.395 ;
        RECT 155.555 -217.085 155.885 -216.755 ;
        RECT 155.555 -218.445 155.885 -218.115 ;
        RECT 155.555 -219.805 155.885 -219.475 ;
        RECT 155.555 -221.165 155.885 -220.835 ;
        RECT 155.555 -222.525 155.885 -222.195 ;
        RECT 155.555 -223.885 155.885 -223.555 ;
        RECT 155.555 -225.245 155.885 -224.915 ;
        RECT 155.555 -226.605 155.885 -226.275 ;
        RECT 155.555 -227.965 155.885 -227.635 ;
        RECT 155.555 -229.325 155.885 -228.995 ;
        RECT 155.555 -230.685 155.885 -230.355 ;
        RECT 155.555 -232.045 155.885 -231.715 ;
        RECT 155.555 -233.405 155.885 -233.075 ;
        RECT 155.555 -234.765 155.885 -234.435 ;
        RECT 155.555 -236.125 155.885 -235.795 ;
        RECT 155.555 -237.485 155.885 -237.155 ;
        RECT 155.555 -238.845 155.885 -238.515 ;
        RECT 155.555 -241.09 155.885 -239.96 ;
        RECT 155.56 -241.205 155.88 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.91 -125.535 156.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 244.04 157.245 245.17 ;
        RECT 156.915 242.595 157.245 242.925 ;
        RECT 156.915 241.235 157.245 241.565 ;
        RECT 156.915 239.875 157.245 240.205 ;
        RECT 156.915 238.515 157.245 238.845 ;
        RECT 156.915 237.155 157.245 237.485 ;
        RECT 156.92 237.155 157.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 -0.845 157.245 -0.515 ;
        RECT 156.915 -2.205 157.245 -1.875 ;
        RECT 156.915 -3.565 157.245 -3.235 ;
        RECT 156.92 -3.565 157.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 244.04 158.605 245.17 ;
        RECT 158.275 242.595 158.605 242.925 ;
        RECT 158.275 241.235 158.605 241.565 ;
        RECT 158.275 239.875 158.605 240.205 ;
        RECT 158.275 238.515 158.605 238.845 ;
        RECT 158.275 237.155 158.605 237.485 ;
        RECT 158.28 237.155 158.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 -0.845 158.605 -0.515 ;
        RECT 158.275 -2.205 158.605 -1.875 ;
        RECT 158.275 -3.565 158.605 -3.235 ;
        RECT 158.28 -3.565 158.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 244.04 159.965 245.17 ;
        RECT 159.635 242.595 159.965 242.925 ;
        RECT 159.635 241.235 159.965 241.565 ;
        RECT 159.635 239.875 159.965 240.205 ;
        RECT 159.635 238.515 159.965 238.845 ;
        RECT 159.635 237.155 159.965 237.485 ;
        RECT 159.64 237.155 159.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -0.845 159.965 -0.515 ;
        RECT 159.635 -2.205 159.965 -1.875 ;
        RECT 159.635 -3.565 159.965 -3.235 ;
        RECT 159.64 -3.565 159.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -123.245 159.965 -122.915 ;
        RECT 159.635 -124.605 159.965 -124.275 ;
        RECT 159.635 -125.965 159.965 -125.635 ;
        RECT 159.635 -127.325 159.965 -126.995 ;
        RECT 159.635 -128.685 159.965 -128.355 ;
        RECT 159.635 -130.045 159.965 -129.715 ;
        RECT 159.635 -131.405 159.965 -131.075 ;
        RECT 159.635 -132.765 159.965 -132.435 ;
        RECT 159.635 -134.125 159.965 -133.795 ;
        RECT 159.635 -135.485 159.965 -135.155 ;
        RECT 159.635 -136.845 159.965 -136.515 ;
        RECT 159.635 -138.205 159.965 -137.875 ;
        RECT 159.635 -139.565 159.965 -139.235 ;
        RECT 159.635 -140.925 159.965 -140.595 ;
        RECT 159.635 -142.285 159.965 -141.955 ;
        RECT 159.635 -143.645 159.965 -143.315 ;
        RECT 159.635 -145.005 159.965 -144.675 ;
        RECT 159.635 -146.365 159.965 -146.035 ;
        RECT 159.635 -147.725 159.965 -147.395 ;
        RECT 159.635 -149.085 159.965 -148.755 ;
        RECT 159.635 -150.445 159.965 -150.115 ;
        RECT 159.635 -151.805 159.965 -151.475 ;
        RECT 159.635 -153.165 159.965 -152.835 ;
        RECT 159.635 -154.525 159.965 -154.195 ;
        RECT 159.635 -155.885 159.965 -155.555 ;
        RECT 159.635 -157.245 159.965 -156.915 ;
        RECT 159.635 -158.605 159.965 -158.275 ;
        RECT 159.635 -159.965 159.965 -159.635 ;
        RECT 159.635 -161.325 159.965 -160.995 ;
        RECT 159.635 -162.685 159.965 -162.355 ;
        RECT 159.635 -164.045 159.965 -163.715 ;
        RECT 159.635 -165.405 159.965 -165.075 ;
        RECT 159.635 -166.765 159.965 -166.435 ;
        RECT 159.635 -168.125 159.965 -167.795 ;
        RECT 159.635 -169.485 159.965 -169.155 ;
        RECT 159.635 -170.845 159.965 -170.515 ;
        RECT 159.635 -172.205 159.965 -171.875 ;
        RECT 159.635 -173.565 159.965 -173.235 ;
        RECT 159.635 -174.925 159.965 -174.595 ;
        RECT 159.635 -176.285 159.965 -175.955 ;
        RECT 159.635 -177.645 159.965 -177.315 ;
        RECT 159.635 -179.005 159.965 -178.675 ;
        RECT 159.635 -180.365 159.965 -180.035 ;
        RECT 159.635 -181.725 159.965 -181.395 ;
        RECT 159.635 -183.085 159.965 -182.755 ;
        RECT 159.635 -184.445 159.965 -184.115 ;
        RECT 159.635 -185.805 159.965 -185.475 ;
        RECT 159.635 -187.165 159.965 -186.835 ;
        RECT 159.635 -188.525 159.965 -188.195 ;
        RECT 159.635 -189.885 159.965 -189.555 ;
        RECT 159.635 -191.245 159.965 -190.915 ;
        RECT 159.635 -192.605 159.965 -192.275 ;
        RECT 159.635 -193.965 159.965 -193.635 ;
        RECT 159.635 -195.325 159.965 -194.995 ;
        RECT 159.635 -196.685 159.965 -196.355 ;
        RECT 159.635 -198.045 159.965 -197.715 ;
        RECT 159.635 -199.405 159.965 -199.075 ;
        RECT 159.635 -200.765 159.965 -200.435 ;
        RECT 159.635 -202.125 159.965 -201.795 ;
        RECT 159.635 -203.485 159.965 -203.155 ;
        RECT 159.635 -204.845 159.965 -204.515 ;
        RECT 159.635 -206.205 159.965 -205.875 ;
        RECT 159.635 -207.565 159.965 -207.235 ;
        RECT 159.635 -208.925 159.965 -208.595 ;
        RECT 159.635 -210.285 159.965 -209.955 ;
        RECT 159.635 -211.645 159.965 -211.315 ;
        RECT 159.635 -213.005 159.965 -212.675 ;
        RECT 159.635 -214.365 159.965 -214.035 ;
        RECT 159.635 -215.725 159.965 -215.395 ;
        RECT 159.635 -217.085 159.965 -216.755 ;
        RECT 159.635 -218.445 159.965 -218.115 ;
        RECT 159.635 -219.805 159.965 -219.475 ;
        RECT 159.635 -221.165 159.965 -220.835 ;
        RECT 159.635 -222.525 159.965 -222.195 ;
        RECT 159.635 -223.885 159.965 -223.555 ;
        RECT 159.635 -225.245 159.965 -224.915 ;
        RECT 159.635 -226.605 159.965 -226.275 ;
        RECT 159.635 -227.965 159.965 -227.635 ;
        RECT 159.635 -229.325 159.965 -228.995 ;
        RECT 159.635 -230.685 159.965 -230.355 ;
        RECT 159.635 -232.045 159.965 -231.715 ;
        RECT 159.635 -233.405 159.965 -233.075 ;
        RECT 159.635 -234.765 159.965 -234.435 ;
        RECT 159.635 -236.125 159.965 -235.795 ;
        RECT 159.635 -237.485 159.965 -237.155 ;
        RECT 159.635 -238.845 159.965 -238.515 ;
        RECT 159.635 -241.09 159.965 -239.96 ;
        RECT 159.64 -241.205 159.96 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 244.04 161.325 245.17 ;
        RECT 160.995 242.595 161.325 242.925 ;
        RECT 160.995 241.235 161.325 241.565 ;
        RECT 160.995 239.875 161.325 240.205 ;
        RECT 160.995 238.515 161.325 238.845 ;
        RECT 160.995 237.155 161.325 237.485 ;
        RECT 161 237.155 161.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 -0.845 161.325 -0.515 ;
        RECT 160.995 -2.205 161.325 -1.875 ;
        RECT 160.995 -3.565 161.325 -3.235 ;
        RECT 161 -3.565 161.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 -123.245 161.325 -122.915 ;
        RECT 160.995 -124.605 161.325 -124.275 ;
        RECT 160.995 -125.965 161.325 -125.635 ;
        RECT 160.995 -127.325 161.325 -126.995 ;
        RECT 160.995 -128.685 161.325 -128.355 ;
        RECT 160.995 -130.045 161.325 -129.715 ;
        RECT 160.995 -131.405 161.325 -131.075 ;
        RECT 160.995 -132.765 161.325 -132.435 ;
        RECT 160.995 -134.125 161.325 -133.795 ;
        RECT 160.995 -135.485 161.325 -135.155 ;
        RECT 160.995 -136.845 161.325 -136.515 ;
        RECT 160.995 -138.205 161.325 -137.875 ;
        RECT 160.995 -139.565 161.325 -139.235 ;
        RECT 160.995 -140.925 161.325 -140.595 ;
        RECT 160.995 -142.285 161.325 -141.955 ;
        RECT 160.995 -143.645 161.325 -143.315 ;
        RECT 160.995 -145.005 161.325 -144.675 ;
        RECT 160.995 -146.365 161.325 -146.035 ;
        RECT 160.995 -147.725 161.325 -147.395 ;
        RECT 160.995 -149.085 161.325 -148.755 ;
        RECT 160.995 -150.445 161.325 -150.115 ;
        RECT 160.995 -151.805 161.325 -151.475 ;
        RECT 160.995 -153.165 161.325 -152.835 ;
        RECT 160.995 -154.525 161.325 -154.195 ;
        RECT 160.995 -155.885 161.325 -155.555 ;
        RECT 160.995 -157.245 161.325 -156.915 ;
        RECT 160.995 -158.605 161.325 -158.275 ;
        RECT 160.995 -159.965 161.325 -159.635 ;
        RECT 160.995 -161.325 161.325 -160.995 ;
        RECT 160.995 -162.685 161.325 -162.355 ;
        RECT 160.995 -164.045 161.325 -163.715 ;
        RECT 160.995 -165.405 161.325 -165.075 ;
        RECT 160.995 -166.765 161.325 -166.435 ;
        RECT 160.995 -168.125 161.325 -167.795 ;
        RECT 160.995 -169.485 161.325 -169.155 ;
        RECT 160.995 -170.845 161.325 -170.515 ;
        RECT 160.995 -172.205 161.325 -171.875 ;
        RECT 160.995 -173.565 161.325 -173.235 ;
        RECT 160.995 -174.925 161.325 -174.595 ;
        RECT 160.995 -176.285 161.325 -175.955 ;
        RECT 160.995 -177.645 161.325 -177.315 ;
        RECT 160.995 -179.005 161.325 -178.675 ;
        RECT 160.995 -180.365 161.325 -180.035 ;
        RECT 160.995 -181.725 161.325 -181.395 ;
        RECT 160.995 -183.085 161.325 -182.755 ;
        RECT 160.995 -184.445 161.325 -184.115 ;
        RECT 160.995 -185.805 161.325 -185.475 ;
        RECT 160.995 -187.165 161.325 -186.835 ;
        RECT 160.995 -188.525 161.325 -188.195 ;
        RECT 160.995 -189.885 161.325 -189.555 ;
        RECT 160.995 -191.245 161.325 -190.915 ;
        RECT 160.995 -192.605 161.325 -192.275 ;
        RECT 160.995 -193.965 161.325 -193.635 ;
        RECT 160.995 -195.325 161.325 -194.995 ;
        RECT 160.995 -196.685 161.325 -196.355 ;
        RECT 160.995 -198.045 161.325 -197.715 ;
        RECT 160.995 -199.405 161.325 -199.075 ;
        RECT 160.995 -200.765 161.325 -200.435 ;
        RECT 160.995 -202.125 161.325 -201.795 ;
        RECT 160.995 -203.485 161.325 -203.155 ;
        RECT 160.995 -204.845 161.325 -204.515 ;
        RECT 160.995 -206.205 161.325 -205.875 ;
        RECT 160.995 -207.565 161.325 -207.235 ;
        RECT 160.995 -208.925 161.325 -208.595 ;
        RECT 160.995 -210.285 161.325 -209.955 ;
        RECT 160.995 -211.645 161.325 -211.315 ;
        RECT 160.995 -213.005 161.325 -212.675 ;
        RECT 160.995 -214.365 161.325 -214.035 ;
        RECT 160.995 -215.725 161.325 -215.395 ;
        RECT 160.995 -217.085 161.325 -216.755 ;
        RECT 160.995 -218.445 161.325 -218.115 ;
        RECT 160.995 -219.805 161.325 -219.475 ;
        RECT 160.995 -221.165 161.325 -220.835 ;
        RECT 160.995 -222.525 161.325 -222.195 ;
        RECT 160.995 -223.885 161.325 -223.555 ;
        RECT 160.995 -225.245 161.325 -224.915 ;
        RECT 160.995 -226.605 161.325 -226.275 ;
        RECT 160.995 -227.965 161.325 -227.635 ;
        RECT 160.995 -229.325 161.325 -228.995 ;
        RECT 160.995 -230.685 161.325 -230.355 ;
        RECT 160.995 -232.045 161.325 -231.715 ;
        RECT 160.995 -233.405 161.325 -233.075 ;
        RECT 160.995 -234.765 161.325 -234.435 ;
        RECT 160.995 -236.125 161.325 -235.795 ;
        RECT 160.995 -237.485 161.325 -237.155 ;
        RECT 160.995 -238.845 161.325 -238.515 ;
        RECT 160.995 -241.09 161.325 -239.96 ;
        RECT 161 -241.205 161.32 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 244.04 162.685 245.17 ;
        RECT 162.355 242.595 162.685 242.925 ;
        RECT 162.355 241.235 162.685 241.565 ;
        RECT 162.355 239.875 162.685 240.205 ;
        RECT 162.355 238.515 162.685 238.845 ;
        RECT 162.355 237.155 162.685 237.485 ;
        RECT 162.36 237.155 162.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 -0.845 162.685 -0.515 ;
        RECT 162.355 -2.205 162.685 -1.875 ;
        RECT 162.355 -3.565 162.685 -3.235 ;
        RECT 162.36 -3.565 162.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 -123.245 162.685 -122.915 ;
        RECT 162.355 -124.605 162.685 -124.275 ;
        RECT 162.355 -125.965 162.685 -125.635 ;
        RECT 162.355 -127.325 162.685 -126.995 ;
        RECT 162.355 -128.685 162.685 -128.355 ;
        RECT 162.355 -130.045 162.685 -129.715 ;
        RECT 162.355 -131.405 162.685 -131.075 ;
        RECT 162.355 -132.765 162.685 -132.435 ;
        RECT 162.355 -134.125 162.685 -133.795 ;
        RECT 162.355 -135.485 162.685 -135.155 ;
        RECT 162.355 -136.845 162.685 -136.515 ;
        RECT 162.355 -138.205 162.685 -137.875 ;
        RECT 162.355 -139.565 162.685 -139.235 ;
        RECT 162.355 -140.925 162.685 -140.595 ;
        RECT 162.355 -142.285 162.685 -141.955 ;
        RECT 162.355 -143.645 162.685 -143.315 ;
        RECT 162.355 -145.005 162.685 -144.675 ;
        RECT 162.355 -146.365 162.685 -146.035 ;
        RECT 162.355 -147.725 162.685 -147.395 ;
        RECT 162.355 -149.085 162.685 -148.755 ;
        RECT 162.355 -150.445 162.685 -150.115 ;
        RECT 162.355 -151.805 162.685 -151.475 ;
        RECT 162.355 -153.165 162.685 -152.835 ;
        RECT 162.355 -154.525 162.685 -154.195 ;
        RECT 162.355 -155.885 162.685 -155.555 ;
        RECT 162.355 -157.245 162.685 -156.915 ;
        RECT 162.355 -158.605 162.685 -158.275 ;
        RECT 162.355 -159.965 162.685 -159.635 ;
        RECT 162.355 -161.325 162.685 -160.995 ;
        RECT 162.355 -162.685 162.685 -162.355 ;
        RECT 162.355 -164.045 162.685 -163.715 ;
        RECT 162.355 -165.405 162.685 -165.075 ;
        RECT 162.355 -166.765 162.685 -166.435 ;
        RECT 162.355 -168.125 162.685 -167.795 ;
        RECT 162.355 -169.485 162.685 -169.155 ;
        RECT 162.355 -170.845 162.685 -170.515 ;
        RECT 162.355 -172.205 162.685 -171.875 ;
        RECT 162.355 -173.565 162.685 -173.235 ;
        RECT 162.355 -174.925 162.685 -174.595 ;
        RECT 162.355 -176.285 162.685 -175.955 ;
        RECT 162.355 -177.645 162.685 -177.315 ;
        RECT 162.355 -179.005 162.685 -178.675 ;
        RECT 162.355 -180.365 162.685 -180.035 ;
        RECT 162.355 -181.725 162.685 -181.395 ;
        RECT 162.355 -183.085 162.685 -182.755 ;
        RECT 162.355 -184.445 162.685 -184.115 ;
        RECT 162.355 -185.805 162.685 -185.475 ;
        RECT 162.355 -187.165 162.685 -186.835 ;
        RECT 162.355 -188.525 162.685 -188.195 ;
        RECT 162.355 -189.885 162.685 -189.555 ;
        RECT 162.355 -191.245 162.685 -190.915 ;
        RECT 162.355 -192.605 162.685 -192.275 ;
        RECT 162.355 -193.965 162.685 -193.635 ;
        RECT 162.355 -195.325 162.685 -194.995 ;
        RECT 162.355 -196.685 162.685 -196.355 ;
        RECT 162.355 -198.045 162.685 -197.715 ;
        RECT 162.355 -199.405 162.685 -199.075 ;
        RECT 162.355 -200.765 162.685 -200.435 ;
        RECT 162.355 -202.125 162.685 -201.795 ;
        RECT 162.355 -203.485 162.685 -203.155 ;
        RECT 162.355 -204.845 162.685 -204.515 ;
        RECT 162.355 -206.205 162.685 -205.875 ;
        RECT 162.355 -207.565 162.685 -207.235 ;
        RECT 162.355 -208.925 162.685 -208.595 ;
        RECT 162.355 -210.285 162.685 -209.955 ;
        RECT 162.355 -211.645 162.685 -211.315 ;
        RECT 162.355 -213.005 162.685 -212.675 ;
        RECT 162.355 -214.365 162.685 -214.035 ;
        RECT 162.355 -215.725 162.685 -215.395 ;
        RECT 162.355 -217.085 162.685 -216.755 ;
        RECT 162.355 -218.445 162.685 -218.115 ;
        RECT 162.355 -219.805 162.685 -219.475 ;
        RECT 162.355 -221.165 162.685 -220.835 ;
        RECT 162.355 -222.525 162.685 -222.195 ;
        RECT 162.355 -223.885 162.685 -223.555 ;
        RECT 162.355 -225.245 162.685 -224.915 ;
        RECT 162.355 -226.605 162.685 -226.275 ;
        RECT 162.355 -227.965 162.685 -227.635 ;
        RECT 162.355 -229.325 162.685 -228.995 ;
        RECT 162.355 -230.685 162.685 -230.355 ;
        RECT 162.355 -232.045 162.685 -231.715 ;
        RECT 162.355 -233.405 162.685 -233.075 ;
        RECT 162.355 -234.765 162.685 -234.435 ;
        RECT 162.355 -236.125 162.685 -235.795 ;
        RECT 162.355 -237.485 162.685 -237.155 ;
        RECT 162.355 -238.845 162.685 -238.515 ;
        RECT 162.355 -241.09 162.685 -239.96 ;
        RECT 162.36 -241.205 162.68 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 244.04 164.045 245.17 ;
        RECT 163.715 242.595 164.045 242.925 ;
        RECT 163.715 241.235 164.045 241.565 ;
        RECT 163.715 239.875 164.045 240.205 ;
        RECT 163.715 238.515 164.045 238.845 ;
        RECT 163.715 237.155 164.045 237.485 ;
        RECT 163.72 237.155 164.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 -0.845 164.045 -0.515 ;
        RECT 163.715 -2.205 164.045 -1.875 ;
        RECT 163.715 -3.565 164.045 -3.235 ;
        RECT 163.72 -3.565 164.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 -149.085 164.045 -148.755 ;
        RECT 163.715 -150.445 164.045 -150.115 ;
        RECT 163.715 -151.805 164.045 -151.475 ;
        RECT 163.715 -153.165 164.045 -152.835 ;
        RECT 163.715 -154.525 164.045 -154.195 ;
        RECT 163.715 -155.885 164.045 -155.555 ;
        RECT 163.715 -157.245 164.045 -156.915 ;
        RECT 163.715 -158.605 164.045 -158.275 ;
        RECT 163.715 -159.965 164.045 -159.635 ;
        RECT 163.715 -161.325 164.045 -160.995 ;
        RECT 163.715 -162.685 164.045 -162.355 ;
        RECT 163.715 -164.045 164.045 -163.715 ;
        RECT 163.715 -165.405 164.045 -165.075 ;
        RECT 163.715 -166.765 164.045 -166.435 ;
        RECT 163.715 -168.125 164.045 -167.795 ;
        RECT 163.715 -169.485 164.045 -169.155 ;
        RECT 163.715 -170.845 164.045 -170.515 ;
        RECT 163.715 -172.205 164.045 -171.875 ;
        RECT 163.715 -173.565 164.045 -173.235 ;
        RECT 163.715 -174.925 164.045 -174.595 ;
        RECT 163.715 -176.285 164.045 -175.955 ;
        RECT 163.715 -177.645 164.045 -177.315 ;
        RECT 163.715 -179.005 164.045 -178.675 ;
        RECT 163.715 -180.365 164.045 -180.035 ;
        RECT 163.715 -181.725 164.045 -181.395 ;
        RECT 163.715 -183.085 164.045 -182.755 ;
        RECT 163.715 -184.445 164.045 -184.115 ;
        RECT 163.715 -185.805 164.045 -185.475 ;
        RECT 163.715 -187.165 164.045 -186.835 ;
        RECT 163.715 -188.525 164.045 -188.195 ;
        RECT 163.715 -189.885 164.045 -189.555 ;
        RECT 163.715 -191.245 164.045 -190.915 ;
        RECT 163.715 -192.605 164.045 -192.275 ;
        RECT 163.715 -193.965 164.045 -193.635 ;
        RECT 163.715 -195.325 164.045 -194.995 ;
        RECT 163.715 -196.685 164.045 -196.355 ;
        RECT 163.715 -198.045 164.045 -197.715 ;
        RECT 163.715 -199.405 164.045 -199.075 ;
        RECT 163.715 -200.765 164.045 -200.435 ;
        RECT 163.715 -202.125 164.045 -201.795 ;
        RECT 163.715 -203.485 164.045 -203.155 ;
        RECT 163.715 -204.845 164.045 -204.515 ;
        RECT 163.715 -206.205 164.045 -205.875 ;
        RECT 163.715 -207.565 164.045 -207.235 ;
        RECT 163.715 -208.925 164.045 -208.595 ;
        RECT 163.715 -210.285 164.045 -209.955 ;
        RECT 163.715 -211.645 164.045 -211.315 ;
        RECT 163.715 -213.005 164.045 -212.675 ;
        RECT 163.715 -214.365 164.045 -214.035 ;
        RECT 163.715 -215.725 164.045 -215.395 ;
        RECT 163.715 -217.085 164.045 -216.755 ;
        RECT 163.715 -218.445 164.045 -218.115 ;
        RECT 163.715 -219.805 164.045 -219.475 ;
        RECT 163.715 -221.165 164.045 -220.835 ;
        RECT 163.715 -222.525 164.045 -222.195 ;
        RECT 163.715 -223.885 164.045 -223.555 ;
        RECT 163.715 -225.245 164.045 -224.915 ;
        RECT 163.715 -226.605 164.045 -226.275 ;
        RECT 163.715 -227.965 164.045 -227.635 ;
        RECT 163.715 -229.325 164.045 -228.995 ;
        RECT 163.715 -230.685 164.045 -230.355 ;
        RECT 163.715 -232.045 164.045 -231.715 ;
        RECT 163.715 -233.405 164.045 -233.075 ;
        RECT 163.715 -234.765 164.045 -234.435 ;
        RECT 163.715 -236.125 164.045 -235.795 ;
        RECT 163.715 -237.485 164.045 -237.155 ;
        RECT 163.715 -238.845 164.045 -238.515 ;
        RECT 163.715 -241.09 164.045 -239.96 ;
        RECT 163.72 -241.205 164.04 -122.24 ;
        RECT 163.715 -123.245 164.045 -122.915 ;
        RECT 163.715 -124.605 164.045 -124.275 ;
        RECT 163.715 -125.965 164.045 -125.635 ;
        RECT 163.715 -127.325 164.045 -126.995 ;
        RECT 163.715 -128.685 164.045 -128.355 ;
        RECT 163.715 -130.045 164.045 -129.715 ;
        RECT 163.715 -131.405 164.045 -131.075 ;
        RECT 163.715 -132.765 164.045 -132.435 ;
        RECT 163.715 -134.125 164.045 -133.795 ;
        RECT 163.715 -135.485 164.045 -135.155 ;
        RECT 163.715 -136.845 164.045 -136.515 ;
        RECT 163.715 -138.205 164.045 -137.875 ;
        RECT 163.715 -139.565 164.045 -139.235 ;
        RECT 163.715 -140.925 164.045 -140.595 ;
        RECT 163.715 -142.285 164.045 -141.955 ;
        RECT 163.715 -143.645 164.045 -143.315 ;
        RECT 163.715 -145.005 164.045 -144.675 ;
        RECT 163.715 -146.365 164.045 -146.035 ;
        RECT 163.715 -147.725 164.045 -147.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -123.245 130.045 -122.915 ;
        RECT 129.715 -124.605 130.045 -124.275 ;
        RECT 129.715 -125.965 130.045 -125.635 ;
        RECT 129.715 -127.325 130.045 -126.995 ;
        RECT 129.715 -128.685 130.045 -128.355 ;
        RECT 129.715 -130.045 130.045 -129.715 ;
        RECT 129.715 -131.405 130.045 -131.075 ;
        RECT 129.715 -132.765 130.045 -132.435 ;
        RECT 129.715 -134.125 130.045 -133.795 ;
        RECT 129.715 -135.485 130.045 -135.155 ;
        RECT 129.715 -136.845 130.045 -136.515 ;
        RECT 129.715 -138.205 130.045 -137.875 ;
        RECT 129.715 -139.565 130.045 -139.235 ;
        RECT 129.715 -140.925 130.045 -140.595 ;
        RECT 129.715 -142.285 130.045 -141.955 ;
        RECT 129.715 -143.645 130.045 -143.315 ;
        RECT 129.715 -145.005 130.045 -144.675 ;
        RECT 129.715 -146.365 130.045 -146.035 ;
        RECT 129.715 -147.725 130.045 -147.395 ;
        RECT 129.715 -149.085 130.045 -148.755 ;
        RECT 129.715 -150.445 130.045 -150.115 ;
        RECT 129.715 -151.805 130.045 -151.475 ;
        RECT 129.715 -153.165 130.045 -152.835 ;
        RECT 129.715 -154.525 130.045 -154.195 ;
        RECT 129.715 -155.885 130.045 -155.555 ;
        RECT 129.715 -157.245 130.045 -156.915 ;
        RECT 129.715 -158.605 130.045 -158.275 ;
        RECT 129.715 -159.965 130.045 -159.635 ;
        RECT 129.715 -161.325 130.045 -160.995 ;
        RECT 129.715 -162.685 130.045 -162.355 ;
        RECT 129.715 -164.045 130.045 -163.715 ;
        RECT 129.715 -165.405 130.045 -165.075 ;
        RECT 129.715 -166.765 130.045 -166.435 ;
        RECT 129.715 -168.125 130.045 -167.795 ;
        RECT 129.715 -169.485 130.045 -169.155 ;
        RECT 129.715 -170.845 130.045 -170.515 ;
        RECT 129.715 -172.205 130.045 -171.875 ;
        RECT 129.715 -173.565 130.045 -173.235 ;
        RECT 129.715 -174.925 130.045 -174.595 ;
        RECT 129.715 -176.285 130.045 -175.955 ;
        RECT 129.715 -177.645 130.045 -177.315 ;
        RECT 129.715 -179.005 130.045 -178.675 ;
        RECT 129.715 -180.365 130.045 -180.035 ;
        RECT 129.715 -181.725 130.045 -181.395 ;
        RECT 129.715 -183.085 130.045 -182.755 ;
        RECT 129.715 -184.445 130.045 -184.115 ;
        RECT 129.715 -185.805 130.045 -185.475 ;
        RECT 129.715 -187.165 130.045 -186.835 ;
        RECT 129.715 -188.525 130.045 -188.195 ;
        RECT 129.715 -189.885 130.045 -189.555 ;
        RECT 129.715 -191.245 130.045 -190.915 ;
        RECT 129.715 -192.605 130.045 -192.275 ;
        RECT 129.715 -193.965 130.045 -193.635 ;
        RECT 129.715 -195.325 130.045 -194.995 ;
        RECT 129.715 -196.685 130.045 -196.355 ;
        RECT 129.715 -198.045 130.045 -197.715 ;
        RECT 129.715 -199.405 130.045 -199.075 ;
        RECT 129.715 -200.765 130.045 -200.435 ;
        RECT 129.715 -202.125 130.045 -201.795 ;
        RECT 129.715 -203.485 130.045 -203.155 ;
        RECT 129.715 -204.845 130.045 -204.515 ;
        RECT 129.715 -206.205 130.045 -205.875 ;
        RECT 129.715 -207.565 130.045 -207.235 ;
        RECT 129.715 -208.925 130.045 -208.595 ;
        RECT 129.715 -210.285 130.045 -209.955 ;
        RECT 129.715 -211.645 130.045 -211.315 ;
        RECT 129.715 -213.005 130.045 -212.675 ;
        RECT 129.715 -214.365 130.045 -214.035 ;
        RECT 129.715 -215.725 130.045 -215.395 ;
        RECT 129.715 -217.085 130.045 -216.755 ;
        RECT 129.715 -218.445 130.045 -218.115 ;
        RECT 129.715 -219.805 130.045 -219.475 ;
        RECT 129.715 -221.165 130.045 -220.835 ;
        RECT 129.715 -222.525 130.045 -222.195 ;
        RECT 129.715 -223.885 130.045 -223.555 ;
        RECT 129.715 -225.245 130.045 -224.915 ;
        RECT 129.715 -226.605 130.045 -226.275 ;
        RECT 129.715 -227.965 130.045 -227.635 ;
        RECT 129.715 -229.325 130.045 -228.995 ;
        RECT 129.715 -230.685 130.045 -230.355 ;
        RECT 129.715 -232.045 130.045 -231.715 ;
        RECT 129.715 -233.405 130.045 -233.075 ;
        RECT 129.715 -234.765 130.045 -234.435 ;
        RECT 129.715 -236.125 130.045 -235.795 ;
        RECT 129.715 -237.485 130.045 -237.155 ;
        RECT 129.715 -238.845 130.045 -238.515 ;
        RECT 129.715 -241.09 130.045 -239.96 ;
        RECT 129.72 -241.205 130.04 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 244.04 131.405 245.17 ;
        RECT 131.075 242.595 131.405 242.925 ;
        RECT 131.075 241.235 131.405 241.565 ;
        RECT 131.075 239.875 131.405 240.205 ;
        RECT 131.075 238.515 131.405 238.845 ;
        RECT 131.075 237.155 131.405 237.485 ;
        RECT 131.08 237.155 131.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 -0.845 131.405 -0.515 ;
        RECT 131.075 -2.205 131.405 -1.875 ;
        RECT 131.075 -3.565 131.405 -3.235 ;
        RECT 131.08 -3.565 131.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 -123.245 131.405 -122.915 ;
        RECT 131.075 -124.605 131.405 -124.275 ;
        RECT 131.075 -125.965 131.405 -125.635 ;
        RECT 131.075 -127.325 131.405 -126.995 ;
        RECT 131.075 -128.685 131.405 -128.355 ;
        RECT 131.075 -130.045 131.405 -129.715 ;
        RECT 131.075 -131.405 131.405 -131.075 ;
        RECT 131.075 -132.765 131.405 -132.435 ;
        RECT 131.075 -134.125 131.405 -133.795 ;
        RECT 131.075 -135.485 131.405 -135.155 ;
        RECT 131.075 -136.845 131.405 -136.515 ;
        RECT 131.075 -138.205 131.405 -137.875 ;
        RECT 131.075 -139.565 131.405 -139.235 ;
        RECT 131.075 -140.925 131.405 -140.595 ;
        RECT 131.075 -142.285 131.405 -141.955 ;
        RECT 131.075 -143.645 131.405 -143.315 ;
        RECT 131.075 -145.005 131.405 -144.675 ;
        RECT 131.075 -146.365 131.405 -146.035 ;
        RECT 131.075 -147.725 131.405 -147.395 ;
        RECT 131.075 -149.085 131.405 -148.755 ;
        RECT 131.075 -150.445 131.405 -150.115 ;
        RECT 131.075 -151.805 131.405 -151.475 ;
        RECT 131.075 -153.165 131.405 -152.835 ;
        RECT 131.075 -154.525 131.405 -154.195 ;
        RECT 131.075 -155.885 131.405 -155.555 ;
        RECT 131.075 -157.245 131.405 -156.915 ;
        RECT 131.075 -158.605 131.405 -158.275 ;
        RECT 131.075 -159.965 131.405 -159.635 ;
        RECT 131.075 -161.325 131.405 -160.995 ;
        RECT 131.075 -162.685 131.405 -162.355 ;
        RECT 131.075 -164.045 131.405 -163.715 ;
        RECT 131.075 -165.405 131.405 -165.075 ;
        RECT 131.075 -166.765 131.405 -166.435 ;
        RECT 131.075 -168.125 131.405 -167.795 ;
        RECT 131.075 -169.485 131.405 -169.155 ;
        RECT 131.075 -170.845 131.405 -170.515 ;
        RECT 131.075 -172.205 131.405 -171.875 ;
        RECT 131.075 -173.565 131.405 -173.235 ;
        RECT 131.075 -174.925 131.405 -174.595 ;
        RECT 131.075 -176.285 131.405 -175.955 ;
        RECT 131.075 -177.645 131.405 -177.315 ;
        RECT 131.075 -179.005 131.405 -178.675 ;
        RECT 131.075 -180.365 131.405 -180.035 ;
        RECT 131.075 -181.725 131.405 -181.395 ;
        RECT 131.075 -183.085 131.405 -182.755 ;
        RECT 131.075 -184.445 131.405 -184.115 ;
        RECT 131.075 -185.805 131.405 -185.475 ;
        RECT 131.075 -187.165 131.405 -186.835 ;
        RECT 131.075 -188.525 131.405 -188.195 ;
        RECT 131.075 -189.885 131.405 -189.555 ;
        RECT 131.075 -191.245 131.405 -190.915 ;
        RECT 131.075 -192.605 131.405 -192.275 ;
        RECT 131.075 -193.965 131.405 -193.635 ;
        RECT 131.075 -195.325 131.405 -194.995 ;
        RECT 131.075 -196.685 131.405 -196.355 ;
        RECT 131.075 -198.045 131.405 -197.715 ;
        RECT 131.075 -199.405 131.405 -199.075 ;
        RECT 131.075 -200.765 131.405 -200.435 ;
        RECT 131.075 -202.125 131.405 -201.795 ;
        RECT 131.075 -203.485 131.405 -203.155 ;
        RECT 131.075 -204.845 131.405 -204.515 ;
        RECT 131.075 -206.205 131.405 -205.875 ;
        RECT 131.075 -207.565 131.405 -207.235 ;
        RECT 131.075 -208.925 131.405 -208.595 ;
        RECT 131.075 -210.285 131.405 -209.955 ;
        RECT 131.075 -211.645 131.405 -211.315 ;
        RECT 131.075 -213.005 131.405 -212.675 ;
        RECT 131.075 -214.365 131.405 -214.035 ;
        RECT 131.075 -215.725 131.405 -215.395 ;
        RECT 131.075 -217.085 131.405 -216.755 ;
        RECT 131.075 -218.445 131.405 -218.115 ;
        RECT 131.075 -219.805 131.405 -219.475 ;
        RECT 131.075 -221.165 131.405 -220.835 ;
        RECT 131.075 -222.525 131.405 -222.195 ;
        RECT 131.075 -223.885 131.405 -223.555 ;
        RECT 131.075 -225.245 131.405 -224.915 ;
        RECT 131.075 -226.605 131.405 -226.275 ;
        RECT 131.075 -227.965 131.405 -227.635 ;
        RECT 131.075 -229.325 131.405 -228.995 ;
        RECT 131.075 -230.685 131.405 -230.355 ;
        RECT 131.075 -232.045 131.405 -231.715 ;
        RECT 131.075 -233.405 131.405 -233.075 ;
        RECT 131.075 -234.765 131.405 -234.435 ;
        RECT 131.075 -236.125 131.405 -235.795 ;
        RECT 131.075 -237.485 131.405 -237.155 ;
        RECT 131.075 -238.845 131.405 -238.515 ;
        RECT 131.075 -241.09 131.405 -239.96 ;
        RECT 131.08 -241.205 131.4 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 244.04 132.765 245.17 ;
        RECT 132.435 242.595 132.765 242.925 ;
        RECT 132.435 241.235 132.765 241.565 ;
        RECT 132.435 239.875 132.765 240.205 ;
        RECT 132.435 238.515 132.765 238.845 ;
        RECT 132.435 237.155 132.765 237.485 ;
        RECT 132.44 237.155 132.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 -0.845 132.765 -0.515 ;
        RECT 132.435 -2.205 132.765 -1.875 ;
        RECT 132.435 -3.565 132.765 -3.235 ;
        RECT 132.44 -3.565 132.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 -123.245 132.765 -122.915 ;
        RECT 132.435 -124.605 132.765 -124.275 ;
        RECT 132.435 -125.965 132.765 -125.635 ;
        RECT 132.435 -127.325 132.765 -126.995 ;
        RECT 132.435 -128.685 132.765 -128.355 ;
        RECT 132.435 -130.045 132.765 -129.715 ;
        RECT 132.435 -131.405 132.765 -131.075 ;
        RECT 132.435 -132.765 132.765 -132.435 ;
        RECT 132.435 -134.125 132.765 -133.795 ;
        RECT 132.435 -135.485 132.765 -135.155 ;
        RECT 132.435 -136.845 132.765 -136.515 ;
        RECT 132.435 -138.205 132.765 -137.875 ;
        RECT 132.435 -139.565 132.765 -139.235 ;
        RECT 132.435 -140.925 132.765 -140.595 ;
        RECT 132.435 -142.285 132.765 -141.955 ;
        RECT 132.435 -143.645 132.765 -143.315 ;
        RECT 132.435 -145.005 132.765 -144.675 ;
        RECT 132.435 -146.365 132.765 -146.035 ;
        RECT 132.435 -147.725 132.765 -147.395 ;
        RECT 132.435 -149.085 132.765 -148.755 ;
        RECT 132.435 -150.445 132.765 -150.115 ;
        RECT 132.435 -151.805 132.765 -151.475 ;
        RECT 132.435 -153.165 132.765 -152.835 ;
        RECT 132.435 -154.525 132.765 -154.195 ;
        RECT 132.435 -155.885 132.765 -155.555 ;
        RECT 132.435 -157.245 132.765 -156.915 ;
        RECT 132.435 -158.605 132.765 -158.275 ;
        RECT 132.435 -159.965 132.765 -159.635 ;
        RECT 132.435 -161.325 132.765 -160.995 ;
        RECT 132.435 -162.685 132.765 -162.355 ;
        RECT 132.435 -164.045 132.765 -163.715 ;
        RECT 132.435 -165.405 132.765 -165.075 ;
        RECT 132.435 -166.765 132.765 -166.435 ;
        RECT 132.435 -168.125 132.765 -167.795 ;
        RECT 132.435 -169.485 132.765 -169.155 ;
        RECT 132.435 -170.845 132.765 -170.515 ;
        RECT 132.435 -172.205 132.765 -171.875 ;
        RECT 132.435 -173.565 132.765 -173.235 ;
        RECT 132.435 -174.925 132.765 -174.595 ;
        RECT 132.435 -176.285 132.765 -175.955 ;
        RECT 132.435 -177.645 132.765 -177.315 ;
        RECT 132.435 -179.005 132.765 -178.675 ;
        RECT 132.435 -180.365 132.765 -180.035 ;
        RECT 132.435 -181.725 132.765 -181.395 ;
        RECT 132.435 -183.085 132.765 -182.755 ;
        RECT 132.435 -184.445 132.765 -184.115 ;
        RECT 132.435 -185.805 132.765 -185.475 ;
        RECT 132.435 -187.165 132.765 -186.835 ;
        RECT 132.435 -188.525 132.765 -188.195 ;
        RECT 132.435 -189.885 132.765 -189.555 ;
        RECT 132.435 -191.245 132.765 -190.915 ;
        RECT 132.435 -192.605 132.765 -192.275 ;
        RECT 132.435 -193.965 132.765 -193.635 ;
        RECT 132.435 -195.325 132.765 -194.995 ;
        RECT 132.435 -196.685 132.765 -196.355 ;
        RECT 132.435 -198.045 132.765 -197.715 ;
        RECT 132.435 -199.405 132.765 -199.075 ;
        RECT 132.435 -200.765 132.765 -200.435 ;
        RECT 132.435 -202.125 132.765 -201.795 ;
        RECT 132.435 -203.485 132.765 -203.155 ;
        RECT 132.435 -204.845 132.765 -204.515 ;
        RECT 132.435 -206.205 132.765 -205.875 ;
        RECT 132.435 -207.565 132.765 -207.235 ;
        RECT 132.435 -208.925 132.765 -208.595 ;
        RECT 132.435 -210.285 132.765 -209.955 ;
        RECT 132.435 -211.645 132.765 -211.315 ;
        RECT 132.435 -213.005 132.765 -212.675 ;
        RECT 132.435 -214.365 132.765 -214.035 ;
        RECT 132.435 -215.725 132.765 -215.395 ;
        RECT 132.435 -217.085 132.765 -216.755 ;
        RECT 132.435 -218.445 132.765 -218.115 ;
        RECT 132.435 -219.805 132.765 -219.475 ;
        RECT 132.435 -221.165 132.765 -220.835 ;
        RECT 132.435 -222.525 132.765 -222.195 ;
        RECT 132.435 -223.885 132.765 -223.555 ;
        RECT 132.435 -225.245 132.765 -224.915 ;
        RECT 132.435 -226.605 132.765 -226.275 ;
        RECT 132.435 -227.965 132.765 -227.635 ;
        RECT 132.435 -229.325 132.765 -228.995 ;
        RECT 132.435 -230.685 132.765 -230.355 ;
        RECT 132.435 -232.045 132.765 -231.715 ;
        RECT 132.435 -233.405 132.765 -233.075 ;
        RECT 132.435 -234.765 132.765 -234.435 ;
        RECT 132.435 -236.125 132.765 -235.795 ;
        RECT 132.435 -237.485 132.765 -237.155 ;
        RECT 132.435 -238.845 132.765 -238.515 ;
        RECT 132.435 -241.09 132.765 -239.96 ;
        RECT 132.44 -241.205 132.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 244.04 134.125 245.17 ;
        RECT 133.795 242.595 134.125 242.925 ;
        RECT 133.795 241.235 134.125 241.565 ;
        RECT 133.795 239.875 134.125 240.205 ;
        RECT 133.795 238.515 134.125 238.845 ;
        RECT 133.795 237.155 134.125 237.485 ;
        RECT 133.8 237.155 134.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 -127.325 134.125 -126.995 ;
        RECT 133.795 -128.685 134.125 -128.355 ;
        RECT 133.795 -130.045 134.125 -129.715 ;
        RECT 133.795 -131.405 134.125 -131.075 ;
        RECT 133.795 -132.765 134.125 -132.435 ;
        RECT 133.795 -134.125 134.125 -133.795 ;
        RECT 133.795 -135.485 134.125 -135.155 ;
        RECT 133.795 -136.845 134.125 -136.515 ;
        RECT 133.795 -138.205 134.125 -137.875 ;
        RECT 133.795 -139.565 134.125 -139.235 ;
        RECT 133.795 -140.925 134.125 -140.595 ;
        RECT 133.795 -142.285 134.125 -141.955 ;
        RECT 133.795 -143.645 134.125 -143.315 ;
        RECT 133.795 -145.005 134.125 -144.675 ;
        RECT 133.795 -146.365 134.125 -146.035 ;
        RECT 133.795 -147.725 134.125 -147.395 ;
        RECT 133.795 -149.085 134.125 -148.755 ;
        RECT 133.795 -150.445 134.125 -150.115 ;
        RECT 133.795 -151.805 134.125 -151.475 ;
        RECT 133.795 -153.165 134.125 -152.835 ;
        RECT 133.795 -154.525 134.125 -154.195 ;
        RECT 133.795 -155.885 134.125 -155.555 ;
        RECT 133.795 -157.245 134.125 -156.915 ;
        RECT 133.795 -158.605 134.125 -158.275 ;
        RECT 133.795 -159.965 134.125 -159.635 ;
        RECT 133.795 -161.325 134.125 -160.995 ;
        RECT 133.795 -162.685 134.125 -162.355 ;
        RECT 133.795 -164.045 134.125 -163.715 ;
        RECT 133.795 -165.405 134.125 -165.075 ;
        RECT 133.795 -166.765 134.125 -166.435 ;
        RECT 133.795 -168.125 134.125 -167.795 ;
        RECT 133.795 -169.485 134.125 -169.155 ;
        RECT 133.795 -170.845 134.125 -170.515 ;
        RECT 133.795 -172.205 134.125 -171.875 ;
        RECT 133.795 -173.565 134.125 -173.235 ;
        RECT 133.795 -174.925 134.125 -174.595 ;
        RECT 133.795 -176.285 134.125 -175.955 ;
        RECT 133.795 -177.645 134.125 -177.315 ;
        RECT 133.795 -179.005 134.125 -178.675 ;
        RECT 133.795 -180.365 134.125 -180.035 ;
        RECT 133.795 -181.725 134.125 -181.395 ;
        RECT 133.795 -183.085 134.125 -182.755 ;
        RECT 133.795 -184.445 134.125 -184.115 ;
        RECT 133.795 -185.805 134.125 -185.475 ;
        RECT 133.795 -187.165 134.125 -186.835 ;
        RECT 133.795 -188.525 134.125 -188.195 ;
        RECT 133.795 -189.885 134.125 -189.555 ;
        RECT 133.795 -191.245 134.125 -190.915 ;
        RECT 133.795 -192.605 134.125 -192.275 ;
        RECT 133.795 -193.965 134.125 -193.635 ;
        RECT 133.795 -195.325 134.125 -194.995 ;
        RECT 133.795 -196.685 134.125 -196.355 ;
        RECT 133.795 -198.045 134.125 -197.715 ;
        RECT 133.795 -199.405 134.125 -199.075 ;
        RECT 133.795 -200.765 134.125 -200.435 ;
        RECT 133.795 -202.125 134.125 -201.795 ;
        RECT 133.795 -203.485 134.125 -203.155 ;
        RECT 133.795 -204.845 134.125 -204.515 ;
        RECT 133.795 -206.205 134.125 -205.875 ;
        RECT 133.795 -207.565 134.125 -207.235 ;
        RECT 133.795 -208.925 134.125 -208.595 ;
        RECT 133.795 -210.285 134.125 -209.955 ;
        RECT 133.795 -211.645 134.125 -211.315 ;
        RECT 133.795 -213.005 134.125 -212.675 ;
        RECT 133.795 -214.365 134.125 -214.035 ;
        RECT 133.795 -215.725 134.125 -215.395 ;
        RECT 133.795 -217.085 134.125 -216.755 ;
        RECT 133.795 -218.445 134.125 -218.115 ;
        RECT 133.795 -219.805 134.125 -219.475 ;
        RECT 133.795 -221.165 134.125 -220.835 ;
        RECT 133.795 -222.525 134.125 -222.195 ;
        RECT 133.795 -223.885 134.125 -223.555 ;
        RECT 133.795 -225.245 134.125 -224.915 ;
        RECT 133.795 -226.605 134.125 -226.275 ;
        RECT 133.795 -227.965 134.125 -227.635 ;
        RECT 133.795 -229.325 134.125 -228.995 ;
        RECT 133.795 -230.685 134.125 -230.355 ;
        RECT 133.795 -232.045 134.125 -231.715 ;
        RECT 133.795 -233.405 134.125 -233.075 ;
        RECT 133.795 -234.765 134.125 -234.435 ;
        RECT 133.795 -236.125 134.125 -235.795 ;
        RECT 133.795 -237.485 134.125 -237.155 ;
        RECT 133.795 -238.845 134.125 -238.515 ;
        RECT 133.795 -241.09 134.125 -239.96 ;
        RECT 133.8 -241.205 134.12 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.11 -125.535 134.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 244.04 135.485 245.17 ;
        RECT 135.155 242.595 135.485 242.925 ;
        RECT 135.155 241.235 135.485 241.565 ;
        RECT 135.155 239.875 135.485 240.205 ;
        RECT 135.155 238.515 135.485 238.845 ;
        RECT 135.155 237.155 135.485 237.485 ;
        RECT 135.16 237.155 135.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 -0.845 135.485 -0.515 ;
        RECT 135.155 -2.205 135.485 -1.875 ;
        RECT 135.155 -3.565 135.485 -3.235 ;
        RECT 135.16 -3.565 135.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 244.04 136.845 245.17 ;
        RECT 136.515 242.595 136.845 242.925 ;
        RECT 136.515 241.235 136.845 241.565 ;
        RECT 136.515 239.875 136.845 240.205 ;
        RECT 136.515 238.515 136.845 238.845 ;
        RECT 136.515 237.155 136.845 237.485 ;
        RECT 136.52 237.155 136.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 -0.845 136.845 -0.515 ;
        RECT 136.515 -2.205 136.845 -1.875 ;
        RECT 136.515 -3.565 136.845 -3.235 ;
        RECT 136.52 -3.565 136.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 244.04 138.205 245.17 ;
        RECT 137.875 242.595 138.205 242.925 ;
        RECT 137.875 241.235 138.205 241.565 ;
        RECT 137.875 239.875 138.205 240.205 ;
        RECT 137.875 238.515 138.205 238.845 ;
        RECT 137.875 237.155 138.205 237.485 ;
        RECT 137.88 237.155 138.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 -0.845 138.205 -0.515 ;
        RECT 137.875 -2.205 138.205 -1.875 ;
        RECT 137.875 -3.565 138.205 -3.235 ;
        RECT 137.88 -3.565 138.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 -123.245 138.205 -122.915 ;
        RECT 137.875 -124.605 138.205 -124.275 ;
        RECT 137.875 -125.965 138.205 -125.635 ;
        RECT 137.875 -127.325 138.205 -126.995 ;
        RECT 137.875 -128.685 138.205 -128.355 ;
        RECT 137.875 -130.045 138.205 -129.715 ;
        RECT 137.875 -131.405 138.205 -131.075 ;
        RECT 137.875 -132.765 138.205 -132.435 ;
        RECT 137.875 -134.125 138.205 -133.795 ;
        RECT 137.875 -135.485 138.205 -135.155 ;
        RECT 137.875 -136.845 138.205 -136.515 ;
        RECT 137.875 -138.205 138.205 -137.875 ;
        RECT 137.875 -139.565 138.205 -139.235 ;
        RECT 137.875 -140.925 138.205 -140.595 ;
        RECT 137.875 -142.285 138.205 -141.955 ;
        RECT 137.875 -143.645 138.205 -143.315 ;
        RECT 137.875 -145.005 138.205 -144.675 ;
        RECT 137.875 -146.365 138.205 -146.035 ;
        RECT 137.875 -147.725 138.205 -147.395 ;
        RECT 137.875 -149.085 138.205 -148.755 ;
        RECT 137.875 -150.445 138.205 -150.115 ;
        RECT 137.875 -151.805 138.205 -151.475 ;
        RECT 137.875 -153.165 138.205 -152.835 ;
        RECT 137.875 -154.525 138.205 -154.195 ;
        RECT 137.875 -155.885 138.205 -155.555 ;
        RECT 137.875 -157.245 138.205 -156.915 ;
        RECT 137.875 -158.605 138.205 -158.275 ;
        RECT 137.875 -159.965 138.205 -159.635 ;
        RECT 137.875 -161.325 138.205 -160.995 ;
        RECT 137.875 -162.685 138.205 -162.355 ;
        RECT 137.875 -164.045 138.205 -163.715 ;
        RECT 137.875 -165.405 138.205 -165.075 ;
        RECT 137.875 -166.765 138.205 -166.435 ;
        RECT 137.875 -168.125 138.205 -167.795 ;
        RECT 137.875 -169.485 138.205 -169.155 ;
        RECT 137.875 -170.845 138.205 -170.515 ;
        RECT 137.875 -172.205 138.205 -171.875 ;
        RECT 137.875 -173.565 138.205 -173.235 ;
        RECT 137.875 -174.925 138.205 -174.595 ;
        RECT 137.875 -176.285 138.205 -175.955 ;
        RECT 137.875 -177.645 138.205 -177.315 ;
        RECT 137.875 -179.005 138.205 -178.675 ;
        RECT 137.875 -180.365 138.205 -180.035 ;
        RECT 137.875 -181.725 138.205 -181.395 ;
        RECT 137.875 -183.085 138.205 -182.755 ;
        RECT 137.875 -184.445 138.205 -184.115 ;
        RECT 137.875 -185.805 138.205 -185.475 ;
        RECT 137.875 -187.165 138.205 -186.835 ;
        RECT 137.875 -188.525 138.205 -188.195 ;
        RECT 137.875 -189.885 138.205 -189.555 ;
        RECT 137.875 -191.245 138.205 -190.915 ;
        RECT 137.875 -192.605 138.205 -192.275 ;
        RECT 137.875 -193.965 138.205 -193.635 ;
        RECT 137.875 -195.325 138.205 -194.995 ;
        RECT 137.875 -196.685 138.205 -196.355 ;
        RECT 137.875 -198.045 138.205 -197.715 ;
        RECT 137.875 -199.405 138.205 -199.075 ;
        RECT 137.875 -200.765 138.205 -200.435 ;
        RECT 137.875 -202.125 138.205 -201.795 ;
        RECT 137.875 -203.485 138.205 -203.155 ;
        RECT 137.875 -204.845 138.205 -204.515 ;
        RECT 137.875 -206.205 138.205 -205.875 ;
        RECT 137.875 -207.565 138.205 -207.235 ;
        RECT 137.875 -208.925 138.205 -208.595 ;
        RECT 137.875 -210.285 138.205 -209.955 ;
        RECT 137.875 -211.645 138.205 -211.315 ;
        RECT 137.875 -213.005 138.205 -212.675 ;
        RECT 137.875 -214.365 138.205 -214.035 ;
        RECT 137.875 -215.725 138.205 -215.395 ;
        RECT 137.875 -217.085 138.205 -216.755 ;
        RECT 137.875 -218.445 138.205 -218.115 ;
        RECT 137.875 -219.805 138.205 -219.475 ;
        RECT 137.875 -221.165 138.205 -220.835 ;
        RECT 137.875 -222.525 138.205 -222.195 ;
        RECT 137.875 -223.885 138.205 -223.555 ;
        RECT 137.875 -225.245 138.205 -224.915 ;
        RECT 137.875 -226.605 138.205 -226.275 ;
        RECT 137.875 -227.965 138.205 -227.635 ;
        RECT 137.875 -229.325 138.205 -228.995 ;
        RECT 137.875 -230.685 138.205 -230.355 ;
        RECT 137.875 -232.045 138.205 -231.715 ;
        RECT 137.875 -233.405 138.205 -233.075 ;
        RECT 137.875 -234.765 138.205 -234.435 ;
        RECT 137.875 -236.125 138.205 -235.795 ;
        RECT 137.875 -237.485 138.205 -237.155 ;
        RECT 137.875 -238.845 138.205 -238.515 ;
        RECT 137.875 -241.09 138.205 -239.96 ;
        RECT 137.88 -241.205 138.2 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 244.04 139.565 245.17 ;
        RECT 139.235 242.595 139.565 242.925 ;
        RECT 139.235 241.235 139.565 241.565 ;
        RECT 139.235 239.875 139.565 240.205 ;
        RECT 139.235 238.515 139.565 238.845 ;
        RECT 139.235 237.155 139.565 237.485 ;
        RECT 139.24 237.155 139.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 -0.845 139.565 -0.515 ;
        RECT 139.235 -2.205 139.565 -1.875 ;
        RECT 139.235 -3.565 139.565 -3.235 ;
        RECT 139.24 -3.565 139.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 -123.245 139.565 -122.915 ;
        RECT 139.235 -124.605 139.565 -124.275 ;
        RECT 139.235 -125.965 139.565 -125.635 ;
        RECT 139.235 -127.325 139.565 -126.995 ;
        RECT 139.235 -128.685 139.565 -128.355 ;
        RECT 139.235 -130.045 139.565 -129.715 ;
        RECT 139.235 -131.405 139.565 -131.075 ;
        RECT 139.235 -132.765 139.565 -132.435 ;
        RECT 139.235 -134.125 139.565 -133.795 ;
        RECT 139.235 -135.485 139.565 -135.155 ;
        RECT 139.235 -136.845 139.565 -136.515 ;
        RECT 139.235 -138.205 139.565 -137.875 ;
        RECT 139.235 -139.565 139.565 -139.235 ;
        RECT 139.235 -140.925 139.565 -140.595 ;
        RECT 139.235 -142.285 139.565 -141.955 ;
        RECT 139.235 -143.645 139.565 -143.315 ;
        RECT 139.235 -145.005 139.565 -144.675 ;
        RECT 139.235 -146.365 139.565 -146.035 ;
        RECT 139.235 -147.725 139.565 -147.395 ;
        RECT 139.235 -149.085 139.565 -148.755 ;
        RECT 139.235 -150.445 139.565 -150.115 ;
        RECT 139.235 -151.805 139.565 -151.475 ;
        RECT 139.235 -153.165 139.565 -152.835 ;
        RECT 139.235 -154.525 139.565 -154.195 ;
        RECT 139.235 -155.885 139.565 -155.555 ;
        RECT 139.235 -157.245 139.565 -156.915 ;
        RECT 139.235 -158.605 139.565 -158.275 ;
        RECT 139.235 -159.965 139.565 -159.635 ;
        RECT 139.235 -161.325 139.565 -160.995 ;
        RECT 139.235 -162.685 139.565 -162.355 ;
        RECT 139.235 -164.045 139.565 -163.715 ;
        RECT 139.235 -165.405 139.565 -165.075 ;
        RECT 139.235 -166.765 139.565 -166.435 ;
        RECT 139.235 -168.125 139.565 -167.795 ;
        RECT 139.235 -169.485 139.565 -169.155 ;
        RECT 139.235 -170.845 139.565 -170.515 ;
        RECT 139.235 -172.205 139.565 -171.875 ;
        RECT 139.235 -173.565 139.565 -173.235 ;
        RECT 139.235 -174.925 139.565 -174.595 ;
        RECT 139.235 -176.285 139.565 -175.955 ;
        RECT 139.235 -177.645 139.565 -177.315 ;
        RECT 139.235 -179.005 139.565 -178.675 ;
        RECT 139.235 -180.365 139.565 -180.035 ;
        RECT 139.235 -181.725 139.565 -181.395 ;
        RECT 139.235 -183.085 139.565 -182.755 ;
        RECT 139.235 -184.445 139.565 -184.115 ;
        RECT 139.235 -185.805 139.565 -185.475 ;
        RECT 139.235 -187.165 139.565 -186.835 ;
        RECT 139.235 -188.525 139.565 -188.195 ;
        RECT 139.235 -189.885 139.565 -189.555 ;
        RECT 139.235 -191.245 139.565 -190.915 ;
        RECT 139.235 -192.605 139.565 -192.275 ;
        RECT 139.235 -193.965 139.565 -193.635 ;
        RECT 139.235 -195.325 139.565 -194.995 ;
        RECT 139.235 -196.685 139.565 -196.355 ;
        RECT 139.235 -198.045 139.565 -197.715 ;
        RECT 139.235 -199.405 139.565 -199.075 ;
        RECT 139.235 -200.765 139.565 -200.435 ;
        RECT 139.235 -202.125 139.565 -201.795 ;
        RECT 139.235 -203.485 139.565 -203.155 ;
        RECT 139.235 -204.845 139.565 -204.515 ;
        RECT 139.235 -206.205 139.565 -205.875 ;
        RECT 139.235 -207.565 139.565 -207.235 ;
        RECT 139.235 -208.925 139.565 -208.595 ;
        RECT 139.235 -210.285 139.565 -209.955 ;
        RECT 139.235 -211.645 139.565 -211.315 ;
        RECT 139.235 -213.005 139.565 -212.675 ;
        RECT 139.235 -214.365 139.565 -214.035 ;
        RECT 139.235 -215.725 139.565 -215.395 ;
        RECT 139.235 -217.085 139.565 -216.755 ;
        RECT 139.235 -218.445 139.565 -218.115 ;
        RECT 139.235 -219.805 139.565 -219.475 ;
        RECT 139.235 -221.165 139.565 -220.835 ;
        RECT 139.235 -222.525 139.565 -222.195 ;
        RECT 139.235 -223.885 139.565 -223.555 ;
        RECT 139.235 -225.245 139.565 -224.915 ;
        RECT 139.235 -226.605 139.565 -226.275 ;
        RECT 139.235 -227.965 139.565 -227.635 ;
        RECT 139.235 -229.325 139.565 -228.995 ;
        RECT 139.235 -230.685 139.565 -230.355 ;
        RECT 139.235 -232.045 139.565 -231.715 ;
        RECT 139.235 -233.405 139.565 -233.075 ;
        RECT 139.235 -234.765 139.565 -234.435 ;
        RECT 139.235 -236.125 139.565 -235.795 ;
        RECT 139.235 -237.485 139.565 -237.155 ;
        RECT 139.235 -238.845 139.565 -238.515 ;
        RECT 139.235 -241.09 139.565 -239.96 ;
        RECT 139.24 -241.205 139.56 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 244.04 140.925 245.17 ;
        RECT 140.595 242.595 140.925 242.925 ;
        RECT 140.595 241.235 140.925 241.565 ;
        RECT 140.595 239.875 140.925 240.205 ;
        RECT 140.595 238.515 140.925 238.845 ;
        RECT 140.595 237.155 140.925 237.485 ;
        RECT 140.6 237.155 140.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -0.845 140.925 -0.515 ;
        RECT 140.595 -2.205 140.925 -1.875 ;
        RECT 140.595 -3.565 140.925 -3.235 ;
        RECT 140.6 -3.565 140.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -123.245 140.925 -122.915 ;
        RECT 140.595 -124.605 140.925 -124.275 ;
        RECT 140.595 -125.965 140.925 -125.635 ;
        RECT 140.595 -127.325 140.925 -126.995 ;
        RECT 140.595 -128.685 140.925 -128.355 ;
        RECT 140.595 -130.045 140.925 -129.715 ;
        RECT 140.595 -131.405 140.925 -131.075 ;
        RECT 140.595 -132.765 140.925 -132.435 ;
        RECT 140.595 -134.125 140.925 -133.795 ;
        RECT 140.595 -135.485 140.925 -135.155 ;
        RECT 140.595 -136.845 140.925 -136.515 ;
        RECT 140.595 -138.205 140.925 -137.875 ;
        RECT 140.595 -139.565 140.925 -139.235 ;
        RECT 140.595 -140.925 140.925 -140.595 ;
        RECT 140.595 -142.285 140.925 -141.955 ;
        RECT 140.595 -143.645 140.925 -143.315 ;
        RECT 140.595 -145.005 140.925 -144.675 ;
        RECT 140.595 -146.365 140.925 -146.035 ;
        RECT 140.595 -147.725 140.925 -147.395 ;
        RECT 140.595 -149.085 140.925 -148.755 ;
        RECT 140.595 -150.445 140.925 -150.115 ;
        RECT 140.595 -151.805 140.925 -151.475 ;
        RECT 140.595 -153.165 140.925 -152.835 ;
        RECT 140.595 -154.525 140.925 -154.195 ;
        RECT 140.595 -155.885 140.925 -155.555 ;
        RECT 140.595 -157.245 140.925 -156.915 ;
        RECT 140.595 -158.605 140.925 -158.275 ;
        RECT 140.595 -159.965 140.925 -159.635 ;
        RECT 140.595 -161.325 140.925 -160.995 ;
        RECT 140.595 -162.685 140.925 -162.355 ;
        RECT 140.595 -164.045 140.925 -163.715 ;
        RECT 140.595 -165.405 140.925 -165.075 ;
        RECT 140.595 -166.765 140.925 -166.435 ;
        RECT 140.595 -168.125 140.925 -167.795 ;
        RECT 140.595 -169.485 140.925 -169.155 ;
        RECT 140.595 -170.845 140.925 -170.515 ;
        RECT 140.595 -172.205 140.925 -171.875 ;
        RECT 140.595 -173.565 140.925 -173.235 ;
        RECT 140.595 -174.925 140.925 -174.595 ;
        RECT 140.595 -176.285 140.925 -175.955 ;
        RECT 140.595 -177.645 140.925 -177.315 ;
        RECT 140.595 -179.005 140.925 -178.675 ;
        RECT 140.595 -180.365 140.925 -180.035 ;
        RECT 140.595 -181.725 140.925 -181.395 ;
        RECT 140.595 -183.085 140.925 -182.755 ;
        RECT 140.595 -184.445 140.925 -184.115 ;
        RECT 140.595 -185.805 140.925 -185.475 ;
        RECT 140.595 -187.165 140.925 -186.835 ;
        RECT 140.595 -188.525 140.925 -188.195 ;
        RECT 140.595 -189.885 140.925 -189.555 ;
        RECT 140.595 -191.245 140.925 -190.915 ;
        RECT 140.595 -192.605 140.925 -192.275 ;
        RECT 140.595 -193.965 140.925 -193.635 ;
        RECT 140.595 -195.325 140.925 -194.995 ;
        RECT 140.595 -196.685 140.925 -196.355 ;
        RECT 140.595 -198.045 140.925 -197.715 ;
        RECT 140.595 -199.405 140.925 -199.075 ;
        RECT 140.595 -200.765 140.925 -200.435 ;
        RECT 140.595 -202.125 140.925 -201.795 ;
        RECT 140.595 -203.485 140.925 -203.155 ;
        RECT 140.595 -204.845 140.925 -204.515 ;
        RECT 140.595 -206.205 140.925 -205.875 ;
        RECT 140.595 -207.565 140.925 -207.235 ;
        RECT 140.595 -208.925 140.925 -208.595 ;
        RECT 140.595 -210.285 140.925 -209.955 ;
        RECT 140.595 -211.645 140.925 -211.315 ;
        RECT 140.595 -213.005 140.925 -212.675 ;
        RECT 140.595 -214.365 140.925 -214.035 ;
        RECT 140.595 -215.725 140.925 -215.395 ;
        RECT 140.595 -217.085 140.925 -216.755 ;
        RECT 140.595 -218.445 140.925 -218.115 ;
        RECT 140.595 -219.805 140.925 -219.475 ;
        RECT 140.595 -221.165 140.925 -220.835 ;
        RECT 140.595 -222.525 140.925 -222.195 ;
        RECT 140.595 -223.885 140.925 -223.555 ;
        RECT 140.595 -225.245 140.925 -224.915 ;
        RECT 140.595 -226.605 140.925 -226.275 ;
        RECT 140.595 -227.965 140.925 -227.635 ;
        RECT 140.595 -229.325 140.925 -228.995 ;
        RECT 140.595 -230.685 140.925 -230.355 ;
        RECT 140.595 -232.045 140.925 -231.715 ;
        RECT 140.595 -233.405 140.925 -233.075 ;
        RECT 140.595 -234.765 140.925 -234.435 ;
        RECT 140.595 -236.125 140.925 -235.795 ;
        RECT 140.595 -237.485 140.925 -237.155 ;
        RECT 140.595 -238.845 140.925 -238.515 ;
        RECT 140.595 -241.09 140.925 -239.96 ;
        RECT 140.6 -241.205 140.92 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 244.04 142.285 245.17 ;
        RECT 141.955 242.595 142.285 242.925 ;
        RECT 141.955 241.235 142.285 241.565 ;
        RECT 141.955 239.875 142.285 240.205 ;
        RECT 141.955 238.515 142.285 238.845 ;
        RECT 141.955 237.155 142.285 237.485 ;
        RECT 141.96 237.155 142.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -0.845 142.285 -0.515 ;
        RECT 141.955 -2.205 142.285 -1.875 ;
        RECT 141.955 -3.565 142.285 -3.235 ;
        RECT 141.96 -3.565 142.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -123.245 142.285 -122.915 ;
        RECT 141.955 -124.605 142.285 -124.275 ;
        RECT 141.955 -125.965 142.285 -125.635 ;
        RECT 141.955 -127.325 142.285 -126.995 ;
        RECT 141.955 -128.685 142.285 -128.355 ;
        RECT 141.955 -130.045 142.285 -129.715 ;
        RECT 141.955 -131.405 142.285 -131.075 ;
        RECT 141.955 -132.765 142.285 -132.435 ;
        RECT 141.955 -134.125 142.285 -133.795 ;
        RECT 141.955 -135.485 142.285 -135.155 ;
        RECT 141.955 -136.845 142.285 -136.515 ;
        RECT 141.955 -138.205 142.285 -137.875 ;
        RECT 141.955 -139.565 142.285 -139.235 ;
        RECT 141.955 -140.925 142.285 -140.595 ;
        RECT 141.955 -142.285 142.285 -141.955 ;
        RECT 141.955 -143.645 142.285 -143.315 ;
        RECT 141.955 -145.005 142.285 -144.675 ;
        RECT 141.955 -146.365 142.285 -146.035 ;
        RECT 141.955 -147.725 142.285 -147.395 ;
        RECT 141.955 -149.085 142.285 -148.755 ;
        RECT 141.955 -150.445 142.285 -150.115 ;
        RECT 141.955 -151.805 142.285 -151.475 ;
        RECT 141.955 -153.165 142.285 -152.835 ;
        RECT 141.955 -154.525 142.285 -154.195 ;
        RECT 141.955 -155.885 142.285 -155.555 ;
        RECT 141.955 -157.245 142.285 -156.915 ;
        RECT 141.955 -158.605 142.285 -158.275 ;
        RECT 141.955 -159.965 142.285 -159.635 ;
        RECT 141.955 -161.325 142.285 -160.995 ;
        RECT 141.955 -162.685 142.285 -162.355 ;
        RECT 141.955 -164.045 142.285 -163.715 ;
        RECT 141.955 -165.405 142.285 -165.075 ;
        RECT 141.955 -166.765 142.285 -166.435 ;
        RECT 141.955 -168.125 142.285 -167.795 ;
        RECT 141.955 -169.485 142.285 -169.155 ;
        RECT 141.955 -170.845 142.285 -170.515 ;
        RECT 141.955 -172.205 142.285 -171.875 ;
        RECT 141.955 -173.565 142.285 -173.235 ;
        RECT 141.955 -174.925 142.285 -174.595 ;
        RECT 141.955 -176.285 142.285 -175.955 ;
        RECT 141.955 -177.645 142.285 -177.315 ;
        RECT 141.955 -179.005 142.285 -178.675 ;
        RECT 141.955 -180.365 142.285 -180.035 ;
        RECT 141.955 -181.725 142.285 -181.395 ;
        RECT 141.955 -183.085 142.285 -182.755 ;
        RECT 141.955 -184.445 142.285 -184.115 ;
        RECT 141.955 -185.805 142.285 -185.475 ;
        RECT 141.955 -187.165 142.285 -186.835 ;
        RECT 141.955 -188.525 142.285 -188.195 ;
        RECT 141.955 -189.885 142.285 -189.555 ;
        RECT 141.955 -191.245 142.285 -190.915 ;
        RECT 141.955 -192.605 142.285 -192.275 ;
        RECT 141.955 -193.965 142.285 -193.635 ;
        RECT 141.955 -195.325 142.285 -194.995 ;
        RECT 141.955 -196.685 142.285 -196.355 ;
        RECT 141.955 -198.045 142.285 -197.715 ;
        RECT 141.955 -199.405 142.285 -199.075 ;
        RECT 141.955 -200.765 142.285 -200.435 ;
        RECT 141.955 -202.125 142.285 -201.795 ;
        RECT 141.955 -203.485 142.285 -203.155 ;
        RECT 141.955 -204.845 142.285 -204.515 ;
        RECT 141.955 -206.205 142.285 -205.875 ;
        RECT 141.955 -207.565 142.285 -207.235 ;
        RECT 141.955 -208.925 142.285 -208.595 ;
        RECT 141.955 -210.285 142.285 -209.955 ;
        RECT 141.955 -211.645 142.285 -211.315 ;
        RECT 141.955 -213.005 142.285 -212.675 ;
        RECT 141.955 -214.365 142.285 -214.035 ;
        RECT 141.955 -215.725 142.285 -215.395 ;
        RECT 141.955 -217.085 142.285 -216.755 ;
        RECT 141.955 -218.445 142.285 -218.115 ;
        RECT 141.955 -219.805 142.285 -219.475 ;
        RECT 141.955 -221.165 142.285 -220.835 ;
        RECT 141.955 -222.525 142.285 -222.195 ;
        RECT 141.955 -223.885 142.285 -223.555 ;
        RECT 141.955 -225.245 142.285 -224.915 ;
        RECT 141.955 -226.605 142.285 -226.275 ;
        RECT 141.955 -227.965 142.285 -227.635 ;
        RECT 141.955 -229.325 142.285 -228.995 ;
        RECT 141.955 -230.685 142.285 -230.355 ;
        RECT 141.955 -232.045 142.285 -231.715 ;
        RECT 141.955 -233.405 142.285 -233.075 ;
        RECT 141.955 -234.765 142.285 -234.435 ;
        RECT 141.955 -236.125 142.285 -235.795 ;
        RECT 141.955 -237.485 142.285 -237.155 ;
        RECT 141.955 -238.845 142.285 -238.515 ;
        RECT 141.955 -241.09 142.285 -239.96 ;
        RECT 141.96 -241.205 142.28 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 244.04 143.645 245.17 ;
        RECT 143.315 242.595 143.645 242.925 ;
        RECT 143.315 241.235 143.645 241.565 ;
        RECT 143.315 239.875 143.645 240.205 ;
        RECT 143.315 238.515 143.645 238.845 ;
        RECT 143.315 237.155 143.645 237.485 ;
        RECT 143.32 237.155 143.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 -0.845 143.645 -0.515 ;
        RECT 143.315 -2.205 143.645 -1.875 ;
        RECT 143.315 -3.565 143.645 -3.235 ;
        RECT 143.32 -3.565 143.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 -123.245 143.645 -122.915 ;
        RECT 143.315 -124.605 143.645 -124.275 ;
        RECT 143.315 -125.965 143.645 -125.635 ;
        RECT 143.315 -127.325 143.645 -126.995 ;
        RECT 143.315 -128.685 143.645 -128.355 ;
        RECT 143.315 -130.045 143.645 -129.715 ;
        RECT 143.315 -131.405 143.645 -131.075 ;
        RECT 143.315 -132.765 143.645 -132.435 ;
        RECT 143.315 -134.125 143.645 -133.795 ;
        RECT 143.315 -135.485 143.645 -135.155 ;
        RECT 143.315 -136.845 143.645 -136.515 ;
        RECT 143.315 -138.205 143.645 -137.875 ;
        RECT 143.315 -139.565 143.645 -139.235 ;
        RECT 143.315 -140.925 143.645 -140.595 ;
        RECT 143.315 -142.285 143.645 -141.955 ;
        RECT 143.315 -143.645 143.645 -143.315 ;
        RECT 143.315 -145.005 143.645 -144.675 ;
        RECT 143.315 -146.365 143.645 -146.035 ;
        RECT 143.315 -147.725 143.645 -147.395 ;
        RECT 143.315 -149.085 143.645 -148.755 ;
        RECT 143.315 -150.445 143.645 -150.115 ;
        RECT 143.315 -151.805 143.645 -151.475 ;
        RECT 143.315 -153.165 143.645 -152.835 ;
        RECT 143.315 -154.525 143.645 -154.195 ;
        RECT 143.315 -155.885 143.645 -155.555 ;
        RECT 143.315 -157.245 143.645 -156.915 ;
        RECT 143.315 -158.605 143.645 -158.275 ;
        RECT 143.315 -159.965 143.645 -159.635 ;
        RECT 143.315 -161.325 143.645 -160.995 ;
        RECT 143.315 -162.685 143.645 -162.355 ;
        RECT 143.315 -164.045 143.645 -163.715 ;
        RECT 143.315 -165.405 143.645 -165.075 ;
        RECT 143.315 -166.765 143.645 -166.435 ;
        RECT 143.315 -168.125 143.645 -167.795 ;
        RECT 143.315 -169.485 143.645 -169.155 ;
        RECT 143.315 -170.845 143.645 -170.515 ;
        RECT 143.315 -172.205 143.645 -171.875 ;
        RECT 143.315 -173.565 143.645 -173.235 ;
        RECT 143.315 -174.925 143.645 -174.595 ;
        RECT 143.315 -176.285 143.645 -175.955 ;
        RECT 143.315 -177.645 143.645 -177.315 ;
        RECT 143.315 -179.005 143.645 -178.675 ;
        RECT 143.315 -180.365 143.645 -180.035 ;
        RECT 143.315 -181.725 143.645 -181.395 ;
        RECT 143.315 -183.085 143.645 -182.755 ;
        RECT 143.315 -184.445 143.645 -184.115 ;
        RECT 143.315 -185.805 143.645 -185.475 ;
        RECT 143.315 -187.165 143.645 -186.835 ;
        RECT 143.315 -188.525 143.645 -188.195 ;
        RECT 143.315 -189.885 143.645 -189.555 ;
        RECT 143.315 -191.245 143.645 -190.915 ;
        RECT 143.315 -192.605 143.645 -192.275 ;
        RECT 143.315 -193.965 143.645 -193.635 ;
        RECT 143.315 -195.325 143.645 -194.995 ;
        RECT 143.315 -196.685 143.645 -196.355 ;
        RECT 143.315 -198.045 143.645 -197.715 ;
        RECT 143.315 -199.405 143.645 -199.075 ;
        RECT 143.315 -200.765 143.645 -200.435 ;
        RECT 143.315 -202.125 143.645 -201.795 ;
        RECT 143.315 -203.485 143.645 -203.155 ;
        RECT 143.315 -204.845 143.645 -204.515 ;
        RECT 143.315 -206.205 143.645 -205.875 ;
        RECT 143.315 -207.565 143.645 -207.235 ;
        RECT 143.315 -208.925 143.645 -208.595 ;
        RECT 143.315 -210.285 143.645 -209.955 ;
        RECT 143.315 -211.645 143.645 -211.315 ;
        RECT 143.315 -213.005 143.645 -212.675 ;
        RECT 143.315 -214.365 143.645 -214.035 ;
        RECT 143.315 -215.725 143.645 -215.395 ;
        RECT 143.315 -217.085 143.645 -216.755 ;
        RECT 143.315 -218.445 143.645 -218.115 ;
        RECT 143.315 -219.805 143.645 -219.475 ;
        RECT 143.315 -221.165 143.645 -220.835 ;
        RECT 143.315 -222.525 143.645 -222.195 ;
        RECT 143.315 -223.885 143.645 -223.555 ;
        RECT 143.315 -225.245 143.645 -224.915 ;
        RECT 143.315 -226.605 143.645 -226.275 ;
        RECT 143.315 -227.965 143.645 -227.635 ;
        RECT 143.315 -229.325 143.645 -228.995 ;
        RECT 143.315 -230.685 143.645 -230.355 ;
        RECT 143.315 -232.045 143.645 -231.715 ;
        RECT 143.315 -233.405 143.645 -233.075 ;
        RECT 143.315 -234.765 143.645 -234.435 ;
        RECT 143.315 -236.125 143.645 -235.795 ;
        RECT 143.315 -237.485 143.645 -237.155 ;
        RECT 143.315 -238.845 143.645 -238.515 ;
        RECT 143.315 -241.09 143.645 -239.96 ;
        RECT 143.32 -241.205 143.64 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 244.04 145.005 245.17 ;
        RECT 144.675 242.595 145.005 242.925 ;
        RECT 144.675 241.235 145.005 241.565 ;
        RECT 144.675 239.875 145.005 240.205 ;
        RECT 144.675 238.515 145.005 238.845 ;
        RECT 144.675 237.155 145.005 237.485 ;
        RECT 144.68 237.155 145 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 -127.325 145.005 -126.995 ;
        RECT 144.675 -128.685 145.005 -128.355 ;
        RECT 144.675 -130.045 145.005 -129.715 ;
        RECT 144.675 -131.405 145.005 -131.075 ;
        RECT 144.675 -132.765 145.005 -132.435 ;
        RECT 144.675 -134.125 145.005 -133.795 ;
        RECT 144.675 -135.485 145.005 -135.155 ;
        RECT 144.675 -136.845 145.005 -136.515 ;
        RECT 144.675 -138.205 145.005 -137.875 ;
        RECT 144.675 -139.565 145.005 -139.235 ;
        RECT 144.675 -140.925 145.005 -140.595 ;
        RECT 144.675 -142.285 145.005 -141.955 ;
        RECT 144.675 -143.645 145.005 -143.315 ;
        RECT 144.675 -145.005 145.005 -144.675 ;
        RECT 144.675 -146.365 145.005 -146.035 ;
        RECT 144.675 -147.725 145.005 -147.395 ;
        RECT 144.675 -149.085 145.005 -148.755 ;
        RECT 144.675 -150.445 145.005 -150.115 ;
        RECT 144.675 -151.805 145.005 -151.475 ;
        RECT 144.675 -153.165 145.005 -152.835 ;
        RECT 144.675 -154.525 145.005 -154.195 ;
        RECT 144.675 -155.885 145.005 -155.555 ;
        RECT 144.675 -157.245 145.005 -156.915 ;
        RECT 144.675 -158.605 145.005 -158.275 ;
        RECT 144.675 -159.965 145.005 -159.635 ;
        RECT 144.675 -161.325 145.005 -160.995 ;
        RECT 144.675 -162.685 145.005 -162.355 ;
        RECT 144.675 -164.045 145.005 -163.715 ;
        RECT 144.675 -165.405 145.005 -165.075 ;
        RECT 144.675 -166.765 145.005 -166.435 ;
        RECT 144.675 -168.125 145.005 -167.795 ;
        RECT 144.675 -169.485 145.005 -169.155 ;
        RECT 144.675 -170.845 145.005 -170.515 ;
        RECT 144.675 -172.205 145.005 -171.875 ;
        RECT 144.675 -173.565 145.005 -173.235 ;
        RECT 144.675 -174.925 145.005 -174.595 ;
        RECT 144.675 -176.285 145.005 -175.955 ;
        RECT 144.675 -177.645 145.005 -177.315 ;
        RECT 144.675 -179.005 145.005 -178.675 ;
        RECT 144.675 -180.365 145.005 -180.035 ;
        RECT 144.675 -181.725 145.005 -181.395 ;
        RECT 144.675 -183.085 145.005 -182.755 ;
        RECT 144.675 -184.445 145.005 -184.115 ;
        RECT 144.675 -185.805 145.005 -185.475 ;
        RECT 144.675 -187.165 145.005 -186.835 ;
        RECT 144.675 -188.525 145.005 -188.195 ;
        RECT 144.675 -189.885 145.005 -189.555 ;
        RECT 144.675 -191.245 145.005 -190.915 ;
        RECT 144.675 -192.605 145.005 -192.275 ;
        RECT 144.675 -193.965 145.005 -193.635 ;
        RECT 144.675 -195.325 145.005 -194.995 ;
        RECT 144.675 -196.685 145.005 -196.355 ;
        RECT 144.675 -198.045 145.005 -197.715 ;
        RECT 144.675 -199.405 145.005 -199.075 ;
        RECT 144.675 -200.765 145.005 -200.435 ;
        RECT 144.675 -202.125 145.005 -201.795 ;
        RECT 144.675 -203.485 145.005 -203.155 ;
        RECT 144.675 -204.845 145.005 -204.515 ;
        RECT 144.675 -206.205 145.005 -205.875 ;
        RECT 144.675 -207.565 145.005 -207.235 ;
        RECT 144.675 -208.925 145.005 -208.595 ;
        RECT 144.675 -210.285 145.005 -209.955 ;
        RECT 144.675 -211.645 145.005 -211.315 ;
        RECT 144.675 -213.005 145.005 -212.675 ;
        RECT 144.675 -214.365 145.005 -214.035 ;
        RECT 144.675 -215.725 145.005 -215.395 ;
        RECT 144.675 -217.085 145.005 -216.755 ;
        RECT 144.675 -218.445 145.005 -218.115 ;
        RECT 144.675 -219.805 145.005 -219.475 ;
        RECT 144.675 -221.165 145.005 -220.835 ;
        RECT 144.675 -222.525 145.005 -222.195 ;
        RECT 144.675 -223.885 145.005 -223.555 ;
        RECT 144.675 -225.245 145.005 -224.915 ;
        RECT 144.675 -226.605 145.005 -226.275 ;
        RECT 144.675 -227.965 145.005 -227.635 ;
        RECT 144.675 -229.325 145.005 -228.995 ;
        RECT 144.675 -230.685 145.005 -230.355 ;
        RECT 144.675 -232.045 145.005 -231.715 ;
        RECT 144.675 -233.405 145.005 -233.075 ;
        RECT 144.675 -234.765 145.005 -234.435 ;
        RECT 144.675 -236.125 145.005 -235.795 ;
        RECT 144.675 -237.485 145.005 -237.155 ;
        RECT 144.675 -238.845 145.005 -238.515 ;
        RECT 144.675 -241.09 145.005 -239.96 ;
        RECT 144.68 -241.205 145 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.01 -125.535 145.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 244.04 146.365 245.17 ;
        RECT 146.035 242.595 146.365 242.925 ;
        RECT 146.035 241.235 146.365 241.565 ;
        RECT 146.035 239.875 146.365 240.205 ;
        RECT 146.035 238.515 146.365 238.845 ;
        RECT 146.035 237.155 146.365 237.485 ;
        RECT 146.04 237.155 146.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 -3.565 146.365 -3.235 ;
        RECT 146.04 -3.565 146.36 -0.515 ;
        RECT 146.035 -0.845 146.365 -0.515 ;
        RECT 146.035 -2.205 146.365 -1.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 244.04 112.365 245.17 ;
        RECT 112.035 242.595 112.365 242.925 ;
        RECT 112.035 241.235 112.365 241.565 ;
        RECT 112.035 239.875 112.365 240.205 ;
        RECT 112.035 238.515 112.365 238.845 ;
        RECT 112.035 237.155 112.365 237.485 ;
        RECT 112.04 237.155 112.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 -127.325 112.365 -126.995 ;
        RECT 112.035 -128.685 112.365 -128.355 ;
        RECT 112.035 -130.045 112.365 -129.715 ;
        RECT 112.035 -131.405 112.365 -131.075 ;
        RECT 112.035 -132.765 112.365 -132.435 ;
        RECT 112.035 -134.125 112.365 -133.795 ;
        RECT 112.035 -135.485 112.365 -135.155 ;
        RECT 112.035 -136.845 112.365 -136.515 ;
        RECT 112.035 -138.205 112.365 -137.875 ;
        RECT 112.035 -139.565 112.365 -139.235 ;
        RECT 112.035 -140.925 112.365 -140.595 ;
        RECT 112.035 -142.285 112.365 -141.955 ;
        RECT 112.035 -143.645 112.365 -143.315 ;
        RECT 112.035 -145.005 112.365 -144.675 ;
        RECT 112.035 -146.365 112.365 -146.035 ;
        RECT 112.035 -147.725 112.365 -147.395 ;
        RECT 112.035 -149.085 112.365 -148.755 ;
        RECT 112.035 -150.445 112.365 -150.115 ;
        RECT 112.035 -151.805 112.365 -151.475 ;
        RECT 112.035 -153.165 112.365 -152.835 ;
        RECT 112.035 -154.525 112.365 -154.195 ;
        RECT 112.035 -155.885 112.365 -155.555 ;
        RECT 112.035 -157.245 112.365 -156.915 ;
        RECT 112.035 -158.605 112.365 -158.275 ;
        RECT 112.035 -159.965 112.365 -159.635 ;
        RECT 112.035 -161.325 112.365 -160.995 ;
        RECT 112.035 -162.685 112.365 -162.355 ;
        RECT 112.035 -164.045 112.365 -163.715 ;
        RECT 112.035 -165.405 112.365 -165.075 ;
        RECT 112.035 -166.765 112.365 -166.435 ;
        RECT 112.035 -168.125 112.365 -167.795 ;
        RECT 112.035 -169.485 112.365 -169.155 ;
        RECT 112.035 -170.845 112.365 -170.515 ;
        RECT 112.035 -172.205 112.365 -171.875 ;
        RECT 112.035 -173.565 112.365 -173.235 ;
        RECT 112.035 -174.925 112.365 -174.595 ;
        RECT 112.035 -176.285 112.365 -175.955 ;
        RECT 112.035 -177.645 112.365 -177.315 ;
        RECT 112.035 -179.005 112.365 -178.675 ;
        RECT 112.035 -180.365 112.365 -180.035 ;
        RECT 112.035 -181.725 112.365 -181.395 ;
        RECT 112.035 -183.085 112.365 -182.755 ;
        RECT 112.035 -184.445 112.365 -184.115 ;
        RECT 112.035 -185.805 112.365 -185.475 ;
        RECT 112.035 -187.165 112.365 -186.835 ;
        RECT 112.035 -188.525 112.365 -188.195 ;
        RECT 112.035 -189.885 112.365 -189.555 ;
        RECT 112.035 -191.245 112.365 -190.915 ;
        RECT 112.035 -192.605 112.365 -192.275 ;
        RECT 112.035 -193.965 112.365 -193.635 ;
        RECT 112.035 -195.325 112.365 -194.995 ;
        RECT 112.035 -196.685 112.365 -196.355 ;
        RECT 112.035 -198.045 112.365 -197.715 ;
        RECT 112.035 -199.405 112.365 -199.075 ;
        RECT 112.035 -200.765 112.365 -200.435 ;
        RECT 112.035 -202.125 112.365 -201.795 ;
        RECT 112.035 -203.485 112.365 -203.155 ;
        RECT 112.035 -204.845 112.365 -204.515 ;
        RECT 112.035 -206.205 112.365 -205.875 ;
        RECT 112.035 -207.565 112.365 -207.235 ;
        RECT 112.035 -208.925 112.365 -208.595 ;
        RECT 112.035 -210.285 112.365 -209.955 ;
        RECT 112.035 -211.645 112.365 -211.315 ;
        RECT 112.035 -213.005 112.365 -212.675 ;
        RECT 112.035 -214.365 112.365 -214.035 ;
        RECT 112.035 -215.725 112.365 -215.395 ;
        RECT 112.035 -217.085 112.365 -216.755 ;
        RECT 112.035 -218.445 112.365 -218.115 ;
        RECT 112.035 -219.805 112.365 -219.475 ;
        RECT 112.035 -221.165 112.365 -220.835 ;
        RECT 112.035 -222.525 112.365 -222.195 ;
        RECT 112.035 -223.885 112.365 -223.555 ;
        RECT 112.035 -225.245 112.365 -224.915 ;
        RECT 112.035 -226.605 112.365 -226.275 ;
        RECT 112.035 -227.965 112.365 -227.635 ;
        RECT 112.035 -229.325 112.365 -228.995 ;
        RECT 112.035 -230.685 112.365 -230.355 ;
        RECT 112.035 -232.045 112.365 -231.715 ;
        RECT 112.035 -233.405 112.365 -233.075 ;
        RECT 112.035 -234.765 112.365 -234.435 ;
        RECT 112.035 -236.125 112.365 -235.795 ;
        RECT 112.035 -237.485 112.365 -237.155 ;
        RECT 112.035 -238.845 112.365 -238.515 ;
        RECT 112.035 -241.09 112.365 -239.96 ;
        RECT 112.04 -241.205 112.36 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.31 -125.535 112.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 244.04 113.725 245.17 ;
        RECT 113.395 242.595 113.725 242.925 ;
        RECT 113.395 241.235 113.725 241.565 ;
        RECT 113.395 239.875 113.725 240.205 ;
        RECT 113.395 238.515 113.725 238.845 ;
        RECT 113.395 237.155 113.725 237.485 ;
        RECT 113.4 237.155 113.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 -0.845 113.725 -0.515 ;
        RECT 113.395 -2.205 113.725 -1.875 ;
        RECT 113.395 -3.565 113.725 -3.235 ;
        RECT 113.4 -3.565 113.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 244.04 115.085 245.17 ;
        RECT 114.755 242.595 115.085 242.925 ;
        RECT 114.755 241.235 115.085 241.565 ;
        RECT 114.755 239.875 115.085 240.205 ;
        RECT 114.755 238.515 115.085 238.845 ;
        RECT 114.755 237.155 115.085 237.485 ;
        RECT 114.76 237.155 115.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 -0.845 115.085 -0.515 ;
        RECT 114.755 -2.205 115.085 -1.875 ;
        RECT 114.755 -3.565 115.085 -3.235 ;
        RECT 114.76 -3.565 115.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 244.04 116.445 245.17 ;
        RECT 116.115 242.595 116.445 242.925 ;
        RECT 116.115 241.235 116.445 241.565 ;
        RECT 116.115 239.875 116.445 240.205 ;
        RECT 116.115 238.515 116.445 238.845 ;
        RECT 116.115 237.155 116.445 237.485 ;
        RECT 116.12 237.155 116.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 -0.845 116.445 -0.515 ;
        RECT 116.115 -2.205 116.445 -1.875 ;
        RECT 116.115 -3.565 116.445 -3.235 ;
        RECT 116.12 -3.565 116.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 -123.245 116.445 -122.915 ;
        RECT 116.115 -124.605 116.445 -124.275 ;
        RECT 116.115 -125.965 116.445 -125.635 ;
        RECT 116.115 -127.325 116.445 -126.995 ;
        RECT 116.115 -128.685 116.445 -128.355 ;
        RECT 116.115 -130.045 116.445 -129.715 ;
        RECT 116.115 -131.405 116.445 -131.075 ;
        RECT 116.115 -132.765 116.445 -132.435 ;
        RECT 116.115 -134.125 116.445 -133.795 ;
        RECT 116.115 -135.485 116.445 -135.155 ;
        RECT 116.115 -136.845 116.445 -136.515 ;
        RECT 116.115 -138.205 116.445 -137.875 ;
        RECT 116.115 -139.565 116.445 -139.235 ;
        RECT 116.115 -140.925 116.445 -140.595 ;
        RECT 116.115 -142.285 116.445 -141.955 ;
        RECT 116.115 -143.645 116.445 -143.315 ;
        RECT 116.115 -145.005 116.445 -144.675 ;
        RECT 116.115 -146.365 116.445 -146.035 ;
        RECT 116.115 -147.725 116.445 -147.395 ;
        RECT 116.115 -149.085 116.445 -148.755 ;
        RECT 116.115 -150.445 116.445 -150.115 ;
        RECT 116.115 -151.805 116.445 -151.475 ;
        RECT 116.115 -153.165 116.445 -152.835 ;
        RECT 116.115 -154.525 116.445 -154.195 ;
        RECT 116.115 -155.885 116.445 -155.555 ;
        RECT 116.115 -157.245 116.445 -156.915 ;
        RECT 116.115 -158.605 116.445 -158.275 ;
        RECT 116.115 -159.965 116.445 -159.635 ;
        RECT 116.115 -161.325 116.445 -160.995 ;
        RECT 116.115 -162.685 116.445 -162.355 ;
        RECT 116.115 -164.045 116.445 -163.715 ;
        RECT 116.115 -165.405 116.445 -165.075 ;
        RECT 116.115 -166.765 116.445 -166.435 ;
        RECT 116.115 -168.125 116.445 -167.795 ;
        RECT 116.115 -169.485 116.445 -169.155 ;
        RECT 116.115 -170.845 116.445 -170.515 ;
        RECT 116.115 -172.205 116.445 -171.875 ;
        RECT 116.115 -173.565 116.445 -173.235 ;
        RECT 116.115 -174.925 116.445 -174.595 ;
        RECT 116.115 -176.285 116.445 -175.955 ;
        RECT 116.115 -177.645 116.445 -177.315 ;
        RECT 116.115 -179.005 116.445 -178.675 ;
        RECT 116.115 -180.365 116.445 -180.035 ;
        RECT 116.115 -181.725 116.445 -181.395 ;
        RECT 116.115 -183.085 116.445 -182.755 ;
        RECT 116.115 -184.445 116.445 -184.115 ;
        RECT 116.115 -185.805 116.445 -185.475 ;
        RECT 116.115 -187.165 116.445 -186.835 ;
        RECT 116.115 -188.525 116.445 -188.195 ;
        RECT 116.115 -189.885 116.445 -189.555 ;
        RECT 116.115 -191.245 116.445 -190.915 ;
        RECT 116.115 -192.605 116.445 -192.275 ;
        RECT 116.115 -193.965 116.445 -193.635 ;
        RECT 116.115 -195.325 116.445 -194.995 ;
        RECT 116.115 -196.685 116.445 -196.355 ;
        RECT 116.115 -198.045 116.445 -197.715 ;
        RECT 116.115 -199.405 116.445 -199.075 ;
        RECT 116.115 -200.765 116.445 -200.435 ;
        RECT 116.115 -202.125 116.445 -201.795 ;
        RECT 116.115 -203.485 116.445 -203.155 ;
        RECT 116.115 -204.845 116.445 -204.515 ;
        RECT 116.115 -206.205 116.445 -205.875 ;
        RECT 116.115 -207.565 116.445 -207.235 ;
        RECT 116.115 -208.925 116.445 -208.595 ;
        RECT 116.115 -210.285 116.445 -209.955 ;
        RECT 116.115 -211.645 116.445 -211.315 ;
        RECT 116.115 -213.005 116.445 -212.675 ;
        RECT 116.115 -214.365 116.445 -214.035 ;
        RECT 116.115 -215.725 116.445 -215.395 ;
        RECT 116.115 -217.085 116.445 -216.755 ;
        RECT 116.115 -218.445 116.445 -218.115 ;
        RECT 116.115 -219.805 116.445 -219.475 ;
        RECT 116.115 -221.165 116.445 -220.835 ;
        RECT 116.115 -222.525 116.445 -222.195 ;
        RECT 116.115 -223.885 116.445 -223.555 ;
        RECT 116.115 -225.245 116.445 -224.915 ;
        RECT 116.115 -226.605 116.445 -226.275 ;
        RECT 116.115 -227.965 116.445 -227.635 ;
        RECT 116.115 -229.325 116.445 -228.995 ;
        RECT 116.115 -230.685 116.445 -230.355 ;
        RECT 116.115 -232.045 116.445 -231.715 ;
        RECT 116.115 -233.405 116.445 -233.075 ;
        RECT 116.115 -234.765 116.445 -234.435 ;
        RECT 116.115 -236.125 116.445 -235.795 ;
        RECT 116.115 -237.485 116.445 -237.155 ;
        RECT 116.115 -238.845 116.445 -238.515 ;
        RECT 116.115 -241.09 116.445 -239.96 ;
        RECT 116.12 -241.205 116.44 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 244.04 117.805 245.17 ;
        RECT 117.475 242.595 117.805 242.925 ;
        RECT 117.475 241.235 117.805 241.565 ;
        RECT 117.475 239.875 117.805 240.205 ;
        RECT 117.475 238.515 117.805 238.845 ;
        RECT 117.475 237.155 117.805 237.485 ;
        RECT 117.48 237.155 117.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -0.845 117.805 -0.515 ;
        RECT 117.475 -2.205 117.805 -1.875 ;
        RECT 117.475 -3.565 117.805 -3.235 ;
        RECT 117.48 -3.565 117.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -123.245 117.805 -122.915 ;
        RECT 117.475 -124.605 117.805 -124.275 ;
        RECT 117.475 -125.965 117.805 -125.635 ;
        RECT 117.475 -127.325 117.805 -126.995 ;
        RECT 117.475 -128.685 117.805 -128.355 ;
        RECT 117.475 -130.045 117.805 -129.715 ;
        RECT 117.475 -131.405 117.805 -131.075 ;
        RECT 117.475 -132.765 117.805 -132.435 ;
        RECT 117.475 -134.125 117.805 -133.795 ;
        RECT 117.475 -135.485 117.805 -135.155 ;
        RECT 117.475 -136.845 117.805 -136.515 ;
        RECT 117.475 -138.205 117.805 -137.875 ;
        RECT 117.475 -139.565 117.805 -139.235 ;
        RECT 117.475 -140.925 117.805 -140.595 ;
        RECT 117.475 -142.285 117.805 -141.955 ;
        RECT 117.475 -143.645 117.805 -143.315 ;
        RECT 117.475 -145.005 117.805 -144.675 ;
        RECT 117.475 -146.365 117.805 -146.035 ;
        RECT 117.475 -147.725 117.805 -147.395 ;
        RECT 117.475 -149.085 117.805 -148.755 ;
        RECT 117.475 -150.445 117.805 -150.115 ;
        RECT 117.475 -151.805 117.805 -151.475 ;
        RECT 117.475 -153.165 117.805 -152.835 ;
        RECT 117.475 -154.525 117.805 -154.195 ;
        RECT 117.475 -155.885 117.805 -155.555 ;
        RECT 117.475 -157.245 117.805 -156.915 ;
        RECT 117.475 -158.605 117.805 -158.275 ;
        RECT 117.475 -159.965 117.805 -159.635 ;
        RECT 117.475 -161.325 117.805 -160.995 ;
        RECT 117.475 -162.685 117.805 -162.355 ;
        RECT 117.475 -164.045 117.805 -163.715 ;
        RECT 117.475 -165.405 117.805 -165.075 ;
        RECT 117.475 -166.765 117.805 -166.435 ;
        RECT 117.475 -168.125 117.805 -167.795 ;
        RECT 117.475 -169.485 117.805 -169.155 ;
        RECT 117.475 -170.845 117.805 -170.515 ;
        RECT 117.475 -172.205 117.805 -171.875 ;
        RECT 117.475 -173.565 117.805 -173.235 ;
        RECT 117.475 -174.925 117.805 -174.595 ;
        RECT 117.475 -176.285 117.805 -175.955 ;
        RECT 117.475 -177.645 117.805 -177.315 ;
        RECT 117.475 -179.005 117.805 -178.675 ;
        RECT 117.475 -180.365 117.805 -180.035 ;
        RECT 117.475 -181.725 117.805 -181.395 ;
        RECT 117.475 -183.085 117.805 -182.755 ;
        RECT 117.475 -184.445 117.805 -184.115 ;
        RECT 117.475 -185.805 117.805 -185.475 ;
        RECT 117.475 -187.165 117.805 -186.835 ;
        RECT 117.475 -188.525 117.805 -188.195 ;
        RECT 117.475 -189.885 117.805 -189.555 ;
        RECT 117.475 -191.245 117.805 -190.915 ;
        RECT 117.475 -192.605 117.805 -192.275 ;
        RECT 117.475 -193.965 117.805 -193.635 ;
        RECT 117.475 -195.325 117.805 -194.995 ;
        RECT 117.475 -196.685 117.805 -196.355 ;
        RECT 117.475 -198.045 117.805 -197.715 ;
        RECT 117.475 -199.405 117.805 -199.075 ;
        RECT 117.475 -200.765 117.805 -200.435 ;
        RECT 117.475 -202.125 117.805 -201.795 ;
        RECT 117.475 -203.485 117.805 -203.155 ;
        RECT 117.475 -204.845 117.805 -204.515 ;
        RECT 117.475 -206.205 117.805 -205.875 ;
        RECT 117.475 -207.565 117.805 -207.235 ;
        RECT 117.475 -208.925 117.805 -208.595 ;
        RECT 117.475 -210.285 117.805 -209.955 ;
        RECT 117.475 -211.645 117.805 -211.315 ;
        RECT 117.475 -213.005 117.805 -212.675 ;
        RECT 117.475 -214.365 117.805 -214.035 ;
        RECT 117.475 -215.725 117.805 -215.395 ;
        RECT 117.475 -217.085 117.805 -216.755 ;
        RECT 117.475 -218.445 117.805 -218.115 ;
        RECT 117.475 -219.805 117.805 -219.475 ;
        RECT 117.475 -221.165 117.805 -220.835 ;
        RECT 117.475 -222.525 117.805 -222.195 ;
        RECT 117.475 -223.885 117.805 -223.555 ;
        RECT 117.475 -225.245 117.805 -224.915 ;
        RECT 117.475 -226.605 117.805 -226.275 ;
        RECT 117.475 -227.965 117.805 -227.635 ;
        RECT 117.475 -229.325 117.805 -228.995 ;
        RECT 117.475 -230.685 117.805 -230.355 ;
        RECT 117.475 -232.045 117.805 -231.715 ;
        RECT 117.475 -233.405 117.805 -233.075 ;
        RECT 117.475 -234.765 117.805 -234.435 ;
        RECT 117.475 -236.125 117.805 -235.795 ;
        RECT 117.475 -237.485 117.805 -237.155 ;
        RECT 117.475 -238.845 117.805 -238.515 ;
        RECT 117.475 -241.09 117.805 -239.96 ;
        RECT 117.48 -241.205 117.8 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 244.04 119.165 245.17 ;
        RECT 118.835 242.595 119.165 242.925 ;
        RECT 118.835 241.235 119.165 241.565 ;
        RECT 118.835 239.875 119.165 240.205 ;
        RECT 118.835 238.515 119.165 238.845 ;
        RECT 118.835 237.155 119.165 237.485 ;
        RECT 118.84 237.155 119.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 -0.845 119.165 -0.515 ;
        RECT 118.835 -2.205 119.165 -1.875 ;
        RECT 118.835 -3.565 119.165 -3.235 ;
        RECT 118.84 -3.565 119.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 -123.245 119.165 -122.915 ;
        RECT 118.835 -124.605 119.165 -124.275 ;
        RECT 118.835 -125.965 119.165 -125.635 ;
        RECT 118.835 -127.325 119.165 -126.995 ;
        RECT 118.835 -128.685 119.165 -128.355 ;
        RECT 118.835 -130.045 119.165 -129.715 ;
        RECT 118.835 -131.405 119.165 -131.075 ;
        RECT 118.835 -132.765 119.165 -132.435 ;
        RECT 118.835 -134.125 119.165 -133.795 ;
        RECT 118.835 -135.485 119.165 -135.155 ;
        RECT 118.835 -136.845 119.165 -136.515 ;
        RECT 118.835 -138.205 119.165 -137.875 ;
        RECT 118.835 -139.565 119.165 -139.235 ;
        RECT 118.835 -140.925 119.165 -140.595 ;
        RECT 118.835 -142.285 119.165 -141.955 ;
        RECT 118.835 -143.645 119.165 -143.315 ;
        RECT 118.835 -145.005 119.165 -144.675 ;
        RECT 118.835 -146.365 119.165 -146.035 ;
        RECT 118.835 -147.725 119.165 -147.395 ;
        RECT 118.835 -149.085 119.165 -148.755 ;
        RECT 118.835 -150.445 119.165 -150.115 ;
        RECT 118.835 -151.805 119.165 -151.475 ;
        RECT 118.835 -153.165 119.165 -152.835 ;
        RECT 118.835 -154.525 119.165 -154.195 ;
        RECT 118.835 -155.885 119.165 -155.555 ;
        RECT 118.835 -157.245 119.165 -156.915 ;
        RECT 118.835 -158.605 119.165 -158.275 ;
        RECT 118.835 -159.965 119.165 -159.635 ;
        RECT 118.835 -161.325 119.165 -160.995 ;
        RECT 118.835 -162.685 119.165 -162.355 ;
        RECT 118.835 -164.045 119.165 -163.715 ;
        RECT 118.835 -165.405 119.165 -165.075 ;
        RECT 118.835 -166.765 119.165 -166.435 ;
        RECT 118.835 -168.125 119.165 -167.795 ;
        RECT 118.835 -169.485 119.165 -169.155 ;
        RECT 118.835 -170.845 119.165 -170.515 ;
        RECT 118.835 -172.205 119.165 -171.875 ;
        RECT 118.835 -173.565 119.165 -173.235 ;
        RECT 118.835 -174.925 119.165 -174.595 ;
        RECT 118.835 -176.285 119.165 -175.955 ;
        RECT 118.835 -177.645 119.165 -177.315 ;
        RECT 118.835 -179.005 119.165 -178.675 ;
        RECT 118.835 -180.365 119.165 -180.035 ;
        RECT 118.835 -181.725 119.165 -181.395 ;
        RECT 118.835 -183.085 119.165 -182.755 ;
        RECT 118.835 -184.445 119.165 -184.115 ;
        RECT 118.835 -185.805 119.165 -185.475 ;
        RECT 118.835 -187.165 119.165 -186.835 ;
        RECT 118.835 -188.525 119.165 -188.195 ;
        RECT 118.835 -189.885 119.165 -189.555 ;
        RECT 118.835 -191.245 119.165 -190.915 ;
        RECT 118.835 -192.605 119.165 -192.275 ;
        RECT 118.835 -193.965 119.165 -193.635 ;
        RECT 118.835 -195.325 119.165 -194.995 ;
        RECT 118.835 -196.685 119.165 -196.355 ;
        RECT 118.835 -198.045 119.165 -197.715 ;
        RECT 118.835 -199.405 119.165 -199.075 ;
        RECT 118.835 -200.765 119.165 -200.435 ;
        RECT 118.835 -202.125 119.165 -201.795 ;
        RECT 118.835 -203.485 119.165 -203.155 ;
        RECT 118.835 -204.845 119.165 -204.515 ;
        RECT 118.835 -206.205 119.165 -205.875 ;
        RECT 118.835 -207.565 119.165 -207.235 ;
        RECT 118.835 -208.925 119.165 -208.595 ;
        RECT 118.835 -210.285 119.165 -209.955 ;
        RECT 118.835 -211.645 119.165 -211.315 ;
        RECT 118.835 -213.005 119.165 -212.675 ;
        RECT 118.835 -214.365 119.165 -214.035 ;
        RECT 118.835 -215.725 119.165 -215.395 ;
        RECT 118.835 -217.085 119.165 -216.755 ;
        RECT 118.835 -218.445 119.165 -218.115 ;
        RECT 118.835 -219.805 119.165 -219.475 ;
        RECT 118.835 -221.165 119.165 -220.835 ;
        RECT 118.835 -222.525 119.165 -222.195 ;
        RECT 118.835 -223.885 119.165 -223.555 ;
        RECT 118.835 -225.245 119.165 -224.915 ;
        RECT 118.835 -226.605 119.165 -226.275 ;
        RECT 118.835 -227.965 119.165 -227.635 ;
        RECT 118.835 -229.325 119.165 -228.995 ;
        RECT 118.835 -230.685 119.165 -230.355 ;
        RECT 118.835 -232.045 119.165 -231.715 ;
        RECT 118.835 -233.405 119.165 -233.075 ;
        RECT 118.835 -234.765 119.165 -234.435 ;
        RECT 118.835 -236.125 119.165 -235.795 ;
        RECT 118.835 -237.485 119.165 -237.155 ;
        RECT 118.835 -238.845 119.165 -238.515 ;
        RECT 118.835 -241.09 119.165 -239.96 ;
        RECT 118.84 -241.205 119.16 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 244.04 120.525 245.17 ;
        RECT 120.195 242.595 120.525 242.925 ;
        RECT 120.195 241.235 120.525 241.565 ;
        RECT 120.195 239.875 120.525 240.205 ;
        RECT 120.195 238.515 120.525 238.845 ;
        RECT 120.195 237.155 120.525 237.485 ;
        RECT 120.2 237.155 120.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 -0.845 120.525 -0.515 ;
        RECT 120.195 -2.205 120.525 -1.875 ;
        RECT 120.195 -3.565 120.525 -3.235 ;
        RECT 120.2 -3.565 120.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 -123.245 120.525 -122.915 ;
        RECT 120.195 -124.605 120.525 -124.275 ;
        RECT 120.195 -125.965 120.525 -125.635 ;
        RECT 120.195 -127.325 120.525 -126.995 ;
        RECT 120.195 -128.685 120.525 -128.355 ;
        RECT 120.195 -130.045 120.525 -129.715 ;
        RECT 120.195 -131.405 120.525 -131.075 ;
        RECT 120.195 -132.765 120.525 -132.435 ;
        RECT 120.195 -134.125 120.525 -133.795 ;
        RECT 120.195 -135.485 120.525 -135.155 ;
        RECT 120.195 -136.845 120.525 -136.515 ;
        RECT 120.195 -138.205 120.525 -137.875 ;
        RECT 120.195 -139.565 120.525 -139.235 ;
        RECT 120.195 -140.925 120.525 -140.595 ;
        RECT 120.195 -142.285 120.525 -141.955 ;
        RECT 120.195 -143.645 120.525 -143.315 ;
        RECT 120.195 -145.005 120.525 -144.675 ;
        RECT 120.195 -146.365 120.525 -146.035 ;
        RECT 120.195 -147.725 120.525 -147.395 ;
        RECT 120.195 -149.085 120.525 -148.755 ;
        RECT 120.195 -150.445 120.525 -150.115 ;
        RECT 120.195 -151.805 120.525 -151.475 ;
        RECT 120.195 -153.165 120.525 -152.835 ;
        RECT 120.195 -154.525 120.525 -154.195 ;
        RECT 120.195 -155.885 120.525 -155.555 ;
        RECT 120.195 -157.245 120.525 -156.915 ;
        RECT 120.195 -158.605 120.525 -158.275 ;
        RECT 120.195 -159.965 120.525 -159.635 ;
        RECT 120.195 -161.325 120.525 -160.995 ;
        RECT 120.195 -162.685 120.525 -162.355 ;
        RECT 120.195 -164.045 120.525 -163.715 ;
        RECT 120.195 -165.405 120.525 -165.075 ;
        RECT 120.195 -166.765 120.525 -166.435 ;
        RECT 120.195 -168.125 120.525 -167.795 ;
        RECT 120.195 -169.485 120.525 -169.155 ;
        RECT 120.195 -170.845 120.525 -170.515 ;
        RECT 120.195 -172.205 120.525 -171.875 ;
        RECT 120.195 -173.565 120.525 -173.235 ;
        RECT 120.195 -174.925 120.525 -174.595 ;
        RECT 120.195 -176.285 120.525 -175.955 ;
        RECT 120.195 -177.645 120.525 -177.315 ;
        RECT 120.195 -179.005 120.525 -178.675 ;
        RECT 120.195 -180.365 120.525 -180.035 ;
        RECT 120.195 -181.725 120.525 -181.395 ;
        RECT 120.195 -183.085 120.525 -182.755 ;
        RECT 120.195 -184.445 120.525 -184.115 ;
        RECT 120.195 -185.805 120.525 -185.475 ;
        RECT 120.195 -187.165 120.525 -186.835 ;
        RECT 120.195 -188.525 120.525 -188.195 ;
        RECT 120.195 -189.885 120.525 -189.555 ;
        RECT 120.195 -191.245 120.525 -190.915 ;
        RECT 120.195 -192.605 120.525 -192.275 ;
        RECT 120.195 -193.965 120.525 -193.635 ;
        RECT 120.195 -195.325 120.525 -194.995 ;
        RECT 120.195 -196.685 120.525 -196.355 ;
        RECT 120.195 -198.045 120.525 -197.715 ;
        RECT 120.195 -199.405 120.525 -199.075 ;
        RECT 120.195 -200.765 120.525 -200.435 ;
        RECT 120.195 -202.125 120.525 -201.795 ;
        RECT 120.195 -203.485 120.525 -203.155 ;
        RECT 120.195 -204.845 120.525 -204.515 ;
        RECT 120.195 -206.205 120.525 -205.875 ;
        RECT 120.195 -207.565 120.525 -207.235 ;
        RECT 120.195 -208.925 120.525 -208.595 ;
        RECT 120.195 -210.285 120.525 -209.955 ;
        RECT 120.195 -211.645 120.525 -211.315 ;
        RECT 120.195 -213.005 120.525 -212.675 ;
        RECT 120.195 -214.365 120.525 -214.035 ;
        RECT 120.195 -215.725 120.525 -215.395 ;
        RECT 120.195 -217.085 120.525 -216.755 ;
        RECT 120.195 -218.445 120.525 -218.115 ;
        RECT 120.195 -219.805 120.525 -219.475 ;
        RECT 120.195 -221.165 120.525 -220.835 ;
        RECT 120.195 -222.525 120.525 -222.195 ;
        RECT 120.195 -223.885 120.525 -223.555 ;
        RECT 120.195 -225.245 120.525 -224.915 ;
        RECT 120.195 -226.605 120.525 -226.275 ;
        RECT 120.195 -227.965 120.525 -227.635 ;
        RECT 120.195 -229.325 120.525 -228.995 ;
        RECT 120.195 -230.685 120.525 -230.355 ;
        RECT 120.195 -232.045 120.525 -231.715 ;
        RECT 120.195 -233.405 120.525 -233.075 ;
        RECT 120.195 -234.765 120.525 -234.435 ;
        RECT 120.195 -236.125 120.525 -235.795 ;
        RECT 120.195 -237.485 120.525 -237.155 ;
        RECT 120.195 -238.845 120.525 -238.515 ;
        RECT 120.195 -241.09 120.525 -239.96 ;
        RECT 120.2 -241.205 120.52 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 244.04 121.885 245.17 ;
        RECT 121.555 242.595 121.885 242.925 ;
        RECT 121.555 241.235 121.885 241.565 ;
        RECT 121.555 239.875 121.885 240.205 ;
        RECT 121.555 238.515 121.885 238.845 ;
        RECT 121.555 237.155 121.885 237.485 ;
        RECT 121.56 237.155 121.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 -0.845 121.885 -0.515 ;
        RECT 121.555 -2.205 121.885 -1.875 ;
        RECT 121.555 -3.565 121.885 -3.235 ;
        RECT 121.56 -3.565 121.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 -123.245 121.885 -122.915 ;
        RECT 121.555 -124.605 121.885 -124.275 ;
        RECT 121.555 -125.965 121.885 -125.635 ;
        RECT 121.555 -127.325 121.885 -126.995 ;
        RECT 121.555 -128.685 121.885 -128.355 ;
        RECT 121.555 -130.045 121.885 -129.715 ;
        RECT 121.555 -131.405 121.885 -131.075 ;
        RECT 121.555 -132.765 121.885 -132.435 ;
        RECT 121.555 -134.125 121.885 -133.795 ;
        RECT 121.555 -135.485 121.885 -135.155 ;
        RECT 121.555 -136.845 121.885 -136.515 ;
        RECT 121.555 -138.205 121.885 -137.875 ;
        RECT 121.555 -139.565 121.885 -139.235 ;
        RECT 121.555 -140.925 121.885 -140.595 ;
        RECT 121.555 -142.285 121.885 -141.955 ;
        RECT 121.555 -143.645 121.885 -143.315 ;
        RECT 121.555 -145.005 121.885 -144.675 ;
        RECT 121.555 -146.365 121.885 -146.035 ;
        RECT 121.555 -147.725 121.885 -147.395 ;
        RECT 121.555 -149.085 121.885 -148.755 ;
        RECT 121.555 -150.445 121.885 -150.115 ;
        RECT 121.555 -151.805 121.885 -151.475 ;
        RECT 121.555 -153.165 121.885 -152.835 ;
        RECT 121.555 -154.525 121.885 -154.195 ;
        RECT 121.555 -155.885 121.885 -155.555 ;
        RECT 121.555 -157.245 121.885 -156.915 ;
        RECT 121.555 -158.605 121.885 -158.275 ;
        RECT 121.555 -159.965 121.885 -159.635 ;
        RECT 121.555 -161.325 121.885 -160.995 ;
        RECT 121.555 -162.685 121.885 -162.355 ;
        RECT 121.555 -164.045 121.885 -163.715 ;
        RECT 121.555 -165.405 121.885 -165.075 ;
        RECT 121.555 -166.765 121.885 -166.435 ;
        RECT 121.555 -168.125 121.885 -167.795 ;
        RECT 121.555 -169.485 121.885 -169.155 ;
        RECT 121.555 -170.845 121.885 -170.515 ;
        RECT 121.555 -172.205 121.885 -171.875 ;
        RECT 121.555 -173.565 121.885 -173.235 ;
        RECT 121.555 -174.925 121.885 -174.595 ;
        RECT 121.555 -176.285 121.885 -175.955 ;
        RECT 121.555 -177.645 121.885 -177.315 ;
        RECT 121.555 -179.005 121.885 -178.675 ;
        RECT 121.555 -180.365 121.885 -180.035 ;
        RECT 121.555 -181.725 121.885 -181.395 ;
        RECT 121.555 -183.085 121.885 -182.755 ;
        RECT 121.555 -184.445 121.885 -184.115 ;
        RECT 121.555 -185.805 121.885 -185.475 ;
        RECT 121.555 -187.165 121.885 -186.835 ;
        RECT 121.555 -188.525 121.885 -188.195 ;
        RECT 121.555 -189.885 121.885 -189.555 ;
        RECT 121.555 -191.245 121.885 -190.915 ;
        RECT 121.555 -192.605 121.885 -192.275 ;
        RECT 121.555 -193.965 121.885 -193.635 ;
        RECT 121.555 -195.325 121.885 -194.995 ;
        RECT 121.555 -196.685 121.885 -196.355 ;
        RECT 121.555 -198.045 121.885 -197.715 ;
        RECT 121.555 -199.405 121.885 -199.075 ;
        RECT 121.555 -200.765 121.885 -200.435 ;
        RECT 121.555 -202.125 121.885 -201.795 ;
        RECT 121.555 -203.485 121.885 -203.155 ;
        RECT 121.555 -204.845 121.885 -204.515 ;
        RECT 121.555 -206.205 121.885 -205.875 ;
        RECT 121.555 -207.565 121.885 -207.235 ;
        RECT 121.555 -208.925 121.885 -208.595 ;
        RECT 121.555 -210.285 121.885 -209.955 ;
        RECT 121.555 -211.645 121.885 -211.315 ;
        RECT 121.555 -213.005 121.885 -212.675 ;
        RECT 121.555 -214.365 121.885 -214.035 ;
        RECT 121.555 -215.725 121.885 -215.395 ;
        RECT 121.555 -217.085 121.885 -216.755 ;
        RECT 121.555 -218.445 121.885 -218.115 ;
        RECT 121.555 -219.805 121.885 -219.475 ;
        RECT 121.555 -221.165 121.885 -220.835 ;
        RECT 121.555 -222.525 121.885 -222.195 ;
        RECT 121.555 -223.885 121.885 -223.555 ;
        RECT 121.555 -225.245 121.885 -224.915 ;
        RECT 121.555 -226.605 121.885 -226.275 ;
        RECT 121.555 -227.965 121.885 -227.635 ;
        RECT 121.555 -229.325 121.885 -228.995 ;
        RECT 121.555 -230.685 121.885 -230.355 ;
        RECT 121.555 -232.045 121.885 -231.715 ;
        RECT 121.555 -233.405 121.885 -233.075 ;
        RECT 121.555 -234.765 121.885 -234.435 ;
        RECT 121.555 -236.125 121.885 -235.795 ;
        RECT 121.555 -237.485 121.885 -237.155 ;
        RECT 121.555 -238.845 121.885 -238.515 ;
        RECT 121.555 -241.09 121.885 -239.96 ;
        RECT 121.56 -241.205 121.88 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 244.04 123.245 245.17 ;
        RECT 122.915 242.595 123.245 242.925 ;
        RECT 122.915 241.235 123.245 241.565 ;
        RECT 122.915 239.875 123.245 240.205 ;
        RECT 122.915 238.515 123.245 238.845 ;
        RECT 122.915 237.155 123.245 237.485 ;
        RECT 122.92 237.155 123.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -127.325 123.245 -126.995 ;
        RECT 122.915 -128.685 123.245 -128.355 ;
        RECT 122.915 -130.045 123.245 -129.715 ;
        RECT 122.915 -131.405 123.245 -131.075 ;
        RECT 122.915 -132.765 123.245 -132.435 ;
        RECT 122.915 -134.125 123.245 -133.795 ;
        RECT 122.915 -135.485 123.245 -135.155 ;
        RECT 122.915 -136.845 123.245 -136.515 ;
        RECT 122.915 -138.205 123.245 -137.875 ;
        RECT 122.915 -139.565 123.245 -139.235 ;
        RECT 122.915 -140.925 123.245 -140.595 ;
        RECT 122.915 -142.285 123.245 -141.955 ;
        RECT 122.915 -143.645 123.245 -143.315 ;
        RECT 122.915 -145.005 123.245 -144.675 ;
        RECT 122.915 -146.365 123.245 -146.035 ;
        RECT 122.915 -147.725 123.245 -147.395 ;
        RECT 122.915 -149.085 123.245 -148.755 ;
        RECT 122.915 -150.445 123.245 -150.115 ;
        RECT 122.915 -151.805 123.245 -151.475 ;
        RECT 122.915 -153.165 123.245 -152.835 ;
        RECT 122.915 -154.525 123.245 -154.195 ;
        RECT 122.915 -155.885 123.245 -155.555 ;
        RECT 122.915 -157.245 123.245 -156.915 ;
        RECT 122.915 -158.605 123.245 -158.275 ;
        RECT 122.915 -159.965 123.245 -159.635 ;
        RECT 122.915 -161.325 123.245 -160.995 ;
        RECT 122.915 -162.685 123.245 -162.355 ;
        RECT 122.915 -164.045 123.245 -163.715 ;
        RECT 122.915 -165.405 123.245 -165.075 ;
        RECT 122.915 -166.765 123.245 -166.435 ;
        RECT 122.915 -168.125 123.245 -167.795 ;
        RECT 122.915 -169.485 123.245 -169.155 ;
        RECT 122.915 -170.845 123.245 -170.515 ;
        RECT 122.915 -172.205 123.245 -171.875 ;
        RECT 122.915 -173.565 123.245 -173.235 ;
        RECT 122.915 -174.925 123.245 -174.595 ;
        RECT 122.915 -176.285 123.245 -175.955 ;
        RECT 122.915 -177.645 123.245 -177.315 ;
        RECT 122.915 -179.005 123.245 -178.675 ;
        RECT 122.915 -180.365 123.245 -180.035 ;
        RECT 122.915 -181.725 123.245 -181.395 ;
        RECT 122.915 -183.085 123.245 -182.755 ;
        RECT 122.915 -184.445 123.245 -184.115 ;
        RECT 122.915 -185.805 123.245 -185.475 ;
        RECT 122.915 -187.165 123.245 -186.835 ;
        RECT 122.915 -188.525 123.245 -188.195 ;
        RECT 122.915 -189.885 123.245 -189.555 ;
        RECT 122.915 -191.245 123.245 -190.915 ;
        RECT 122.915 -192.605 123.245 -192.275 ;
        RECT 122.915 -193.965 123.245 -193.635 ;
        RECT 122.915 -195.325 123.245 -194.995 ;
        RECT 122.915 -196.685 123.245 -196.355 ;
        RECT 122.915 -198.045 123.245 -197.715 ;
        RECT 122.915 -199.405 123.245 -199.075 ;
        RECT 122.915 -200.765 123.245 -200.435 ;
        RECT 122.915 -202.125 123.245 -201.795 ;
        RECT 122.915 -203.485 123.245 -203.155 ;
        RECT 122.915 -204.845 123.245 -204.515 ;
        RECT 122.915 -206.205 123.245 -205.875 ;
        RECT 122.915 -207.565 123.245 -207.235 ;
        RECT 122.915 -208.925 123.245 -208.595 ;
        RECT 122.915 -210.285 123.245 -209.955 ;
        RECT 122.915 -211.645 123.245 -211.315 ;
        RECT 122.915 -213.005 123.245 -212.675 ;
        RECT 122.915 -214.365 123.245 -214.035 ;
        RECT 122.915 -215.725 123.245 -215.395 ;
        RECT 122.915 -217.085 123.245 -216.755 ;
        RECT 122.915 -218.445 123.245 -218.115 ;
        RECT 122.915 -219.805 123.245 -219.475 ;
        RECT 122.915 -221.165 123.245 -220.835 ;
        RECT 122.915 -222.525 123.245 -222.195 ;
        RECT 122.915 -223.885 123.245 -223.555 ;
        RECT 122.915 -225.245 123.245 -224.915 ;
        RECT 122.915 -226.605 123.245 -226.275 ;
        RECT 122.915 -227.965 123.245 -227.635 ;
        RECT 122.915 -229.325 123.245 -228.995 ;
        RECT 122.915 -230.685 123.245 -230.355 ;
        RECT 122.915 -232.045 123.245 -231.715 ;
        RECT 122.915 -233.405 123.245 -233.075 ;
        RECT 122.915 -234.765 123.245 -234.435 ;
        RECT 122.915 -236.125 123.245 -235.795 ;
        RECT 122.915 -237.485 123.245 -237.155 ;
        RECT 122.915 -238.845 123.245 -238.515 ;
        RECT 122.915 -241.09 123.245 -239.96 ;
        RECT 122.92 -241.205 123.24 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.21 -125.535 123.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 244.04 124.605 245.17 ;
        RECT 124.275 242.595 124.605 242.925 ;
        RECT 124.275 241.235 124.605 241.565 ;
        RECT 124.275 239.875 124.605 240.205 ;
        RECT 124.275 238.515 124.605 238.845 ;
        RECT 124.275 237.155 124.605 237.485 ;
        RECT 124.28 237.155 124.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 -0.845 124.605 -0.515 ;
        RECT 124.275 -2.205 124.605 -1.875 ;
        RECT 124.275 -3.565 124.605 -3.235 ;
        RECT 124.28 -3.565 124.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 244.04 125.965 245.17 ;
        RECT 125.635 242.595 125.965 242.925 ;
        RECT 125.635 241.235 125.965 241.565 ;
        RECT 125.635 239.875 125.965 240.205 ;
        RECT 125.635 238.515 125.965 238.845 ;
        RECT 125.635 237.155 125.965 237.485 ;
        RECT 125.64 237.155 125.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 -0.845 125.965 -0.515 ;
        RECT 125.635 -2.205 125.965 -1.875 ;
        RECT 125.635 -3.565 125.965 -3.235 ;
        RECT 125.64 -3.565 125.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 244.04 127.325 245.17 ;
        RECT 126.995 242.595 127.325 242.925 ;
        RECT 126.995 241.235 127.325 241.565 ;
        RECT 126.995 239.875 127.325 240.205 ;
        RECT 126.995 238.515 127.325 238.845 ;
        RECT 126.995 237.155 127.325 237.485 ;
        RECT 127 237.155 127.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 -0.845 127.325 -0.515 ;
        RECT 126.995 -2.205 127.325 -1.875 ;
        RECT 126.995 -3.565 127.325 -3.235 ;
        RECT 127 -3.565 127.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 -123.245 127.325 -122.915 ;
        RECT 126.995 -124.605 127.325 -124.275 ;
        RECT 126.995 -125.965 127.325 -125.635 ;
        RECT 126.995 -127.325 127.325 -126.995 ;
        RECT 126.995 -128.685 127.325 -128.355 ;
        RECT 126.995 -130.045 127.325 -129.715 ;
        RECT 126.995 -131.405 127.325 -131.075 ;
        RECT 126.995 -132.765 127.325 -132.435 ;
        RECT 126.995 -134.125 127.325 -133.795 ;
        RECT 126.995 -135.485 127.325 -135.155 ;
        RECT 126.995 -136.845 127.325 -136.515 ;
        RECT 126.995 -138.205 127.325 -137.875 ;
        RECT 126.995 -139.565 127.325 -139.235 ;
        RECT 126.995 -140.925 127.325 -140.595 ;
        RECT 126.995 -142.285 127.325 -141.955 ;
        RECT 126.995 -143.645 127.325 -143.315 ;
        RECT 126.995 -145.005 127.325 -144.675 ;
        RECT 126.995 -146.365 127.325 -146.035 ;
        RECT 126.995 -147.725 127.325 -147.395 ;
        RECT 126.995 -149.085 127.325 -148.755 ;
        RECT 126.995 -150.445 127.325 -150.115 ;
        RECT 126.995 -151.805 127.325 -151.475 ;
        RECT 126.995 -153.165 127.325 -152.835 ;
        RECT 126.995 -154.525 127.325 -154.195 ;
        RECT 126.995 -155.885 127.325 -155.555 ;
        RECT 126.995 -157.245 127.325 -156.915 ;
        RECT 126.995 -158.605 127.325 -158.275 ;
        RECT 126.995 -159.965 127.325 -159.635 ;
        RECT 126.995 -161.325 127.325 -160.995 ;
        RECT 126.995 -162.685 127.325 -162.355 ;
        RECT 126.995 -164.045 127.325 -163.715 ;
        RECT 126.995 -165.405 127.325 -165.075 ;
        RECT 126.995 -166.765 127.325 -166.435 ;
        RECT 126.995 -168.125 127.325 -167.795 ;
        RECT 126.995 -169.485 127.325 -169.155 ;
        RECT 126.995 -170.845 127.325 -170.515 ;
        RECT 126.995 -172.205 127.325 -171.875 ;
        RECT 126.995 -173.565 127.325 -173.235 ;
        RECT 126.995 -174.925 127.325 -174.595 ;
        RECT 126.995 -176.285 127.325 -175.955 ;
        RECT 126.995 -177.645 127.325 -177.315 ;
        RECT 126.995 -179.005 127.325 -178.675 ;
        RECT 126.995 -180.365 127.325 -180.035 ;
        RECT 126.995 -181.725 127.325 -181.395 ;
        RECT 126.995 -183.085 127.325 -182.755 ;
        RECT 126.995 -184.445 127.325 -184.115 ;
        RECT 126.995 -185.805 127.325 -185.475 ;
        RECT 126.995 -187.165 127.325 -186.835 ;
        RECT 126.995 -188.525 127.325 -188.195 ;
        RECT 126.995 -189.885 127.325 -189.555 ;
        RECT 126.995 -191.245 127.325 -190.915 ;
        RECT 126.995 -192.605 127.325 -192.275 ;
        RECT 126.995 -193.965 127.325 -193.635 ;
        RECT 126.995 -195.325 127.325 -194.995 ;
        RECT 126.995 -196.685 127.325 -196.355 ;
        RECT 126.995 -198.045 127.325 -197.715 ;
        RECT 126.995 -199.405 127.325 -199.075 ;
        RECT 126.995 -200.765 127.325 -200.435 ;
        RECT 126.995 -202.125 127.325 -201.795 ;
        RECT 126.995 -203.485 127.325 -203.155 ;
        RECT 126.995 -204.845 127.325 -204.515 ;
        RECT 126.995 -206.205 127.325 -205.875 ;
        RECT 126.995 -207.565 127.325 -207.235 ;
        RECT 126.995 -208.925 127.325 -208.595 ;
        RECT 126.995 -210.285 127.325 -209.955 ;
        RECT 126.995 -211.645 127.325 -211.315 ;
        RECT 126.995 -213.005 127.325 -212.675 ;
        RECT 126.995 -214.365 127.325 -214.035 ;
        RECT 126.995 -215.725 127.325 -215.395 ;
        RECT 126.995 -217.085 127.325 -216.755 ;
        RECT 126.995 -218.445 127.325 -218.115 ;
        RECT 126.995 -219.805 127.325 -219.475 ;
        RECT 126.995 -221.165 127.325 -220.835 ;
        RECT 126.995 -222.525 127.325 -222.195 ;
        RECT 126.995 -223.885 127.325 -223.555 ;
        RECT 126.995 -225.245 127.325 -224.915 ;
        RECT 126.995 -226.605 127.325 -226.275 ;
        RECT 126.995 -227.965 127.325 -227.635 ;
        RECT 126.995 -229.325 127.325 -228.995 ;
        RECT 126.995 -230.685 127.325 -230.355 ;
        RECT 126.995 -232.045 127.325 -231.715 ;
        RECT 126.995 -233.405 127.325 -233.075 ;
        RECT 126.995 -234.765 127.325 -234.435 ;
        RECT 126.995 -236.125 127.325 -235.795 ;
        RECT 126.995 -237.485 127.325 -237.155 ;
        RECT 126.995 -238.845 127.325 -238.515 ;
        RECT 126.995 -241.09 127.325 -239.96 ;
        RECT 127 -241.205 127.32 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 244.04 128.685 245.17 ;
        RECT 128.355 242.595 128.685 242.925 ;
        RECT 128.355 241.235 128.685 241.565 ;
        RECT 128.355 239.875 128.685 240.205 ;
        RECT 128.355 238.515 128.685 238.845 ;
        RECT 128.355 237.155 128.685 237.485 ;
        RECT 128.36 237.155 128.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -0.845 128.685 -0.515 ;
        RECT 128.355 -2.205 128.685 -1.875 ;
        RECT 128.355 -3.565 128.685 -3.235 ;
        RECT 128.36 -3.565 128.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -123.245 128.685 -122.915 ;
        RECT 128.355 -124.605 128.685 -124.275 ;
        RECT 128.355 -125.965 128.685 -125.635 ;
        RECT 128.355 -127.325 128.685 -126.995 ;
        RECT 128.355 -128.685 128.685 -128.355 ;
        RECT 128.355 -130.045 128.685 -129.715 ;
        RECT 128.355 -131.405 128.685 -131.075 ;
        RECT 128.355 -132.765 128.685 -132.435 ;
        RECT 128.355 -134.125 128.685 -133.795 ;
        RECT 128.355 -135.485 128.685 -135.155 ;
        RECT 128.355 -136.845 128.685 -136.515 ;
        RECT 128.355 -138.205 128.685 -137.875 ;
        RECT 128.355 -139.565 128.685 -139.235 ;
        RECT 128.355 -140.925 128.685 -140.595 ;
        RECT 128.355 -142.285 128.685 -141.955 ;
        RECT 128.355 -143.645 128.685 -143.315 ;
        RECT 128.355 -145.005 128.685 -144.675 ;
        RECT 128.355 -146.365 128.685 -146.035 ;
        RECT 128.355 -147.725 128.685 -147.395 ;
        RECT 128.355 -149.085 128.685 -148.755 ;
        RECT 128.355 -150.445 128.685 -150.115 ;
        RECT 128.355 -151.805 128.685 -151.475 ;
        RECT 128.355 -153.165 128.685 -152.835 ;
        RECT 128.355 -154.525 128.685 -154.195 ;
        RECT 128.355 -155.885 128.685 -155.555 ;
        RECT 128.355 -157.245 128.685 -156.915 ;
        RECT 128.355 -158.605 128.685 -158.275 ;
        RECT 128.355 -159.965 128.685 -159.635 ;
        RECT 128.355 -161.325 128.685 -160.995 ;
        RECT 128.355 -162.685 128.685 -162.355 ;
        RECT 128.355 -164.045 128.685 -163.715 ;
        RECT 128.355 -165.405 128.685 -165.075 ;
        RECT 128.355 -166.765 128.685 -166.435 ;
        RECT 128.355 -168.125 128.685 -167.795 ;
        RECT 128.355 -169.485 128.685 -169.155 ;
        RECT 128.355 -170.845 128.685 -170.515 ;
        RECT 128.355 -172.205 128.685 -171.875 ;
        RECT 128.355 -173.565 128.685 -173.235 ;
        RECT 128.355 -174.925 128.685 -174.595 ;
        RECT 128.355 -176.285 128.685 -175.955 ;
        RECT 128.355 -177.645 128.685 -177.315 ;
        RECT 128.355 -179.005 128.685 -178.675 ;
        RECT 128.355 -180.365 128.685 -180.035 ;
        RECT 128.355 -181.725 128.685 -181.395 ;
        RECT 128.355 -183.085 128.685 -182.755 ;
        RECT 128.355 -184.445 128.685 -184.115 ;
        RECT 128.355 -185.805 128.685 -185.475 ;
        RECT 128.355 -187.165 128.685 -186.835 ;
        RECT 128.355 -188.525 128.685 -188.195 ;
        RECT 128.355 -189.885 128.685 -189.555 ;
        RECT 128.355 -191.245 128.685 -190.915 ;
        RECT 128.355 -192.605 128.685 -192.275 ;
        RECT 128.355 -193.965 128.685 -193.635 ;
        RECT 128.355 -195.325 128.685 -194.995 ;
        RECT 128.355 -196.685 128.685 -196.355 ;
        RECT 128.355 -198.045 128.685 -197.715 ;
        RECT 128.355 -199.405 128.685 -199.075 ;
        RECT 128.355 -200.765 128.685 -200.435 ;
        RECT 128.355 -202.125 128.685 -201.795 ;
        RECT 128.355 -203.485 128.685 -203.155 ;
        RECT 128.355 -204.845 128.685 -204.515 ;
        RECT 128.355 -206.205 128.685 -205.875 ;
        RECT 128.355 -207.565 128.685 -207.235 ;
        RECT 128.355 -208.925 128.685 -208.595 ;
        RECT 128.355 -210.285 128.685 -209.955 ;
        RECT 128.355 -211.645 128.685 -211.315 ;
        RECT 128.355 -213.005 128.685 -212.675 ;
        RECT 128.355 -214.365 128.685 -214.035 ;
        RECT 128.355 -215.725 128.685 -215.395 ;
        RECT 128.355 -217.085 128.685 -216.755 ;
        RECT 128.355 -218.445 128.685 -218.115 ;
        RECT 128.355 -219.805 128.685 -219.475 ;
        RECT 128.355 -221.165 128.685 -220.835 ;
        RECT 128.355 -222.525 128.685 -222.195 ;
        RECT 128.355 -223.885 128.685 -223.555 ;
        RECT 128.355 -225.245 128.685 -224.915 ;
        RECT 128.355 -226.605 128.685 -226.275 ;
        RECT 128.355 -227.965 128.685 -227.635 ;
        RECT 128.355 -229.325 128.685 -228.995 ;
        RECT 128.355 -230.685 128.685 -230.355 ;
        RECT 128.355 -232.045 128.685 -231.715 ;
        RECT 128.355 -233.405 128.685 -233.075 ;
        RECT 128.355 -234.765 128.685 -234.435 ;
        RECT 128.355 -236.125 128.685 -235.795 ;
        RECT 128.355 -237.485 128.685 -237.155 ;
        RECT 128.355 -238.845 128.685 -238.515 ;
        RECT 128.355 -241.09 128.685 -239.96 ;
        RECT 128.36 -241.205 128.68 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 244.04 130.045 245.17 ;
        RECT 129.715 242.595 130.045 242.925 ;
        RECT 129.715 241.235 130.045 241.565 ;
        RECT 129.715 239.875 130.045 240.205 ;
        RECT 129.715 238.515 130.045 238.845 ;
        RECT 129.715 237.155 130.045 237.485 ;
        RECT 129.72 237.155 130.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -3.565 130.045 -3.235 ;
        RECT 129.72 -3.565 130.04 -0.515 ;
        RECT 129.715 -0.845 130.045 -0.515 ;
        RECT 129.715 -2.205 130.045 -1.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 244.04 96.045 245.17 ;
        RECT 95.715 242.595 96.045 242.925 ;
        RECT 95.715 241.235 96.045 241.565 ;
        RECT 95.715 239.875 96.045 240.205 ;
        RECT 95.715 238.515 96.045 238.845 ;
        RECT 95.715 237.155 96.045 237.485 ;
        RECT 95.72 237.155 96.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 -0.845 96.045 -0.515 ;
        RECT 95.715 -2.205 96.045 -1.875 ;
        RECT 95.715 -3.565 96.045 -3.235 ;
        RECT 95.72 -3.565 96.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 -123.245 96.045 -122.915 ;
        RECT 95.715 -124.605 96.045 -124.275 ;
        RECT 95.715 -125.965 96.045 -125.635 ;
        RECT 95.715 -127.325 96.045 -126.995 ;
        RECT 95.715 -128.685 96.045 -128.355 ;
        RECT 95.715 -130.045 96.045 -129.715 ;
        RECT 95.715 -131.405 96.045 -131.075 ;
        RECT 95.715 -132.765 96.045 -132.435 ;
        RECT 95.715 -134.125 96.045 -133.795 ;
        RECT 95.715 -135.485 96.045 -135.155 ;
        RECT 95.715 -136.845 96.045 -136.515 ;
        RECT 95.715 -138.205 96.045 -137.875 ;
        RECT 95.715 -139.565 96.045 -139.235 ;
        RECT 95.715 -140.925 96.045 -140.595 ;
        RECT 95.715 -142.285 96.045 -141.955 ;
        RECT 95.715 -143.645 96.045 -143.315 ;
        RECT 95.715 -145.005 96.045 -144.675 ;
        RECT 95.715 -146.365 96.045 -146.035 ;
        RECT 95.715 -147.725 96.045 -147.395 ;
        RECT 95.715 -149.085 96.045 -148.755 ;
        RECT 95.715 -150.445 96.045 -150.115 ;
        RECT 95.715 -151.805 96.045 -151.475 ;
        RECT 95.715 -153.165 96.045 -152.835 ;
        RECT 95.715 -154.525 96.045 -154.195 ;
        RECT 95.715 -155.885 96.045 -155.555 ;
        RECT 95.715 -157.245 96.045 -156.915 ;
        RECT 95.715 -158.605 96.045 -158.275 ;
        RECT 95.715 -159.965 96.045 -159.635 ;
        RECT 95.715 -161.325 96.045 -160.995 ;
        RECT 95.715 -162.685 96.045 -162.355 ;
        RECT 95.715 -164.045 96.045 -163.715 ;
        RECT 95.715 -165.405 96.045 -165.075 ;
        RECT 95.715 -166.765 96.045 -166.435 ;
        RECT 95.715 -168.125 96.045 -167.795 ;
        RECT 95.715 -169.485 96.045 -169.155 ;
        RECT 95.715 -170.845 96.045 -170.515 ;
        RECT 95.715 -172.205 96.045 -171.875 ;
        RECT 95.715 -173.565 96.045 -173.235 ;
        RECT 95.715 -174.925 96.045 -174.595 ;
        RECT 95.715 -176.285 96.045 -175.955 ;
        RECT 95.715 -177.645 96.045 -177.315 ;
        RECT 95.715 -179.005 96.045 -178.675 ;
        RECT 95.715 -180.365 96.045 -180.035 ;
        RECT 95.715 -181.725 96.045 -181.395 ;
        RECT 95.715 -183.085 96.045 -182.755 ;
        RECT 95.715 -184.445 96.045 -184.115 ;
        RECT 95.715 -185.805 96.045 -185.475 ;
        RECT 95.715 -187.165 96.045 -186.835 ;
        RECT 95.715 -188.525 96.045 -188.195 ;
        RECT 95.715 -189.885 96.045 -189.555 ;
        RECT 95.715 -191.245 96.045 -190.915 ;
        RECT 95.715 -192.605 96.045 -192.275 ;
        RECT 95.715 -193.965 96.045 -193.635 ;
        RECT 95.715 -195.325 96.045 -194.995 ;
        RECT 95.715 -196.685 96.045 -196.355 ;
        RECT 95.715 -198.045 96.045 -197.715 ;
        RECT 95.715 -199.405 96.045 -199.075 ;
        RECT 95.715 -200.765 96.045 -200.435 ;
        RECT 95.715 -202.125 96.045 -201.795 ;
        RECT 95.715 -203.485 96.045 -203.155 ;
        RECT 95.715 -204.845 96.045 -204.515 ;
        RECT 95.715 -206.205 96.045 -205.875 ;
        RECT 95.715 -207.565 96.045 -207.235 ;
        RECT 95.715 -208.925 96.045 -208.595 ;
        RECT 95.715 -210.285 96.045 -209.955 ;
        RECT 95.715 -211.645 96.045 -211.315 ;
        RECT 95.715 -213.005 96.045 -212.675 ;
        RECT 95.715 -214.365 96.045 -214.035 ;
        RECT 95.715 -215.725 96.045 -215.395 ;
        RECT 95.715 -217.085 96.045 -216.755 ;
        RECT 95.715 -218.445 96.045 -218.115 ;
        RECT 95.715 -219.805 96.045 -219.475 ;
        RECT 95.715 -221.165 96.045 -220.835 ;
        RECT 95.715 -222.525 96.045 -222.195 ;
        RECT 95.715 -223.885 96.045 -223.555 ;
        RECT 95.715 -225.245 96.045 -224.915 ;
        RECT 95.715 -226.605 96.045 -226.275 ;
        RECT 95.715 -227.965 96.045 -227.635 ;
        RECT 95.715 -229.325 96.045 -228.995 ;
        RECT 95.715 -230.685 96.045 -230.355 ;
        RECT 95.715 -232.045 96.045 -231.715 ;
        RECT 95.715 -233.405 96.045 -233.075 ;
        RECT 95.715 -234.765 96.045 -234.435 ;
        RECT 95.715 -236.125 96.045 -235.795 ;
        RECT 95.715 -237.485 96.045 -237.155 ;
        RECT 95.715 -238.845 96.045 -238.515 ;
        RECT 95.715 -241.09 96.045 -239.96 ;
        RECT 95.72 -241.205 96.04 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 244.04 97.405 245.17 ;
        RECT 97.075 242.595 97.405 242.925 ;
        RECT 97.075 241.235 97.405 241.565 ;
        RECT 97.075 239.875 97.405 240.205 ;
        RECT 97.075 238.515 97.405 238.845 ;
        RECT 97.075 237.155 97.405 237.485 ;
        RECT 97.08 237.155 97.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 -0.845 97.405 -0.515 ;
        RECT 97.075 -2.205 97.405 -1.875 ;
        RECT 97.075 -3.565 97.405 -3.235 ;
        RECT 97.08 -3.565 97.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 -123.245 97.405 -122.915 ;
        RECT 97.075 -124.605 97.405 -124.275 ;
        RECT 97.075 -125.965 97.405 -125.635 ;
        RECT 97.075 -127.325 97.405 -126.995 ;
        RECT 97.075 -128.685 97.405 -128.355 ;
        RECT 97.075 -130.045 97.405 -129.715 ;
        RECT 97.075 -131.405 97.405 -131.075 ;
        RECT 97.075 -132.765 97.405 -132.435 ;
        RECT 97.075 -134.125 97.405 -133.795 ;
        RECT 97.075 -135.485 97.405 -135.155 ;
        RECT 97.075 -136.845 97.405 -136.515 ;
        RECT 97.075 -138.205 97.405 -137.875 ;
        RECT 97.075 -139.565 97.405 -139.235 ;
        RECT 97.075 -140.925 97.405 -140.595 ;
        RECT 97.075 -142.285 97.405 -141.955 ;
        RECT 97.075 -143.645 97.405 -143.315 ;
        RECT 97.075 -145.005 97.405 -144.675 ;
        RECT 97.075 -146.365 97.405 -146.035 ;
        RECT 97.075 -147.725 97.405 -147.395 ;
        RECT 97.075 -149.085 97.405 -148.755 ;
        RECT 97.075 -150.445 97.405 -150.115 ;
        RECT 97.075 -151.805 97.405 -151.475 ;
        RECT 97.075 -153.165 97.405 -152.835 ;
        RECT 97.075 -154.525 97.405 -154.195 ;
        RECT 97.075 -155.885 97.405 -155.555 ;
        RECT 97.075 -157.245 97.405 -156.915 ;
        RECT 97.075 -158.605 97.405 -158.275 ;
        RECT 97.075 -159.965 97.405 -159.635 ;
        RECT 97.075 -161.325 97.405 -160.995 ;
        RECT 97.075 -162.685 97.405 -162.355 ;
        RECT 97.075 -164.045 97.405 -163.715 ;
        RECT 97.075 -165.405 97.405 -165.075 ;
        RECT 97.075 -166.765 97.405 -166.435 ;
        RECT 97.075 -168.125 97.405 -167.795 ;
        RECT 97.075 -169.485 97.405 -169.155 ;
        RECT 97.075 -170.845 97.405 -170.515 ;
        RECT 97.075 -172.205 97.405 -171.875 ;
        RECT 97.075 -173.565 97.405 -173.235 ;
        RECT 97.075 -174.925 97.405 -174.595 ;
        RECT 97.075 -176.285 97.405 -175.955 ;
        RECT 97.075 -177.645 97.405 -177.315 ;
        RECT 97.075 -179.005 97.405 -178.675 ;
        RECT 97.075 -180.365 97.405 -180.035 ;
        RECT 97.075 -181.725 97.405 -181.395 ;
        RECT 97.075 -183.085 97.405 -182.755 ;
        RECT 97.075 -184.445 97.405 -184.115 ;
        RECT 97.075 -185.805 97.405 -185.475 ;
        RECT 97.075 -187.165 97.405 -186.835 ;
        RECT 97.075 -188.525 97.405 -188.195 ;
        RECT 97.075 -189.885 97.405 -189.555 ;
        RECT 97.075 -191.245 97.405 -190.915 ;
        RECT 97.075 -192.605 97.405 -192.275 ;
        RECT 97.075 -193.965 97.405 -193.635 ;
        RECT 97.075 -195.325 97.405 -194.995 ;
        RECT 97.075 -196.685 97.405 -196.355 ;
        RECT 97.075 -198.045 97.405 -197.715 ;
        RECT 97.075 -199.405 97.405 -199.075 ;
        RECT 97.075 -200.765 97.405 -200.435 ;
        RECT 97.075 -202.125 97.405 -201.795 ;
        RECT 97.075 -203.485 97.405 -203.155 ;
        RECT 97.075 -204.845 97.405 -204.515 ;
        RECT 97.075 -206.205 97.405 -205.875 ;
        RECT 97.075 -207.565 97.405 -207.235 ;
        RECT 97.075 -208.925 97.405 -208.595 ;
        RECT 97.075 -210.285 97.405 -209.955 ;
        RECT 97.075 -211.645 97.405 -211.315 ;
        RECT 97.075 -213.005 97.405 -212.675 ;
        RECT 97.075 -214.365 97.405 -214.035 ;
        RECT 97.075 -215.725 97.405 -215.395 ;
        RECT 97.075 -217.085 97.405 -216.755 ;
        RECT 97.075 -218.445 97.405 -218.115 ;
        RECT 97.075 -219.805 97.405 -219.475 ;
        RECT 97.075 -221.165 97.405 -220.835 ;
        RECT 97.075 -222.525 97.405 -222.195 ;
        RECT 97.075 -223.885 97.405 -223.555 ;
        RECT 97.075 -225.245 97.405 -224.915 ;
        RECT 97.075 -226.605 97.405 -226.275 ;
        RECT 97.075 -227.965 97.405 -227.635 ;
        RECT 97.075 -229.325 97.405 -228.995 ;
        RECT 97.075 -230.685 97.405 -230.355 ;
        RECT 97.075 -232.045 97.405 -231.715 ;
        RECT 97.075 -233.405 97.405 -233.075 ;
        RECT 97.075 -234.765 97.405 -234.435 ;
        RECT 97.075 -236.125 97.405 -235.795 ;
        RECT 97.075 -237.485 97.405 -237.155 ;
        RECT 97.075 -238.845 97.405 -238.515 ;
        RECT 97.075 -241.09 97.405 -239.96 ;
        RECT 97.08 -241.205 97.4 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 244.04 98.765 245.17 ;
        RECT 98.435 242.595 98.765 242.925 ;
        RECT 98.435 241.235 98.765 241.565 ;
        RECT 98.435 239.875 98.765 240.205 ;
        RECT 98.435 238.515 98.765 238.845 ;
        RECT 98.435 237.155 98.765 237.485 ;
        RECT 98.44 237.155 98.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -0.845 98.765 -0.515 ;
        RECT 98.435 -2.205 98.765 -1.875 ;
        RECT 98.435 -3.565 98.765 -3.235 ;
        RECT 98.44 -3.565 98.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -123.245 98.765 -122.915 ;
        RECT 98.435 -124.605 98.765 -124.275 ;
        RECT 98.435 -125.965 98.765 -125.635 ;
        RECT 98.435 -127.325 98.765 -126.995 ;
        RECT 98.435 -128.685 98.765 -128.355 ;
        RECT 98.435 -130.045 98.765 -129.715 ;
        RECT 98.435 -131.405 98.765 -131.075 ;
        RECT 98.435 -132.765 98.765 -132.435 ;
        RECT 98.435 -134.125 98.765 -133.795 ;
        RECT 98.435 -135.485 98.765 -135.155 ;
        RECT 98.435 -136.845 98.765 -136.515 ;
        RECT 98.435 -138.205 98.765 -137.875 ;
        RECT 98.435 -139.565 98.765 -139.235 ;
        RECT 98.435 -140.925 98.765 -140.595 ;
        RECT 98.435 -142.285 98.765 -141.955 ;
        RECT 98.435 -143.645 98.765 -143.315 ;
        RECT 98.435 -145.005 98.765 -144.675 ;
        RECT 98.435 -146.365 98.765 -146.035 ;
        RECT 98.435 -147.725 98.765 -147.395 ;
        RECT 98.435 -149.085 98.765 -148.755 ;
        RECT 98.435 -150.445 98.765 -150.115 ;
        RECT 98.435 -151.805 98.765 -151.475 ;
        RECT 98.435 -153.165 98.765 -152.835 ;
        RECT 98.435 -154.525 98.765 -154.195 ;
        RECT 98.435 -155.885 98.765 -155.555 ;
        RECT 98.435 -157.245 98.765 -156.915 ;
        RECT 98.435 -158.605 98.765 -158.275 ;
        RECT 98.435 -159.965 98.765 -159.635 ;
        RECT 98.435 -161.325 98.765 -160.995 ;
        RECT 98.435 -162.685 98.765 -162.355 ;
        RECT 98.435 -164.045 98.765 -163.715 ;
        RECT 98.435 -165.405 98.765 -165.075 ;
        RECT 98.435 -166.765 98.765 -166.435 ;
        RECT 98.435 -168.125 98.765 -167.795 ;
        RECT 98.435 -169.485 98.765 -169.155 ;
        RECT 98.435 -170.845 98.765 -170.515 ;
        RECT 98.435 -172.205 98.765 -171.875 ;
        RECT 98.435 -173.565 98.765 -173.235 ;
        RECT 98.435 -174.925 98.765 -174.595 ;
        RECT 98.435 -176.285 98.765 -175.955 ;
        RECT 98.435 -177.645 98.765 -177.315 ;
        RECT 98.435 -179.005 98.765 -178.675 ;
        RECT 98.435 -180.365 98.765 -180.035 ;
        RECT 98.435 -181.725 98.765 -181.395 ;
        RECT 98.435 -183.085 98.765 -182.755 ;
        RECT 98.435 -184.445 98.765 -184.115 ;
        RECT 98.435 -185.805 98.765 -185.475 ;
        RECT 98.435 -187.165 98.765 -186.835 ;
        RECT 98.435 -188.525 98.765 -188.195 ;
        RECT 98.435 -189.885 98.765 -189.555 ;
        RECT 98.435 -191.245 98.765 -190.915 ;
        RECT 98.435 -192.605 98.765 -192.275 ;
        RECT 98.435 -193.965 98.765 -193.635 ;
        RECT 98.435 -195.325 98.765 -194.995 ;
        RECT 98.435 -196.685 98.765 -196.355 ;
        RECT 98.435 -198.045 98.765 -197.715 ;
        RECT 98.435 -199.405 98.765 -199.075 ;
        RECT 98.435 -200.765 98.765 -200.435 ;
        RECT 98.435 -202.125 98.765 -201.795 ;
        RECT 98.435 -203.485 98.765 -203.155 ;
        RECT 98.435 -204.845 98.765 -204.515 ;
        RECT 98.435 -206.205 98.765 -205.875 ;
        RECT 98.435 -207.565 98.765 -207.235 ;
        RECT 98.435 -208.925 98.765 -208.595 ;
        RECT 98.435 -210.285 98.765 -209.955 ;
        RECT 98.435 -211.645 98.765 -211.315 ;
        RECT 98.435 -213.005 98.765 -212.675 ;
        RECT 98.435 -214.365 98.765 -214.035 ;
        RECT 98.435 -215.725 98.765 -215.395 ;
        RECT 98.435 -217.085 98.765 -216.755 ;
        RECT 98.435 -218.445 98.765 -218.115 ;
        RECT 98.435 -219.805 98.765 -219.475 ;
        RECT 98.435 -221.165 98.765 -220.835 ;
        RECT 98.435 -222.525 98.765 -222.195 ;
        RECT 98.435 -223.885 98.765 -223.555 ;
        RECT 98.435 -225.245 98.765 -224.915 ;
        RECT 98.435 -226.605 98.765 -226.275 ;
        RECT 98.435 -227.965 98.765 -227.635 ;
        RECT 98.435 -229.325 98.765 -228.995 ;
        RECT 98.435 -230.685 98.765 -230.355 ;
        RECT 98.435 -232.045 98.765 -231.715 ;
        RECT 98.435 -233.405 98.765 -233.075 ;
        RECT 98.435 -234.765 98.765 -234.435 ;
        RECT 98.435 -236.125 98.765 -235.795 ;
        RECT 98.435 -237.485 98.765 -237.155 ;
        RECT 98.435 -238.845 98.765 -238.515 ;
        RECT 98.435 -241.09 98.765 -239.96 ;
        RECT 98.44 -241.205 98.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 244.04 100.125 245.17 ;
        RECT 99.795 242.595 100.125 242.925 ;
        RECT 99.795 241.235 100.125 241.565 ;
        RECT 99.795 239.875 100.125 240.205 ;
        RECT 99.795 238.515 100.125 238.845 ;
        RECT 99.795 237.155 100.125 237.485 ;
        RECT 99.8 237.155 100.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 -0.845 100.125 -0.515 ;
        RECT 99.795 -2.205 100.125 -1.875 ;
        RECT 99.795 -3.565 100.125 -3.235 ;
        RECT 99.8 -3.565 100.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 -123.245 100.125 -122.915 ;
        RECT 99.795 -124.605 100.125 -124.275 ;
        RECT 99.795 -125.965 100.125 -125.635 ;
        RECT 99.795 -127.325 100.125 -126.995 ;
        RECT 99.795 -128.685 100.125 -128.355 ;
        RECT 99.795 -130.045 100.125 -129.715 ;
        RECT 99.795 -131.405 100.125 -131.075 ;
        RECT 99.795 -132.765 100.125 -132.435 ;
        RECT 99.795 -134.125 100.125 -133.795 ;
        RECT 99.795 -135.485 100.125 -135.155 ;
        RECT 99.795 -136.845 100.125 -136.515 ;
        RECT 99.795 -138.205 100.125 -137.875 ;
        RECT 99.795 -139.565 100.125 -139.235 ;
        RECT 99.795 -140.925 100.125 -140.595 ;
        RECT 99.795 -142.285 100.125 -141.955 ;
        RECT 99.795 -143.645 100.125 -143.315 ;
        RECT 99.795 -145.005 100.125 -144.675 ;
        RECT 99.795 -146.365 100.125 -146.035 ;
        RECT 99.795 -147.725 100.125 -147.395 ;
        RECT 99.795 -149.085 100.125 -148.755 ;
        RECT 99.795 -150.445 100.125 -150.115 ;
        RECT 99.795 -151.805 100.125 -151.475 ;
        RECT 99.795 -153.165 100.125 -152.835 ;
        RECT 99.795 -154.525 100.125 -154.195 ;
        RECT 99.795 -155.885 100.125 -155.555 ;
        RECT 99.795 -157.245 100.125 -156.915 ;
        RECT 99.795 -158.605 100.125 -158.275 ;
        RECT 99.795 -159.965 100.125 -159.635 ;
        RECT 99.795 -161.325 100.125 -160.995 ;
        RECT 99.795 -162.685 100.125 -162.355 ;
        RECT 99.795 -164.045 100.125 -163.715 ;
        RECT 99.795 -165.405 100.125 -165.075 ;
        RECT 99.795 -166.765 100.125 -166.435 ;
        RECT 99.795 -168.125 100.125 -167.795 ;
        RECT 99.795 -169.485 100.125 -169.155 ;
        RECT 99.795 -170.845 100.125 -170.515 ;
        RECT 99.795 -172.205 100.125 -171.875 ;
        RECT 99.795 -173.565 100.125 -173.235 ;
        RECT 99.795 -174.925 100.125 -174.595 ;
        RECT 99.795 -176.285 100.125 -175.955 ;
        RECT 99.795 -177.645 100.125 -177.315 ;
        RECT 99.795 -179.005 100.125 -178.675 ;
        RECT 99.795 -180.365 100.125 -180.035 ;
        RECT 99.795 -181.725 100.125 -181.395 ;
        RECT 99.795 -183.085 100.125 -182.755 ;
        RECT 99.795 -184.445 100.125 -184.115 ;
        RECT 99.795 -185.805 100.125 -185.475 ;
        RECT 99.795 -187.165 100.125 -186.835 ;
        RECT 99.795 -188.525 100.125 -188.195 ;
        RECT 99.795 -189.885 100.125 -189.555 ;
        RECT 99.795 -191.245 100.125 -190.915 ;
        RECT 99.795 -192.605 100.125 -192.275 ;
        RECT 99.795 -193.965 100.125 -193.635 ;
        RECT 99.795 -195.325 100.125 -194.995 ;
        RECT 99.795 -196.685 100.125 -196.355 ;
        RECT 99.795 -198.045 100.125 -197.715 ;
        RECT 99.795 -199.405 100.125 -199.075 ;
        RECT 99.795 -200.765 100.125 -200.435 ;
        RECT 99.795 -202.125 100.125 -201.795 ;
        RECT 99.795 -203.485 100.125 -203.155 ;
        RECT 99.795 -204.845 100.125 -204.515 ;
        RECT 99.795 -206.205 100.125 -205.875 ;
        RECT 99.795 -207.565 100.125 -207.235 ;
        RECT 99.795 -208.925 100.125 -208.595 ;
        RECT 99.795 -210.285 100.125 -209.955 ;
        RECT 99.795 -211.645 100.125 -211.315 ;
        RECT 99.795 -213.005 100.125 -212.675 ;
        RECT 99.795 -214.365 100.125 -214.035 ;
        RECT 99.795 -215.725 100.125 -215.395 ;
        RECT 99.795 -217.085 100.125 -216.755 ;
        RECT 99.795 -218.445 100.125 -218.115 ;
        RECT 99.795 -219.805 100.125 -219.475 ;
        RECT 99.795 -221.165 100.125 -220.835 ;
        RECT 99.795 -222.525 100.125 -222.195 ;
        RECT 99.795 -223.885 100.125 -223.555 ;
        RECT 99.795 -225.245 100.125 -224.915 ;
        RECT 99.795 -226.605 100.125 -226.275 ;
        RECT 99.795 -227.965 100.125 -227.635 ;
        RECT 99.795 -229.325 100.125 -228.995 ;
        RECT 99.795 -230.685 100.125 -230.355 ;
        RECT 99.795 -232.045 100.125 -231.715 ;
        RECT 99.795 -233.405 100.125 -233.075 ;
        RECT 99.795 -234.765 100.125 -234.435 ;
        RECT 99.795 -236.125 100.125 -235.795 ;
        RECT 99.795 -237.485 100.125 -237.155 ;
        RECT 99.795 -238.845 100.125 -238.515 ;
        RECT 99.795 -241.09 100.125 -239.96 ;
        RECT 99.8 -241.205 100.12 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 244.04 101.485 245.17 ;
        RECT 101.155 242.595 101.485 242.925 ;
        RECT 101.155 241.235 101.485 241.565 ;
        RECT 101.155 239.875 101.485 240.205 ;
        RECT 101.155 238.515 101.485 238.845 ;
        RECT 101.155 237.155 101.485 237.485 ;
        RECT 101.16 237.155 101.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 -127.325 101.485 -126.995 ;
        RECT 101.155 -128.685 101.485 -128.355 ;
        RECT 101.155 -130.045 101.485 -129.715 ;
        RECT 101.155 -131.405 101.485 -131.075 ;
        RECT 101.155 -132.765 101.485 -132.435 ;
        RECT 101.155 -134.125 101.485 -133.795 ;
        RECT 101.155 -135.485 101.485 -135.155 ;
        RECT 101.155 -136.845 101.485 -136.515 ;
        RECT 101.155 -138.205 101.485 -137.875 ;
        RECT 101.155 -139.565 101.485 -139.235 ;
        RECT 101.155 -140.925 101.485 -140.595 ;
        RECT 101.155 -142.285 101.485 -141.955 ;
        RECT 101.155 -143.645 101.485 -143.315 ;
        RECT 101.155 -145.005 101.485 -144.675 ;
        RECT 101.155 -146.365 101.485 -146.035 ;
        RECT 101.155 -147.725 101.485 -147.395 ;
        RECT 101.155 -149.085 101.485 -148.755 ;
        RECT 101.155 -150.445 101.485 -150.115 ;
        RECT 101.155 -151.805 101.485 -151.475 ;
        RECT 101.155 -153.165 101.485 -152.835 ;
        RECT 101.155 -154.525 101.485 -154.195 ;
        RECT 101.155 -155.885 101.485 -155.555 ;
        RECT 101.155 -157.245 101.485 -156.915 ;
        RECT 101.155 -158.605 101.485 -158.275 ;
        RECT 101.155 -159.965 101.485 -159.635 ;
        RECT 101.155 -161.325 101.485 -160.995 ;
        RECT 101.155 -162.685 101.485 -162.355 ;
        RECT 101.155 -164.045 101.485 -163.715 ;
        RECT 101.155 -165.405 101.485 -165.075 ;
        RECT 101.155 -166.765 101.485 -166.435 ;
        RECT 101.155 -168.125 101.485 -167.795 ;
        RECT 101.155 -169.485 101.485 -169.155 ;
        RECT 101.155 -170.845 101.485 -170.515 ;
        RECT 101.155 -172.205 101.485 -171.875 ;
        RECT 101.155 -173.565 101.485 -173.235 ;
        RECT 101.155 -174.925 101.485 -174.595 ;
        RECT 101.155 -176.285 101.485 -175.955 ;
        RECT 101.155 -177.645 101.485 -177.315 ;
        RECT 101.155 -179.005 101.485 -178.675 ;
        RECT 101.155 -180.365 101.485 -180.035 ;
        RECT 101.155 -181.725 101.485 -181.395 ;
        RECT 101.155 -183.085 101.485 -182.755 ;
        RECT 101.155 -184.445 101.485 -184.115 ;
        RECT 101.155 -185.805 101.485 -185.475 ;
        RECT 101.155 -187.165 101.485 -186.835 ;
        RECT 101.155 -188.525 101.485 -188.195 ;
        RECT 101.155 -189.885 101.485 -189.555 ;
        RECT 101.155 -191.245 101.485 -190.915 ;
        RECT 101.155 -192.605 101.485 -192.275 ;
        RECT 101.155 -193.965 101.485 -193.635 ;
        RECT 101.155 -195.325 101.485 -194.995 ;
        RECT 101.155 -196.685 101.485 -196.355 ;
        RECT 101.155 -198.045 101.485 -197.715 ;
        RECT 101.155 -199.405 101.485 -199.075 ;
        RECT 101.155 -200.765 101.485 -200.435 ;
        RECT 101.155 -202.125 101.485 -201.795 ;
        RECT 101.155 -203.485 101.485 -203.155 ;
        RECT 101.155 -204.845 101.485 -204.515 ;
        RECT 101.155 -206.205 101.485 -205.875 ;
        RECT 101.155 -207.565 101.485 -207.235 ;
        RECT 101.155 -208.925 101.485 -208.595 ;
        RECT 101.155 -210.285 101.485 -209.955 ;
        RECT 101.155 -211.645 101.485 -211.315 ;
        RECT 101.155 -213.005 101.485 -212.675 ;
        RECT 101.155 -214.365 101.485 -214.035 ;
        RECT 101.155 -215.725 101.485 -215.395 ;
        RECT 101.155 -217.085 101.485 -216.755 ;
        RECT 101.155 -218.445 101.485 -218.115 ;
        RECT 101.155 -219.805 101.485 -219.475 ;
        RECT 101.155 -221.165 101.485 -220.835 ;
        RECT 101.155 -222.525 101.485 -222.195 ;
        RECT 101.155 -223.885 101.485 -223.555 ;
        RECT 101.155 -225.245 101.485 -224.915 ;
        RECT 101.155 -226.605 101.485 -226.275 ;
        RECT 101.155 -227.965 101.485 -227.635 ;
        RECT 101.155 -229.325 101.485 -228.995 ;
        RECT 101.155 -230.685 101.485 -230.355 ;
        RECT 101.155 -232.045 101.485 -231.715 ;
        RECT 101.155 -233.405 101.485 -233.075 ;
        RECT 101.155 -234.765 101.485 -234.435 ;
        RECT 101.155 -236.125 101.485 -235.795 ;
        RECT 101.155 -237.485 101.485 -237.155 ;
        RECT 101.155 -238.845 101.485 -238.515 ;
        RECT 101.155 -241.09 101.485 -239.96 ;
        RECT 101.16 -241.205 101.48 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.41 -125.535 101.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 244.04 102.845 245.17 ;
        RECT 102.515 242.595 102.845 242.925 ;
        RECT 102.515 241.235 102.845 241.565 ;
        RECT 102.515 239.875 102.845 240.205 ;
        RECT 102.515 238.515 102.845 238.845 ;
        RECT 102.515 237.155 102.845 237.485 ;
        RECT 102.52 237.155 102.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 -0.845 102.845 -0.515 ;
        RECT 102.515 -2.205 102.845 -1.875 ;
        RECT 102.515 -3.565 102.845 -3.235 ;
        RECT 102.52 -3.565 102.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 244.04 104.205 245.17 ;
        RECT 103.875 242.595 104.205 242.925 ;
        RECT 103.875 241.235 104.205 241.565 ;
        RECT 103.875 239.875 104.205 240.205 ;
        RECT 103.875 238.515 104.205 238.845 ;
        RECT 103.875 237.155 104.205 237.485 ;
        RECT 103.88 237.155 104.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 -0.845 104.205 -0.515 ;
        RECT 103.875 -2.205 104.205 -1.875 ;
        RECT 103.875 -3.565 104.205 -3.235 ;
        RECT 103.88 -3.565 104.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 244.04 105.565 245.17 ;
        RECT 105.235 242.595 105.565 242.925 ;
        RECT 105.235 241.235 105.565 241.565 ;
        RECT 105.235 239.875 105.565 240.205 ;
        RECT 105.235 238.515 105.565 238.845 ;
        RECT 105.235 237.155 105.565 237.485 ;
        RECT 105.24 237.155 105.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -0.845 105.565 -0.515 ;
        RECT 105.235 -2.205 105.565 -1.875 ;
        RECT 105.235 -3.565 105.565 -3.235 ;
        RECT 105.24 -3.565 105.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -123.245 105.565 -122.915 ;
        RECT 105.235 -124.605 105.565 -124.275 ;
        RECT 105.235 -125.965 105.565 -125.635 ;
        RECT 105.235 -127.325 105.565 -126.995 ;
        RECT 105.235 -128.685 105.565 -128.355 ;
        RECT 105.235 -130.045 105.565 -129.715 ;
        RECT 105.235 -131.405 105.565 -131.075 ;
        RECT 105.235 -132.765 105.565 -132.435 ;
        RECT 105.235 -134.125 105.565 -133.795 ;
        RECT 105.235 -135.485 105.565 -135.155 ;
        RECT 105.235 -136.845 105.565 -136.515 ;
        RECT 105.235 -138.205 105.565 -137.875 ;
        RECT 105.235 -139.565 105.565 -139.235 ;
        RECT 105.235 -140.925 105.565 -140.595 ;
        RECT 105.235 -142.285 105.565 -141.955 ;
        RECT 105.235 -143.645 105.565 -143.315 ;
        RECT 105.235 -145.005 105.565 -144.675 ;
        RECT 105.235 -146.365 105.565 -146.035 ;
        RECT 105.235 -147.725 105.565 -147.395 ;
        RECT 105.235 -149.085 105.565 -148.755 ;
        RECT 105.235 -150.445 105.565 -150.115 ;
        RECT 105.235 -151.805 105.565 -151.475 ;
        RECT 105.235 -153.165 105.565 -152.835 ;
        RECT 105.235 -154.525 105.565 -154.195 ;
        RECT 105.235 -155.885 105.565 -155.555 ;
        RECT 105.235 -157.245 105.565 -156.915 ;
        RECT 105.235 -158.605 105.565 -158.275 ;
        RECT 105.235 -159.965 105.565 -159.635 ;
        RECT 105.235 -161.325 105.565 -160.995 ;
        RECT 105.235 -162.685 105.565 -162.355 ;
        RECT 105.235 -164.045 105.565 -163.715 ;
        RECT 105.235 -165.405 105.565 -165.075 ;
        RECT 105.235 -166.765 105.565 -166.435 ;
        RECT 105.235 -168.125 105.565 -167.795 ;
        RECT 105.235 -169.485 105.565 -169.155 ;
        RECT 105.235 -170.845 105.565 -170.515 ;
        RECT 105.235 -172.205 105.565 -171.875 ;
        RECT 105.235 -173.565 105.565 -173.235 ;
        RECT 105.235 -174.925 105.565 -174.595 ;
        RECT 105.235 -176.285 105.565 -175.955 ;
        RECT 105.235 -177.645 105.565 -177.315 ;
        RECT 105.235 -179.005 105.565 -178.675 ;
        RECT 105.235 -180.365 105.565 -180.035 ;
        RECT 105.235 -181.725 105.565 -181.395 ;
        RECT 105.235 -183.085 105.565 -182.755 ;
        RECT 105.235 -184.445 105.565 -184.115 ;
        RECT 105.235 -185.805 105.565 -185.475 ;
        RECT 105.235 -187.165 105.565 -186.835 ;
        RECT 105.235 -188.525 105.565 -188.195 ;
        RECT 105.235 -189.885 105.565 -189.555 ;
        RECT 105.235 -191.245 105.565 -190.915 ;
        RECT 105.235 -192.605 105.565 -192.275 ;
        RECT 105.235 -193.965 105.565 -193.635 ;
        RECT 105.235 -195.325 105.565 -194.995 ;
        RECT 105.235 -196.685 105.565 -196.355 ;
        RECT 105.235 -198.045 105.565 -197.715 ;
        RECT 105.235 -199.405 105.565 -199.075 ;
        RECT 105.235 -200.765 105.565 -200.435 ;
        RECT 105.235 -202.125 105.565 -201.795 ;
        RECT 105.235 -203.485 105.565 -203.155 ;
        RECT 105.235 -204.845 105.565 -204.515 ;
        RECT 105.235 -206.205 105.565 -205.875 ;
        RECT 105.235 -207.565 105.565 -207.235 ;
        RECT 105.235 -208.925 105.565 -208.595 ;
        RECT 105.235 -210.285 105.565 -209.955 ;
        RECT 105.235 -211.645 105.565 -211.315 ;
        RECT 105.235 -213.005 105.565 -212.675 ;
        RECT 105.235 -214.365 105.565 -214.035 ;
        RECT 105.235 -215.725 105.565 -215.395 ;
        RECT 105.235 -217.085 105.565 -216.755 ;
        RECT 105.235 -218.445 105.565 -218.115 ;
        RECT 105.235 -219.805 105.565 -219.475 ;
        RECT 105.235 -221.165 105.565 -220.835 ;
        RECT 105.235 -222.525 105.565 -222.195 ;
        RECT 105.235 -223.885 105.565 -223.555 ;
        RECT 105.235 -225.245 105.565 -224.915 ;
        RECT 105.235 -226.605 105.565 -226.275 ;
        RECT 105.235 -227.965 105.565 -227.635 ;
        RECT 105.235 -229.325 105.565 -228.995 ;
        RECT 105.235 -230.685 105.565 -230.355 ;
        RECT 105.235 -232.045 105.565 -231.715 ;
        RECT 105.235 -233.405 105.565 -233.075 ;
        RECT 105.235 -234.765 105.565 -234.435 ;
        RECT 105.235 -236.125 105.565 -235.795 ;
        RECT 105.235 -237.485 105.565 -237.155 ;
        RECT 105.235 -238.845 105.565 -238.515 ;
        RECT 105.235 -241.09 105.565 -239.96 ;
        RECT 105.24 -241.205 105.56 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 244.04 106.925 245.17 ;
        RECT 106.595 242.595 106.925 242.925 ;
        RECT 106.595 241.235 106.925 241.565 ;
        RECT 106.595 239.875 106.925 240.205 ;
        RECT 106.595 238.515 106.925 238.845 ;
        RECT 106.595 237.155 106.925 237.485 ;
        RECT 106.6 237.155 106.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 -0.845 106.925 -0.515 ;
        RECT 106.595 -2.205 106.925 -1.875 ;
        RECT 106.595 -3.565 106.925 -3.235 ;
        RECT 106.6 -3.565 106.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 -123.245 106.925 -122.915 ;
        RECT 106.595 -124.605 106.925 -124.275 ;
        RECT 106.595 -125.965 106.925 -125.635 ;
        RECT 106.595 -127.325 106.925 -126.995 ;
        RECT 106.595 -128.685 106.925 -128.355 ;
        RECT 106.595 -130.045 106.925 -129.715 ;
        RECT 106.595 -131.405 106.925 -131.075 ;
        RECT 106.595 -132.765 106.925 -132.435 ;
        RECT 106.595 -134.125 106.925 -133.795 ;
        RECT 106.595 -135.485 106.925 -135.155 ;
        RECT 106.595 -136.845 106.925 -136.515 ;
        RECT 106.595 -138.205 106.925 -137.875 ;
        RECT 106.595 -139.565 106.925 -139.235 ;
        RECT 106.595 -140.925 106.925 -140.595 ;
        RECT 106.595 -142.285 106.925 -141.955 ;
        RECT 106.595 -143.645 106.925 -143.315 ;
        RECT 106.595 -145.005 106.925 -144.675 ;
        RECT 106.595 -146.365 106.925 -146.035 ;
        RECT 106.595 -147.725 106.925 -147.395 ;
        RECT 106.595 -149.085 106.925 -148.755 ;
        RECT 106.595 -150.445 106.925 -150.115 ;
        RECT 106.595 -151.805 106.925 -151.475 ;
        RECT 106.595 -153.165 106.925 -152.835 ;
        RECT 106.595 -154.525 106.925 -154.195 ;
        RECT 106.595 -155.885 106.925 -155.555 ;
        RECT 106.595 -157.245 106.925 -156.915 ;
        RECT 106.595 -158.605 106.925 -158.275 ;
        RECT 106.595 -159.965 106.925 -159.635 ;
        RECT 106.595 -161.325 106.925 -160.995 ;
        RECT 106.595 -162.685 106.925 -162.355 ;
        RECT 106.595 -164.045 106.925 -163.715 ;
        RECT 106.595 -165.405 106.925 -165.075 ;
        RECT 106.595 -166.765 106.925 -166.435 ;
        RECT 106.595 -168.125 106.925 -167.795 ;
        RECT 106.595 -169.485 106.925 -169.155 ;
        RECT 106.595 -170.845 106.925 -170.515 ;
        RECT 106.595 -172.205 106.925 -171.875 ;
        RECT 106.595 -173.565 106.925 -173.235 ;
        RECT 106.595 -174.925 106.925 -174.595 ;
        RECT 106.595 -176.285 106.925 -175.955 ;
        RECT 106.595 -177.645 106.925 -177.315 ;
        RECT 106.595 -179.005 106.925 -178.675 ;
        RECT 106.595 -180.365 106.925 -180.035 ;
        RECT 106.595 -181.725 106.925 -181.395 ;
        RECT 106.595 -183.085 106.925 -182.755 ;
        RECT 106.595 -184.445 106.925 -184.115 ;
        RECT 106.595 -185.805 106.925 -185.475 ;
        RECT 106.595 -187.165 106.925 -186.835 ;
        RECT 106.595 -188.525 106.925 -188.195 ;
        RECT 106.595 -189.885 106.925 -189.555 ;
        RECT 106.595 -191.245 106.925 -190.915 ;
        RECT 106.595 -192.605 106.925 -192.275 ;
        RECT 106.595 -193.965 106.925 -193.635 ;
        RECT 106.595 -195.325 106.925 -194.995 ;
        RECT 106.595 -196.685 106.925 -196.355 ;
        RECT 106.595 -198.045 106.925 -197.715 ;
        RECT 106.595 -199.405 106.925 -199.075 ;
        RECT 106.595 -200.765 106.925 -200.435 ;
        RECT 106.595 -202.125 106.925 -201.795 ;
        RECT 106.595 -203.485 106.925 -203.155 ;
        RECT 106.595 -204.845 106.925 -204.515 ;
        RECT 106.595 -206.205 106.925 -205.875 ;
        RECT 106.595 -207.565 106.925 -207.235 ;
        RECT 106.595 -208.925 106.925 -208.595 ;
        RECT 106.595 -210.285 106.925 -209.955 ;
        RECT 106.595 -211.645 106.925 -211.315 ;
        RECT 106.595 -213.005 106.925 -212.675 ;
        RECT 106.595 -214.365 106.925 -214.035 ;
        RECT 106.595 -215.725 106.925 -215.395 ;
        RECT 106.595 -217.085 106.925 -216.755 ;
        RECT 106.595 -218.445 106.925 -218.115 ;
        RECT 106.595 -219.805 106.925 -219.475 ;
        RECT 106.595 -221.165 106.925 -220.835 ;
        RECT 106.595 -222.525 106.925 -222.195 ;
        RECT 106.595 -223.885 106.925 -223.555 ;
        RECT 106.595 -225.245 106.925 -224.915 ;
        RECT 106.595 -226.605 106.925 -226.275 ;
        RECT 106.595 -227.965 106.925 -227.635 ;
        RECT 106.595 -229.325 106.925 -228.995 ;
        RECT 106.595 -230.685 106.925 -230.355 ;
        RECT 106.595 -232.045 106.925 -231.715 ;
        RECT 106.595 -233.405 106.925 -233.075 ;
        RECT 106.595 -234.765 106.925 -234.435 ;
        RECT 106.595 -236.125 106.925 -235.795 ;
        RECT 106.595 -237.485 106.925 -237.155 ;
        RECT 106.595 -238.845 106.925 -238.515 ;
        RECT 106.595 -241.09 106.925 -239.96 ;
        RECT 106.6 -241.205 106.92 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 244.04 108.285 245.17 ;
        RECT 107.955 242.595 108.285 242.925 ;
        RECT 107.955 241.235 108.285 241.565 ;
        RECT 107.955 239.875 108.285 240.205 ;
        RECT 107.955 238.515 108.285 238.845 ;
        RECT 107.955 237.155 108.285 237.485 ;
        RECT 107.96 237.155 108.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 -0.845 108.285 -0.515 ;
        RECT 107.955 -2.205 108.285 -1.875 ;
        RECT 107.955 -3.565 108.285 -3.235 ;
        RECT 107.96 -3.565 108.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 -123.245 108.285 -122.915 ;
        RECT 107.955 -124.605 108.285 -124.275 ;
        RECT 107.955 -125.965 108.285 -125.635 ;
        RECT 107.955 -127.325 108.285 -126.995 ;
        RECT 107.955 -128.685 108.285 -128.355 ;
        RECT 107.955 -130.045 108.285 -129.715 ;
        RECT 107.955 -131.405 108.285 -131.075 ;
        RECT 107.955 -132.765 108.285 -132.435 ;
        RECT 107.955 -134.125 108.285 -133.795 ;
        RECT 107.955 -135.485 108.285 -135.155 ;
        RECT 107.955 -136.845 108.285 -136.515 ;
        RECT 107.955 -138.205 108.285 -137.875 ;
        RECT 107.955 -139.565 108.285 -139.235 ;
        RECT 107.955 -140.925 108.285 -140.595 ;
        RECT 107.955 -142.285 108.285 -141.955 ;
        RECT 107.955 -143.645 108.285 -143.315 ;
        RECT 107.955 -145.005 108.285 -144.675 ;
        RECT 107.955 -146.365 108.285 -146.035 ;
        RECT 107.955 -147.725 108.285 -147.395 ;
        RECT 107.955 -149.085 108.285 -148.755 ;
        RECT 107.955 -150.445 108.285 -150.115 ;
        RECT 107.955 -151.805 108.285 -151.475 ;
        RECT 107.955 -153.165 108.285 -152.835 ;
        RECT 107.955 -154.525 108.285 -154.195 ;
        RECT 107.955 -155.885 108.285 -155.555 ;
        RECT 107.955 -157.245 108.285 -156.915 ;
        RECT 107.955 -158.605 108.285 -158.275 ;
        RECT 107.955 -159.965 108.285 -159.635 ;
        RECT 107.955 -161.325 108.285 -160.995 ;
        RECT 107.955 -162.685 108.285 -162.355 ;
        RECT 107.955 -164.045 108.285 -163.715 ;
        RECT 107.955 -165.405 108.285 -165.075 ;
        RECT 107.955 -166.765 108.285 -166.435 ;
        RECT 107.955 -168.125 108.285 -167.795 ;
        RECT 107.955 -169.485 108.285 -169.155 ;
        RECT 107.955 -170.845 108.285 -170.515 ;
        RECT 107.955 -172.205 108.285 -171.875 ;
        RECT 107.955 -173.565 108.285 -173.235 ;
        RECT 107.955 -174.925 108.285 -174.595 ;
        RECT 107.955 -176.285 108.285 -175.955 ;
        RECT 107.955 -177.645 108.285 -177.315 ;
        RECT 107.955 -179.005 108.285 -178.675 ;
        RECT 107.955 -180.365 108.285 -180.035 ;
        RECT 107.955 -181.725 108.285 -181.395 ;
        RECT 107.955 -183.085 108.285 -182.755 ;
        RECT 107.955 -184.445 108.285 -184.115 ;
        RECT 107.955 -185.805 108.285 -185.475 ;
        RECT 107.955 -187.165 108.285 -186.835 ;
        RECT 107.955 -188.525 108.285 -188.195 ;
        RECT 107.955 -189.885 108.285 -189.555 ;
        RECT 107.955 -191.245 108.285 -190.915 ;
        RECT 107.955 -192.605 108.285 -192.275 ;
        RECT 107.955 -193.965 108.285 -193.635 ;
        RECT 107.955 -195.325 108.285 -194.995 ;
        RECT 107.955 -196.685 108.285 -196.355 ;
        RECT 107.955 -198.045 108.285 -197.715 ;
        RECT 107.955 -199.405 108.285 -199.075 ;
        RECT 107.955 -200.765 108.285 -200.435 ;
        RECT 107.955 -202.125 108.285 -201.795 ;
        RECT 107.955 -203.485 108.285 -203.155 ;
        RECT 107.955 -204.845 108.285 -204.515 ;
        RECT 107.955 -206.205 108.285 -205.875 ;
        RECT 107.955 -207.565 108.285 -207.235 ;
        RECT 107.955 -208.925 108.285 -208.595 ;
        RECT 107.955 -210.285 108.285 -209.955 ;
        RECT 107.955 -211.645 108.285 -211.315 ;
        RECT 107.955 -213.005 108.285 -212.675 ;
        RECT 107.955 -214.365 108.285 -214.035 ;
        RECT 107.955 -215.725 108.285 -215.395 ;
        RECT 107.955 -217.085 108.285 -216.755 ;
        RECT 107.955 -218.445 108.285 -218.115 ;
        RECT 107.955 -219.805 108.285 -219.475 ;
        RECT 107.955 -221.165 108.285 -220.835 ;
        RECT 107.955 -222.525 108.285 -222.195 ;
        RECT 107.955 -223.885 108.285 -223.555 ;
        RECT 107.955 -225.245 108.285 -224.915 ;
        RECT 107.955 -226.605 108.285 -226.275 ;
        RECT 107.955 -227.965 108.285 -227.635 ;
        RECT 107.955 -229.325 108.285 -228.995 ;
        RECT 107.955 -230.685 108.285 -230.355 ;
        RECT 107.955 -232.045 108.285 -231.715 ;
        RECT 107.955 -233.405 108.285 -233.075 ;
        RECT 107.955 -234.765 108.285 -234.435 ;
        RECT 107.955 -236.125 108.285 -235.795 ;
        RECT 107.955 -237.485 108.285 -237.155 ;
        RECT 107.955 -238.845 108.285 -238.515 ;
        RECT 107.955 -241.09 108.285 -239.96 ;
        RECT 107.96 -241.205 108.28 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 244.04 109.645 245.17 ;
        RECT 109.315 242.595 109.645 242.925 ;
        RECT 109.315 241.235 109.645 241.565 ;
        RECT 109.315 239.875 109.645 240.205 ;
        RECT 109.315 238.515 109.645 238.845 ;
        RECT 109.315 237.155 109.645 237.485 ;
        RECT 109.32 237.155 109.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 -0.845 109.645 -0.515 ;
        RECT 109.315 -2.205 109.645 -1.875 ;
        RECT 109.315 -3.565 109.645 -3.235 ;
        RECT 109.32 -3.565 109.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 -123.245 109.645 -122.915 ;
        RECT 109.315 -124.605 109.645 -124.275 ;
        RECT 109.315 -125.965 109.645 -125.635 ;
        RECT 109.315 -127.325 109.645 -126.995 ;
        RECT 109.315 -128.685 109.645 -128.355 ;
        RECT 109.315 -130.045 109.645 -129.715 ;
        RECT 109.315 -131.405 109.645 -131.075 ;
        RECT 109.315 -132.765 109.645 -132.435 ;
        RECT 109.315 -134.125 109.645 -133.795 ;
        RECT 109.315 -135.485 109.645 -135.155 ;
        RECT 109.315 -136.845 109.645 -136.515 ;
        RECT 109.315 -138.205 109.645 -137.875 ;
        RECT 109.315 -139.565 109.645 -139.235 ;
        RECT 109.315 -140.925 109.645 -140.595 ;
        RECT 109.315 -142.285 109.645 -141.955 ;
        RECT 109.315 -143.645 109.645 -143.315 ;
        RECT 109.315 -145.005 109.645 -144.675 ;
        RECT 109.315 -146.365 109.645 -146.035 ;
        RECT 109.315 -147.725 109.645 -147.395 ;
        RECT 109.315 -149.085 109.645 -148.755 ;
        RECT 109.315 -150.445 109.645 -150.115 ;
        RECT 109.315 -151.805 109.645 -151.475 ;
        RECT 109.315 -153.165 109.645 -152.835 ;
        RECT 109.315 -154.525 109.645 -154.195 ;
        RECT 109.315 -155.885 109.645 -155.555 ;
        RECT 109.315 -157.245 109.645 -156.915 ;
        RECT 109.315 -158.605 109.645 -158.275 ;
        RECT 109.315 -159.965 109.645 -159.635 ;
        RECT 109.315 -161.325 109.645 -160.995 ;
        RECT 109.315 -162.685 109.645 -162.355 ;
        RECT 109.315 -164.045 109.645 -163.715 ;
        RECT 109.315 -165.405 109.645 -165.075 ;
        RECT 109.315 -166.765 109.645 -166.435 ;
        RECT 109.315 -168.125 109.645 -167.795 ;
        RECT 109.315 -169.485 109.645 -169.155 ;
        RECT 109.315 -170.845 109.645 -170.515 ;
        RECT 109.315 -172.205 109.645 -171.875 ;
        RECT 109.315 -173.565 109.645 -173.235 ;
        RECT 109.315 -174.925 109.645 -174.595 ;
        RECT 109.315 -176.285 109.645 -175.955 ;
        RECT 109.315 -177.645 109.645 -177.315 ;
        RECT 109.315 -179.005 109.645 -178.675 ;
        RECT 109.315 -180.365 109.645 -180.035 ;
        RECT 109.315 -181.725 109.645 -181.395 ;
        RECT 109.315 -183.085 109.645 -182.755 ;
        RECT 109.315 -184.445 109.645 -184.115 ;
        RECT 109.315 -185.805 109.645 -185.475 ;
        RECT 109.315 -187.165 109.645 -186.835 ;
        RECT 109.315 -188.525 109.645 -188.195 ;
        RECT 109.315 -189.885 109.645 -189.555 ;
        RECT 109.315 -191.245 109.645 -190.915 ;
        RECT 109.315 -192.605 109.645 -192.275 ;
        RECT 109.315 -193.965 109.645 -193.635 ;
        RECT 109.315 -195.325 109.645 -194.995 ;
        RECT 109.315 -196.685 109.645 -196.355 ;
        RECT 109.315 -198.045 109.645 -197.715 ;
        RECT 109.315 -199.405 109.645 -199.075 ;
        RECT 109.315 -200.765 109.645 -200.435 ;
        RECT 109.315 -202.125 109.645 -201.795 ;
        RECT 109.315 -203.485 109.645 -203.155 ;
        RECT 109.315 -204.845 109.645 -204.515 ;
        RECT 109.315 -206.205 109.645 -205.875 ;
        RECT 109.315 -207.565 109.645 -207.235 ;
        RECT 109.315 -208.925 109.645 -208.595 ;
        RECT 109.315 -210.285 109.645 -209.955 ;
        RECT 109.315 -211.645 109.645 -211.315 ;
        RECT 109.315 -213.005 109.645 -212.675 ;
        RECT 109.315 -214.365 109.645 -214.035 ;
        RECT 109.315 -215.725 109.645 -215.395 ;
        RECT 109.315 -217.085 109.645 -216.755 ;
        RECT 109.315 -218.445 109.645 -218.115 ;
        RECT 109.315 -219.805 109.645 -219.475 ;
        RECT 109.315 -221.165 109.645 -220.835 ;
        RECT 109.315 -222.525 109.645 -222.195 ;
        RECT 109.315 -223.885 109.645 -223.555 ;
        RECT 109.315 -225.245 109.645 -224.915 ;
        RECT 109.315 -226.605 109.645 -226.275 ;
        RECT 109.315 -227.965 109.645 -227.635 ;
        RECT 109.315 -229.325 109.645 -228.995 ;
        RECT 109.315 -230.685 109.645 -230.355 ;
        RECT 109.315 -232.045 109.645 -231.715 ;
        RECT 109.315 -233.405 109.645 -233.075 ;
        RECT 109.315 -234.765 109.645 -234.435 ;
        RECT 109.315 -236.125 109.645 -235.795 ;
        RECT 109.315 -237.485 109.645 -237.155 ;
        RECT 109.315 -238.845 109.645 -238.515 ;
        RECT 109.315 -241.09 109.645 -239.96 ;
        RECT 109.32 -241.205 109.64 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 244.04 111.005 245.17 ;
        RECT 110.675 242.595 111.005 242.925 ;
        RECT 110.675 241.235 111.005 241.565 ;
        RECT 110.675 239.875 111.005 240.205 ;
        RECT 110.675 238.515 111.005 238.845 ;
        RECT 110.675 237.155 111.005 237.485 ;
        RECT 110.68 237.155 111 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -0.845 111.005 -0.515 ;
        RECT 110.675 -2.205 111.005 -1.875 ;
        RECT 110.675 -3.565 111.005 -3.235 ;
        RECT 110.68 -3.565 111 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -215.725 111.005 -215.395 ;
        RECT 110.675 -217.085 111.005 -216.755 ;
        RECT 110.675 -218.445 111.005 -218.115 ;
        RECT 110.675 -219.805 111.005 -219.475 ;
        RECT 110.675 -221.165 111.005 -220.835 ;
        RECT 110.675 -222.525 111.005 -222.195 ;
        RECT 110.675 -223.885 111.005 -223.555 ;
        RECT 110.675 -225.245 111.005 -224.915 ;
        RECT 110.675 -226.605 111.005 -226.275 ;
        RECT 110.675 -227.965 111.005 -227.635 ;
        RECT 110.675 -229.325 111.005 -228.995 ;
        RECT 110.675 -230.685 111.005 -230.355 ;
        RECT 110.675 -232.045 111.005 -231.715 ;
        RECT 110.675 -233.405 111.005 -233.075 ;
        RECT 110.675 -234.765 111.005 -234.435 ;
        RECT 110.675 -236.125 111.005 -235.795 ;
        RECT 110.675 -237.485 111.005 -237.155 ;
        RECT 110.675 -238.845 111.005 -238.515 ;
        RECT 110.675 -241.09 111.005 -239.96 ;
        RECT 110.68 -241.205 111 -122.24 ;
        RECT 110.675 -123.245 111.005 -122.915 ;
        RECT 110.675 -124.605 111.005 -124.275 ;
        RECT 110.675 -125.965 111.005 -125.635 ;
        RECT 110.675 -127.325 111.005 -126.995 ;
        RECT 110.675 -128.685 111.005 -128.355 ;
        RECT 110.675 -130.045 111.005 -129.715 ;
        RECT 110.675 -131.405 111.005 -131.075 ;
        RECT 110.675 -132.765 111.005 -132.435 ;
        RECT 110.675 -134.125 111.005 -133.795 ;
        RECT 110.675 -135.485 111.005 -135.155 ;
        RECT 110.675 -136.845 111.005 -136.515 ;
        RECT 110.675 -138.205 111.005 -137.875 ;
        RECT 110.675 -139.565 111.005 -139.235 ;
        RECT 110.675 -140.925 111.005 -140.595 ;
        RECT 110.675 -142.285 111.005 -141.955 ;
        RECT 110.675 -143.645 111.005 -143.315 ;
        RECT 110.675 -145.005 111.005 -144.675 ;
        RECT 110.675 -146.365 111.005 -146.035 ;
        RECT 110.675 -147.725 111.005 -147.395 ;
        RECT 110.675 -149.085 111.005 -148.755 ;
        RECT 110.675 -150.445 111.005 -150.115 ;
        RECT 110.675 -151.805 111.005 -151.475 ;
        RECT 110.675 -153.165 111.005 -152.835 ;
        RECT 110.675 -154.525 111.005 -154.195 ;
        RECT 110.675 -155.885 111.005 -155.555 ;
        RECT 110.675 -157.245 111.005 -156.915 ;
        RECT 110.675 -158.605 111.005 -158.275 ;
        RECT 110.675 -159.965 111.005 -159.635 ;
        RECT 110.675 -161.325 111.005 -160.995 ;
        RECT 110.675 -162.685 111.005 -162.355 ;
        RECT 110.675 -164.045 111.005 -163.715 ;
        RECT 110.675 -165.405 111.005 -165.075 ;
        RECT 110.675 -166.765 111.005 -166.435 ;
        RECT 110.675 -168.125 111.005 -167.795 ;
        RECT 110.675 -169.485 111.005 -169.155 ;
        RECT 110.675 -170.845 111.005 -170.515 ;
        RECT 110.675 -172.205 111.005 -171.875 ;
        RECT 110.675 -173.565 111.005 -173.235 ;
        RECT 110.675 -174.925 111.005 -174.595 ;
        RECT 110.675 -176.285 111.005 -175.955 ;
        RECT 110.675 -177.645 111.005 -177.315 ;
        RECT 110.675 -179.005 111.005 -178.675 ;
        RECT 110.675 -180.365 111.005 -180.035 ;
        RECT 110.675 -181.725 111.005 -181.395 ;
        RECT 110.675 -183.085 111.005 -182.755 ;
        RECT 110.675 -184.445 111.005 -184.115 ;
        RECT 110.675 -185.805 111.005 -185.475 ;
        RECT 110.675 -187.165 111.005 -186.835 ;
        RECT 110.675 -188.525 111.005 -188.195 ;
        RECT 110.675 -189.885 111.005 -189.555 ;
        RECT 110.675 -191.245 111.005 -190.915 ;
        RECT 110.675 -192.605 111.005 -192.275 ;
        RECT 110.675 -193.965 111.005 -193.635 ;
        RECT 110.675 -195.325 111.005 -194.995 ;
        RECT 110.675 -196.685 111.005 -196.355 ;
        RECT 110.675 -198.045 111.005 -197.715 ;
        RECT 110.675 -199.405 111.005 -199.075 ;
        RECT 110.675 -200.765 111.005 -200.435 ;
        RECT 110.675 -202.125 111.005 -201.795 ;
        RECT 110.675 -203.485 111.005 -203.155 ;
        RECT 110.675 -204.845 111.005 -204.515 ;
        RECT 110.675 -206.205 111.005 -205.875 ;
        RECT 110.675 -207.565 111.005 -207.235 ;
        RECT 110.675 -208.925 111.005 -208.595 ;
        RECT 110.675 -210.285 111.005 -209.955 ;
        RECT 110.675 -211.645 111.005 -211.315 ;
        RECT 110.675 -213.005 111.005 -212.675 ;
        RECT 110.675 -214.365 111.005 -214.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 244.04 77.005 245.17 ;
        RECT 76.675 242.595 77.005 242.925 ;
        RECT 76.675 241.235 77.005 241.565 ;
        RECT 76.675 239.875 77.005 240.205 ;
        RECT 76.675 238.515 77.005 238.845 ;
        RECT 76.675 237.155 77.005 237.485 ;
        RECT 76.68 237.155 77 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 -0.845 77.005 -0.515 ;
        RECT 76.675 -2.205 77.005 -1.875 ;
        RECT 76.675 -3.565 77.005 -3.235 ;
        RECT 76.68 -3.565 77 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 -123.245 77.005 -122.915 ;
        RECT 76.675 -124.605 77.005 -124.275 ;
        RECT 76.675 -125.965 77.005 -125.635 ;
        RECT 76.675 -127.325 77.005 -126.995 ;
        RECT 76.675 -128.685 77.005 -128.355 ;
        RECT 76.675 -130.045 77.005 -129.715 ;
        RECT 76.675 -131.405 77.005 -131.075 ;
        RECT 76.675 -132.765 77.005 -132.435 ;
        RECT 76.675 -134.125 77.005 -133.795 ;
        RECT 76.675 -135.485 77.005 -135.155 ;
        RECT 76.675 -136.845 77.005 -136.515 ;
        RECT 76.675 -138.205 77.005 -137.875 ;
        RECT 76.675 -139.565 77.005 -139.235 ;
        RECT 76.675 -140.925 77.005 -140.595 ;
        RECT 76.675 -142.285 77.005 -141.955 ;
        RECT 76.675 -143.645 77.005 -143.315 ;
        RECT 76.675 -145.005 77.005 -144.675 ;
        RECT 76.675 -146.365 77.005 -146.035 ;
        RECT 76.675 -147.725 77.005 -147.395 ;
        RECT 76.675 -149.085 77.005 -148.755 ;
        RECT 76.675 -150.445 77.005 -150.115 ;
        RECT 76.675 -151.805 77.005 -151.475 ;
        RECT 76.675 -153.165 77.005 -152.835 ;
        RECT 76.675 -154.525 77.005 -154.195 ;
        RECT 76.675 -155.885 77.005 -155.555 ;
        RECT 76.675 -157.245 77.005 -156.915 ;
        RECT 76.675 -158.605 77.005 -158.275 ;
        RECT 76.675 -159.965 77.005 -159.635 ;
        RECT 76.675 -161.325 77.005 -160.995 ;
        RECT 76.675 -162.685 77.005 -162.355 ;
        RECT 76.675 -164.045 77.005 -163.715 ;
        RECT 76.675 -165.405 77.005 -165.075 ;
        RECT 76.675 -166.765 77.005 -166.435 ;
        RECT 76.675 -168.125 77.005 -167.795 ;
        RECT 76.675 -169.485 77.005 -169.155 ;
        RECT 76.675 -170.845 77.005 -170.515 ;
        RECT 76.675 -172.205 77.005 -171.875 ;
        RECT 76.675 -173.565 77.005 -173.235 ;
        RECT 76.675 -174.925 77.005 -174.595 ;
        RECT 76.675 -176.285 77.005 -175.955 ;
        RECT 76.675 -177.645 77.005 -177.315 ;
        RECT 76.675 -179.005 77.005 -178.675 ;
        RECT 76.675 -180.365 77.005 -180.035 ;
        RECT 76.675 -181.725 77.005 -181.395 ;
        RECT 76.675 -183.085 77.005 -182.755 ;
        RECT 76.675 -184.445 77.005 -184.115 ;
        RECT 76.675 -185.805 77.005 -185.475 ;
        RECT 76.675 -187.165 77.005 -186.835 ;
        RECT 76.675 -188.525 77.005 -188.195 ;
        RECT 76.675 -189.885 77.005 -189.555 ;
        RECT 76.675 -191.245 77.005 -190.915 ;
        RECT 76.675 -192.605 77.005 -192.275 ;
        RECT 76.675 -193.965 77.005 -193.635 ;
        RECT 76.675 -195.325 77.005 -194.995 ;
        RECT 76.675 -196.685 77.005 -196.355 ;
        RECT 76.675 -198.045 77.005 -197.715 ;
        RECT 76.675 -199.405 77.005 -199.075 ;
        RECT 76.675 -200.765 77.005 -200.435 ;
        RECT 76.675 -202.125 77.005 -201.795 ;
        RECT 76.675 -203.485 77.005 -203.155 ;
        RECT 76.675 -204.845 77.005 -204.515 ;
        RECT 76.675 -206.205 77.005 -205.875 ;
        RECT 76.675 -207.565 77.005 -207.235 ;
        RECT 76.675 -208.925 77.005 -208.595 ;
        RECT 76.675 -210.285 77.005 -209.955 ;
        RECT 76.675 -211.645 77.005 -211.315 ;
        RECT 76.675 -213.005 77.005 -212.675 ;
        RECT 76.675 -214.365 77.005 -214.035 ;
        RECT 76.675 -215.725 77.005 -215.395 ;
        RECT 76.675 -217.085 77.005 -216.755 ;
        RECT 76.675 -218.445 77.005 -218.115 ;
        RECT 76.675 -219.805 77.005 -219.475 ;
        RECT 76.675 -221.165 77.005 -220.835 ;
        RECT 76.675 -222.525 77.005 -222.195 ;
        RECT 76.675 -223.885 77.005 -223.555 ;
        RECT 76.675 -225.245 77.005 -224.915 ;
        RECT 76.675 -226.605 77.005 -226.275 ;
        RECT 76.675 -227.965 77.005 -227.635 ;
        RECT 76.675 -229.325 77.005 -228.995 ;
        RECT 76.675 -230.685 77.005 -230.355 ;
        RECT 76.675 -232.045 77.005 -231.715 ;
        RECT 76.675 -233.405 77.005 -233.075 ;
        RECT 76.675 -234.765 77.005 -234.435 ;
        RECT 76.675 -236.125 77.005 -235.795 ;
        RECT 76.675 -237.485 77.005 -237.155 ;
        RECT 76.675 -238.845 77.005 -238.515 ;
        RECT 76.675 -241.09 77.005 -239.96 ;
        RECT 76.68 -241.205 77 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 244.04 78.365 245.17 ;
        RECT 78.035 242.595 78.365 242.925 ;
        RECT 78.035 241.235 78.365 241.565 ;
        RECT 78.035 239.875 78.365 240.205 ;
        RECT 78.035 238.515 78.365 238.845 ;
        RECT 78.035 237.155 78.365 237.485 ;
        RECT 78.04 237.155 78.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -0.845 78.365 -0.515 ;
        RECT 78.035 -2.205 78.365 -1.875 ;
        RECT 78.035 -3.565 78.365 -3.235 ;
        RECT 78.04 -3.565 78.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -123.245 78.365 -122.915 ;
        RECT 78.035 -124.605 78.365 -124.275 ;
        RECT 78.035 -125.965 78.365 -125.635 ;
        RECT 78.035 -127.325 78.365 -126.995 ;
        RECT 78.035 -128.685 78.365 -128.355 ;
        RECT 78.035 -130.045 78.365 -129.715 ;
        RECT 78.035 -131.405 78.365 -131.075 ;
        RECT 78.035 -132.765 78.365 -132.435 ;
        RECT 78.035 -134.125 78.365 -133.795 ;
        RECT 78.035 -135.485 78.365 -135.155 ;
        RECT 78.035 -136.845 78.365 -136.515 ;
        RECT 78.035 -138.205 78.365 -137.875 ;
        RECT 78.035 -139.565 78.365 -139.235 ;
        RECT 78.035 -140.925 78.365 -140.595 ;
        RECT 78.035 -142.285 78.365 -141.955 ;
        RECT 78.035 -143.645 78.365 -143.315 ;
        RECT 78.035 -145.005 78.365 -144.675 ;
        RECT 78.035 -146.365 78.365 -146.035 ;
        RECT 78.035 -147.725 78.365 -147.395 ;
        RECT 78.035 -149.085 78.365 -148.755 ;
        RECT 78.035 -150.445 78.365 -150.115 ;
        RECT 78.035 -151.805 78.365 -151.475 ;
        RECT 78.035 -153.165 78.365 -152.835 ;
        RECT 78.035 -154.525 78.365 -154.195 ;
        RECT 78.035 -155.885 78.365 -155.555 ;
        RECT 78.035 -157.245 78.365 -156.915 ;
        RECT 78.035 -158.605 78.365 -158.275 ;
        RECT 78.035 -159.965 78.365 -159.635 ;
        RECT 78.035 -161.325 78.365 -160.995 ;
        RECT 78.035 -162.685 78.365 -162.355 ;
        RECT 78.035 -164.045 78.365 -163.715 ;
        RECT 78.035 -165.405 78.365 -165.075 ;
        RECT 78.035 -166.765 78.365 -166.435 ;
        RECT 78.035 -168.125 78.365 -167.795 ;
        RECT 78.035 -169.485 78.365 -169.155 ;
        RECT 78.035 -170.845 78.365 -170.515 ;
        RECT 78.035 -172.205 78.365 -171.875 ;
        RECT 78.035 -173.565 78.365 -173.235 ;
        RECT 78.035 -174.925 78.365 -174.595 ;
        RECT 78.035 -176.285 78.365 -175.955 ;
        RECT 78.035 -177.645 78.365 -177.315 ;
        RECT 78.035 -179.005 78.365 -178.675 ;
        RECT 78.035 -180.365 78.365 -180.035 ;
        RECT 78.035 -181.725 78.365 -181.395 ;
        RECT 78.035 -183.085 78.365 -182.755 ;
        RECT 78.035 -184.445 78.365 -184.115 ;
        RECT 78.035 -185.805 78.365 -185.475 ;
        RECT 78.035 -187.165 78.365 -186.835 ;
        RECT 78.035 -188.525 78.365 -188.195 ;
        RECT 78.035 -189.885 78.365 -189.555 ;
        RECT 78.035 -191.245 78.365 -190.915 ;
        RECT 78.035 -192.605 78.365 -192.275 ;
        RECT 78.035 -193.965 78.365 -193.635 ;
        RECT 78.035 -195.325 78.365 -194.995 ;
        RECT 78.035 -196.685 78.365 -196.355 ;
        RECT 78.035 -198.045 78.365 -197.715 ;
        RECT 78.035 -199.405 78.365 -199.075 ;
        RECT 78.035 -200.765 78.365 -200.435 ;
        RECT 78.035 -202.125 78.365 -201.795 ;
        RECT 78.035 -203.485 78.365 -203.155 ;
        RECT 78.035 -204.845 78.365 -204.515 ;
        RECT 78.035 -206.205 78.365 -205.875 ;
        RECT 78.035 -207.565 78.365 -207.235 ;
        RECT 78.035 -208.925 78.365 -208.595 ;
        RECT 78.035 -210.285 78.365 -209.955 ;
        RECT 78.035 -211.645 78.365 -211.315 ;
        RECT 78.035 -213.005 78.365 -212.675 ;
        RECT 78.035 -214.365 78.365 -214.035 ;
        RECT 78.035 -215.725 78.365 -215.395 ;
        RECT 78.035 -217.085 78.365 -216.755 ;
        RECT 78.035 -218.445 78.365 -218.115 ;
        RECT 78.035 -219.805 78.365 -219.475 ;
        RECT 78.035 -221.165 78.365 -220.835 ;
        RECT 78.035 -222.525 78.365 -222.195 ;
        RECT 78.035 -223.885 78.365 -223.555 ;
        RECT 78.035 -225.245 78.365 -224.915 ;
        RECT 78.035 -226.605 78.365 -226.275 ;
        RECT 78.035 -227.965 78.365 -227.635 ;
        RECT 78.035 -229.325 78.365 -228.995 ;
        RECT 78.035 -230.685 78.365 -230.355 ;
        RECT 78.035 -232.045 78.365 -231.715 ;
        RECT 78.035 -233.405 78.365 -233.075 ;
        RECT 78.035 -234.765 78.365 -234.435 ;
        RECT 78.035 -236.125 78.365 -235.795 ;
        RECT 78.035 -237.485 78.365 -237.155 ;
        RECT 78.035 -238.845 78.365 -238.515 ;
        RECT 78.035 -241.09 78.365 -239.96 ;
        RECT 78.04 -241.205 78.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 244.04 79.725 245.17 ;
        RECT 79.395 242.595 79.725 242.925 ;
        RECT 79.395 241.235 79.725 241.565 ;
        RECT 79.395 239.875 79.725 240.205 ;
        RECT 79.395 238.515 79.725 238.845 ;
        RECT 79.395 237.155 79.725 237.485 ;
        RECT 79.4 237.155 79.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 -127.325 79.725 -126.995 ;
        RECT 79.395 -128.685 79.725 -128.355 ;
        RECT 79.395 -130.045 79.725 -129.715 ;
        RECT 79.395 -131.405 79.725 -131.075 ;
        RECT 79.395 -132.765 79.725 -132.435 ;
        RECT 79.395 -134.125 79.725 -133.795 ;
        RECT 79.395 -135.485 79.725 -135.155 ;
        RECT 79.395 -136.845 79.725 -136.515 ;
        RECT 79.395 -138.205 79.725 -137.875 ;
        RECT 79.395 -139.565 79.725 -139.235 ;
        RECT 79.395 -140.925 79.725 -140.595 ;
        RECT 79.395 -142.285 79.725 -141.955 ;
        RECT 79.395 -143.645 79.725 -143.315 ;
        RECT 79.395 -145.005 79.725 -144.675 ;
        RECT 79.395 -146.365 79.725 -146.035 ;
        RECT 79.395 -147.725 79.725 -147.395 ;
        RECT 79.395 -149.085 79.725 -148.755 ;
        RECT 79.395 -150.445 79.725 -150.115 ;
        RECT 79.395 -151.805 79.725 -151.475 ;
        RECT 79.395 -153.165 79.725 -152.835 ;
        RECT 79.395 -154.525 79.725 -154.195 ;
        RECT 79.395 -155.885 79.725 -155.555 ;
        RECT 79.395 -157.245 79.725 -156.915 ;
        RECT 79.395 -158.605 79.725 -158.275 ;
        RECT 79.395 -159.965 79.725 -159.635 ;
        RECT 79.395 -161.325 79.725 -160.995 ;
        RECT 79.395 -162.685 79.725 -162.355 ;
        RECT 79.395 -164.045 79.725 -163.715 ;
        RECT 79.395 -165.405 79.725 -165.075 ;
        RECT 79.395 -166.765 79.725 -166.435 ;
        RECT 79.395 -168.125 79.725 -167.795 ;
        RECT 79.395 -169.485 79.725 -169.155 ;
        RECT 79.395 -170.845 79.725 -170.515 ;
        RECT 79.395 -172.205 79.725 -171.875 ;
        RECT 79.395 -173.565 79.725 -173.235 ;
        RECT 79.395 -174.925 79.725 -174.595 ;
        RECT 79.395 -176.285 79.725 -175.955 ;
        RECT 79.395 -177.645 79.725 -177.315 ;
        RECT 79.395 -179.005 79.725 -178.675 ;
        RECT 79.395 -180.365 79.725 -180.035 ;
        RECT 79.395 -181.725 79.725 -181.395 ;
        RECT 79.395 -183.085 79.725 -182.755 ;
        RECT 79.395 -184.445 79.725 -184.115 ;
        RECT 79.395 -185.805 79.725 -185.475 ;
        RECT 79.395 -187.165 79.725 -186.835 ;
        RECT 79.395 -188.525 79.725 -188.195 ;
        RECT 79.395 -189.885 79.725 -189.555 ;
        RECT 79.395 -191.245 79.725 -190.915 ;
        RECT 79.395 -192.605 79.725 -192.275 ;
        RECT 79.395 -193.965 79.725 -193.635 ;
        RECT 79.395 -195.325 79.725 -194.995 ;
        RECT 79.395 -196.685 79.725 -196.355 ;
        RECT 79.395 -198.045 79.725 -197.715 ;
        RECT 79.395 -199.405 79.725 -199.075 ;
        RECT 79.395 -200.765 79.725 -200.435 ;
        RECT 79.395 -202.125 79.725 -201.795 ;
        RECT 79.395 -203.485 79.725 -203.155 ;
        RECT 79.395 -204.845 79.725 -204.515 ;
        RECT 79.395 -206.205 79.725 -205.875 ;
        RECT 79.395 -207.565 79.725 -207.235 ;
        RECT 79.395 -208.925 79.725 -208.595 ;
        RECT 79.395 -210.285 79.725 -209.955 ;
        RECT 79.395 -211.645 79.725 -211.315 ;
        RECT 79.395 -213.005 79.725 -212.675 ;
        RECT 79.395 -214.365 79.725 -214.035 ;
        RECT 79.395 -215.725 79.725 -215.395 ;
        RECT 79.395 -217.085 79.725 -216.755 ;
        RECT 79.395 -218.445 79.725 -218.115 ;
        RECT 79.395 -219.805 79.725 -219.475 ;
        RECT 79.395 -221.165 79.725 -220.835 ;
        RECT 79.395 -222.525 79.725 -222.195 ;
        RECT 79.395 -223.885 79.725 -223.555 ;
        RECT 79.395 -225.245 79.725 -224.915 ;
        RECT 79.395 -226.605 79.725 -226.275 ;
        RECT 79.395 -227.965 79.725 -227.635 ;
        RECT 79.395 -229.325 79.725 -228.995 ;
        RECT 79.395 -230.685 79.725 -230.355 ;
        RECT 79.395 -232.045 79.725 -231.715 ;
        RECT 79.395 -233.405 79.725 -233.075 ;
        RECT 79.395 -234.765 79.725 -234.435 ;
        RECT 79.395 -236.125 79.725 -235.795 ;
        RECT 79.395 -237.485 79.725 -237.155 ;
        RECT 79.395 -238.845 79.725 -238.515 ;
        RECT 79.395 -241.09 79.725 -239.96 ;
        RECT 79.4 -241.205 79.72 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.61 -125.535 79.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 244.04 81.085 245.17 ;
        RECT 80.755 242.595 81.085 242.925 ;
        RECT 80.755 241.235 81.085 241.565 ;
        RECT 80.755 239.875 81.085 240.205 ;
        RECT 80.755 238.515 81.085 238.845 ;
        RECT 80.755 237.155 81.085 237.485 ;
        RECT 80.76 237.155 81.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 -0.845 81.085 -0.515 ;
        RECT 80.755 -2.205 81.085 -1.875 ;
        RECT 80.755 -3.565 81.085 -3.235 ;
        RECT 80.76 -3.565 81.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 244.04 82.445 245.17 ;
        RECT 82.115 242.595 82.445 242.925 ;
        RECT 82.115 241.235 82.445 241.565 ;
        RECT 82.115 239.875 82.445 240.205 ;
        RECT 82.115 238.515 82.445 238.845 ;
        RECT 82.115 237.155 82.445 237.485 ;
        RECT 82.12 237.155 82.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 -0.845 82.445 -0.515 ;
        RECT 82.115 -2.205 82.445 -1.875 ;
        RECT 82.115 -3.565 82.445 -3.235 ;
        RECT 82.12 -3.565 82.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 244.04 83.805 245.17 ;
        RECT 83.475 242.595 83.805 242.925 ;
        RECT 83.475 241.235 83.805 241.565 ;
        RECT 83.475 239.875 83.805 240.205 ;
        RECT 83.475 238.515 83.805 238.845 ;
        RECT 83.475 237.155 83.805 237.485 ;
        RECT 83.48 237.155 83.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 -0.845 83.805 -0.515 ;
        RECT 83.475 -2.205 83.805 -1.875 ;
        RECT 83.475 -3.565 83.805 -3.235 ;
        RECT 83.48 -3.565 83.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 -123.245 83.805 -122.915 ;
        RECT 83.475 -124.605 83.805 -124.275 ;
        RECT 83.475 -125.965 83.805 -125.635 ;
        RECT 83.475 -127.325 83.805 -126.995 ;
        RECT 83.475 -128.685 83.805 -128.355 ;
        RECT 83.475 -130.045 83.805 -129.715 ;
        RECT 83.475 -131.405 83.805 -131.075 ;
        RECT 83.475 -132.765 83.805 -132.435 ;
        RECT 83.475 -134.125 83.805 -133.795 ;
        RECT 83.475 -135.485 83.805 -135.155 ;
        RECT 83.475 -136.845 83.805 -136.515 ;
        RECT 83.475 -138.205 83.805 -137.875 ;
        RECT 83.475 -139.565 83.805 -139.235 ;
        RECT 83.475 -140.925 83.805 -140.595 ;
        RECT 83.475 -142.285 83.805 -141.955 ;
        RECT 83.475 -143.645 83.805 -143.315 ;
        RECT 83.475 -145.005 83.805 -144.675 ;
        RECT 83.475 -146.365 83.805 -146.035 ;
        RECT 83.475 -147.725 83.805 -147.395 ;
        RECT 83.475 -149.085 83.805 -148.755 ;
        RECT 83.475 -150.445 83.805 -150.115 ;
        RECT 83.475 -151.805 83.805 -151.475 ;
        RECT 83.475 -153.165 83.805 -152.835 ;
        RECT 83.475 -154.525 83.805 -154.195 ;
        RECT 83.475 -155.885 83.805 -155.555 ;
        RECT 83.475 -157.245 83.805 -156.915 ;
        RECT 83.475 -158.605 83.805 -158.275 ;
        RECT 83.475 -159.965 83.805 -159.635 ;
        RECT 83.475 -161.325 83.805 -160.995 ;
        RECT 83.475 -162.685 83.805 -162.355 ;
        RECT 83.475 -164.045 83.805 -163.715 ;
        RECT 83.475 -165.405 83.805 -165.075 ;
        RECT 83.475 -166.765 83.805 -166.435 ;
        RECT 83.475 -168.125 83.805 -167.795 ;
        RECT 83.475 -169.485 83.805 -169.155 ;
        RECT 83.475 -170.845 83.805 -170.515 ;
        RECT 83.475 -172.205 83.805 -171.875 ;
        RECT 83.475 -173.565 83.805 -173.235 ;
        RECT 83.475 -174.925 83.805 -174.595 ;
        RECT 83.475 -176.285 83.805 -175.955 ;
        RECT 83.475 -177.645 83.805 -177.315 ;
        RECT 83.475 -179.005 83.805 -178.675 ;
        RECT 83.475 -180.365 83.805 -180.035 ;
        RECT 83.475 -181.725 83.805 -181.395 ;
        RECT 83.475 -183.085 83.805 -182.755 ;
        RECT 83.475 -184.445 83.805 -184.115 ;
        RECT 83.475 -185.805 83.805 -185.475 ;
        RECT 83.475 -187.165 83.805 -186.835 ;
        RECT 83.475 -188.525 83.805 -188.195 ;
        RECT 83.475 -189.885 83.805 -189.555 ;
        RECT 83.475 -191.245 83.805 -190.915 ;
        RECT 83.475 -192.605 83.805 -192.275 ;
        RECT 83.475 -193.965 83.805 -193.635 ;
        RECT 83.475 -195.325 83.805 -194.995 ;
        RECT 83.475 -196.685 83.805 -196.355 ;
        RECT 83.475 -198.045 83.805 -197.715 ;
        RECT 83.475 -199.405 83.805 -199.075 ;
        RECT 83.475 -200.765 83.805 -200.435 ;
        RECT 83.475 -202.125 83.805 -201.795 ;
        RECT 83.475 -203.485 83.805 -203.155 ;
        RECT 83.475 -204.845 83.805 -204.515 ;
        RECT 83.475 -206.205 83.805 -205.875 ;
        RECT 83.475 -207.565 83.805 -207.235 ;
        RECT 83.475 -208.925 83.805 -208.595 ;
        RECT 83.475 -210.285 83.805 -209.955 ;
        RECT 83.475 -211.645 83.805 -211.315 ;
        RECT 83.475 -213.005 83.805 -212.675 ;
        RECT 83.475 -214.365 83.805 -214.035 ;
        RECT 83.475 -215.725 83.805 -215.395 ;
        RECT 83.475 -217.085 83.805 -216.755 ;
        RECT 83.475 -218.445 83.805 -218.115 ;
        RECT 83.475 -219.805 83.805 -219.475 ;
        RECT 83.475 -221.165 83.805 -220.835 ;
        RECT 83.475 -222.525 83.805 -222.195 ;
        RECT 83.475 -223.885 83.805 -223.555 ;
        RECT 83.475 -225.245 83.805 -224.915 ;
        RECT 83.475 -226.605 83.805 -226.275 ;
        RECT 83.475 -227.965 83.805 -227.635 ;
        RECT 83.475 -229.325 83.805 -228.995 ;
        RECT 83.475 -230.685 83.805 -230.355 ;
        RECT 83.475 -232.045 83.805 -231.715 ;
        RECT 83.475 -233.405 83.805 -233.075 ;
        RECT 83.475 -234.765 83.805 -234.435 ;
        RECT 83.475 -236.125 83.805 -235.795 ;
        RECT 83.475 -237.485 83.805 -237.155 ;
        RECT 83.475 -238.845 83.805 -238.515 ;
        RECT 83.475 -241.09 83.805 -239.96 ;
        RECT 83.48 -241.205 83.8 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 244.04 85.165 245.17 ;
        RECT 84.835 242.595 85.165 242.925 ;
        RECT 84.835 241.235 85.165 241.565 ;
        RECT 84.835 239.875 85.165 240.205 ;
        RECT 84.835 238.515 85.165 238.845 ;
        RECT 84.835 237.155 85.165 237.485 ;
        RECT 84.84 237.155 85.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 -0.845 85.165 -0.515 ;
        RECT 84.835 -2.205 85.165 -1.875 ;
        RECT 84.835 -3.565 85.165 -3.235 ;
        RECT 84.84 -3.565 85.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 -123.245 85.165 -122.915 ;
        RECT 84.835 -124.605 85.165 -124.275 ;
        RECT 84.835 -125.965 85.165 -125.635 ;
        RECT 84.835 -127.325 85.165 -126.995 ;
        RECT 84.835 -128.685 85.165 -128.355 ;
        RECT 84.835 -130.045 85.165 -129.715 ;
        RECT 84.835 -131.405 85.165 -131.075 ;
        RECT 84.835 -132.765 85.165 -132.435 ;
        RECT 84.835 -134.125 85.165 -133.795 ;
        RECT 84.835 -135.485 85.165 -135.155 ;
        RECT 84.835 -136.845 85.165 -136.515 ;
        RECT 84.835 -138.205 85.165 -137.875 ;
        RECT 84.835 -139.565 85.165 -139.235 ;
        RECT 84.835 -140.925 85.165 -140.595 ;
        RECT 84.835 -142.285 85.165 -141.955 ;
        RECT 84.835 -143.645 85.165 -143.315 ;
        RECT 84.835 -145.005 85.165 -144.675 ;
        RECT 84.835 -146.365 85.165 -146.035 ;
        RECT 84.835 -147.725 85.165 -147.395 ;
        RECT 84.835 -149.085 85.165 -148.755 ;
        RECT 84.835 -150.445 85.165 -150.115 ;
        RECT 84.835 -151.805 85.165 -151.475 ;
        RECT 84.835 -153.165 85.165 -152.835 ;
        RECT 84.835 -154.525 85.165 -154.195 ;
        RECT 84.835 -155.885 85.165 -155.555 ;
        RECT 84.835 -157.245 85.165 -156.915 ;
        RECT 84.835 -158.605 85.165 -158.275 ;
        RECT 84.835 -159.965 85.165 -159.635 ;
        RECT 84.835 -161.325 85.165 -160.995 ;
        RECT 84.835 -162.685 85.165 -162.355 ;
        RECT 84.835 -164.045 85.165 -163.715 ;
        RECT 84.835 -165.405 85.165 -165.075 ;
        RECT 84.835 -166.765 85.165 -166.435 ;
        RECT 84.835 -168.125 85.165 -167.795 ;
        RECT 84.835 -169.485 85.165 -169.155 ;
        RECT 84.835 -170.845 85.165 -170.515 ;
        RECT 84.835 -172.205 85.165 -171.875 ;
        RECT 84.835 -173.565 85.165 -173.235 ;
        RECT 84.835 -174.925 85.165 -174.595 ;
        RECT 84.835 -176.285 85.165 -175.955 ;
        RECT 84.835 -177.645 85.165 -177.315 ;
        RECT 84.835 -179.005 85.165 -178.675 ;
        RECT 84.835 -180.365 85.165 -180.035 ;
        RECT 84.835 -181.725 85.165 -181.395 ;
        RECT 84.835 -183.085 85.165 -182.755 ;
        RECT 84.835 -184.445 85.165 -184.115 ;
        RECT 84.835 -185.805 85.165 -185.475 ;
        RECT 84.835 -187.165 85.165 -186.835 ;
        RECT 84.835 -188.525 85.165 -188.195 ;
        RECT 84.835 -189.885 85.165 -189.555 ;
        RECT 84.835 -191.245 85.165 -190.915 ;
        RECT 84.835 -192.605 85.165 -192.275 ;
        RECT 84.835 -193.965 85.165 -193.635 ;
        RECT 84.835 -195.325 85.165 -194.995 ;
        RECT 84.835 -196.685 85.165 -196.355 ;
        RECT 84.835 -198.045 85.165 -197.715 ;
        RECT 84.835 -199.405 85.165 -199.075 ;
        RECT 84.835 -200.765 85.165 -200.435 ;
        RECT 84.835 -202.125 85.165 -201.795 ;
        RECT 84.835 -203.485 85.165 -203.155 ;
        RECT 84.835 -204.845 85.165 -204.515 ;
        RECT 84.835 -206.205 85.165 -205.875 ;
        RECT 84.835 -207.565 85.165 -207.235 ;
        RECT 84.835 -208.925 85.165 -208.595 ;
        RECT 84.835 -210.285 85.165 -209.955 ;
        RECT 84.835 -211.645 85.165 -211.315 ;
        RECT 84.835 -213.005 85.165 -212.675 ;
        RECT 84.835 -214.365 85.165 -214.035 ;
        RECT 84.835 -215.725 85.165 -215.395 ;
        RECT 84.835 -217.085 85.165 -216.755 ;
        RECT 84.835 -218.445 85.165 -218.115 ;
        RECT 84.835 -219.805 85.165 -219.475 ;
        RECT 84.835 -221.165 85.165 -220.835 ;
        RECT 84.835 -222.525 85.165 -222.195 ;
        RECT 84.835 -223.885 85.165 -223.555 ;
        RECT 84.835 -225.245 85.165 -224.915 ;
        RECT 84.835 -226.605 85.165 -226.275 ;
        RECT 84.835 -227.965 85.165 -227.635 ;
        RECT 84.835 -229.325 85.165 -228.995 ;
        RECT 84.835 -230.685 85.165 -230.355 ;
        RECT 84.835 -232.045 85.165 -231.715 ;
        RECT 84.835 -233.405 85.165 -233.075 ;
        RECT 84.835 -234.765 85.165 -234.435 ;
        RECT 84.835 -236.125 85.165 -235.795 ;
        RECT 84.835 -237.485 85.165 -237.155 ;
        RECT 84.835 -238.845 85.165 -238.515 ;
        RECT 84.835 -241.09 85.165 -239.96 ;
        RECT 84.84 -241.205 85.16 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 244.04 86.525 245.17 ;
        RECT 86.195 242.595 86.525 242.925 ;
        RECT 86.195 241.235 86.525 241.565 ;
        RECT 86.195 239.875 86.525 240.205 ;
        RECT 86.195 238.515 86.525 238.845 ;
        RECT 86.195 237.155 86.525 237.485 ;
        RECT 86.2 237.155 86.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -0.845 86.525 -0.515 ;
        RECT 86.195 -2.205 86.525 -1.875 ;
        RECT 86.195 -3.565 86.525 -3.235 ;
        RECT 86.2 -3.565 86.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -123.245 86.525 -122.915 ;
        RECT 86.195 -124.605 86.525 -124.275 ;
        RECT 86.195 -125.965 86.525 -125.635 ;
        RECT 86.195 -127.325 86.525 -126.995 ;
        RECT 86.195 -128.685 86.525 -128.355 ;
        RECT 86.195 -130.045 86.525 -129.715 ;
        RECT 86.195 -131.405 86.525 -131.075 ;
        RECT 86.195 -132.765 86.525 -132.435 ;
        RECT 86.195 -134.125 86.525 -133.795 ;
        RECT 86.195 -135.485 86.525 -135.155 ;
        RECT 86.195 -136.845 86.525 -136.515 ;
        RECT 86.195 -138.205 86.525 -137.875 ;
        RECT 86.195 -139.565 86.525 -139.235 ;
        RECT 86.195 -140.925 86.525 -140.595 ;
        RECT 86.195 -142.285 86.525 -141.955 ;
        RECT 86.195 -143.645 86.525 -143.315 ;
        RECT 86.195 -145.005 86.525 -144.675 ;
        RECT 86.195 -146.365 86.525 -146.035 ;
        RECT 86.195 -147.725 86.525 -147.395 ;
        RECT 86.195 -149.085 86.525 -148.755 ;
        RECT 86.195 -150.445 86.525 -150.115 ;
        RECT 86.195 -151.805 86.525 -151.475 ;
        RECT 86.195 -153.165 86.525 -152.835 ;
        RECT 86.195 -154.525 86.525 -154.195 ;
        RECT 86.195 -155.885 86.525 -155.555 ;
        RECT 86.195 -157.245 86.525 -156.915 ;
        RECT 86.195 -158.605 86.525 -158.275 ;
        RECT 86.195 -159.965 86.525 -159.635 ;
        RECT 86.195 -161.325 86.525 -160.995 ;
        RECT 86.195 -162.685 86.525 -162.355 ;
        RECT 86.195 -164.045 86.525 -163.715 ;
        RECT 86.195 -165.405 86.525 -165.075 ;
        RECT 86.195 -166.765 86.525 -166.435 ;
        RECT 86.195 -168.125 86.525 -167.795 ;
        RECT 86.195 -169.485 86.525 -169.155 ;
        RECT 86.195 -170.845 86.525 -170.515 ;
        RECT 86.195 -172.205 86.525 -171.875 ;
        RECT 86.195 -173.565 86.525 -173.235 ;
        RECT 86.195 -174.925 86.525 -174.595 ;
        RECT 86.195 -176.285 86.525 -175.955 ;
        RECT 86.195 -177.645 86.525 -177.315 ;
        RECT 86.195 -179.005 86.525 -178.675 ;
        RECT 86.195 -180.365 86.525 -180.035 ;
        RECT 86.195 -181.725 86.525 -181.395 ;
        RECT 86.195 -183.085 86.525 -182.755 ;
        RECT 86.195 -184.445 86.525 -184.115 ;
        RECT 86.195 -185.805 86.525 -185.475 ;
        RECT 86.195 -187.165 86.525 -186.835 ;
        RECT 86.195 -188.525 86.525 -188.195 ;
        RECT 86.195 -189.885 86.525 -189.555 ;
        RECT 86.195 -191.245 86.525 -190.915 ;
        RECT 86.195 -192.605 86.525 -192.275 ;
        RECT 86.195 -193.965 86.525 -193.635 ;
        RECT 86.195 -195.325 86.525 -194.995 ;
        RECT 86.195 -196.685 86.525 -196.355 ;
        RECT 86.195 -198.045 86.525 -197.715 ;
        RECT 86.195 -199.405 86.525 -199.075 ;
        RECT 86.195 -200.765 86.525 -200.435 ;
        RECT 86.195 -202.125 86.525 -201.795 ;
        RECT 86.195 -203.485 86.525 -203.155 ;
        RECT 86.195 -204.845 86.525 -204.515 ;
        RECT 86.195 -206.205 86.525 -205.875 ;
        RECT 86.195 -207.565 86.525 -207.235 ;
        RECT 86.195 -208.925 86.525 -208.595 ;
        RECT 86.195 -210.285 86.525 -209.955 ;
        RECT 86.195 -211.645 86.525 -211.315 ;
        RECT 86.195 -213.005 86.525 -212.675 ;
        RECT 86.195 -214.365 86.525 -214.035 ;
        RECT 86.195 -215.725 86.525 -215.395 ;
        RECT 86.195 -217.085 86.525 -216.755 ;
        RECT 86.195 -218.445 86.525 -218.115 ;
        RECT 86.195 -219.805 86.525 -219.475 ;
        RECT 86.195 -221.165 86.525 -220.835 ;
        RECT 86.195 -222.525 86.525 -222.195 ;
        RECT 86.195 -223.885 86.525 -223.555 ;
        RECT 86.195 -225.245 86.525 -224.915 ;
        RECT 86.195 -226.605 86.525 -226.275 ;
        RECT 86.195 -227.965 86.525 -227.635 ;
        RECT 86.195 -229.325 86.525 -228.995 ;
        RECT 86.195 -230.685 86.525 -230.355 ;
        RECT 86.195 -232.045 86.525 -231.715 ;
        RECT 86.195 -233.405 86.525 -233.075 ;
        RECT 86.195 -234.765 86.525 -234.435 ;
        RECT 86.195 -236.125 86.525 -235.795 ;
        RECT 86.195 -237.485 86.525 -237.155 ;
        RECT 86.195 -238.845 86.525 -238.515 ;
        RECT 86.195 -241.09 86.525 -239.96 ;
        RECT 86.2 -241.205 86.52 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 244.04 87.885 245.17 ;
        RECT 87.555 242.595 87.885 242.925 ;
        RECT 87.555 241.235 87.885 241.565 ;
        RECT 87.555 239.875 87.885 240.205 ;
        RECT 87.555 238.515 87.885 238.845 ;
        RECT 87.555 237.155 87.885 237.485 ;
        RECT 87.56 237.155 87.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 -0.845 87.885 -0.515 ;
        RECT 87.555 -2.205 87.885 -1.875 ;
        RECT 87.555 -3.565 87.885 -3.235 ;
        RECT 87.56 -3.565 87.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 -123.245 87.885 -122.915 ;
        RECT 87.555 -124.605 87.885 -124.275 ;
        RECT 87.555 -125.965 87.885 -125.635 ;
        RECT 87.555 -127.325 87.885 -126.995 ;
        RECT 87.555 -128.685 87.885 -128.355 ;
        RECT 87.555 -130.045 87.885 -129.715 ;
        RECT 87.555 -131.405 87.885 -131.075 ;
        RECT 87.555 -132.765 87.885 -132.435 ;
        RECT 87.555 -134.125 87.885 -133.795 ;
        RECT 87.555 -135.485 87.885 -135.155 ;
        RECT 87.555 -136.845 87.885 -136.515 ;
        RECT 87.555 -138.205 87.885 -137.875 ;
        RECT 87.555 -139.565 87.885 -139.235 ;
        RECT 87.555 -140.925 87.885 -140.595 ;
        RECT 87.555 -142.285 87.885 -141.955 ;
        RECT 87.555 -143.645 87.885 -143.315 ;
        RECT 87.555 -145.005 87.885 -144.675 ;
        RECT 87.555 -146.365 87.885 -146.035 ;
        RECT 87.555 -147.725 87.885 -147.395 ;
        RECT 87.555 -149.085 87.885 -148.755 ;
        RECT 87.555 -150.445 87.885 -150.115 ;
        RECT 87.555 -151.805 87.885 -151.475 ;
        RECT 87.555 -153.165 87.885 -152.835 ;
        RECT 87.555 -154.525 87.885 -154.195 ;
        RECT 87.555 -155.885 87.885 -155.555 ;
        RECT 87.555 -157.245 87.885 -156.915 ;
        RECT 87.555 -158.605 87.885 -158.275 ;
        RECT 87.555 -159.965 87.885 -159.635 ;
        RECT 87.555 -161.325 87.885 -160.995 ;
        RECT 87.555 -162.685 87.885 -162.355 ;
        RECT 87.555 -164.045 87.885 -163.715 ;
        RECT 87.555 -165.405 87.885 -165.075 ;
        RECT 87.555 -166.765 87.885 -166.435 ;
        RECT 87.555 -168.125 87.885 -167.795 ;
        RECT 87.555 -169.485 87.885 -169.155 ;
        RECT 87.555 -170.845 87.885 -170.515 ;
        RECT 87.555 -172.205 87.885 -171.875 ;
        RECT 87.555 -173.565 87.885 -173.235 ;
        RECT 87.555 -174.925 87.885 -174.595 ;
        RECT 87.555 -176.285 87.885 -175.955 ;
        RECT 87.555 -177.645 87.885 -177.315 ;
        RECT 87.555 -179.005 87.885 -178.675 ;
        RECT 87.555 -180.365 87.885 -180.035 ;
        RECT 87.555 -181.725 87.885 -181.395 ;
        RECT 87.555 -183.085 87.885 -182.755 ;
        RECT 87.555 -184.445 87.885 -184.115 ;
        RECT 87.555 -185.805 87.885 -185.475 ;
        RECT 87.555 -187.165 87.885 -186.835 ;
        RECT 87.555 -188.525 87.885 -188.195 ;
        RECT 87.555 -189.885 87.885 -189.555 ;
        RECT 87.555 -191.245 87.885 -190.915 ;
        RECT 87.555 -192.605 87.885 -192.275 ;
        RECT 87.555 -193.965 87.885 -193.635 ;
        RECT 87.555 -195.325 87.885 -194.995 ;
        RECT 87.555 -196.685 87.885 -196.355 ;
        RECT 87.555 -198.045 87.885 -197.715 ;
        RECT 87.555 -199.405 87.885 -199.075 ;
        RECT 87.555 -200.765 87.885 -200.435 ;
        RECT 87.555 -202.125 87.885 -201.795 ;
        RECT 87.555 -203.485 87.885 -203.155 ;
        RECT 87.555 -204.845 87.885 -204.515 ;
        RECT 87.555 -206.205 87.885 -205.875 ;
        RECT 87.555 -207.565 87.885 -207.235 ;
        RECT 87.555 -208.925 87.885 -208.595 ;
        RECT 87.555 -210.285 87.885 -209.955 ;
        RECT 87.555 -211.645 87.885 -211.315 ;
        RECT 87.555 -213.005 87.885 -212.675 ;
        RECT 87.555 -214.365 87.885 -214.035 ;
        RECT 87.555 -215.725 87.885 -215.395 ;
        RECT 87.555 -217.085 87.885 -216.755 ;
        RECT 87.555 -218.445 87.885 -218.115 ;
        RECT 87.555 -219.805 87.885 -219.475 ;
        RECT 87.555 -221.165 87.885 -220.835 ;
        RECT 87.555 -222.525 87.885 -222.195 ;
        RECT 87.555 -223.885 87.885 -223.555 ;
        RECT 87.555 -225.245 87.885 -224.915 ;
        RECT 87.555 -226.605 87.885 -226.275 ;
        RECT 87.555 -227.965 87.885 -227.635 ;
        RECT 87.555 -229.325 87.885 -228.995 ;
        RECT 87.555 -230.685 87.885 -230.355 ;
        RECT 87.555 -232.045 87.885 -231.715 ;
        RECT 87.555 -233.405 87.885 -233.075 ;
        RECT 87.555 -234.765 87.885 -234.435 ;
        RECT 87.555 -236.125 87.885 -235.795 ;
        RECT 87.555 -237.485 87.885 -237.155 ;
        RECT 87.555 -238.845 87.885 -238.515 ;
        RECT 87.555 -241.09 87.885 -239.96 ;
        RECT 87.56 -241.205 87.88 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 244.04 89.245 245.17 ;
        RECT 88.915 242.595 89.245 242.925 ;
        RECT 88.915 241.235 89.245 241.565 ;
        RECT 88.915 239.875 89.245 240.205 ;
        RECT 88.915 238.515 89.245 238.845 ;
        RECT 88.915 237.155 89.245 237.485 ;
        RECT 88.92 237.155 89.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 -0.845 89.245 -0.515 ;
        RECT 88.915 -2.205 89.245 -1.875 ;
        RECT 88.915 -3.565 89.245 -3.235 ;
        RECT 88.92 -3.565 89.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 -123.245 89.245 -122.915 ;
        RECT 88.915 -124.605 89.245 -124.275 ;
        RECT 88.915 -125.965 89.245 -125.635 ;
        RECT 88.915 -127.325 89.245 -126.995 ;
        RECT 88.915 -128.685 89.245 -128.355 ;
        RECT 88.915 -130.045 89.245 -129.715 ;
        RECT 88.915 -131.405 89.245 -131.075 ;
        RECT 88.915 -132.765 89.245 -132.435 ;
        RECT 88.915 -134.125 89.245 -133.795 ;
        RECT 88.915 -135.485 89.245 -135.155 ;
        RECT 88.915 -136.845 89.245 -136.515 ;
        RECT 88.915 -138.205 89.245 -137.875 ;
        RECT 88.915 -139.565 89.245 -139.235 ;
        RECT 88.915 -140.925 89.245 -140.595 ;
        RECT 88.915 -142.285 89.245 -141.955 ;
        RECT 88.915 -143.645 89.245 -143.315 ;
        RECT 88.915 -145.005 89.245 -144.675 ;
        RECT 88.915 -146.365 89.245 -146.035 ;
        RECT 88.915 -147.725 89.245 -147.395 ;
        RECT 88.915 -149.085 89.245 -148.755 ;
        RECT 88.915 -150.445 89.245 -150.115 ;
        RECT 88.915 -151.805 89.245 -151.475 ;
        RECT 88.915 -153.165 89.245 -152.835 ;
        RECT 88.915 -154.525 89.245 -154.195 ;
        RECT 88.915 -155.885 89.245 -155.555 ;
        RECT 88.915 -157.245 89.245 -156.915 ;
        RECT 88.915 -158.605 89.245 -158.275 ;
        RECT 88.915 -159.965 89.245 -159.635 ;
        RECT 88.915 -161.325 89.245 -160.995 ;
        RECT 88.915 -162.685 89.245 -162.355 ;
        RECT 88.915 -164.045 89.245 -163.715 ;
        RECT 88.915 -165.405 89.245 -165.075 ;
        RECT 88.915 -166.765 89.245 -166.435 ;
        RECT 88.915 -168.125 89.245 -167.795 ;
        RECT 88.915 -169.485 89.245 -169.155 ;
        RECT 88.915 -170.845 89.245 -170.515 ;
        RECT 88.915 -172.205 89.245 -171.875 ;
        RECT 88.915 -173.565 89.245 -173.235 ;
        RECT 88.915 -174.925 89.245 -174.595 ;
        RECT 88.915 -176.285 89.245 -175.955 ;
        RECT 88.915 -177.645 89.245 -177.315 ;
        RECT 88.915 -179.005 89.245 -178.675 ;
        RECT 88.915 -180.365 89.245 -180.035 ;
        RECT 88.915 -181.725 89.245 -181.395 ;
        RECT 88.915 -183.085 89.245 -182.755 ;
        RECT 88.915 -184.445 89.245 -184.115 ;
        RECT 88.915 -185.805 89.245 -185.475 ;
        RECT 88.915 -187.165 89.245 -186.835 ;
        RECT 88.915 -188.525 89.245 -188.195 ;
        RECT 88.915 -189.885 89.245 -189.555 ;
        RECT 88.915 -191.245 89.245 -190.915 ;
        RECT 88.915 -192.605 89.245 -192.275 ;
        RECT 88.915 -193.965 89.245 -193.635 ;
        RECT 88.915 -195.325 89.245 -194.995 ;
        RECT 88.915 -196.685 89.245 -196.355 ;
        RECT 88.915 -198.045 89.245 -197.715 ;
        RECT 88.915 -199.405 89.245 -199.075 ;
        RECT 88.915 -200.765 89.245 -200.435 ;
        RECT 88.915 -202.125 89.245 -201.795 ;
        RECT 88.915 -203.485 89.245 -203.155 ;
        RECT 88.915 -204.845 89.245 -204.515 ;
        RECT 88.915 -206.205 89.245 -205.875 ;
        RECT 88.915 -207.565 89.245 -207.235 ;
        RECT 88.915 -208.925 89.245 -208.595 ;
        RECT 88.915 -210.285 89.245 -209.955 ;
        RECT 88.915 -211.645 89.245 -211.315 ;
        RECT 88.915 -213.005 89.245 -212.675 ;
        RECT 88.915 -214.365 89.245 -214.035 ;
        RECT 88.915 -215.725 89.245 -215.395 ;
        RECT 88.915 -217.085 89.245 -216.755 ;
        RECT 88.915 -218.445 89.245 -218.115 ;
        RECT 88.915 -219.805 89.245 -219.475 ;
        RECT 88.915 -221.165 89.245 -220.835 ;
        RECT 88.915 -222.525 89.245 -222.195 ;
        RECT 88.915 -223.885 89.245 -223.555 ;
        RECT 88.915 -225.245 89.245 -224.915 ;
        RECT 88.915 -226.605 89.245 -226.275 ;
        RECT 88.915 -227.965 89.245 -227.635 ;
        RECT 88.915 -229.325 89.245 -228.995 ;
        RECT 88.915 -230.685 89.245 -230.355 ;
        RECT 88.915 -232.045 89.245 -231.715 ;
        RECT 88.915 -233.405 89.245 -233.075 ;
        RECT 88.915 -234.765 89.245 -234.435 ;
        RECT 88.915 -236.125 89.245 -235.795 ;
        RECT 88.915 -237.485 89.245 -237.155 ;
        RECT 88.915 -238.845 89.245 -238.515 ;
        RECT 88.915 -241.09 89.245 -239.96 ;
        RECT 88.92 -241.205 89.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 244.04 90.605 245.17 ;
        RECT 90.275 242.595 90.605 242.925 ;
        RECT 90.275 241.235 90.605 241.565 ;
        RECT 90.275 239.875 90.605 240.205 ;
        RECT 90.275 238.515 90.605 238.845 ;
        RECT 90.275 237.155 90.605 237.485 ;
        RECT 90.28 237.155 90.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 -127.325 90.605 -126.995 ;
        RECT 90.275 -128.685 90.605 -128.355 ;
        RECT 90.275 -130.045 90.605 -129.715 ;
        RECT 90.275 -131.405 90.605 -131.075 ;
        RECT 90.275 -132.765 90.605 -132.435 ;
        RECT 90.275 -134.125 90.605 -133.795 ;
        RECT 90.275 -135.485 90.605 -135.155 ;
        RECT 90.275 -136.845 90.605 -136.515 ;
        RECT 90.275 -138.205 90.605 -137.875 ;
        RECT 90.275 -139.565 90.605 -139.235 ;
        RECT 90.275 -140.925 90.605 -140.595 ;
        RECT 90.275 -142.285 90.605 -141.955 ;
        RECT 90.275 -143.645 90.605 -143.315 ;
        RECT 90.275 -145.005 90.605 -144.675 ;
        RECT 90.275 -146.365 90.605 -146.035 ;
        RECT 90.275 -147.725 90.605 -147.395 ;
        RECT 90.275 -149.085 90.605 -148.755 ;
        RECT 90.275 -150.445 90.605 -150.115 ;
        RECT 90.275 -151.805 90.605 -151.475 ;
        RECT 90.275 -153.165 90.605 -152.835 ;
        RECT 90.275 -154.525 90.605 -154.195 ;
        RECT 90.275 -155.885 90.605 -155.555 ;
        RECT 90.275 -157.245 90.605 -156.915 ;
        RECT 90.275 -158.605 90.605 -158.275 ;
        RECT 90.275 -159.965 90.605 -159.635 ;
        RECT 90.275 -161.325 90.605 -160.995 ;
        RECT 90.275 -162.685 90.605 -162.355 ;
        RECT 90.275 -164.045 90.605 -163.715 ;
        RECT 90.275 -165.405 90.605 -165.075 ;
        RECT 90.275 -166.765 90.605 -166.435 ;
        RECT 90.275 -168.125 90.605 -167.795 ;
        RECT 90.275 -169.485 90.605 -169.155 ;
        RECT 90.275 -170.845 90.605 -170.515 ;
        RECT 90.275 -172.205 90.605 -171.875 ;
        RECT 90.275 -173.565 90.605 -173.235 ;
        RECT 90.275 -174.925 90.605 -174.595 ;
        RECT 90.275 -176.285 90.605 -175.955 ;
        RECT 90.275 -177.645 90.605 -177.315 ;
        RECT 90.275 -179.005 90.605 -178.675 ;
        RECT 90.275 -180.365 90.605 -180.035 ;
        RECT 90.275 -181.725 90.605 -181.395 ;
        RECT 90.275 -183.085 90.605 -182.755 ;
        RECT 90.275 -184.445 90.605 -184.115 ;
        RECT 90.275 -185.805 90.605 -185.475 ;
        RECT 90.275 -187.165 90.605 -186.835 ;
        RECT 90.275 -188.525 90.605 -188.195 ;
        RECT 90.275 -189.885 90.605 -189.555 ;
        RECT 90.275 -191.245 90.605 -190.915 ;
        RECT 90.275 -192.605 90.605 -192.275 ;
        RECT 90.275 -193.965 90.605 -193.635 ;
        RECT 90.275 -195.325 90.605 -194.995 ;
        RECT 90.275 -196.685 90.605 -196.355 ;
        RECT 90.275 -198.045 90.605 -197.715 ;
        RECT 90.275 -199.405 90.605 -199.075 ;
        RECT 90.275 -200.765 90.605 -200.435 ;
        RECT 90.275 -202.125 90.605 -201.795 ;
        RECT 90.275 -203.485 90.605 -203.155 ;
        RECT 90.275 -204.845 90.605 -204.515 ;
        RECT 90.275 -206.205 90.605 -205.875 ;
        RECT 90.275 -207.565 90.605 -207.235 ;
        RECT 90.275 -208.925 90.605 -208.595 ;
        RECT 90.275 -210.285 90.605 -209.955 ;
        RECT 90.275 -211.645 90.605 -211.315 ;
        RECT 90.275 -213.005 90.605 -212.675 ;
        RECT 90.275 -214.365 90.605 -214.035 ;
        RECT 90.275 -215.725 90.605 -215.395 ;
        RECT 90.275 -217.085 90.605 -216.755 ;
        RECT 90.275 -218.445 90.605 -218.115 ;
        RECT 90.275 -219.805 90.605 -219.475 ;
        RECT 90.275 -221.165 90.605 -220.835 ;
        RECT 90.275 -222.525 90.605 -222.195 ;
        RECT 90.275 -223.885 90.605 -223.555 ;
        RECT 90.275 -225.245 90.605 -224.915 ;
        RECT 90.275 -226.605 90.605 -226.275 ;
        RECT 90.275 -227.965 90.605 -227.635 ;
        RECT 90.275 -229.325 90.605 -228.995 ;
        RECT 90.275 -230.685 90.605 -230.355 ;
        RECT 90.275 -232.045 90.605 -231.715 ;
        RECT 90.275 -233.405 90.605 -233.075 ;
        RECT 90.275 -234.765 90.605 -234.435 ;
        RECT 90.275 -236.125 90.605 -235.795 ;
        RECT 90.275 -237.485 90.605 -237.155 ;
        RECT 90.275 -238.845 90.605 -238.515 ;
        RECT 90.275 -241.09 90.605 -239.96 ;
        RECT 90.28 -241.205 90.6 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.51 -125.535 90.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 244.04 91.965 245.17 ;
        RECT 91.635 242.595 91.965 242.925 ;
        RECT 91.635 241.235 91.965 241.565 ;
        RECT 91.635 239.875 91.965 240.205 ;
        RECT 91.635 238.515 91.965 238.845 ;
        RECT 91.635 237.155 91.965 237.485 ;
        RECT 91.64 237.155 91.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 -0.845 91.965 -0.515 ;
        RECT 91.635 -2.205 91.965 -1.875 ;
        RECT 91.635 -3.565 91.965 -3.235 ;
        RECT 91.64 -3.565 91.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 244.04 93.325 245.17 ;
        RECT 92.995 242.595 93.325 242.925 ;
        RECT 92.995 241.235 93.325 241.565 ;
        RECT 92.995 239.875 93.325 240.205 ;
        RECT 92.995 238.515 93.325 238.845 ;
        RECT 92.995 237.155 93.325 237.485 ;
        RECT 93 237.155 93.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 -0.845 93.325 -0.515 ;
        RECT 92.995 -2.205 93.325 -1.875 ;
        RECT 92.995 -3.565 93.325 -3.235 ;
        RECT 93 -3.565 93.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 244.04 94.685 245.17 ;
        RECT 94.355 242.595 94.685 242.925 ;
        RECT 94.355 241.235 94.685 241.565 ;
        RECT 94.355 239.875 94.685 240.205 ;
        RECT 94.355 238.515 94.685 238.845 ;
        RECT 94.355 237.155 94.685 237.485 ;
        RECT 94.36 237.155 94.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 -0.845 94.685 -0.515 ;
        RECT 94.355 -2.205 94.685 -1.875 ;
        RECT 94.355 -3.565 94.685 -3.235 ;
        RECT 94.36 -3.565 94.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 -207.565 94.685 -207.235 ;
        RECT 94.355 -208.925 94.685 -208.595 ;
        RECT 94.355 -210.285 94.685 -209.955 ;
        RECT 94.355 -211.645 94.685 -211.315 ;
        RECT 94.355 -213.005 94.685 -212.675 ;
        RECT 94.355 -214.365 94.685 -214.035 ;
        RECT 94.355 -215.725 94.685 -215.395 ;
        RECT 94.355 -217.085 94.685 -216.755 ;
        RECT 94.355 -218.445 94.685 -218.115 ;
        RECT 94.355 -219.805 94.685 -219.475 ;
        RECT 94.355 -221.165 94.685 -220.835 ;
        RECT 94.355 -222.525 94.685 -222.195 ;
        RECT 94.355 -223.885 94.685 -223.555 ;
        RECT 94.355 -225.245 94.685 -224.915 ;
        RECT 94.355 -226.605 94.685 -226.275 ;
        RECT 94.355 -227.965 94.685 -227.635 ;
        RECT 94.355 -229.325 94.685 -228.995 ;
        RECT 94.355 -230.685 94.685 -230.355 ;
        RECT 94.355 -232.045 94.685 -231.715 ;
        RECT 94.355 -233.405 94.685 -233.075 ;
        RECT 94.355 -234.765 94.685 -234.435 ;
        RECT 94.355 -236.125 94.685 -235.795 ;
        RECT 94.355 -237.485 94.685 -237.155 ;
        RECT 94.355 -238.845 94.685 -238.515 ;
        RECT 94.355 -241.09 94.685 -239.96 ;
        RECT 94.36 -241.205 94.68 -122.24 ;
        RECT 94.355 -123.245 94.685 -122.915 ;
        RECT 94.355 -124.605 94.685 -124.275 ;
        RECT 94.355 -125.965 94.685 -125.635 ;
        RECT 94.355 -127.325 94.685 -126.995 ;
        RECT 94.355 -128.685 94.685 -128.355 ;
        RECT 94.355 -130.045 94.685 -129.715 ;
        RECT 94.355 -131.405 94.685 -131.075 ;
        RECT 94.355 -132.765 94.685 -132.435 ;
        RECT 94.355 -134.125 94.685 -133.795 ;
        RECT 94.355 -135.485 94.685 -135.155 ;
        RECT 94.355 -136.845 94.685 -136.515 ;
        RECT 94.355 -138.205 94.685 -137.875 ;
        RECT 94.355 -139.565 94.685 -139.235 ;
        RECT 94.355 -140.925 94.685 -140.595 ;
        RECT 94.355 -142.285 94.685 -141.955 ;
        RECT 94.355 -143.645 94.685 -143.315 ;
        RECT 94.355 -145.005 94.685 -144.675 ;
        RECT 94.355 -146.365 94.685 -146.035 ;
        RECT 94.355 -147.725 94.685 -147.395 ;
        RECT 94.355 -149.085 94.685 -148.755 ;
        RECT 94.355 -150.445 94.685 -150.115 ;
        RECT 94.355 -151.805 94.685 -151.475 ;
        RECT 94.355 -153.165 94.685 -152.835 ;
        RECT 94.355 -154.525 94.685 -154.195 ;
        RECT 94.355 -155.885 94.685 -155.555 ;
        RECT 94.355 -157.245 94.685 -156.915 ;
        RECT 94.355 -158.605 94.685 -158.275 ;
        RECT 94.355 -159.965 94.685 -159.635 ;
        RECT 94.355 -161.325 94.685 -160.995 ;
        RECT 94.355 -162.685 94.685 -162.355 ;
        RECT 94.355 -164.045 94.685 -163.715 ;
        RECT 94.355 -165.405 94.685 -165.075 ;
        RECT 94.355 -166.765 94.685 -166.435 ;
        RECT 94.355 -168.125 94.685 -167.795 ;
        RECT 94.355 -169.485 94.685 -169.155 ;
        RECT 94.355 -170.845 94.685 -170.515 ;
        RECT 94.355 -172.205 94.685 -171.875 ;
        RECT 94.355 -173.565 94.685 -173.235 ;
        RECT 94.355 -174.925 94.685 -174.595 ;
        RECT 94.355 -176.285 94.685 -175.955 ;
        RECT 94.355 -177.645 94.685 -177.315 ;
        RECT 94.355 -179.005 94.685 -178.675 ;
        RECT 94.355 -180.365 94.685 -180.035 ;
        RECT 94.355 -181.725 94.685 -181.395 ;
        RECT 94.355 -183.085 94.685 -182.755 ;
        RECT 94.355 -184.445 94.685 -184.115 ;
        RECT 94.355 -185.805 94.685 -185.475 ;
        RECT 94.355 -187.165 94.685 -186.835 ;
        RECT 94.355 -188.525 94.685 -188.195 ;
        RECT 94.355 -189.885 94.685 -189.555 ;
        RECT 94.355 -191.245 94.685 -190.915 ;
        RECT 94.355 -192.605 94.685 -192.275 ;
        RECT 94.355 -193.965 94.685 -193.635 ;
        RECT 94.355 -195.325 94.685 -194.995 ;
        RECT 94.355 -196.685 94.685 -196.355 ;
        RECT 94.355 -198.045 94.685 -197.715 ;
        RECT 94.355 -199.405 94.685 -199.075 ;
        RECT 94.355 -200.765 94.685 -200.435 ;
        RECT 94.355 -202.125 94.685 -201.795 ;
        RECT 94.355 -203.485 94.685 -203.155 ;
        RECT 94.355 -204.845 94.685 -204.515 ;
        RECT 94.355 -206.205 94.685 -205.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 244.04 57.965 245.17 ;
        RECT 57.635 242.595 57.965 242.925 ;
        RECT 57.635 241.235 57.965 241.565 ;
        RECT 57.635 239.875 57.965 240.205 ;
        RECT 57.635 238.515 57.965 238.845 ;
        RECT 57.635 237.155 57.965 237.485 ;
        RECT 57.64 237.155 57.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 -127.325 57.965 -126.995 ;
        RECT 57.635 -128.685 57.965 -128.355 ;
        RECT 57.635 -130.045 57.965 -129.715 ;
        RECT 57.635 -131.405 57.965 -131.075 ;
        RECT 57.635 -132.765 57.965 -132.435 ;
        RECT 57.635 -134.125 57.965 -133.795 ;
        RECT 57.635 -135.485 57.965 -135.155 ;
        RECT 57.635 -136.845 57.965 -136.515 ;
        RECT 57.635 -138.205 57.965 -137.875 ;
        RECT 57.635 -139.565 57.965 -139.235 ;
        RECT 57.635 -140.925 57.965 -140.595 ;
        RECT 57.635 -142.285 57.965 -141.955 ;
        RECT 57.635 -143.645 57.965 -143.315 ;
        RECT 57.635 -145.005 57.965 -144.675 ;
        RECT 57.635 -146.365 57.965 -146.035 ;
        RECT 57.635 -147.725 57.965 -147.395 ;
        RECT 57.635 -149.085 57.965 -148.755 ;
        RECT 57.635 -150.445 57.965 -150.115 ;
        RECT 57.635 -151.805 57.965 -151.475 ;
        RECT 57.635 -153.165 57.965 -152.835 ;
        RECT 57.635 -154.525 57.965 -154.195 ;
        RECT 57.635 -155.885 57.965 -155.555 ;
        RECT 57.635 -157.245 57.965 -156.915 ;
        RECT 57.635 -158.605 57.965 -158.275 ;
        RECT 57.635 -159.965 57.965 -159.635 ;
        RECT 57.635 -161.325 57.965 -160.995 ;
        RECT 57.635 -162.685 57.965 -162.355 ;
        RECT 57.635 -164.045 57.965 -163.715 ;
        RECT 57.635 -165.405 57.965 -165.075 ;
        RECT 57.635 -166.765 57.965 -166.435 ;
        RECT 57.635 -168.125 57.965 -167.795 ;
        RECT 57.635 -169.485 57.965 -169.155 ;
        RECT 57.635 -170.845 57.965 -170.515 ;
        RECT 57.635 -172.205 57.965 -171.875 ;
        RECT 57.635 -173.565 57.965 -173.235 ;
        RECT 57.635 -174.925 57.965 -174.595 ;
        RECT 57.635 -176.285 57.965 -175.955 ;
        RECT 57.635 -177.645 57.965 -177.315 ;
        RECT 57.635 -179.005 57.965 -178.675 ;
        RECT 57.635 -180.365 57.965 -180.035 ;
        RECT 57.635 -181.725 57.965 -181.395 ;
        RECT 57.635 -183.085 57.965 -182.755 ;
        RECT 57.635 -184.445 57.965 -184.115 ;
        RECT 57.635 -185.805 57.965 -185.475 ;
        RECT 57.635 -187.165 57.965 -186.835 ;
        RECT 57.635 -188.525 57.965 -188.195 ;
        RECT 57.635 -189.885 57.965 -189.555 ;
        RECT 57.635 -191.245 57.965 -190.915 ;
        RECT 57.635 -192.605 57.965 -192.275 ;
        RECT 57.635 -193.965 57.965 -193.635 ;
        RECT 57.635 -195.325 57.965 -194.995 ;
        RECT 57.635 -196.685 57.965 -196.355 ;
        RECT 57.635 -198.045 57.965 -197.715 ;
        RECT 57.635 -199.405 57.965 -199.075 ;
        RECT 57.635 -200.765 57.965 -200.435 ;
        RECT 57.635 -202.125 57.965 -201.795 ;
        RECT 57.635 -203.485 57.965 -203.155 ;
        RECT 57.635 -204.845 57.965 -204.515 ;
        RECT 57.635 -206.205 57.965 -205.875 ;
        RECT 57.635 -207.565 57.965 -207.235 ;
        RECT 57.635 -208.925 57.965 -208.595 ;
        RECT 57.635 -210.285 57.965 -209.955 ;
        RECT 57.635 -211.645 57.965 -211.315 ;
        RECT 57.635 -213.005 57.965 -212.675 ;
        RECT 57.635 -214.365 57.965 -214.035 ;
        RECT 57.635 -215.725 57.965 -215.395 ;
        RECT 57.635 -217.085 57.965 -216.755 ;
        RECT 57.635 -218.445 57.965 -218.115 ;
        RECT 57.635 -219.805 57.965 -219.475 ;
        RECT 57.635 -221.165 57.965 -220.835 ;
        RECT 57.635 -222.525 57.965 -222.195 ;
        RECT 57.635 -223.885 57.965 -223.555 ;
        RECT 57.635 -225.245 57.965 -224.915 ;
        RECT 57.635 -226.605 57.965 -226.275 ;
        RECT 57.635 -227.965 57.965 -227.635 ;
        RECT 57.635 -229.325 57.965 -228.995 ;
        RECT 57.635 -230.685 57.965 -230.355 ;
        RECT 57.635 -232.045 57.965 -231.715 ;
        RECT 57.635 -233.405 57.965 -233.075 ;
        RECT 57.635 -234.765 57.965 -234.435 ;
        RECT 57.635 -236.125 57.965 -235.795 ;
        RECT 57.635 -237.485 57.965 -237.155 ;
        RECT 57.635 -238.845 57.965 -238.515 ;
        RECT 57.635 -241.09 57.965 -239.96 ;
        RECT 57.64 -241.205 57.96 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.81 -125.535 58.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 244.04 59.325 245.17 ;
        RECT 58.995 242.595 59.325 242.925 ;
        RECT 58.995 241.235 59.325 241.565 ;
        RECT 58.995 239.875 59.325 240.205 ;
        RECT 58.995 238.515 59.325 238.845 ;
        RECT 58.995 237.155 59.325 237.485 ;
        RECT 59 237.155 59.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 -0.845 59.325 -0.515 ;
        RECT 58.995 -2.205 59.325 -1.875 ;
        RECT 58.995 -3.565 59.325 -3.235 ;
        RECT 59 -3.565 59.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 244.04 60.685 245.17 ;
        RECT 60.355 242.595 60.685 242.925 ;
        RECT 60.355 241.235 60.685 241.565 ;
        RECT 60.355 239.875 60.685 240.205 ;
        RECT 60.355 238.515 60.685 238.845 ;
        RECT 60.355 237.155 60.685 237.485 ;
        RECT 60.36 237.155 60.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 -0.845 60.685 -0.515 ;
        RECT 60.355 -2.205 60.685 -1.875 ;
        RECT 60.355 -3.565 60.685 -3.235 ;
        RECT 60.36 -3.565 60.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 244.04 62.045 245.17 ;
        RECT 61.715 242.595 62.045 242.925 ;
        RECT 61.715 241.235 62.045 241.565 ;
        RECT 61.715 239.875 62.045 240.205 ;
        RECT 61.715 238.515 62.045 238.845 ;
        RECT 61.715 237.155 62.045 237.485 ;
        RECT 61.72 237.155 62.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -0.845 62.045 -0.515 ;
        RECT 61.715 -2.205 62.045 -1.875 ;
        RECT 61.715 -3.565 62.045 -3.235 ;
        RECT 61.72 -3.565 62.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -123.245 62.045 -122.915 ;
        RECT 61.715 -124.605 62.045 -124.275 ;
        RECT 61.715 -125.965 62.045 -125.635 ;
        RECT 61.715 -127.325 62.045 -126.995 ;
        RECT 61.715 -128.685 62.045 -128.355 ;
        RECT 61.715 -130.045 62.045 -129.715 ;
        RECT 61.715 -131.405 62.045 -131.075 ;
        RECT 61.715 -132.765 62.045 -132.435 ;
        RECT 61.715 -134.125 62.045 -133.795 ;
        RECT 61.715 -135.485 62.045 -135.155 ;
        RECT 61.715 -136.845 62.045 -136.515 ;
        RECT 61.715 -138.205 62.045 -137.875 ;
        RECT 61.715 -139.565 62.045 -139.235 ;
        RECT 61.715 -140.925 62.045 -140.595 ;
        RECT 61.715 -142.285 62.045 -141.955 ;
        RECT 61.715 -143.645 62.045 -143.315 ;
        RECT 61.715 -145.005 62.045 -144.675 ;
        RECT 61.715 -146.365 62.045 -146.035 ;
        RECT 61.715 -147.725 62.045 -147.395 ;
        RECT 61.715 -149.085 62.045 -148.755 ;
        RECT 61.715 -150.445 62.045 -150.115 ;
        RECT 61.715 -151.805 62.045 -151.475 ;
        RECT 61.715 -153.165 62.045 -152.835 ;
        RECT 61.715 -154.525 62.045 -154.195 ;
        RECT 61.715 -155.885 62.045 -155.555 ;
        RECT 61.715 -157.245 62.045 -156.915 ;
        RECT 61.715 -158.605 62.045 -158.275 ;
        RECT 61.715 -159.965 62.045 -159.635 ;
        RECT 61.715 -161.325 62.045 -160.995 ;
        RECT 61.715 -162.685 62.045 -162.355 ;
        RECT 61.715 -164.045 62.045 -163.715 ;
        RECT 61.715 -165.405 62.045 -165.075 ;
        RECT 61.715 -166.765 62.045 -166.435 ;
        RECT 61.715 -168.125 62.045 -167.795 ;
        RECT 61.715 -169.485 62.045 -169.155 ;
        RECT 61.715 -170.845 62.045 -170.515 ;
        RECT 61.715 -172.205 62.045 -171.875 ;
        RECT 61.715 -173.565 62.045 -173.235 ;
        RECT 61.715 -174.925 62.045 -174.595 ;
        RECT 61.715 -176.285 62.045 -175.955 ;
        RECT 61.715 -177.645 62.045 -177.315 ;
        RECT 61.715 -179.005 62.045 -178.675 ;
        RECT 61.715 -180.365 62.045 -180.035 ;
        RECT 61.715 -181.725 62.045 -181.395 ;
        RECT 61.715 -183.085 62.045 -182.755 ;
        RECT 61.715 -184.445 62.045 -184.115 ;
        RECT 61.715 -185.805 62.045 -185.475 ;
        RECT 61.715 -187.165 62.045 -186.835 ;
        RECT 61.715 -188.525 62.045 -188.195 ;
        RECT 61.715 -189.885 62.045 -189.555 ;
        RECT 61.715 -191.245 62.045 -190.915 ;
        RECT 61.715 -192.605 62.045 -192.275 ;
        RECT 61.715 -193.965 62.045 -193.635 ;
        RECT 61.715 -195.325 62.045 -194.995 ;
        RECT 61.715 -196.685 62.045 -196.355 ;
        RECT 61.715 -198.045 62.045 -197.715 ;
        RECT 61.715 -199.405 62.045 -199.075 ;
        RECT 61.715 -200.765 62.045 -200.435 ;
        RECT 61.715 -202.125 62.045 -201.795 ;
        RECT 61.715 -203.485 62.045 -203.155 ;
        RECT 61.715 -204.845 62.045 -204.515 ;
        RECT 61.715 -206.205 62.045 -205.875 ;
        RECT 61.715 -207.565 62.045 -207.235 ;
        RECT 61.715 -208.925 62.045 -208.595 ;
        RECT 61.715 -210.285 62.045 -209.955 ;
        RECT 61.715 -211.645 62.045 -211.315 ;
        RECT 61.715 -213.005 62.045 -212.675 ;
        RECT 61.715 -214.365 62.045 -214.035 ;
        RECT 61.715 -215.725 62.045 -215.395 ;
        RECT 61.715 -217.085 62.045 -216.755 ;
        RECT 61.715 -218.445 62.045 -218.115 ;
        RECT 61.715 -219.805 62.045 -219.475 ;
        RECT 61.715 -221.165 62.045 -220.835 ;
        RECT 61.715 -222.525 62.045 -222.195 ;
        RECT 61.715 -223.885 62.045 -223.555 ;
        RECT 61.715 -225.245 62.045 -224.915 ;
        RECT 61.715 -226.605 62.045 -226.275 ;
        RECT 61.715 -227.965 62.045 -227.635 ;
        RECT 61.715 -229.325 62.045 -228.995 ;
        RECT 61.715 -230.685 62.045 -230.355 ;
        RECT 61.715 -232.045 62.045 -231.715 ;
        RECT 61.715 -233.405 62.045 -233.075 ;
        RECT 61.715 -234.765 62.045 -234.435 ;
        RECT 61.715 -236.125 62.045 -235.795 ;
        RECT 61.715 -237.485 62.045 -237.155 ;
        RECT 61.715 -238.845 62.045 -238.515 ;
        RECT 61.715 -241.09 62.045 -239.96 ;
        RECT 61.72 -241.205 62.04 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 244.04 63.405 245.17 ;
        RECT 63.075 242.595 63.405 242.925 ;
        RECT 63.075 241.235 63.405 241.565 ;
        RECT 63.075 239.875 63.405 240.205 ;
        RECT 63.075 238.515 63.405 238.845 ;
        RECT 63.075 237.155 63.405 237.485 ;
        RECT 63.08 237.155 63.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 -0.845 63.405 -0.515 ;
        RECT 63.075 -2.205 63.405 -1.875 ;
        RECT 63.075 -3.565 63.405 -3.235 ;
        RECT 63.08 -3.565 63.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 -123.245 63.405 -122.915 ;
        RECT 63.075 -124.605 63.405 -124.275 ;
        RECT 63.075 -125.965 63.405 -125.635 ;
        RECT 63.075 -127.325 63.405 -126.995 ;
        RECT 63.075 -128.685 63.405 -128.355 ;
        RECT 63.075 -130.045 63.405 -129.715 ;
        RECT 63.075 -131.405 63.405 -131.075 ;
        RECT 63.075 -132.765 63.405 -132.435 ;
        RECT 63.075 -134.125 63.405 -133.795 ;
        RECT 63.075 -135.485 63.405 -135.155 ;
        RECT 63.075 -136.845 63.405 -136.515 ;
        RECT 63.075 -138.205 63.405 -137.875 ;
        RECT 63.075 -139.565 63.405 -139.235 ;
        RECT 63.075 -140.925 63.405 -140.595 ;
        RECT 63.075 -142.285 63.405 -141.955 ;
        RECT 63.075 -143.645 63.405 -143.315 ;
        RECT 63.075 -145.005 63.405 -144.675 ;
        RECT 63.075 -146.365 63.405 -146.035 ;
        RECT 63.075 -147.725 63.405 -147.395 ;
        RECT 63.075 -149.085 63.405 -148.755 ;
        RECT 63.075 -150.445 63.405 -150.115 ;
        RECT 63.075 -151.805 63.405 -151.475 ;
        RECT 63.075 -153.165 63.405 -152.835 ;
        RECT 63.075 -154.525 63.405 -154.195 ;
        RECT 63.075 -155.885 63.405 -155.555 ;
        RECT 63.075 -157.245 63.405 -156.915 ;
        RECT 63.075 -158.605 63.405 -158.275 ;
        RECT 63.075 -159.965 63.405 -159.635 ;
        RECT 63.075 -161.325 63.405 -160.995 ;
        RECT 63.075 -162.685 63.405 -162.355 ;
        RECT 63.075 -164.045 63.405 -163.715 ;
        RECT 63.075 -165.405 63.405 -165.075 ;
        RECT 63.075 -166.765 63.405 -166.435 ;
        RECT 63.075 -168.125 63.405 -167.795 ;
        RECT 63.075 -169.485 63.405 -169.155 ;
        RECT 63.075 -170.845 63.405 -170.515 ;
        RECT 63.075 -172.205 63.405 -171.875 ;
        RECT 63.075 -173.565 63.405 -173.235 ;
        RECT 63.075 -174.925 63.405 -174.595 ;
        RECT 63.075 -176.285 63.405 -175.955 ;
        RECT 63.075 -177.645 63.405 -177.315 ;
        RECT 63.075 -179.005 63.405 -178.675 ;
        RECT 63.075 -180.365 63.405 -180.035 ;
        RECT 63.075 -181.725 63.405 -181.395 ;
        RECT 63.075 -183.085 63.405 -182.755 ;
        RECT 63.075 -184.445 63.405 -184.115 ;
        RECT 63.075 -185.805 63.405 -185.475 ;
        RECT 63.075 -187.165 63.405 -186.835 ;
        RECT 63.075 -188.525 63.405 -188.195 ;
        RECT 63.075 -189.885 63.405 -189.555 ;
        RECT 63.075 -191.245 63.405 -190.915 ;
        RECT 63.075 -192.605 63.405 -192.275 ;
        RECT 63.075 -193.965 63.405 -193.635 ;
        RECT 63.075 -195.325 63.405 -194.995 ;
        RECT 63.075 -196.685 63.405 -196.355 ;
        RECT 63.075 -198.045 63.405 -197.715 ;
        RECT 63.075 -199.405 63.405 -199.075 ;
        RECT 63.075 -200.765 63.405 -200.435 ;
        RECT 63.075 -202.125 63.405 -201.795 ;
        RECT 63.075 -203.485 63.405 -203.155 ;
        RECT 63.075 -204.845 63.405 -204.515 ;
        RECT 63.075 -206.205 63.405 -205.875 ;
        RECT 63.075 -207.565 63.405 -207.235 ;
        RECT 63.075 -208.925 63.405 -208.595 ;
        RECT 63.075 -210.285 63.405 -209.955 ;
        RECT 63.075 -211.645 63.405 -211.315 ;
        RECT 63.075 -213.005 63.405 -212.675 ;
        RECT 63.075 -214.365 63.405 -214.035 ;
        RECT 63.075 -215.725 63.405 -215.395 ;
        RECT 63.075 -217.085 63.405 -216.755 ;
        RECT 63.075 -218.445 63.405 -218.115 ;
        RECT 63.075 -219.805 63.405 -219.475 ;
        RECT 63.075 -221.165 63.405 -220.835 ;
        RECT 63.075 -222.525 63.405 -222.195 ;
        RECT 63.075 -223.885 63.405 -223.555 ;
        RECT 63.075 -225.245 63.405 -224.915 ;
        RECT 63.075 -226.605 63.405 -226.275 ;
        RECT 63.075 -227.965 63.405 -227.635 ;
        RECT 63.075 -229.325 63.405 -228.995 ;
        RECT 63.075 -230.685 63.405 -230.355 ;
        RECT 63.075 -232.045 63.405 -231.715 ;
        RECT 63.075 -233.405 63.405 -233.075 ;
        RECT 63.075 -234.765 63.405 -234.435 ;
        RECT 63.075 -236.125 63.405 -235.795 ;
        RECT 63.075 -237.485 63.405 -237.155 ;
        RECT 63.075 -238.845 63.405 -238.515 ;
        RECT 63.075 -241.09 63.405 -239.96 ;
        RECT 63.08 -241.205 63.4 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 244.04 64.765 245.17 ;
        RECT 64.435 242.595 64.765 242.925 ;
        RECT 64.435 241.235 64.765 241.565 ;
        RECT 64.435 239.875 64.765 240.205 ;
        RECT 64.435 238.515 64.765 238.845 ;
        RECT 64.435 237.155 64.765 237.485 ;
        RECT 64.44 237.155 64.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 -0.845 64.765 -0.515 ;
        RECT 64.435 -2.205 64.765 -1.875 ;
        RECT 64.435 -3.565 64.765 -3.235 ;
        RECT 64.44 -3.565 64.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 -123.245 64.765 -122.915 ;
        RECT 64.435 -124.605 64.765 -124.275 ;
        RECT 64.435 -125.965 64.765 -125.635 ;
        RECT 64.435 -127.325 64.765 -126.995 ;
        RECT 64.435 -128.685 64.765 -128.355 ;
        RECT 64.435 -130.045 64.765 -129.715 ;
        RECT 64.435 -131.405 64.765 -131.075 ;
        RECT 64.435 -132.765 64.765 -132.435 ;
        RECT 64.435 -134.125 64.765 -133.795 ;
        RECT 64.435 -135.485 64.765 -135.155 ;
        RECT 64.435 -136.845 64.765 -136.515 ;
        RECT 64.435 -138.205 64.765 -137.875 ;
        RECT 64.435 -139.565 64.765 -139.235 ;
        RECT 64.435 -140.925 64.765 -140.595 ;
        RECT 64.435 -142.285 64.765 -141.955 ;
        RECT 64.435 -143.645 64.765 -143.315 ;
        RECT 64.435 -145.005 64.765 -144.675 ;
        RECT 64.435 -146.365 64.765 -146.035 ;
        RECT 64.435 -147.725 64.765 -147.395 ;
        RECT 64.435 -149.085 64.765 -148.755 ;
        RECT 64.435 -150.445 64.765 -150.115 ;
        RECT 64.435 -151.805 64.765 -151.475 ;
        RECT 64.435 -153.165 64.765 -152.835 ;
        RECT 64.435 -154.525 64.765 -154.195 ;
        RECT 64.435 -155.885 64.765 -155.555 ;
        RECT 64.435 -157.245 64.765 -156.915 ;
        RECT 64.435 -158.605 64.765 -158.275 ;
        RECT 64.435 -159.965 64.765 -159.635 ;
        RECT 64.435 -161.325 64.765 -160.995 ;
        RECT 64.435 -162.685 64.765 -162.355 ;
        RECT 64.435 -164.045 64.765 -163.715 ;
        RECT 64.435 -165.405 64.765 -165.075 ;
        RECT 64.435 -166.765 64.765 -166.435 ;
        RECT 64.435 -168.125 64.765 -167.795 ;
        RECT 64.435 -169.485 64.765 -169.155 ;
        RECT 64.435 -170.845 64.765 -170.515 ;
        RECT 64.435 -172.205 64.765 -171.875 ;
        RECT 64.435 -173.565 64.765 -173.235 ;
        RECT 64.435 -174.925 64.765 -174.595 ;
        RECT 64.435 -176.285 64.765 -175.955 ;
        RECT 64.435 -177.645 64.765 -177.315 ;
        RECT 64.435 -179.005 64.765 -178.675 ;
        RECT 64.435 -180.365 64.765 -180.035 ;
        RECT 64.435 -181.725 64.765 -181.395 ;
        RECT 64.435 -183.085 64.765 -182.755 ;
        RECT 64.435 -184.445 64.765 -184.115 ;
        RECT 64.435 -185.805 64.765 -185.475 ;
        RECT 64.435 -187.165 64.765 -186.835 ;
        RECT 64.435 -188.525 64.765 -188.195 ;
        RECT 64.435 -189.885 64.765 -189.555 ;
        RECT 64.435 -191.245 64.765 -190.915 ;
        RECT 64.435 -192.605 64.765 -192.275 ;
        RECT 64.435 -193.965 64.765 -193.635 ;
        RECT 64.435 -195.325 64.765 -194.995 ;
        RECT 64.435 -196.685 64.765 -196.355 ;
        RECT 64.435 -198.045 64.765 -197.715 ;
        RECT 64.435 -199.405 64.765 -199.075 ;
        RECT 64.435 -200.765 64.765 -200.435 ;
        RECT 64.435 -202.125 64.765 -201.795 ;
        RECT 64.435 -203.485 64.765 -203.155 ;
        RECT 64.435 -204.845 64.765 -204.515 ;
        RECT 64.435 -206.205 64.765 -205.875 ;
        RECT 64.435 -207.565 64.765 -207.235 ;
        RECT 64.435 -208.925 64.765 -208.595 ;
        RECT 64.435 -210.285 64.765 -209.955 ;
        RECT 64.435 -211.645 64.765 -211.315 ;
        RECT 64.435 -213.005 64.765 -212.675 ;
        RECT 64.435 -214.365 64.765 -214.035 ;
        RECT 64.435 -215.725 64.765 -215.395 ;
        RECT 64.435 -217.085 64.765 -216.755 ;
        RECT 64.435 -218.445 64.765 -218.115 ;
        RECT 64.435 -219.805 64.765 -219.475 ;
        RECT 64.435 -221.165 64.765 -220.835 ;
        RECT 64.435 -222.525 64.765 -222.195 ;
        RECT 64.435 -223.885 64.765 -223.555 ;
        RECT 64.435 -225.245 64.765 -224.915 ;
        RECT 64.435 -226.605 64.765 -226.275 ;
        RECT 64.435 -227.965 64.765 -227.635 ;
        RECT 64.435 -229.325 64.765 -228.995 ;
        RECT 64.435 -230.685 64.765 -230.355 ;
        RECT 64.435 -232.045 64.765 -231.715 ;
        RECT 64.435 -233.405 64.765 -233.075 ;
        RECT 64.435 -234.765 64.765 -234.435 ;
        RECT 64.435 -236.125 64.765 -235.795 ;
        RECT 64.435 -237.485 64.765 -237.155 ;
        RECT 64.435 -238.845 64.765 -238.515 ;
        RECT 64.435 -241.09 64.765 -239.96 ;
        RECT 64.44 -241.205 64.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 244.04 66.125 245.17 ;
        RECT 65.795 242.595 66.125 242.925 ;
        RECT 65.795 241.235 66.125 241.565 ;
        RECT 65.795 239.875 66.125 240.205 ;
        RECT 65.795 238.515 66.125 238.845 ;
        RECT 65.795 237.155 66.125 237.485 ;
        RECT 65.8 237.155 66.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -0.845 66.125 -0.515 ;
        RECT 65.795 -2.205 66.125 -1.875 ;
        RECT 65.795 -3.565 66.125 -3.235 ;
        RECT 65.8 -3.565 66.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -123.245 66.125 -122.915 ;
        RECT 65.795 -124.605 66.125 -124.275 ;
        RECT 65.795 -125.965 66.125 -125.635 ;
        RECT 65.795 -127.325 66.125 -126.995 ;
        RECT 65.795 -128.685 66.125 -128.355 ;
        RECT 65.795 -130.045 66.125 -129.715 ;
        RECT 65.795 -131.405 66.125 -131.075 ;
        RECT 65.795 -132.765 66.125 -132.435 ;
        RECT 65.795 -134.125 66.125 -133.795 ;
        RECT 65.795 -135.485 66.125 -135.155 ;
        RECT 65.795 -136.845 66.125 -136.515 ;
        RECT 65.795 -138.205 66.125 -137.875 ;
        RECT 65.795 -139.565 66.125 -139.235 ;
        RECT 65.795 -140.925 66.125 -140.595 ;
        RECT 65.795 -142.285 66.125 -141.955 ;
        RECT 65.795 -143.645 66.125 -143.315 ;
        RECT 65.795 -145.005 66.125 -144.675 ;
        RECT 65.795 -146.365 66.125 -146.035 ;
        RECT 65.795 -147.725 66.125 -147.395 ;
        RECT 65.795 -149.085 66.125 -148.755 ;
        RECT 65.795 -150.445 66.125 -150.115 ;
        RECT 65.795 -151.805 66.125 -151.475 ;
        RECT 65.795 -153.165 66.125 -152.835 ;
        RECT 65.795 -154.525 66.125 -154.195 ;
        RECT 65.795 -155.885 66.125 -155.555 ;
        RECT 65.795 -157.245 66.125 -156.915 ;
        RECT 65.795 -158.605 66.125 -158.275 ;
        RECT 65.795 -159.965 66.125 -159.635 ;
        RECT 65.795 -161.325 66.125 -160.995 ;
        RECT 65.795 -162.685 66.125 -162.355 ;
        RECT 65.795 -164.045 66.125 -163.715 ;
        RECT 65.795 -165.405 66.125 -165.075 ;
        RECT 65.795 -166.765 66.125 -166.435 ;
        RECT 65.795 -168.125 66.125 -167.795 ;
        RECT 65.795 -169.485 66.125 -169.155 ;
        RECT 65.795 -170.845 66.125 -170.515 ;
        RECT 65.795 -172.205 66.125 -171.875 ;
        RECT 65.795 -173.565 66.125 -173.235 ;
        RECT 65.795 -174.925 66.125 -174.595 ;
        RECT 65.795 -176.285 66.125 -175.955 ;
        RECT 65.795 -177.645 66.125 -177.315 ;
        RECT 65.795 -179.005 66.125 -178.675 ;
        RECT 65.795 -180.365 66.125 -180.035 ;
        RECT 65.795 -181.725 66.125 -181.395 ;
        RECT 65.795 -183.085 66.125 -182.755 ;
        RECT 65.795 -184.445 66.125 -184.115 ;
        RECT 65.795 -185.805 66.125 -185.475 ;
        RECT 65.795 -187.165 66.125 -186.835 ;
        RECT 65.795 -188.525 66.125 -188.195 ;
        RECT 65.795 -189.885 66.125 -189.555 ;
        RECT 65.795 -191.245 66.125 -190.915 ;
        RECT 65.795 -192.605 66.125 -192.275 ;
        RECT 65.795 -193.965 66.125 -193.635 ;
        RECT 65.795 -195.325 66.125 -194.995 ;
        RECT 65.795 -196.685 66.125 -196.355 ;
        RECT 65.795 -198.045 66.125 -197.715 ;
        RECT 65.795 -199.405 66.125 -199.075 ;
        RECT 65.795 -200.765 66.125 -200.435 ;
        RECT 65.795 -202.125 66.125 -201.795 ;
        RECT 65.795 -203.485 66.125 -203.155 ;
        RECT 65.795 -204.845 66.125 -204.515 ;
        RECT 65.795 -206.205 66.125 -205.875 ;
        RECT 65.795 -207.565 66.125 -207.235 ;
        RECT 65.795 -208.925 66.125 -208.595 ;
        RECT 65.795 -210.285 66.125 -209.955 ;
        RECT 65.795 -211.645 66.125 -211.315 ;
        RECT 65.795 -213.005 66.125 -212.675 ;
        RECT 65.795 -214.365 66.125 -214.035 ;
        RECT 65.795 -215.725 66.125 -215.395 ;
        RECT 65.795 -217.085 66.125 -216.755 ;
        RECT 65.795 -218.445 66.125 -218.115 ;
        RECT 65.795 -219.805 66.125 -219.475 ;
        RECT 65.795 -221.165 66.125 -220.835 ;
        RECT 65.795 -222.525 66.125 -222.195 ;
        RECT 65.795 -223.885 66.125 -223.555 ;
        RECT 65.795 -225.245 66.125 -224.915 ;
        RECT 65.795 -226.605 66.125 -226.275 ;
        RECT 65.795 -227.965 66.125 -227.635 ;
        RECT 65.795 -229.325 66.125 -228.995 ;
        RECT 65.795 -230.685 66.125 -230.355 ;
        RECT 65.795 -232.045 66.125 -231.715 ;
        RECT 65.795 -233.405 66.125 -233.075 ;
        RECT 65.795 -234.765 66.125 -234.435 ;
        RECT 65.795 -236.125 66.125 -235.795 ;
        RECT 65.795 -237.485 66.125 -237.155 ;
        RECT 65.795 -238.845 66.125 -238.515 ;
        RECT 65.795 -241.09 66.125 -239.96 ;
        RECT 65.8 -241.205 66.12 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 244.04 67.485 245.17 ;
        RECT 67.155 242.595 67.485 242.925 ;
        RECT 67.155 241.235 67.485 241.565 ;
        RECT 67.155 239.875 67.485 240.205 ;
        RECT 67.155 238.515 67.485 238.845 ;
        RECT 67.155 237.155 67.485 237.485 ;
        RECT 67.16 237.155 67.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 -0.845 67.485 -0.515 ;
        RECT 67.155 -2.205 67.485 -1.875 ;
        RECT 67.155 -3.565 67.485 -3.235 ;
        RECT 67.16 -3.565 67.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 -123.245 67.485 -122.915 ;
        RECT 67.155 -124.605 67.485 -124.275 ;
        RECT 67.155 -125.965 67.485 -125.635 ;
        RECT 67.155 -127.325 67.485 -126.995 ;
        RECT 67.155 -128.685 67.485 -128.355 ;
        RECT 67.155 -130.045 67.485 -129.715 ;
        RECT 67.155 -131.405 67.485 -131.075 ;
        RECT 67.155 -132.765 67.485 -132.435 ;
        RECT 67.155 -134.125 67.485 -133.795 ;
        RECT 67.155 -135.485 67.485 -135.155 ;
        RECT 67.155 -136.845 67.485 -136.515 ;
        RECT 67.155 -138.205 67.485 -137.875 ;
        RECT 67.155 -139.565 67.485 -139.235 ;
        RECT 67.155 -140.925 67.485 -140.595 ;
        RECT 67.155 -142.285 67.485 -141.955 ;
        RECT 67.155 -143.645 67.485 -143.315 ;
        RECT 67.155 -145.005 67.485 -144.675 ;
        RECT 67.155 -146.365 67.485 -146.035 ;
        RECT 67.155 -147.725 67.485 -147.395 ;
        RECT 67.155 -149.085 67.485 -148.755 ;
        RECT 67.155 -150.445 67.485 -150.115 ;
        RECT 67.155 -151.805 67.485 -151.475 ;
        RECT 67.155 -153.165 67.485 -152.835 ;
        RECT 67.155 -154.525 67.485 -154.195 ;
        RECT 67.155 -155.885 67.485 -155.555 ;
        RECT 67.155 -157.245 67.485 -156.915 ;
        RECT 67.155 -158.605 67.485 -158.275 ;
        RECT 67.155 -159.965 67.485 -159.635 ;
        RECT 67.155 -161.325 67.485 -160.995 ;
        RECT 67.155 -162.685 67.485 -162.355 ;
        RECT 67.155 -164.045 67.485 -163.715 ;
        RECT 67.155 -165.405 67.485 -165.075 ;
        RECT 67.155 -166.765 67.485 -166.435 ;
        RECT 67.155 -168.125 67.485 -167.795 ;
        RECT 67.155 -169.485 67.485 -169.155 ;
        RECT 67.155 -170.845 67.485 -170.515 ;
        RECT 67.155 -172.205 67.485 -171.875 ;
        RECT 67.155 -173.565 67.485 -173.235 ;
        RECT 67.155 -174.925 67.485 -174.595 ;
        RECT 67.155 -176.285 67.485 -175.955 ;
        RECT 67.155 -177.645 67.485 -177.315 ;
        RECT 67.155 -179.005 67.485 -178.675 ;
        RECT 67.155 -180.365 67.485 -180.035 ;
        RECT 67.155 -181.725 67.485 -181.395 ;
        RECT 67.155 -183.085 67.485 -182.755 ;
        RECT 67.155 -184.445 67.485 -184.115 ;
        RECT 67.155 -185.805 67.485 -185.475 ;
        RECT 67.155 -187.165 67.485 -186.835 ;
        RECT 67.155 -188.525 67.485 -188.195 ;
        RECT 67.155 -189.885 67.485 -189.555 ;
        RECT 67.155 -191.245 67.485 -190.915 ;
        RECT 67.155 -192.605 67.485 -192.275 ;
        RECT 67.155 -193.965 67.485 -193.635 ;
        RECT 67.155 -195.325 67.485 -194.995 ;
        RECT 67.155 -196.685 67.485 -196.355 ;
        RECT 67.155 -198.045 67.485 -197.715 ;
        RECT 67.155 -199.405 67.485 -199.075 ;
        RECT 67.155 -200.765 67.485 -200.435 ;
        RECT 67.155 -202.125 67.485 -201.795 ;
        RECT 67.155 -203.485 67.485 -203.155 ;
        RECT 67.155 -204.845 67.485 -204.515 ;
        RECT 67.155 -206.205 67.485 -205.875 ;
        RECT 67.155 -207.565 67.485 -207.235 ;
        RECT 67.155 -208.925 67.485 -208.595 ;
        RECT 67.155 -210.285 67.485 -209.955 ;
        RECT 67.155 -211.645 67.485 -211.315 ;
        RECT 67.155 -213.005 67.485 -212.675 ;
        RECT 67.155 -214.365 67.485 -214.035 ;
        RECT 67.155 -215.725 67.485 -215.395 ;
        RECT 67.155 -217.085 67.485 -216.755 ;
        RECT 67.155 -218.445 67.485 -218.115 ;
        RECT 67.155 -219.805 67.485 -219.475 ;
        RECT 67.155 -221.165 67.485 -220.835 ;
        RECT 67.155 -222.525 67.485 -222.195 ;
        RECT 67.155 -223.885 67.485 -223.555 ;
        RECT 67.155 -225.245 67.485 -224.915 ;
        RECT 67.155 -226.605 67.485 -226.275 ;
        RECT 67.155 -227.965 67.485 -227.635 ;
        RECT 67.155 -229.325 67.485 -228.995 ;
        RECT 67.155 -230.685 67.485 -230.355 ;
        RECT 67.155 -232.045 67.485 -231.715 ;
        RECT 67.155 -233.405 67.485 -233.075 ;
        RECT 67.155 -234.765 67.485 -234.435 ;
        RECT 67.155 -236.125 67.485 -235.795 ;
        RECT 67.155 -237.485 67.485 -237.155 ;
        RECT 67.155 -238.845 67.485 -238.515 ;
        RECT 67.155 -241.09 67.485 -239.96 ;
        RECT 67.16 -241.205 67.48 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 244.04 68.845 245.17 ;
        RECT 68.515 242.595 68.845 242.925 ;
        RECT 68.515 241.235 68.845 241.565 ;
        RECT 68.515 239.875 68.845 240.205 ;
        RECT 68.515 238.515 68.845 238.845 ;
        RECT 68.515 237.155 68.845 237.485 ;
        RECT 68.52 237.155 68.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 -127.325 68.845 -126.995 ;
        RECT 68.515 -128.685 68.845 -128.355 ;
        RECT 68.515 -130.045 68.845 -129.715 ;
        RECT 68.515 -131.405 68.845 -131.075 ;
        RECT 68.515 -132.765 68.845 -132.435 ;
        RECT 68.515 -134.125 68.845 -133.795 ;
        RECT 68.515 -135.485 68.845 -135.155 ;
        RECT 68.515 -136.845 68.845 -136.515 ;
        RECT 68.515 -138.205 68.845 -137.875 ;
        RECT 68.515 -139.565 68.845 -139.235 ;
        RECT 68.515 -140.925 68.845 -140.595 ;
        RECT 68.515 -142.285 68.845 -141.955 ;
        RECT 68.515 -143.645 68.845 -143.315 ;
        RECT 68.515 -145.005 68.845 -144.675 ;
        RECT 68.515 -146.365 68.845 -146.035 ;
        RECT 68.515 -147.725 68.845 -147.395 ;
        RECT 68.515 -149.085 68.845 -148.755 ;
        RECT 68.515 -150.445 68.845 -150.115 ;
        RECT 68.515 -151.805 68.845 -151.475 ;
        RECT 68.515 -153.165 68.845 -152.835 ;
        RECT 68.515 -154.525 68.845 -154.195 ;
        RECT 68.515 -155.885 68.845 -155.555 ;
        RECT 68.515 -157.245 68.845 -156.915 ;
        RECT 68.515 -158.605 68.845 -158.275 ;
        RECT 68.515 -159.965 68.845 -159.635 ;
        RECT 68.515 -161.325 68.845 -160.995 ;
        RECT 68.515 -162.685 68.845 -162.355 ;
        RECT 68.515 -164.045 68.845 -163.715 ;
        RECT 68.515 -165.405 68.845 -165.075 ;
        RECT 68.515 -166.765 68.845 -166.435 ;
        RECT 68.515 -168.125 68.845 -167.795 ;
        RECT 68.515 -169.485 68.845 -169.155 ;
        RECT 68.515 -170.845 68.845 -170.515 ;
        RECT 68.515 -172.205 68.845 -171.875 ;
        RECT 68.515 -173.565 68.845 -173.235 ;
        RECT 68.515 -174.925 68.845 -174.595 ;
        RECT 68.515 -176.285 68.845 -175.955 ;
        RECT 68.515 -177.645 68.845 -177.315 ;
        RECT 68.515 -179.005 68.845 -178.675 ;
        RECT 68.515 -180.365 68.845 -180.035 ;
        RECT 68.515 -181.725 68.845 -181.395 ;
        RECT 68.515 -183.085 68.845 -182.755 ;
        RECT 68.515 -184.445 68.845 -184.115 ;
        RECT 68.515 -185.805 68.845 -185.475 ;
        RECT 68.515 -187.165 68.845 -186.835 ;
        RECT 68.515 -188.525 68.845 -188.195 ;
        RECT 68.515 -189.885 68.845 -189.555 ;
        RECT 68.515 -191.245 68.845 -190.915 ;
        RECT 68.515 -192.605 68.845 -192.275 ;
        RECT 68.515 -193.965 68.845 -193.635 ;
        RECT 68.515 -195.325 68.845 -194.995 ;
        RECT 68.515 -196.685 68.845 -196.355 ;
        RECT 68.515 -198.045 68.845 -197.715 ;
        RECT 68.515 -199.405 68.845 -199.075 ;
        RECT 68.515 -200.765 68.845 -200.435 ;
        RECT 68.515 -202.125 68.845 -201.795 ;
        RECT 68.515 -203.485 68.845 -203.155 ;
        RECT 68.515 -204.845 68.845 -204.515 ;
        RECT 68.515 -206.205 68.845 -205.875 ;
        RECT 68.515 -207.565 68.845 -207.235 ;
        RECT 68.515 -208.925 68.845 -208.595 ;
        RECT 68.515 -210.285 68.845 -209.955 ;
        RECT 68.515 -211.645 68.845 -211.315 ;
        RECT 68.515 -213.005 68.845 -212.675 ;
        RECT 68.515 -214.365 68.845 -214.035 ;
        RECT 68.515 -215.725 68.845 -215.395 ;
        RECT 68.515 -217.085 68.845 -216.755 ;
        RECT 68.515 -218.445 68.845 -218.115 ;
        RECT 68.515 -219.805 68.845 -219.475 ;
        RECT 68.515 -221.165 68.845 -220.835 ;
        RECT 68.515 -222.525 68.845 -222.195 ;
        RECT 68.515 -223.885 68.845 -223.555 ;
        RECT 68.515 -225.245 68.845 -224.915 ;
        RECT 68.515 -226.605 68.845 -226.275 ;
        RECT 68.515 -227.965 68.845 -227.635 ;
        RECT 68.515 -229.325 68.845 -228.995 ;
        RECT 68.515 -230.685 68.845 -230.355 ;
        RECT 68.515 -232.045 68.845 -231.715 ;
        RECT 68.515 -233.405 68.845 -233.075 ;
        RECT 68.515 -234.765 68.845 -234.435 ;
        RECT 68.515 -236.125 68.845 -235.795 ;
        RECT 68.515 -237.485 68.845 -237.155 ;
        RECT 68.515 -238.845 68.845 -238.515 ;
        RECT 68.515 -241.09 68.845 -239.96 ;
        RECT 68.52 -241.205 68.84 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.71 -125.535 69.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 244.04 70.205 245.17 ;
        RECT 69.875 242.595 70.205 242.925 ;
        RECT 69.875 241.235 70.205 241.565 ;
        RECT 69.875 239.875 70.205 240.205 ;
        RECT 69.875 238.515 70.205 238.845 ;
        RECT 69.875 237.155 70.205 237.485 ;
        RECT 69.88 237.155 70.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 -0.845 70.205 -0.515 ;
        RECT 69.875 -2.205 70.205 -1.875 ;
        RECT 69.875 -3.565 70.205 -3.235 ;
        RECT 69.88 -3.565 70.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 244.04 71.565 245.17 ;
        RECT 71.235 242.595 71.565 242.925 ;
        RECT 71.235 241.235 71.565 241.565 ;
        RECT 71.235 239.875 71.565 240.205 ;
        RECT 71.235 238.515 71.565 238.845 ;
        RECT 71.235 237.155 71.565 237.485 ;
        RECT 71.24 237.155 71.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 -0.845 71.565 -0.515 ;
        RECT 71.235 -2.205 71.565 -1.875 ;
        RECT 71.235 -3.565 71.565 -3.235 ;
        RECT 71.24 -3.565 71.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 244.04 72.925 245.17 ;
        RECT 72.595 242.595 72.925 242.925 ;
        RECT 72.595 241.235 72.925 241.565 ;
        RECT 72.595 239.875 72.925 240.205 ;
        RECT 72.595 238.515 72.925 238.845 ;
        RECT 72.595 237.155 72.925 237.485 ;
        RECT 72.6 237.155 72.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 -0.845 72.925 -0.515 ;
        RECT 72.595 -2.205 72.925 -1.875 ;
        RECT 72.595 -3.565 72.925 -3.235 ;
        RECT 72.6 -3.565 72.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 -123.245 72.925 -122.915 ;
        RECT 72.595 -124.605 72.925 -124.275 ;
        RECT 72.595 -125.965 72.925 -125.635 ;
        RECT 72.595 -127.325 72.925 -126.995 ;
        RECT 72.595 -128.685 72.925 -128.355 ;
        RECT 72.595 -130.045 72.925 -129.715 ;
        RECT 72.595 -131.405 72.925 -131.075 ;
        RECT 72.595 -132.765 72.925 -132.435 ;
        RECT 72.595 -134.125 72.925 -133.795 ;
        RECT 72.595 -135.485 72.925 -135.155 ;
        RECT 72.595 -136.845 72.925 -136.515 ;
        RECT 72.595 -138.205 72.925 -137.875 ;
        RECT 72.595 -139.565 72.925 -139.235 ;
        RECT 72.595 -140.925 72.925 -140.595 ;
        RECT 72.595 -142.285 72.925 -141.955 ;
        RECT 72.595 -143.645 72.925 -143.315 ;
        RECT 72.595 -145.005 72.925 -144.675 ;
        RECT 72.595 -146.365 72.925 -146.035 ;
        RECT 72.595 -147.725 72.925 -147.395 ;
        RECT 72.595 -149.085 72.925 -148.755 ;
        RECT 72.595 -150.445 72.925 -150.115 ;
        RECT 72.595 -151.805 72.925 -151.475 ;
        RECT 72.595 -153.165 72.925 -152.835 ;
        RECT 72.595 -154.525 72.925 -154.195 ;
        RECT 72.595 -155.885 72.925 -155.555 ;
        RECT 72.595 -157.245 72.925 -156.915 ;
        RECT 72.595 -158.605 72.925 -158.275 ;
        RECT 72.595 -159.965 72.925 -159.635 ;
        RECT 72.595 -161.325 72.925 -160.995 ;
        RECT 72.595 -162.685 72.925 -162.355 ;
        RECT 72.595 -164.045 72.925 -163.715 ;
        RECT 72.595 -165.405 72.925 -165.075 ;
        RECT 72.595 -166.765 72.925 -166.435 ;
        RECT 72.595 -168.125 72.925 -167.795 ;
        RECT 72.595 -169.485 72.925 -169.155 ;
        RECT 72.595 -170.845 72.925 -170.515 ;
        RECT 72.595 -172.205 72.925 -171.875 ;
        RECT 72.595 -173.565 72.925 -173.235 ;
        RECT 72.595 -174.925 72.925 -174.595 ;
        RECT 72.595 -176.285 72.925 -175.955 ;
        RECT 72.595 -177.645 72.925 -177.315 ;
        RECT 72.595 -179.005 72.925 -178.675 ;
        RECT 72.595 -180.365 72.925 -180.035 ;
        RECT 72.595 -181.725 72.925 -181.395 ;
        RECT 72.595 -183.085 72.925 -182.755 ;
        RECT 72.595 -184.445 72.925 -184.115 ;
        RECT 72.595 -185.805 72.925 -185.475 ;
        RECT 72.595 -187.165 72.925 -186.835 ;
        RECT 72.595 -188.525 72.925 -188.195 ;
        RECT 72.595 -189.885 72.925 -189.555 ;
        RECT 72.595 -191.245 72.925 -190.915 ;
        RECT 72.595 -192.605 72.925 -192.275 ;
        RECT 72.595 -193.965 72.925 -193.635 ;
        RECT 72.595 -195.325 72.925 -194.995 ;
        RECT 72.595 -196.685 72.925 -196.355 ;
        RECT 72.595 -198.045 72.925 -197.715 ;
        RECT 72.595 -199.405 72.925 -199.075 ;
        RECT 72.595 -200.765 72.925 -200.435 ;
        RECT 72.595 -202.125 72.925 -201.795 ;
        RECT 72.595 -203.485 72.925 -203.155 ;
        RECT 72.595 -204.845 72.925 -204.515 ;
        RECT 72.595 -206.205 72.925 -205.875 ;
        RECT 72.595 -207.565 72.925 -207.235 ;
        RECT 72.595 -208.925 72.925 -208.595 ;
        RECT 72.595 -210.285 72.925 -209.955 ;
        RECT 72.595 -211.645 72.925 -211.315 ;
        RECT 72.595 -213.005 72.925 -212.675 ;
        RECT 72.595 -214.365 72.925 -214.035 ;
        RECT 72.595 -215.725 72.925 -215.395 ;
        RECT 72.595 -217.085 72.925 -216.755 ;
        RECT 72.595 -218.445 72.925 -218.115 ;
        RECT 72.595 -219.805 72.925 -219.475 ;
        RECT 72.595 -221.165 72.925 -220.835 ;
        RECT 72.595 -222.525 72.925 -222.195 ;
        RECT 72.595 -223.885 72.925 -223.555 ;
        RECT 72.595 -225.245 72.925 -224.915 ;
        RECT 72.595 -226.605 72.925 -226.275 ;
        RECT 72.595 -227.965 72.925 -227.635 ;
        RECT 72.595 -229.325 72.925 -228.995 ;
        RECT 72.595 -230.685 72.925 -230.355 ;
        RECT 72.595 -232.045 72.925 -231.715 ;
        RECT 72.595 -233.405 72.925 -233.075 ;
        RECT 72.595 -234.765 72.925 -234.435 ;
        RECT 72.595 -236.125 72.925 -235.795 ;
        RECT 72.595 -237.485 72.925 -237.155 ;
        RECT 72.595 -238.845 72.925 -238.515 ;
        RECT 72.595 -241.09 72.925 -239.96 ;
        RECT 72.6 -241.205 72.92 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 244.04 74.285 245.17 ;
        RECT 73.955 242.595 74.285 242.925 ;
        RECT 73.955 241.235 74.285 241.565 ;
        RECT 73.955 239.875 74.285 240.205 ;
        RECT 73.955 238.515 74.285 238.845 ;
        RECT 73.955 237.155 74.285 237.485 ;
        RECT 73.96 237.155 74.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -0.845 74.285 -0.515 ;
        RECT 73.955 -2.205 74.285 -1.875 ;
        RECT 73.955 -3.565 74.285 -3.235 ;
        RECT 73.96 -3.565 74.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -123.245 74.285 -122.915 ;
        RECT 73.955 -124.605 74.285 -124.275 ;
        RECT 73.955 -125.965 74.285 -125.635 ;
        RECT 73.955 -127.325 74.285 -126.995 ;
        RECT 73.955 -128.685 74.285 -128.355 ;
        RECT 73.955 -130.045 74.285 -129.715 ;
        RECT 73.955 -131.405 74.285 -131.075 ;
        RECT 73.955 -132.765 74.285 -132.435 ;
        RECT 73.955 -134.125 74.285 -133.795 ;
        RECT 73.955 -135.485 74.285 -135.155 ;
        RECT 73.955 -136.845 74.285 -136.515 ;
        RECT 73.955 -138.205 74.285 -137.875 ;
        RECT 73.955 -139.565 74.285 -139.235 ;
        RECT 73.955 -140.925 74.285 -140.595 ;
        RECT 73.955 -142.285 74.285 -141.955 ;
        RECT 73.955 -143.645 74.285 -143.315 ;
        RECT 73.955 -145.005 74.285 -144.675 ;
        RECT 73.955 -146.365 74.285 -146.035 ;
        RECT 73.955 -147.725 74.285 -147.395 ;
        RECT 73.955 -149.085 74.285 -148.755 ;
        RECT 73.955 -150.445 74.285 -150.115 ;
        RECT 73.955 -151.805 74.285 -151.475 ;
        RECT 73.955 -153.165 74.285 -152.835 ;
        RECT 73.955 -154.525 74.285 -154.195 ;
        RECT 73.955 -155.885 74.285 -155.555 ;
        RECT 73.955 -157.245 74.285 -156.915 ;
        RECT 73.955 -158.605 74.285 -158.275 ;
        RECT 73.955 -159.965 74.285 -159.635 ;
        RECT 73.955 -161.325 74.285 -160.995 ;
        RECT 73.955 -162.685 74.285 -162.355 ;
        RECT 73.955 -164.045 74.285 -163.715 ;
        RECT 73.955 -165.405 74.285 -165.075 ;
        RECT 73.955 -166.765 74.285 -166.435 ;
        RECT 73.955 -168.125 74.285 -167.795 ;
        RECT 73.955 -169.485 74.285 -169.155 ;
        RECT 73.955 -170.845 74.285 -170.515 ;
        RECT 73.955 -172.205 74.285 -171.875 ;
        RECT 73.955 -173.565 74.285 -173.235 ;
        RECT 73.955 -174.925 74.285 -174.595 ;
        RECT 73.955 -176.285 74.285 -175.955 ;
        RECT 73.955 -177.645 74.285 -177.315 ;
        RECT 73.955 -179.005 74.285 -178.675 ;
        RECT 73.955 -180.365 74.285 -180.035 ;
        RECT 73.955 -181.725 74.285 -181.395 ;
        RECT 73.955 -183.085 74.285 -182.755 ;
        RECT 73.955 -184.445 74.285 -184.115 ;
        RECT 73.955 -185.805 74.285 -185.475 ;
        RECT 73.955 -187.165 74.285 -186.835 ;
        RECT 73.955 -188.525 74.285 -188.195 ;
        RECT 73.955 -189.885 74.285 -189.555 ;
        RECT 73.955 -191.245 74.285 -190.915 ;
        RECT 73.955 -192.605 74.285 -192.275 ;
        RECT 73.955 -193.965 74.285 -193.635 ;
        RECT 73.955 -195.325 74.285 -194.995 ;
        RECT 73.955 -196.685 74.285 -196.355 ;
        RECT 73.955 -198.045 74.285 -197.715 ;
        RECT 73.955 -199.405 74.285 -199.075 ;
        RECT 73.955 -200.765 74.285 -200.435 ;
        RECT 73.955 -202.125 74.285 -201.795 ;
        RECT 73.955 -203.485 74.285 -203.155 ;
        RECT 73.955 -204.845 74.285 -204.515 ;
        RECT 73.955 -206.205 74.285 -205.875 ;
        RECT 73.955 -207.565 74.285 -207.235 ;
        RECT 73.955 -208.925 74.285 -208.595 ;
        RECT 73.955 -210.285 74.285 -209.955 ;
        RECT 73.955 -211.645 74.285 -211.315 ;
        RECT 73.955 -213.005 74.285 -212.675 ;
        RECT 73.955 -214.365 74.285 -214.035 ;
        RECT 73.955 -215.725 74.285 -215.395 ;
        RECT 73.955 -217.085 74.285 -216.755 ;
        RECT 73.955 -218.445 74.285 -218.115 ;
        RECT 73.955 -219.805 74.285 -219.475 ;
        RECT 73.955 -221.165 74.285 -220.835 ;
        RECT 73.955 -222.525 74.285 -222.195 ;
        RECT 73.955 -223.885 74.285 -223.555 ;
        RECT 73.955 -225.245 74.285 -224.915 ;
        RECT 73.955 -226.605 74.285 -226.275 ;
        RECT 73.955 -227.965 74.285 -227.635 ;
        RECT 73.955 -229.325 74.285 -228.995 ;
        RECT 73.955 -230.685 74.285 -230.355 ;
        RECT 73.955 -232.045 74.285 -231.715 ;
        RECT 73.955 -233.405 74.285 -233.075 ;
        RECT 73.955 -234.765 74.285 -234.435 ;
        RECT 73.955 -236.125 74.285 -235.795 ;
        RECT 73.955 -237.485 74.285 -237.155 ;
        RECT 73.955 -238.845 74.285 -238.515 ;
        RECT 73.955 -241.09 74.285 -239.96 ;
        RECT 73.96 -241.205 74.28 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 244.04 75.645 245.17 ;
        RECT 75.315 242.595 75.645 242.925 ;
        RECT 75.315 241.235 75.645 241.565 ;
        RECT 75.315 239.875 75.645 240.205 ;
        RECT 75.315 238.515 75.645 238.845 ;
        RECT 75.315 237.155 75.645 237.485 ;
        RECT 75.32 237.155 75.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 -0.845 75.645 -0.515 ;
        RECT 75.315 -2.205 75.645 -1.875 ;
        RECT 75.315 -3.565 75.645 -3.235 ;
        RECT 75.32 -3.565 75.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 -177.645 75.645 -177.315 ;
        RECT 75.315 -179.005 75.645 -178.675 ;
        RECT 75.315 -180.365 75.645 -180.035 ;
        RECT 75.315 -181.725 75.645 -181.395 ;
        RECT 75.315 -183.085 75.645 -182.755 ;
        RECT 75.315 -184.445 75.645 -184.115 ;
        RECT 75.315 -185.805 75.645 -185.475 ;
        RECT 75.315 -187.165 75.645 -186.835 ;
        RECT 75.315 -188.525 75.645 -188.195 ;
        RECT 75.315 -189.885 75.645 -189.555 ;
        RECT 75.315 -191.245 75.645 -190.915 ;
        RECT 75.315 -192.605 75.645 -192.275 ;
        RECT 75.315 -193.965 75.645 -193.635 ;
        RECT 75.315 -195.325 75.645 -194.995 ;
        RECT 75.315 -196.685 75.645 -196.355 ;
        RECT 75.315 -198.045 75.645 -197.715 ;
        RECT 75.315 -199.405 75.645 -199.075 ;
        RECT 75.315 -200.765 75.645 -200.435 ;
        RECT 75.315 -202.125 75.645 -201.795 ;
        RECT 75.315 -203.485 75.645 -203.155 ;
        RECT 75.315 -204.845 75.645 -204.515 ;
        RECT 75.315 -206.205 75.645 -205.875 ;
        RECT 75.315 -207.565 75.645 -207.235 ;
        RECT 75.315 -208.925 75.645 -208.595 ;
        RECT 75.315 -210.285 75.645 -209.955 ;
        RECT 75.315 -211.645 75.645 -211.315 ;
        RECT 75.315 -213.005 75.645 -212.675 ;
        RECT 75.315 -214.365 75.645 -214.035 ;
        RECT 75.315 -215.725 75.645 -215.395 ;
        RECT 75.315 -217.085 75.645 -216.755 ;
        RECT 75.315 -218.445 75.645 -218.115 ;
        RECT 75.315 -219.805 75.645 -219.475 ;
        RECT 75.315 -221.165 75.645 -220.835 ;
        RECT 75.315 -222.525 75.645 -222.195 ;
        RECT 75.315 -223.885 75.645 -223.555 ;
        RECT 75.315 -225.245 75.645 -224.915 ;
        RECT 75.315 -226.605 75.645 -226.275 ;
        RECT 75.315 -227.965 75.645 -227.635 ;
        RECT 75.315 -229.325 75.645 -228.995 ;
        RECT 75.315 -230.685 75.645 -230.355 ;
        RECT 75.315 -232.045 75.645 -231.715 ;
        RECT 75.315 -233.405 75.645 -233.075 ;
        RECT 75.315 -234.765 75.645 -234.435 ;
        RECT 75.315 -236.125 75.645 -235.795 ;
        RECT 75.315 -237.485 75.645 -237.155 ;
        RECT 75.315 -238.845 75.645 -238.515 ;
        RECT 75.315 -241.09 75.645 -239.96 ;
        RECT 75.32 -241.205 75.64 -122.24 ;
        RECT 75.315 -123.245 75.645 -122.915 ;
        RECT 75.315 -124.605 75.645 -124.275 ;
        RECT 75.315 -125.965 75.645 -125.635 ;
        RECT 75.315 -127.325 75.645 -126.995 ;
        RECT 75.315 -128.685 75.645 -128.355 ;
        RECT 75.315 -130.045 75.645 -129.715 ;
        RECT 75.315 -131.405 75.645 -131.075 ;
        RECT 75.315 -132.765 75.645 -132.435 ;
        RECT 75.315 -134.125 75.645 -133.795 ;
        RECT 75.315 -135.485 75.645 -135.155 ;
        RECT 75.315 -136.845 75.645 -136.515 ;
        RECT 75.315 -138.205 75.645 -137.875 ;
        RECT 75.315 -139.565 75.645 -139.235 ;
        RECT 75.315 -140.925 75.645 -140.595 ;
        RECT 75.315 -142.285 75.645 -141.955 ;
        RECT 75.315 -143.645 75.645 -143.315 ;
        RECT 75.315 -145.005 75.645 -144.675 ;
        RECT 75.315 -146.365 75.645 -146.035 ;
        RECT 75.315 -147.725 75.645 -147.395 ;
        RECT 75.315 -149.085 75.645 -148.755 ;
        RECT 75.315 -150.445 75.645 -150.115 ;
        RECT 75.315 -151.805 75.645 -151.475 ;
        RECT 75.315 -153.165 75.645 -152.835 ;
        RECT 75.315 -154.525 75.645 -154.195 ;
        RECT 75.315 -155.885 75.645 -155.555 ;
        RECT 75.315 -157.245 75.645 -156.915 ;
        RECT 75.315 -158.605 75.645 -158.275 ;
        RECT 75.315 -159.965 75.645 -159.635 ;
        RECT 75.315 -161.325 75.645 -160.995 ;
        RECT 75.315 -162.685 75.645 -162.355 ;
        RECT 75.315 -164.045 75.645 -163.715 ;
        RECT 75.315 -165.405 75.645 -165.075 ;
        RECT 75.315 -166.765 75.645 -166.435 ;
        RECT 75.315 -168.125 75.645 -167.795 ;
        RECT 75.315 -169.485 75.645 -169.155 ;
        RECT 75.315 -170.845 75.645 -170.515 ;
        RECT 75.315 -172.205 75.645 -171.875 ;
        RECT 75.315 -173.565 75.645 -173.235 ;
        RECT 75.315 -174.925 75.645 -174.595 ;
        RECT 75.315 -176.285 75.645 -175.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 244.04 41.645 245.17 ;
        RECT 41.315 242.595 41.645 242.925 ;
        RECT 41.315 241.235 41.645 241.565 ;
        RECT 41.315 239.875 41.645 240.205 ;
        RECT 41.315 238.515 41.645 238.845 ;
        RECT 41.315 237.155 41.645 237.485 ;
        RECT 41.32 237.155 41.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 -0.845 41.645 -0.515 ;
        RECT 41.315 -2.205 41.645 -1.875 ;
        RECT 41.315 -3.565 41.645 -3.235 ;
        RECT 41.32 -3.565 41.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 -123.245 41.645 -122.915 ;
        RECT 41.315 -124.605 41.645 -124.275 ;
        RECT 41.315 -125.965 41.645 -125.635 ;
        RECT 41.315 -127.325 41.645 -126.995 ;
        RECT 41.315 -128.685 41.645 -128.355 ;
        RECT 41.315 -130.045 41.645 -129.715 ;
        RECT 41.315 -131.405 41.645 -131.075 ;
        RECT 41.315 -132.765 41.645 -132.435 ;
        RECT 41.315 -134.125 41.645 -133.795 ;
        RECT 41.315 -135.485 41.645 -135.155 ;
        RECT 41.315 -136.845 41.645 -136.515 ;
        RECT 41.315 -138.205 41.645 -137.875 ;
        RECT 41.315 -139.565 41.645 -139.235 ;
        RECT 41.315 -140.925 41.645 -140.595 ;
        RECT 41.315 -142.285 41.645 -141.955 ;
        RECT 41.315 -143.645 41.645 -143.315 ;
        RECT 41.315 -145.005 41.645 -144.675 ;
        RECT 41.315 -146.365 41.645 -146.035 ;
        RECT 41.315 -147.725 41.645 -147.395 ;
        RECT 41.315 -149.085 41.645 -148.755 ;
        RECT 41.315 -150.445 41.645 -150.115 ;
        RECT 41.315 -151.805 41.645 -151.475 ;
        RECT 41.315 -153.165 41.645 -152.835 ;
        RECT 41.315 -154.525 41.645 -154.195 ;
        RECT 41.315 -155.885 41.645 -155.555 ;
        RECT 41.315 -157.245 41.645 -156.915 ;
        RECT 41.315 -158.605 41.645 -158.275 ;
        RECT 41.315 -159.965 41.645 -159.635 ;
        RECT 41.315 -161.325 41.645 -160.995 ;
        RECT 41.315 -162.685 41.645 -162.355 ;
        RECT 41.315 -164.045 41.645 -163.715 ;
        RECT 41.315 -165.405 41.645 -165.075 ;
        RECT 41.315 -166.765 41.645 -166.435 ;
        RECT 41.315 -168.125 41.645 -167.795 ;
        RECT 41.315 -169.485 41.645 -169.155 ;
        RECT 41.315 -170.845 41.645 -170.515 ;
        RECT 41.315 -172.205 41.645 -171.875 ;
        RECT 41.315 -173.565 41.645 -173.235 ;
        RECT 41.315 -174.925 41.645 -174.595 ;
        RECT 41.315 -176.285 41.645 -175.955 ;
        RECT 41.315 -177.645 41.645 -177.315 ;
        RECT 41.315 -179.005 41.645 -178.675 ;
        RECT 41.315 -180.365 41.645 -180.035 ;
        RECT 41.315 -181.725 41.645 -181.395 ;
        RECT 41.315 -183.085 41.645 -182.755 ;
        RECT 41.315 -184.445 41.645 -184.115 ;
        RECT 41.315 -185.805 41.645 -185.475 ;
        RECT 41.315 -187.165 41.645 -186.835 ;
        RECT 41.315 -188.525 41.645 -188.195 ;
        RECT 41.315 -189.885 41.645 -189.555 ;
        RECT 41.315 -191.245 41.645 -190.915 ;
        RECT 41.315 -192.605 41.645 -192.275 ;
        RECT 41.315 -193.965 41.645 -193.635 ;
        RECT 41.315 -195.325 41.645 -194.995 ;
        RECT 41.315 -196.685 41.645 -196.355 ;
        RECT 41.315 -198.045 41.645 -197.715 ;
        RECT 41.315 -199.405 41.645 -199.075 ;
        RECT 41.315 -200.765 41.645 -200.435 ;
        RECT 41.315 -202.125 41.645 -201.795 ;
        RECT 41.315 -203.485 41.645 -203.155 ;
        RECT 41.315 -204.845 41.645 -204.515 ;
        RECT 41.315 -206.205 41.645 -205.875 ;
        RECT 41.315 -207.565 41.645 -207.235 ;
        RECT 41.315 -208.925 41.645 -208.595 ;
        RECT 41.315 -210.285 41.645 -209.955 ;
        RECT 41.315 -211.645 41.645 -211.315 ;
        RECT 41.315 -213.005 41.645 -212.675 ;
        RECT 41.315 -214.365 41.645 -214.035 ;
        RECT 41.315 -215.725 41.645 -215.395 ;
        RECT 41.315 -217.085 41.645 -216.755 ;
        RECT 41.315 -218.445 41.645 -218.115 ;
        RECT 41.315 -219.805 41.645 -219.475 ;
        RECT 41.315 -221.165 41.645 -220.835 ;
        RECT 41.315 -222.525 41.645 -222.195 ;
        RECT 41.315 -223.885 41.645 -223.555 ;
        RECT 41.315 -225.245 41.645 -224.915 ;
        RECT 41.315 -226.605 41.645 -226.275 ;
        RECT 41.315 -227.965 41.645 -227.635 ;
        RECT 41.315 -229.325 41.645 -228.995 ;
        RECT 41.315 -230.685 41.645 -230.355 ;
        RECT 41.315 -232.045 41.645 -231.715 ;
        RECT 41.315 -233.405 41.645 -233.075 ;
        RECT 41.315 -234.765 41.645 -234.435 ;
        RECT 41.315 -236.125 41.645 -235.795 ;
        RECT 41.315 -237.485 41.645 -237.155 ;
        RECT 41.315 -238.845 41.645 -238.515 ;
        RECT 41.315 -241.09 41.645 -239.96 ;
        RECT 41.32 -241.205 41.64 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 244.04 43.005 245.17 ;
        RECT 42.675 242.595 43.005 242.925 ;
        RECT 42.675 241.235 43.005 241.565 ;
        RECT 42.675 239.875 43.005 240.205 ;
        RECT 42.675 238.515 43.005 238.845 ;
        RECT 42.675 237.155 43.005 237.485 ;
        RECT 42.68 237.155 43 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 -0.845 43.005 -0.515 ;
        RECT 42.675 -2.205 43.005 -1.875 ;
        RECT 42.675 -3.565 43.005 -3.235 ;
        RECT 42.68 -3.565 43 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 -123.245 43.005 -122.915 ;
        RECT 42.675 -124.605 43.005 -124.275 ;
        RECT 42.675 -125.965 43.005 -125.635 ;
        RECT 42.675 -127.325 43.005 -126.995 ;
        RECT 42.675 -128.685 43.005 -128.355 ;
        RECT 42.675 -130.045 43.005 -129.715 ;
        RECT 42.675 -131.405 43.005 -131.075 ;
        RECT 42.675 -132.765 43.005 -132.435 ;
        RECT 42.675 -134.125 43.005 -133.795 ;
        RECT 42.675 -135.485 43.005 -135.155 ;
        RECT 42.675 -136.845 43.005 -136.515 ;
        RECT 42.675 -138.205 43.005 -137.875 ;
        RECT 42.675 -139.565 43.005 -139.235 ;
        RECT 42.675 -140.925 43.005 -140.595 ;
        RECT 42.675 -142.285 43.005 -141.955 ;
        RECT 42.675 -143.645 43.005 -143.315 ;
        RECT 42.675 -145.005 43.005 -144.675 ;
        RECT 42.675 -146.365 43.005 -146.035 ;
        RECT 42.675 -147.725 43.005 -147.395 ;
        RECT 42.675 -149.085 43.005 -148.755 ;
        RECT 42.675 -150.445 43.005 -150.115 ;
        RECT 42.675 -151.805 43.005 -151.475 ;
        RECT 42.675 -153.165 43.005 -152.835 ;
        RECT 42.675 -154.525 43.005 -154.195 ;
        RECT 42.675 -155.885 43.005 -155.555 ;
        RECT 42.675 -157.245 43.005 -156.915 ;
        RECT 42.675 -158.605 43.005 -158.275 ;
        RECT 42.675 -159.965 43.005 -159.635 ;
        RECT 42.675 -161.325 43.005 -160.995 ;
        RECT 42.675 -162.685 43.005 -162.355 ;
        RECT 42.675 -164.045 43.005 -163.715 ;
        RECT 42.675 -165.405 43.005 -165.075 ;
        RECT 42.675 -166.765 43.005 -166.435 ;
        RECT 42.675 -168.125 43.005 -167.795 ;
        RECT 42.675 -169.485 43.005 -169.155 ;
        RECT 42.675 -170.845 43.005 -170.515 ;
        RECT 42.675 -172.205 43.005 -171.875 ;
        RECT 42.675 -173.565 43.005 -173.235 ;
        RECT 42.675 -174.925 43.005 -174.595 ;
        RECT 42.675 -176.285 43.005 -175.955 ;
        RECT 42.675 -177.645 43.005 -177.315 ;
        RECT 42.675 -179.005 43.005 -178.675 ;
        RECT 42.675 -180.365 43.005 -180.035 ;
        RECT 42.675 -181.725 43.005 -181.395 ;
        RECT 42.675 -183.085 43.005 -182.755 ;
        RECT 42.675 -184.445 43.005 -184.115 ;
        RECT 42.675 -185.805 43.005 -185.475 ;
        RECT 42.675 -187.165 43.005 -186.835 ;
        RECT 42.675 -188.525 43.005 -188.195 ;
        RECT 42.675 -189.885 43.005 -189.555 ;
        RECT 42.675 -191.245 43.005 -190.915 ;
        RECT 42.675 -192.605 43.005 -192.275 ;
        RECT 42.675 -193.965 43.005 -193.635 ;
        RECT 42.675 -195.325 43.005 -194.995 ;
        RECT 42.675 -196.685 43.005 -196.355 ;
        RECT 42.675 -198.045 43.005 -197.715 ;
        RECT 42.675 -199.405 43.005 -199.075 ;
        RECT 42.675 -200.765 43.005 -200.435 ;
        RECT 42.675 -202.125 43.005 -201.795 ;
        RECT 42.675 -203.485 43.005 -203.155 ;
        RECT 42.675 -204.845 43.005 -204.515 ;
        RECT 42.675 -206.205 43.005 -205.875 ;
        RECT 42.675 -207.565 43.005 -207.235 ;
        RECT 42.675 -208.925 43.005 -208.595 ;
        RECT 42.675 -210.285 43.005 -209.955 ;
        RECT 42.675 -211.645 43.005 -211.315 ;
        RECT 42.675 -213.005 43.005 -212.675 ;
        RECT 42.675 -214.365 43.005 -214.035 ;
        RECT 42.675 -215.725 43.005 -215.395 ;
        RECT 42.675 -217.085 43.005 -216.755 ;
        RECT 42.675 -218.445 43.005 -218.115 ;
        RECT 42.675 -219.805 43.005 -219.475 ;
        RECT 42.675 -221.165 43.005 -220.835 ;
        RECT 42.675 -222.525 43.005 -222.195 ;
        RECT 42.675 -223.885 43.005 -223.555 ;
        RECT 42.675 -225.245 43.005 -224.915 ;
        RECT 42.675 -226.605 43.005 -226.275 ;
        RECT 42.675 -227.965 43.005 -227.635 ;
        RECT 42.675 -229.325 43.005 -228.995 ;
        RECT 42.675 -230.685 43.005 -230.355 ;
        RECT 42.675 -232.045 43.005 -231.715 ;
        RECT 42.675 -233.405 43.005 -233.075 ;
        RECT 42.675 -234.765 43.005 -234.435 ;
        RECT 42.675 -236.125 43.005 -235.795 ;
        RECT 42.675 -237.485 43.005 -237.155 ;
        RECT 42.675 -238.845 43.005 -238.515 ;
        RECT 42.675 -241.09 43.005 -239.96 ;
        RECT 42.68 -241.205 43 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 244.04 44.365 245.17 ;
        RECT 44.035 242.595 44.365 242.925 ;
        RECT 44.035 241.235 44.365 241.565 ;
        RECT 44.035 239.875 44.365 240.205 ;
        RECT 44.035 238.515 44.365 238.845 ;
        RECT 44.035 237.155 44.365 237.485 ;
        RECT 44.04 237.155 44.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -0.845 44.365 -0.515 ;
        RECT 44.035 -2.205 44.365 -1.875 ;
        RECT 44.035 -3.565 44.365 -3.235 ;
        RECT 44.04 -3.565 44.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -123.245 44.365 -122.915 ;
        RECT 44.035 -124.605 44.365 -124.275 ;
        RECT 44.035 -125.965 44.365 -125.635 ;
        RECT 44.035 -127.325 44.365 -126.995 ;
        RECT 44.035 -128.685 44.365 -128.355 ;
        RECT 44.035 -130.045 44.365 -129.715 ;
        RECT 44.035 -131.405 44.365 -131.075 ;
        RECT 44.035 -132.765 44.365 -132.435 ;
        RECT 44.035 -134.125 44.365 -133.795 ;
        RECT 44.035 -135.485 44.365 -135.155 ;
        RECT 44.035 -136.845 44.365 -136.515 ;
        RECT 44.035 -138.205 44.365 -137.875 ;
        RECT 44.035 -139.565 44.365 -139.235 ;
        RECT 44.035 -140.925 44.365 -140.595 ;
        RECT 44.035 -142.285 44.365 -141.955 ;
        RECT 44.035 -143.645 44.365 -143.315 ;
        RECT 44.035 -145.005 44.365 -144.675 ;
        RECT 44.035 -146.365 44.365 -146.035 ;
        RECT 44.035 -147.725 44.365 -147.395 ;
        RECT 44.035 -149.085 44.365 -148.755 ;
        RECT 44.035 -150.445 44.365 -150.115 ;
        RECT 44.035 -151.805 44.365 -151.475 ;
        RECT 44.035 -153.165 44.365 -152.835 ;
        RECT 44.035 -154.525 44.365 -154.195 ;
        RECT 44.035 -155.885 44.365 -155.555 ;
        RECT 44.035 -157.245 44.365 -156.915 ;
        RECT 44.035 -158.605 44.365 -158.275 ;
        RECT 44.035 -159.965 44.365 -159.635 ;
        RECT 44.035 -161.325 44.365 -160.995 ;
        RECT 44.035 -162.685 44.365 -162.355 ;
        RECT 44.035 -164.045 44.365 -163.715 ;
        RECT 44.035 -165.405 44.365 -165.075 ;
        RECT 44.035 -166.765 44.365 -166.435 ;
        RECT 44.035 -168.125 44.365 -167.795 ;
        RECT 44.035 -169.485 44.365 -169.155 ;
        RECT 44.035 -170.845 44.365 -170.515 ;
        RECT 44.035 -172.205 44.365 -171.875 ;
        RECT 44.035 -173.565 44.365 -173.235 ;
        RECT 44.035 -174.925 44.365 -174.595 ;
        RECT 44.035 -176.285 44.365 -175.955 ;
        RECT 44.035 -177.645 44.365 -177.315 ;
        RECT 44.035 -179.005 44.365 -178.675 ;
        RECT 44.035 -180.365 44.365 -180.035 ;
        RECT 44.035 -181.725 44.365 -181.395 ;
        RECT 44.035 -183.085 44.365 -182.755 ;
        RECT 44.035 -184.445 44.365 -184.115 ;
        RECT 44.035 -185.805 44.365 -185.475 ;
        RECT 44.035 -187.165 44.365 -186.835 ;
        RECT 44.035 -188.525 44.365 -188.195 ;
        RECT 44.035 -189.885 44.365 -189.555 ;
        RECT 44.035 -191.245 44.365 -190.915 ;
        RECT 44.035 -192.605 44.365 -192.275 ;
        RECT 44.035 -193.965 44.365 -193.635 ;
        RECT 44.035 -195.325 44.365 -194.995 ;
        RECT 44.035 -196.685 44.365 -196.355 ;
        RECT 44.035 -198.045 44.365 -197.715 ;
        RECT 44.035 -199.405 44.365 -199.075 ;
        RECT 44.035 -200.765 44.365 -200.435 ;
        RECT 44.035 -202.125 44.365 -201.795 ;
        RECT 44.035 -203.485 44.365 -203.155 ;
        RECT 44.035 -204.845 44.365 -204.515 ;
        RECT 44.035 -206.205 44.365 -205.875 ;
        RECT 44.035 -207.565 44.365 -207.235 ;
        RECT 44.035 -208.925 44.365 -208.595 ;
        RECT 44.035 -210.285 44.365 -209.955 ;
        RECT 44.035 -211.645 44.365 -211.315 ;
        RECT 44.035 -213.005 44.365 -212.675 ;
        RECT 44.035 -214.365 44.365 -214.035 ;
        RECT 44.035 -215.725 44.365 -215.395 ;
        RECT 44.035 -217.085 44.365 -216.755 ;
        RECT 44.035 -218.445 44.365 -218.115 ;
        RECT 44.035 -219.805 44.365 -219.475 ;
        RECT 44.035 -221.165 44.365 -220.835 ;
        RECT 44.035 -222.525 44.365 -222.195 ;
        RECT 44.035 -223.885 44.365 -223.555 ;
        RECT 44.035 -225.245 44.365 -224.915 ;
        RECT 44.035 -226.605 44.365 -226.275 ;
        RECT 44.035 -227.965 44.365 -227.635 ;
        RECT 44.035 -229.325 44.365 -228.995 ;
        RECT 44.035 -230.685 44.365 -230.355 ;
        RECT 44.035 -232.045 44.365 -231.715 ;
        RECT 44.035 -233.405 44.365 -233.075 ;
        RECT 44.035 -234.765 44.365 -234.435 ;
        RECT 44.035 -236.125 44.365 -235.795 ;
        RECT 44.035 -237.485 44.365 -237.155 ;
        RECT 44.035 -238.845 44.365 -238.515 ;
        RECT 44.035 -241.09 44.365 -239.96 ;
        RECT 44.04 -241.205 44.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 244.04 45.725 245.17 ;
        RECT 45.395 242.595 45.725 242.925 ;
        RECT 45.395 241.235 45.725 241.565 ;
        RECT 45.395 239.875 45.725 240.205 ;
        RECT 45.395 238.515 45.725 238.845 ;
        RECT 45.395 237.155 45.725 237.485 ;
        RECT 45.4 237.155 45.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 -0.845 45.725 -0.515 ;
        RECT 45.395 -2.205 45.725 -1.875 ;
        RECT 45.395 -3.565 45.725 -3.235 ;
        RECT 45.4 -3.565 45.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 -123.245 45.725 -122.915 ;
        RECT 45.395 -124.605 45.725 -124.275 ;
        RECT 45.395 -125.965 45.725 -125.635 ;
        RECT 45.395 -127.325 45.725 -126.995 ;
        RECT 45.395 -128.685 45.725 -128.355 ;
        RECT 45.395 -130.045 45.725 -129.715 ;
        RECT 45.395 -131.405 45.725 -131.075 ;
        RECT 45.395 -132.765 45.725 -132.435 ;
        RECT 45.395 -134.125 45.725 -133.795 ;
        RECT 45.395 -135.485 45.725 -135.155 ;
        RECT 45.395 -136.845 45.725 -136.515 ;
        RECT 45.395 -138.205 45.725 -137.875 ;
        RECT 45.395 -139.565 45.725 -139.235 ;
        RECT 45.395 -140.925 45.725 -140.595 ;
        RECT 45.395 -142.285 45.725 -141.955 ;
        RECT 45.395 -143.645 45.725 -143.315 ;
        RECT 45.395 -145.005 45.725 -144.675 ;
        RECT 45.395 -146.365 45.725 -146.035 ;
        RECT 45.395 -147.725 45.725 -147.395 ;
        RECT 45.395 -149.085 45.725 -148.755 ;
        RECT 45.395 -150.445 45.725 -150.115 ;
        RECT 45.395 -151.805 45.725 -151.475 ;
        RECT 45.395 -153.165 45.725 -152.835 ;
        RECT 45.395 -154.525 45.725 -154.195 ;
        RECT 45.395 -155.885 45.725 -155.555 ;
        RECT 45.395 -157.245 45.725 -156.915 ;
        RECT 45.395 -158.605 45.725 -158.275 ;
        RECT 45.395 -159.965 45.725 -159.635 ;
        RECT 45.395 -161.325 45.725 -160.995 ;
        RECT 45.395 -162.685 45.725 -162.355 ;
        RECT 45.395 -164.045 45.725 -163.715 ;
        RECT 45.395 -165.405 45.725 -165.075 ;
        RECT 45.395 -166.765 45.725 -166.435 ;
        RECT 45.395 -168.125 45.725 -167.795 ;
        RECT 45.395 -169.485 45.725 -169.155 ;
        RECT 45.395 -170.845 45.725 -170.515 ;
        RECT 45.395 -172.205 45.725 -171.875 ;
        RECT 45.395 -173.565 45.725 -173.235 ;
        RECT 45.395 -174.925 45.725 -174.595 ;
        RECT 45.395 -176.285 45.725 -175.955 ;
        RECT 45.395 -177.645 45.725 -177.315 ;
        RECT 45.395 -179.005 45.725 -178.675 ;
        RECT 45.395 -180.365 45.725 -180.035 ;
        RECT 45.395 -181.725 45.725 -181.395 ;
        RECT 45.395 -183.085 45.725 -182.755 ;
        RECT 45.395 -184.445 45.725 -184.115 ;
        RECT 45.395 -185.805 45.725 -185.475 ;
        RECT 45.395 -187.165 45.725 -186.835 ;
        RECT 45.395 -188.525 45.725 -188.195 ;
        RECT 45.395 -189.885 45.725 -189.555 ;
        RECT 45.395 -191.245 45.725 -190.915 ;
        RECT 45.395 -192.605 45.725 -192.275 ;
        RECT 45.395 -193.965 45.725 -193.635 ;
        RECT 45.395 -195.325 45.725 -194.995 ;
        RECT 45.395 -196.685 45.725 -196.355 ;
        RECT 45.395 -198.045 45.725 -197.715 ;
        RECT 45.395 -199.405 45.725 -199.075 ;
        RECT 45.395 -200.765 45.725 -200.435 ;
        RECT 45.395 -202.125 45.725 -201.795 ;
        RECT 45.395 -203.485 45.725 -203.155 ;
        RECT 45.395 -204.845 45.725 -204.515 ;
        RECT 45.395 -206.205 45.725 -205.875 ;
        RECT 45.395 -207.565 45.725 -207.235 ;
        RECT 45.395 -208.925 45.725 -208.595 ;
        RECT 45.395 -210.285 45.725 -209.955 ;
        RECT 45.395 -211.645 45.725 -211.315 ;
        RECT 45.395 -213.005 45.725 -212.675 ;
        RECT 45.395 -214.365 45.725 -214.035 ;
        RECT 45.395 -215.725 45.725 -215.395 ;
        RECT 45.395 -217.085 45.725 -216.755 ;
        RECT 45.395 -218.445 45.725 -218.115 ;
        RECT 45.395 -219.805 45.725 -219.475 ;
        RECT 45.395 -221.165 45.725 -220.835 ;
        RECT 45.395 -222.525 45.725 -222.195 ;
        RECT 45.395 -223.885 45.725 -223.555 ;
        RECT 45.395 -225.245 45.725 -224.915 ;
        RECT 45.395 -226.605 45.725 -226.275 ;
        RECT 45.395 -227.965 45.725 -227.635 ;
        RECT 45.395 -229.325 45.725 -228.995 ;
        RECT 45.395 -230.685 45.725 -230.355 ;
        RECT 45.395 -232.045 45.725 -231.715 ;
        RECT 45.395 -233.405 45.725 -233.075 ;
        RECT 45.395 -234.765 45.725 -234.435 ;
        RECT 45.395 -236.125 45.725 -235.795 ;
        RECT 45.395 -237.485 45.725 -237.155 ;
        RECT 45.395 -238.845 45.725 -238.515 ;
        RECT 45.395 -241.09 45.725 -239.96 ;
        RECT 45.4 -241.205 45.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 244.04 47.085 245.17 ;
        RECT 46.755 242.595 47.085 242.925 ;
        RECT 46.755 241.235 47.085 241.565 ;
        RECT 46.755 239.875 47.085 240.205 ;
        RECT 46.755 238.515 47.085 238.845 ;
        RECT 46.755 237.155 47.085 237.485 ;
        RECT 46.76 237.155 47.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 -127.325 47.085 -126.995 ;
        RECT 46.755 -128.685 47.085 -128.355 ;
        RECT 46.755 -130.045 47.085 -129.715 ;
        RECT 46.755 -131.405 47.085 -131.075 ;
        RECT 46.755 -132.765 47.085 -132.435 ;
        RECT 46.755 -134.125 47.085 -133.795 ;
        RECT 46.755 -135.485 47.085 -135.155 ;
        RECT 46.755 -136.845 47.085 -136.515 ;
        RECT 46.755 -138.205 47.085 -137.875 ;
        RECT 46.755 -139.565 47.085 -139.235 ;
        RECT 46.755 -140.925 47.085 -140.595 ;
        RECT 46.755 -142.285 47.085 -141.955 ;
        RECT 46.755 -143.645 47.085 -143.315 ;
        RECT 46.755 -145.005 47.085 -144.675 ;
        RECT 46.755 -146.365 47.085 -146.035 ;
        RECT 46.755 -147.725 47.085 -147.395 ;
        RECT 46.755 -149.085 47.085 -148.755 ;
        RECT 46.755 -150.445 47.085 -150.115 ;
        RECT 46.755 -151.805 47.085 -151.475 ;
        RECT 46.755 -153.165 47.085 -152.835 ;
        RECT 46.755 -154.525 47.085 -154.195 ;
        RECT 46.755 -155.885 47.085 -155.555 ;
        RECT 46.755 -157.245 47.085 -156.915 ;
        RECT 46.755 -158.605 47.085 -158.275 ;
        RECT 46.755 -159.965 47.085 -159.635 ;
        RECT 46.755 -161.325 47.085 -160.995 ;
        RECT 46.755 -162.685 47.085 -162.355 ;
        RECT 46.755 -164.045 47.085 -163.715 ;
        RECT 46.755 -165.405 47.085 -165.075 ;
        RECT 46.755 -166.765 47.085 -166.435 ;
        RECT 46.755 -168.125 47.085 -167.795 ;
        RECT 46.755 -169.485 47.085 -169.155 ;
        RECT 46.755 -170.845 47.085 -170.515 ;
        RECT 46.755 -172.205 47.085 -171.875 ;
        RECT 46.755 -173.565 47.085 -173.235 ;
        RECT 46.755 -174.925 47.085 -174.595 ;
        RECT 46.755 -176.285 47.085 -175.955 ;
        RECT 46.755 -177.645 47.085 -177.315 ;
        RECT 46.755 -179.005 47.085 -178.675 ;
        RECT 46.755 -180.365 47.085 -180.035 ;
        RECT 46.755 -181.725 47.085 -181.395 ;
        RECT 46.755 -183.085 47.085 -182.755 ;
        RECT 46.755 -184.445 47.085 -184.115 ;
        RECT 46.755 -185.805 47.085 -185.475 ;
        RECT 46.755 -187.165 47.085 -186.835 ;
        RECT 46.755 -188.525 47.085 -188.195 ;
        RECT 46.755 -189.885 47.085 -189.555 ;
        RECT 46.755 -191.245 47.085 -190.915 ;
        RECT 46.755 -192.605 47.085 -192.275 ;
        RECT 46.755 -193.965 47.085 -193.635 ;
        RECT 46.755 -195.325 47.085 -194.995 ;
        RECT 46.755 -196.685 47.085 -196.355 ;
        RECT 46.755 -198.045 47.085 -197.715 ;
        RECT 46.755 -199.405 47.085 -199.075 ;
        RECT 46.755 -200.765 47.085 -200.435 ;
        RECT 46.755 -202.125 47.085 -201.795 ;
        RECT 46.755 -203.485 47.085 -203.155 ;
        RECT 46.755 -204.845 47.085 -204.515 ;
        RECT 46.755 -206.205 47.085 -205.875 ;
        RECT 46.755 -207.565 47.085 -207.235 ;
        RECT 46.755 -208.925 47.085 -208.595 ;
        RECT 46.755 -210.285 47.085 -209.955 ;
        RECT 46.755 -211.645 47.085 -211.315 ;
        RECT 46.755 -213.005 47.085 -212.675 ;
        RECT 46.755 -214.365 47.085 -214.035 ;
        RECT 46.755 -215.725 47.085 -215.395 ;
        RECT 46.755 -217.085 47.085 -216.755 ;
        RECT 46.755 -218.445 47.085 -218.115 ;
        RECT 46.755 -219.805 47.085 -219.475 ;
        RECT 46.755 -221.165 47.085 -220.835 ;
        RECT 46.755 -222.525 47.085 -222.195 ;
        RECT 46.755 -223.885 47.085 -223.555 ;
        RECT 46.755 -225.245 47.085 -224.915 ;
        RECT 46.755 -226.605 47.085 -226.275 ;
        RECT 46.755 -227.965 47.085 -227.635 ;
        RECT 46.755 -229.325 47.085 -228.995 ;
        RECT 46.755 -230.685 47.085 -230.355 ;
        RECT 46.755 -232.045 47.085 -231.715 ;
        RECT 46.755 -233.405 47.085 -233.075 ;
        RECT 46.755 -234.765 47.085 -234.435 ;
        RECT 46.755 -236.125 47.085 -235.795 ;
        RECT 46.755 -237.485 47.085 -237.155 ;
        RECT 46.755 -238.845 47.085 -238.515 ;
        RECT 46.755 -241.09 47.085 -239.96 ;
        RECT 46.76 -241.205 47.08 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.91 -125.535 47.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 244.04 48.445 245.17 ;
        RECT 48.115 242.595 48.445 242.925 ;
        RECT 48.115 241.235 48.445 241.565 ;
        RECT 48.115 239.875 48.445 240.205 ;
        RECT 48.115 238.515 48.445 238.845 ;
        RECT 48.115 237.155 48.445 237.485 ;
        RECT 48.12 237.155 48.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 -0.845 48.445 -0.515 ;
        RECT 48.115 -2.205 48.445 -1.875 ;
        RECT 48.115 -3.565 48.445 -3.235 ;
        RECT 48.12 -3.565 48.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 244.04 49.805 245.17 ;
        RECT 49.475 242.595 49.805 242.925 ;
        RECT 49.475 241.235 49.805 241.565 ;
        RECT 49.475 239.875 49.805 240.205 ;
        RECT 49.475 238.515 49.805 238.845 ;
        RECT 49.475 237.155 49.805 237.485 ;
        RECT 49.48 237.155 49.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 -0.845 49.805 -0.515 ;
        RECT 49.475 -2.205 49.805 -1.875 ;
        RECT 49.475 -3.565 49.805 -3.235 ;
        RECT 49.48 -3.565 49.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 244.04 51.165 245.17 ;
        RECT 50.835 242.595 51.165 242.925 ;
        RECT 50.835 241.235 51.165 241.565 ;
        RECT 50.835 239.875 51.165 240.205 ;
        RECT 50.835 238.515 51.165 238.845 ;
        RECT 50.835 237.155 51.165 237.485 ;
        RECT 50.84 237.155 51.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 -0.845 51.165 -0.515 ;
        RECT 50.835 -2.205 51.165 -1.875 ;
        RECT 50.835 -3.565 51.165 -3.235 ;
        RECT 50.84 -3.565 51.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 -123.245 51.165 -122.915 ;
        RECT 50.835 -124.605 51.165 -124.275 ;
        RECT 50.835 -125.965 51.165 -125.635 ;
        RECT 50.835 -127.325 51.165 -126.995 ;
        RECT 50.835 -128.685 51.165 -128.355 ;
        RECT 50.835 -130.045 51.165 -129.715 ;
        RECT 50.835 -131.405 51.165 -131.075 ;
        RECT 50.835 -132.765 51.165 -132.435 ;
        RECT 50.835 -134.125 51.165 -133.795 ;
        RECT 50.835 -135.485 51.165 -135.155 ;
        RECT 50.835 -136.845 51.165 -136.515 ;
        RECT 50.835 -138.205 51.165 -137.875 ;
        RECT 50.835 -139.565 51.165 -139.235 ;
        RECT 50.835 -140.925 51.165 -140.595 ;
        RECT 50.835 -142.285 51.165 -141.955 ;
        RECT 50.835 -143.645 51.165 -143.315 ;
        RECT 50.835 -145.005 51.165 -144.675 ;
        RECT 50.835 -146.365 51.165 -146.035 ;
        RECT 50.835 -147.725 51.165 -147.395 ;
        RECT 50.835 -149.085 51.165 -148.755 ;
        RECT 50.835 -150.445 51.165 -150.115 ;
        RECT 50.835 -151.805 51.165 -151.475 ;
        RECT 50.835 -153.165 51.165 -152.835 ;
        RECT 50.835 -154.525 51.165 -154.195 ;
        RECT 50.835 -155.885 51.165 -155.555 ;
        RECT 50.835 -157.245 51.165 -156.915 ;
        RECT 50.835 -158.605 51.165 -158.275 ;
        RECT 50.835 -159.965 51.165 -159.635 ;
        RECT 50.835 -161.325 51.165 -160.995 ;
        RECT 50.835 -162.685 51.165 -162.355 ;
        RECT 50.835 -164.045 51.165 -163.715 ;
        RECT 50.835 -165.405 51.165 -165.075 ;
        RECT 50.835 -166.765 51.165 -166.435 ;
        RECT 50.835 -168.125 51.165 -167.795 ;
        RECT 50.835 -169.485 51.165 -169.155 ;
        RECT 50.835 -170.845 51.165 -170.515 ;
        RECT 50.835 -172.205 51.165 -171.875 ;
        RECT 50.835 -173.565 51.165 -173.235 ;
        RECT 50.835 -174.925 51.165 -174.595 ;
        RECT 50.835 -176.285 51.165 -175.955 ;
        RECT 50.835 -177.645 51.165 -177.315 ;
        RECT 50.835 -179.005 51.165 -178.675 ;
        RECT 50.835 -180.365 51.165 -180.035 ;
        RECT 50.835 -181.725 51.165 -181.395 ;
        RECT 50.835 -183.085 51.165 -182.755 ;
        RECT 50.835 -184.445 51.165 -184.115 ;
        RECT 50.835 -185.805 51.165 -185.475 ;
        RECT 50.835 -187.165 51.165 -186.835 ;
        RECT 50.835 -188.525 51.165 -188.195 ;
        RECT 50.835 -189.885 51.165 -189.555 ;
        RECT 50.835 -191.245 51.165 -190.915 ;
        RECT 50.835 -192.605 51.165 -192.275 ;
        RECT 50.835 -193.965 51.165 -193.635 ;
        RECT 50.835 -195.325 51.165 -194.995 ;
        RECT 50.835 -196.685 51.165 -196.355 ;
        RECT 50.835 -198.045 51.165 -197.715 ;
        RECT 50.835 -199.405 51.165 -199.075 ;
        RECT 50.835 -200.765 51.165 -200.435 ;
        RECT 50.835 -202.125 51.165 -201.795 ;
        RECT 50.835 -203.485 51.165 -203.155 ;
        RECT 50.835 -204.845 51.165 -204.515 ;
        RECT 50.835 -206.205 51.165 -205.875 ;
        RECT 50.835 -207.565 51.165 -207.235 ;
        RECT 50.835 -208.925 51.165 -208.595 ;
        RECT 50.835 -210.285 51.165 -209.955 ;
        RECT 50.835 -211.645 51.165 -211.315 ;
        RECT 50.835 -213.005 51.165 -212.675 ;
        RECT 50.835 -214.365 51.165 -214.035 ;
        RECT 50.835 -215.725 51.165 -215.395 ;
        RECT 50.835 -217.085 51.165 -216.755 ;
        RECT 50.835 -218.445 51.165 -218.115 ;
        RECT 50.835 -219.805 51.165 -219.475 ;
        RECT 50.835 -221.165 51.165 -220.835 ;
        RECT 50.835 -222.525 51.165 -222.195 ;
        RECT 50.835 -223.885 51.165 -223.555 ;
        RECT 50.835 -225.245 51.165 -224.915 ;
        RECT 50.835 -226.605 51.165 -226.275 ;
        RECT 50.835 -227.965 51.165 -227.635 ;
        RECT 50.835 -229.325 51.165 -228.995 ;
        RECT 50.835 -230.685 51.165 -230.355 ;
        RECT 50.835 -232.045 51.165 -231.715 ;
        RECT 50.835 -233.405 51.165 -233.075 ;
        RECT 50.835 -234.765 51.165 -234.435 ;
        RECT 50.835 -236.125 51.165 -235.795 ;
        RECT 50.835 -237.485 51.165 -237.155 ;
        RECT 50.835 -238.845 51.165 -238.515 ;
        RECT 50.835 -241.09 51.165 -239.96 ;
        RECT 50.84 -241.205 51.16 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 244.04 52.525 245.17 ;
        RECT 52.195 242.595 52.525 242.925 ;
        RECT 52.195 241.235 52.525 241.565 ;
        RECT 52.195 239.875 52.525 240.205 ;
        RECT 52.195 238.515 52.525 238.845 ;
        RECT 52.195 237.155 52.525 237.485 ;
        RECT 52.2 237.155 52.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 -0.845 52.525 -0.515 ;
        RECT 52.195 -2.205 52.525 -1.875 ;
        RECT 52.195 -3.565 52.525 -3.235 ;
        RECT 52.2 -3.565 52.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 -123.245 52.525 -122.915 ;
        RECT 52.195 -124.605 52.525 -124.275 ;
        RECT 52.195 -125.965 52.525 -125.635 ;
        RECT 52.195 -127.325 52.525 -126.995 ;
        RECT 52.195 -128.685 52.525 -128.355 ;
        RECT 52.195 -130.045 52.525 -129.715 ;
        RECT 52.195 -131.405 52.525 -131.075 ;
        RECT 52.195 -132.765 52.525 -132.435 ;
        RECT 52.195 -134.125 52.525 -133.795 ;
        RECT 52.195 -135.485 52.525 -135.155 ;
        RECT 52.195 -136.845 52.525 -136.515 ;
        RECT 52.195 -138.205 52.525 -137.875 ;
        RECT 52.195 -139.565 52.525 -139.235 ;
        RECT 52.195 -140.925 52.525 -140.595 ;
        RECT 52.195 -142.285 52.525 -141.955 ;
        RECT 52.195 -143.645 52.525 -143.315 ;
        RECT 52.195 -145.005 52.525 -144.675 ;
        RECT 52.195 -146.365 52.525 -146.035 ;
        RECT 52.195 -147.725 52.525 -147.395 ;
        RECT 52.195 -149.085 52.525 -148.755 ;
        RECT 52.195 -150.445 52.525 -150.115 ;
        RECT 52.195 -151.805 52.525 -151.475 ;
        RECT 52.195 -153.165 52.525 -152.835 ;
        RECT 52.195 -154.525 52.525 -154.195 ;
        RECT 52.195 -155.885 52.525 -155.555 ;
        RECT 52.195 -157.245 52.525 -156.915 ;
        RECT 52.195 -158.605 52.525 -158.275 ;
        RECT 52.195 -159.965 52.525 -159.635 ;
        RECT 52.195 -161.325 52.525 -160.995 ;
        RECT 52.195 -162.685 52.525 -162.355 ;
        RECT 52.195 -164.045 52.525 -163.715 ;
        RECT 52.195 -165.405 52.525 -165.075 ;
        RECT 52.195 -166.765 52.525 -166.435 ;
        RECT 52.195 -168.125 52.525 -167.795 ;
        RECT 52.195 -169.485 52.525 -169.155 ;
        RECT 52.195 -170.845 52.525 -170.515 ;
        RECT 52.195 -172.205 52.525 -171.875 ;
        RECT 52.195 -173.565 52.525 -173.235 ;
        RECT 52.195 -174.925 52.525 -174.595 ;
        RECT 52.195 -176.285 52.525 -175.955 ;
        RECT 52.195 -177.645 52.525 -177.315 ;
        RECT 52.195 -179.005 52.525 -178.675 ;
        RECT 52.195 -180.365 52.525 -180.035 ;
        RECT 52.195 -181.725 52.525 -181.395 ;
        RECT 52.195 -183.085 52.525 -182.755 ;
        RECT 52.195 -184.445 52.525 -184.115 ;
        RECT 52.195 -185.805 52.525 -185.475 ;
        RECT 52.195 -187.165 52.525 -186.835 ;
        RECT 52.195 -188.525 52.525 -188.195 ;
        RECT 52.195 -189.885 52.525 -189.555 ;
        RECT 52.195 -191.245 52.525 -190.915 ;
        RECT 52.195 -192.605 52.525 -192.275 ;
        RECT 52.195 -193.965 52.525 -193.635 ;
        RECT 52.195 -195.325 52.525 -194.995 ;
        RECT 52.195 -196.685 52.525 -196.355 ;
        RECT 52.195 -198.045 52.525 -197.715 ;
        RECT 52.195 -199.405 52.525 -199.075 ;
        RECT 52.195 -200.765 52.525 -200.435 ;
        RECT 52.195 -202.125 52.525 -201.795 ;
        RECT 52.195 -203.485 52.525 -203.155 ;
        RECT 52.195 -204.845 52.525 -204.515 ;
        RECT 52.195 -206.205 52.525 -205.875 ;
        RECT 52.195 -207.565 52.525 -207.235 ;
        RECT 52.195 -208.925 52.525 -208.595 ;
        RECT 52.195 -210.285 52.525 -209.955 ;
        RECT 52.195 -211.645 52.525 -211.315 ;
        RECT 52.195 -213.005 52.525 -212.675 ;
        RECT 52.195 -214.365 52.525 -214.035 ;
        RECT 52.195 -215.725 52.525 -215.395 ;
        RECT 52.195 -217.085 52.525 -216.755 ;
        RECT 52.195 -218.445 52.525 -218.115 ;
        RECT 52.195 -219.805 52.525 -219.475 ;
        RECT 52.195 -221.165 52.525 -220.835 ;
        RECT 52.195 -222.525 52.525 -222.195 ;
        RECT 52.195 -223.885 52.525 -223.555 ;
        RECT 52.195 -225.245 52.525 -224.915 ;
        RECT 52.195 -226.605 52.525 -226.275 ;
        RECT 52.195 -227.965 52.525 -227.635 ;
        RECT 52.195 -229.325 52.525 -228.995 ;
        RECT 52.195 -230.685 52.525 -230.355 ;
        RECT 52.195 -232.045 52.525 -231.715 ;
        RECT 52.195 -233.405 52.525 -233.075 ;
        RECT 52.195 -234.765 52.525 -234.435 ;
        RECT 52.195 -236.125 52.525 -235.795 ;
        RECT 52.195 -237.485 52.525 -237.155 ;
        RECT 52.195 -238.845 52.525 -238.515 ;
        RECT 52.195 -241.09 52.525 -239.96 ;
        RECT 52.2 -241.205 52.52 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 244.04 53.885 245.17 ;
        RECT 53.555 242.595 53.885 242.925 ;
        RECT 53.555 241.235 53.885 241.565 ;
        RECT 53.555 239.875 53.885 240.205 ;
        RECT 53.555 238.515 53.885 238.845 ;
        RECT 53.555 237.155 53.885 237.485 ;
        RECT 53.56 237.155 53.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -0.845 53.885 -0.515 ;
        RECT 53.555 -2.205 53.885 -1.875 ;
        RECT 53.555 -3.565 53.885 -3.235 ;
        RECT 53.56 -3.565 53.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -123.245 53.885 -122.915 ;
        RECT 53.555 -124.605 53.885 -124.275 ;
        RECT 53.555 -125.965 53.885 -125.635 ;
        RECT 53.555 -127.325 53.885 -126.995 ;
        RECT 53.555 -128.685 53.885 -128.355 ;
        RECT 53.555 -130.045 53.885 -129.715 ;
        RECT 53.555 -131.405 53.885 -131.075 ;
        RECT 53.555 -132.765 53.885 -132.435 ;
        RECT 53.555 -134.125 53.885 -133.795 ;
        RECT 53.555 -135.485 53.885 -135.155 ;
        RECT 53.555 -136.845 53.885 -136.515 ;
        RECT 53.555 -138.205 53.885 -137.875 ;
        RECT 53.555 -139.565 53.885 -139.235 ;
        RECT 53.555 -140.925 53.885 -140.595 ;
        RECT 53.555 -142.285 53.885 -141.955 ;
        RECT 53.555 -143.645 53.885 -143.315 ;
        RECT 53.555 -145.005 53.885 -144.675 ;
        RECT 53.555 -146.365 53.885 -146.035 ;
        RECT 53.555 -147.725 53.885 -147.395 ;
        RECT 53.555 -149.085 53.885 -148.755 ;
        RECT 53.555 -150.445 53.885 -150.115 ;
        RECT 53.555 -151.805 53.885 -151.475 ;
        RECT 53.555 -153.165 53.885 -152.835 ;
        RECT 53.555 -154.525 53.885 -154.195 ;
        RECT 53.555 -155.885 53.885 -155.555 ;
        RECT 53.555 -157.245 53.885 -156.915 ;
        RECT 53.555 -158.605 53.885 -158.275 ;
        RECT 53.555 -159.965 53.885 -159.635 ;
        RECT 53.555 -161.325 53.885 -160.995 ;
        RECT 53.555 -162.685 53.885 -162.355 ;
        RECT 53.555 -164.045 53.885 -163.715 ;
        RECT 53.555 -165.405 53.885 -165.075 ;
        RECT 53.555 -166.765 53.885 -166.435 ;
        RECT 53.555 -168.125 53.885 -167.795 ;
        RECT 53.555 -169.485 53.885 -169.155 ;
        RECT 53.555 -170.845 53.885 -170.515 ;
        RECT 53.555 -172.205 53.885 -171.875 ;
        RECT 53.555 -173.565 53.885 -173.235 ;
        RECT 53.555 -174.925 53.885 -174.595 ;
        RECT 53.555 -176.285 53.885 -175.955 ;
        RECT 53.555 -177.645 53.885 -177.315 ;
        RECT 53.555 -179.005 53.885 -178.675 ;
        RECT 53.555 -180.365 53.885 -180.035 ;
        RECT 53.555 -181.725 53.885 -181.395 ;
        RECT 53.555 -183.085 53.885 -182.755 ;
        RECT 53.555 -184.445 53.885 -184.115 ;
        RECT 53.555 -185.805 53.885 -185.475 ;
        RECT 53.555 -187.165 53.885 -186.835 ;
        RECT 53.555 -188.525 53.885 -188.195 ;
        RECT 53.555 -189.885 53.885 -189.555 ;
        RECT 53.555 -191.245 53.885 -190.915 ;
        RECT 53.555 -192.605 53.885 -192.275 ;
        RECT 53.555 -193.965 53.885 -193.635 ;
        RECT 53.555 -195.325 53.885 -194.995 ;
        RECT 53.555 -196.685 53.885 -196.355 ;
        RECT 53.555 -198.045 53.885 -197.715 ;
        RECT 53.555 -199.405 53.885 -199.075 ;
        RECT 53.555 -200.765 53.885 -200.435 ;
        RECT 53.555 -202.125 53.885 -201.795 ;
        RECT 53.555 -203.485 53.885 -203.155 ;
        RECT 53.555 -204.845 53.885 -204.515 ;
        RECT 53.555 -206.205 53.885 -205.875 ;
        RECT 53.555 -207.565 53.885 -207.235 ;
        RECT 53.555 -208.925 53.885 -208.595 ;
        RECT 53.555 -210.285 53.885 -209.955 ;
        RECT 53.555 -211.645 53.885 -211.315 ;
        RECT 53.555 -213.005 53.885 -212.675 ;
        RECT 53.555 -214.365 53.885 -214.035 ;
        RECT 53.555 -215.725 53.885 -215.395 ;
        RECT 53.555 -217.085 53.885 -216.755 ;
        RECT 53.555 -218.445 53.885 -218.115 ;
        RECT 53.555 -219.805 53.885 -219.475 ;
        RECT 53.555 -221.165 53.885 -220.835 ;
        RECT 53.555 -222.525 53.885 -222.195 ;
        RECT 53.555 -223.885 53.885 -223.555 ;
        RECT 53.555 -225.245 53.885 -224.915 ;
        RECT 53.555 -226.605 53.885 -226.275 ;
        RECT 53.555 -227.965 53.885 -227.635 ;
        RECT 53.555 -229.325 53.885 -228.995 ;
        RECT 53.555 -230.685 53.885 -230.355 ;
        RECT 53.555 -232.045 53.885 -231.715 ;
        RECT 53.555 -233.405 53.885 -233.075 ;
        RECT 53.555 -234.765 53.885 -234.435 ;
        RECT 53.555 -236.125 53.885 -235.795 ;
        RECT 53.555 -237.485 53.885 -237.155 ;
        RECT 53.555 -238.845 53.885 -238.515 ;
        RECT 53.555 -241.09 53.885 -239.96 ;
        RECT 53.56 -241.205 53.88 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 244.04 55.245 245.17 ;
        RECT 54.915 242.595 55.245 242.925 ;
        RECT 54.915 241.235 55.245 241.565 ;
        RECT 54.915 239.875 55.245 240.205 ;
        RECT 54.915 238.515 55.245 238.845 ;
        RECT 54.915 237.155 55.245 237.485 ;
        RECT 54.92 237.155 55.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 -0.845 55.245 -0.515 ;
        RECT 54.915 -2.205 55.245 -1.875 ;
        RECT 54.915 -3.565 55.245 -3.235 ;
        RECT 54.92 -3.565 55.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 -123.245 55.245 -122.915 ;
        RECT 54.915 -124.605 55.245 -124.275 ;
        RECT 54.915 -125.965 55.245 -125.635 ;
        RECT 54.915 -127.325 55.245 -126.995 ;
        RECT 54.915 -128.685 55.245 -128.355 ;
        RECT 54.915 -130.045 55.245 -129.715 ;
        RECT 54.915 -131.405 55.245 -131.075 ;
        RECT 54.915 -132.765 55.245 -132.435 ;
        RECT 54.915 -134.125 55.245 -133.795 ;
        RECT 54.915 -135.485 55.245 -135.155 ;
        RECT 54.915 -136.845 55.245 -136.515 ;
        RECT 54.915 -138.205 55.245 -137.875 ;
        RECT 54.915 -139.565 55.245 -139.235 ;
        RECT 54.915 -140.925 55.245 -140.595 ;
        RECT 54.915 -142.285 55.245 -141.955 ;
        RECT 54.915 -143.645 55.245 -143.315 ;
        RECT 54.915 -145.005 55.245 -144.675 ;
        RECT 54.915 -146.365 55.245 -146.035 ;
        RECT 54.915 -147.725 55.245 -147.395 ;
        RECT 54.915 -149.085 55.245 -148.755 ;
        RECT 54.915 -150.445 55.245 -150.115 ;
        RECT 54.915 -151.805 55.245 -151.475 ;
        RECT 54.915 -153.165 55.245 -152.835 ;
        RECT 54.915 -154.525 55.245 -154.195 ;
        RECT 54.915 -155.885 55.245 -155.555 ;
        RECT 54.915 -157.245 55.245 -156.915 ;
        RECT 54.915 -158.605 55.245 -158.275 ;
        RECT 54.915 -159.965 55.245 -159.635 ;
        RECT 54.915 -161.325 55.245 -160.995 ;
        RECT 54.915 -162.685 55.245 -162.355 ;
        RECT 54.915 -164.045 55.245 -163.715 ;
        RECT 54.915 -165.405 55.245 -165.075 ;
        RECT 54.915 -166.765 55.245 -166.435 ;
        RECT 54.915 -168.125 55.245 -167.795 ;
        RECT 54.915 -169.485 55.245 -169.155 ;
        RECT 54.915 -170.845 55.245 -170.515 ;
        RECT 54.915 -172.205 55.245 -171.875 ;
        RECT 54.915 -173.565 55.245 -173.235 ;
        RECT 54.915 -174.925 55.245 -174.595 ;
        RECT 54.915 -176.285 55.245 -175.955 ;
        RECT 54.915 -177.645 55.245 -177.315 ;
        RECT 54.915 -179.005 55.245 -178.675 ;
        RECT 54.915 -180.365 55.245 -180.035 ;
        RECT 54.915 -181.725 55.245 -181.395 ;
        RECT 54.915 -183.085 55.245 -182.755 ;
        RECT 54.915 -184.445 55.245 -184.115 ;
        RECT 54.915 -185.805 55.245 -185.475 ;
        RECT 54.915 -187.165 55.245 -186.835 ;
        RECT 54.915 -188.525 55.245 -188.195 ;
        RECT 54.915 -189.885 55.245 -189.555 ;
        RECT 54.915 -191.245 55.245 -190.915 ;
        RECT 54.915 -192.605 55.245 -192.275 ;
        RECT 54.915 -193.965 55.245 -193.635 ;
        RECT 54.915 -195.325 55.245 -194.995 ;
        RECT 54.915 -196.685 55.245 -196.355 ;
        RECT 54.915 -198.045 55.245 -197.715 ;
        RECT 54.915 -199.405 55.245 -199.075 ;
        RECT 54.915 -200.765 55.245 -200.435 ;
        RECT 54.915 -202.125 55.245 -201.795 ;
        RECT 54.915 -203.485 55.245 -203.155 ;
        RECT 54.915 -204.845 55.245 -204.515 ;
        RECT 54.915 -206.205 55.245 -205.875 ;
        RECT 54.915 -207.565 55.245 -207.235 ;
        RECT 54.915 -208.925 55.245 -208.595 ;
        RECT 54.915 -210.285 55.245 -209.955 ;
        RECT 54.915 -211.645 55.245 -211.315 ;
        RECT 54.915 -213.005 55.245 -212.675 ;
        RECT 54.915 -214.365 55.245 -214.035 ;
        RECT 54.915 -215.725 55.245 -215.395 ;
        RECT 54.915 -217.085 55.245 -216.755 ;
        RECT 54.915 -218.445 55.245 -218.115 ;
        RECT 54.915 -219.805 55.245 -219.475 ;
        RECT 54.915 -221.165 55.245 -220.835 ;
        RECT 54.915 -222.525 55.245 -222.195 ;
        RECT 54.915 -223.885 55.245 -223.555 ;
        RECT 54.915 -225.245 55.245 -224.915 ;
        RECT 54.915 -226.605 55.245 -226.275 ;
        RECT 54.915 -227.965 55.245 -227.635 ;
        RECT 54.915 -229.325 55.245 -228.995 ;
        RECT 54.915 -230.685 55.245 -230.355 ;
        RECT 54.915 -232.045 55.245 -231.715 ;
        RECT 54.915 -233.405 55.245 -233.075 ;
        RECT 54.915 -234.765 55.245 -234.435 ;
        RECT 54.915 -236.125 55.245 -235.795 ;
        RECT 54.915 -237.485 55.245 -237.155 ;
        RECT 54.915 -238.845 55.245 -238.515 ;
        RECT 54.915 -241.09 55.245 -239.96 ;
        RECT 54.92 -241.205 55.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 244.04 56.605 245.17 ;
        RECT 56.275 242.595 56.605 242.925 ;
        RECT 56.275 241.235 56.605 241.565 ;
        RECT 56.275 239.875 56.605 240.205 ;
        RECT 56.275 238.515 56.605 238.845 ;
        RECT 56.275 237.155 56.605 237.485 ;
        RECT 56.28 237.155 56.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -0.845 56.605 -0.515 ;
        RECT 56.275 -2.205 56.605 -1.875 ;
        RECT 56.275 -3.565 56.605 -3.235 ;
        RECT 56.28 -3.565 56.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -147.725 56.605 -147.395 ;
        RECT 56.275 -149.085 56.605 -148.755 ;
        RECT 56.275 -150.445 56.605 -150.115 ;
        RECT 56.275 -151.805 56.605 -151.475 ;
        RECT 56.275 -153.165 56.605 -152.835 ;
        RECT 56.275 -154.525 56.605 -154.195 ;
        RECT 56.275 -155.885 56.605 -155.555 ;
        RECT 56.275 -157.245 56.605 -156.915 ;
        RECT 56.275 -158.605 56.605 -158.275 ;
        RECT 56.275 -159.965 56.605 -159.635 ;
        RECT 56.275 -161.325 56.605 -160.995 ;
        RECT 56.275 -162.685 56.605 -162.355 ;
        RECT 56.275 -164.045 56.605 -163.715 ;
        RECT 56.275 -165.405 56.605 -165.075 ;
        RECT 56.275 -166.765 56.605 -166.435 ;
        RECT 56.275 -168.125 56.605 -167.795 ;
        RECT 56.275 -169.485 56.605 -169.155 ;
        RECT 56.275 -170.845 56.605 -170.515 ;
        RECT 56.275 -172.205 56.605 -171.875 ;
        RECT 56.275 -173.565 56.605 -173.235 ;
        RECT 56.275 -174.925 56.605 -174.595 ;
        RECT 56.275 -176.285 56.605 -175.955 ;
        RECT 56.275 -177.645 56.605 -177.315 ;
        RECT 56.275 -179.005 56.605 -178.675 ;
        RECT 56.275 -180.365 56.605 -180.035 ;
        RECT 56.275 -181.725 56.605 -181.395 ;
        RECT 56.275 -183.085 56.605 -182.755 ;
        RECT 56.275 -184.445 56.605 -184.115 ;
        RECT 56.275 -185.805 56.605 -185.475 ;
        RECT 56.275 -187.165 56.605 -186.835 ;
        RECT 56.275 -188.525 56.605 -188.195 ;
        RECT 56.275 -189.885 56.605 -189.555 ;
        RECT 56.275 -191.245 56.605 -190.915 ;
        RECT 56.275 -192.605 56.605 -192.275 ;
        RECT 56.275 -193.965 56.605 -193.635 ;
        RECT 56.275 -195.325 56.605 -194.995 ;
        RECT 56.275 -196.685 56.605 -196.355 ;
        RECT 56.275 -198.045 56.605 -197.715 ;
        RECT 56.275 -199.405 56.605 -199.075 ;
        RECT 56.275 -200.765 56.605 -200.435 ;
        RECT 56.275 -202.125 56.605 -201.795 ;
        RECT 56.275 -203.485 56.605 -203.155 ;
        RECT 56.275 -204.845 56.605 -204.515 ;
        RECT 56.275 -206.205 56.605 -205.875 ;
        RECT 56.275 -207.565 56.605 -207.235 ;
        RECT 56.275 -208.925 56.605 -208.595 ;
        RECT 56.275 -210.285 56.605 -209.955 ;
        RECT 56.275 -211.645 56.605 -211.315 ;
        RECT 56.275 -213.005 56.605 -212.675 ;
        RECT 56.275 -214.365 56.605 -214.035 ;
        RECT 56.275 -215.725 56.605 -215.395 ;
        RECT 56.275 -217.085 56.605 -216.755 ;
        RECT 56.275 -218.445 56.605 -218.115 ;
        RECT 56.275 -219.805 56.605 -219.475 ;
        RECT 56.275 -221.165 56.605 -220.835 ;
        RECT 56.275 -222.525 56.605 -222.195 ;
        RECT 56.275 -223.885 56.605 -223.555 ;
        RECT 56.275 -225.245 56.605 -224.915 ;
        RECT 56.275 -226.605 56.605 -226.275 ;
        RECT 56.275 -227.965 56.605 -227.635 ;
        RECT 56.275 -229.325 56.605 -228.995 ;
        RECT 56.275 -230.685 56.605 -230.355 ;
        RECT 56.275 -232.045 56.605 -231.715 ;
        RECT 56.275 -233.405 56.605 -233.075 ;
        RECT 56.275 -234.765 56.605 -234.435 ;
        RECT 56.275 -236.125 56.605 -235.795 ;
        RECT 56.275 -237.485 56.605 -237.155 ;
        RECT 56.275 -238.845 56.605 -238.515 ;
        RECT 56.275 -241.09 56.605 -239.96 ;
        RECT 56.28 -241.205 56.6 -122.24 ;
        RECT 56.275 -123.245 56.605 -122.915 ;
        RECT 56.275 -124.605 56.605 -124.275 ;
        RECT 56.275 -125.965 56.605 -125.635 ;
        RECT 56.275 -127.325 56.605 -126.995 ;
        RECT 56.275 -128.685 56.605 -128.355 ;
        RECT 56.275 -130.045 56.605 -129.715 ;
        RECT 56.275 -131.405 56.605 -131.075 ;
        RECT 56.275 -132.765 56.605 -132.435 ;
        RECT 56.275 -134.125 56.605 -133.795 ;
        RECT 56.275 -135.485 56.605 -135.155 ;
        RECT 56.275 -136.845 56.605 -136.515 ;
        RECT 56.275 -138.205 56.605 -137.875 ;
        RECT 56.275 -139.565 56.605 -139.235 ;
        RECT 56.275 -140.925 56.605 -140.595 ;
        RECT 56.275 -142.285 56.605 -141.955 ;
        RECT 56.275 -143.645 56.605 -143.315 ;
        RECT 56.275 -145.005 56.605 -144.675 ;
        RECT 56.275 -146.365 56.605 -146.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 -123.245 22.605 -122.915 ;
        RECT 22.275 -124.605 22.605 -124.275 ;
        RECT 22.275 -125.965 22.605 -125.635 ;
        RECT 22.275 -127.325 22.605 -126.995 ;
        RECT 22.275 -128.685 22.605 -128.355 ;
        RECT 22.275 -130.045 22.605 -129.715 ;
        RECT 22.275 -131.405 22.605 -131.075 ;
        RECT 22.275 -132.765 22.605 -132.435 ;
        RECT 22.275 -134.125 22.605 -133.795 ;
        RECT 22.275 -135.485 22.605 -135.155 ;
        RECT 22.275 -136.845 22.605 -136.515 ;
        RECT 22.275 -138.205 22.605 -137.875 ;
        RECT 22.275 -139.565 22.605 -139.235 ;
        RECT 22.275 -140.925 22.605 -140.595 ;
        RECT 22.275 -142.285 22.605 -141.955 ;
        RECT 22.275 -143.645 22.605 -143.315 ;
        RECT 22.275 -145.005 22.605 -144.675 ;
        RECT 22.275 -146.365 22.605 -146.035 ;
        RECT 22.275 -147.725 22.605 -147.395 ;
        RECT 22.275 -149.085 22.605 -148.755 ;
        RECT 22.275 -150.445 22.605 -150.115 ;
        RECT 22.275 -151.805 22.605 -151.475 ;
        RECT 22.275 -153.165 22.605 -152.835 ;
        RECT 22.275 -154.525 22.605 -154.195 ;
        RECT 22.275 -155.885 22.605 -155.555 ;
        RECT 22.275 -157.245 22.605 -156.915 ;
        RECT 22.275 -158.605 22.605 -158.275 ;
        RECT 22.275 -159.965 22.605 -159.635 ;
        RECT 22.275 -161.325 22.605 -160.995 ;
        RECT 22.275 -162.685 22.605 -162.355 ;
        RECT 22.275 -164.045 22.605 -163.715 ;
        RECT 22.275 -165.405 22.605 -165.075 ;
        RECT 22.275 -166.765 22.605 -166.435 ;
        RECT 22.275 -168.125 22.605 -167.795 ;
        RECT 22.275 -169.485 22.605 -169.155 ;
        RECT 22.275 -170.845 22.605 -170.515 ;
        RECT 22.275 -172.205 22.605 -171.875 ;
        RECT 22.275 -173.565 22.605 -173.235 ;
        RECT 22.275 -174.925 22.605 -174.595 ;
        RECT 22.275 -176.285 22.605 -175.955 ;
        RECT 22.275 -177.645 22.605 -177.315 ;
        RECT 22.275 -179.005 22.605 -178.675 ;
        RECT 22.275 -180.365 22.605 -180.035 ;
        RECT 22.275 -181.725 22.605 -181.395 ;
        RECT 22.275 -183.085 22.605 -182.755 ;
        RECT 22.275 -184.445 22.605 -184.115 ;
        RECT 22.275 -185.805 22.605 -185.475 ;
        RECT 22.275 -187.165 22.605 -186.835 ;
        RECT 22.275 -188.525 22.605 -188.195 ;
        RECT 22.275 -189.885 22.605 -189.555 ;
        RECT 22.275 -191.245 22.605 -190.915 ;
        RECT 22.275 -192.605 22.605 -192.275 ;
        RECT 22.275 -193.965 22.605 -193.635 ;
        RECT 22.275 -195.325 22.605 -194.995 ;
        RECT 22.275 -196.685 22.605 -196.355 ;
        RECT 22.275 -198.045 22.605 -197.715 ;
        RECT 22.275 -199.405 22.605 -199.075 ;
        RECT 22.275 -200.765 22.605 -200.435 ;
        RECT 22.275 -202.125 22.605 -201.795 ;
        RECT 22.275 -203.485 22.605 -203.155 ;
        RECT 22.275 -204.845 22.605 -204.515 ;
        RECT 22.275 -206.205 22.605 -205.875 ;
        RECT 22.275 -207.565 22.605 -207.235 ;
        RECT 22.275 -208.925 22.605 -208.595 ;
        RECT 22.275 -210.285 22.605 -209.955 ;
        RECT 22.275 -211.645 22.605 -211.315 ;
        RECT 22.275 -213.005 22.605 -212.675 ;
        RECT 22.275 -214.365 22.605 -214.035 ;
        RECT 22.275 -215.725 22.605 -215.395 ;
        RECT 22.275 -217.085 22.605 -216.755 ;
        RECT 22.275 -218.445 22.605 -218.115 ;
        RECT 22.275 -219.805 22.605 -219.475 ;
        RECT 22.275 -221.165 22.605 -220.835 ;
        RECT 22.275 -222.525 22.605 -222.195 ;
        RECT 22.275 -223.885 22.605 -223.555 ;
        RECT 22.275 -225.245 22.605 -224.915 ;
        RECT 22.275 -226.605 22.605 -226.275 ;
        RECT 22.275 -227.965 22.605 -227.635 ;
        RECT 22.275 -229.325 22.605 -228.995 ;
        RECT 22.275 -230.685 22.605 -230.355 ;
        RECT 22.275 -232.045 22.605 -231.715 ;
        RECT 22.275 -233.405 22.605 -233.075 ;
        RECT 22.275 -234.765 22.605 -234.435 ;
        RECT 22.275 -236.125 22.605 -235.795 ;
        RECT 22.275 -237.485 22.605 -237.155 ;
        RECT 22.275 -238.845 22.605 -238.515 ;
        RECT 22.275 -241.09 22.605 -239.96 ;
        RECT 22.28 -241.205 22.6 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 244.04 23.965 245.17 ;
        RECT 23.635 242.595 23.965 242.925 ;
        RECT 23.635 241.235 23.965 241.565 ;
        RECT 23.635 239.875 23.965 240.205 ;
        RECT 23.635 238.515 23.965 238.845 ;
        RECT 23.635 237.155 23.965 237.485 ;
        RECT 23.64 237.155 23.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 -0.845 23.965 -0.515 ;
        RECT 23.635 -2.205 23.965 -1.875 ;
        RECT 23.635 -3.565 23.965 -3.235 ;
        RECT 23.64 -3.565 23.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 -123.245 23.965 -122.915 ;
        RECT 23.635 -124.605 23.965 -124.275 ;
        RECT 23.635 -125.965 23.965 -125.635 ;
        RECT 23.635 -127.325 23.965 -126.995 ;
        RECT 23.635 -128.685 23.965 -128.355 ;
        RECT 23.635 -130.045 23.965 -129.715 ;
        RECT 23.635 -131.405 23.965 -131.075 ;
        RECT 23.635 -132.765 23.965 -132.435 ;
        RECT 23.635 -134.125 23.965 -133.795 ;
        RECT 23.635 -135.485 23.965 -135.155 ;
        RECT 23.635 -136.845 23.965 -136.515 ;
        RECT 23.635 -138.205 23.965 -137.875 ;
        RECT 23.635 -139.565 23.965 -139.235 ;
        RECT 23.635 -140.925 23.965 -140.595 ;
        RECT 23.635 -142.285 23.965 -141.955 ;
        RECT 23.635 -143.645 23.965 -143.315 ;
        RECT 23.635 -145.005 23.965 -144.675 ;
        RECT 23.635 -146.365 23.965 -146.035 ;
        RECT 23.635 -147.725 23.965 -147.395 ;
        RECT 23.635 -149.085 23.965 -148.755 ;
        RECT 23.635 -150.445 23.965 -150.115 ;
        RECT 23.635 -151.805 23.965 -151.475 ;
        RECT 23.635 -153.165 23.965 -152.835 ;
        RECT 23.635 -154.525 23.965 -154.195 ;
        RECT 23.635 -155.885 23.965 -155.555 ;
        RECT 23.635 -157.245 23.965 -156.915 ;
        RECT 23.635 -158.605 23.965 -158.275 ;
        RECT 23.635 -159.965 23.965 -159.635 ;
        RECT 23.635 -161.325 23.965 -160.995 ;
        RECT 23.635 -162.685 23.965 -162.355 ;
        RECT 23.635 -164.045 23.965 -163.715 ;
        RECT 23.635 -165.405 23.965 -165.075 ;
        RECT 23.635 -166.765 23.965 -166.435 ;
        RECT 23.635 -168.125 23.965 -167.795 ;
        RECT 23.635 -169.485 23.965 -169.155 ;
        RECT 23.635 -170.845 23.965 -170.515 ;
        RECT 23.635 -172.205 23.965 -171.875 ;
        RECT 23.635 -173.565 23.965 -173.235 ;
        RECT 23.635 -174.925 23.965 -174.595 ;
        RECT 23.635 -176.285 23.965 -175.955 ;
        RECT 23.635 -177.645 23.965 -177.315 ;
        RECT 23.635 -179.005 23.965 -178.675 ;
        RECT 23.635 -180.365 23.965 -180.035 ;
        RECT 23.635 -181.725 23.965 -181.395 ;
        RECT 23.635 -183.085 23.965 -182.755 ;
        RECT 23.635 -184.445 23.965 -184.115 ;
        RECT 23.635 -185.805 23.965 -185.475 ;
        RECT 23.635 -187.165 23.965 -186.835 ;
        RECT 23.635 -188.525 23.965 -188.195 ;
        RECT 23.635 -189.885 23.965 -189.555 ;
        RECT 23.635 -191.245 23.965 -190.915 ;
        RECT 23.635 -192.605 23.965 -192.275 ;
        RECT 23.635 -193.965 23.965 -193.635 ;
        RECT 23.635 -195.325 23.965 -194.995 ;
        RECT 23.635 -196.685 23.965 -196.355 ;
        RECT 23.635 -198.045 23.965 -197.715 ;
        RECT 23.635 -199.405 23.965 -199.075 ;
        RECT 23.635 -200.765 23.965 -200.435 ;
        RECT 23.635 -202.125 23.965 -201.795 ;
        RECT 23.635 -203.485 23.965 -203.155 ;
        RECT 23.635 -204.845 23.965 -204.515 ;
        RECT 23.635 -206.205 23.965 -205.875 ;
        RECT 23.635 -207.565 23.965 -207.235 ;
        RECT 23.635 -208.925 23.965 -208.595 ;
        RECT 23.635 -210.285 23.965 -209.955 ;
        RECT 23.635 -211.645 23.965 -211.315 ;
        RECT 23.635 -213.005 23.965 -212.675 ;
        RECT 23.635 -214.365 23.965 -214.035 ;
        RECT 23.635 -215.725 23.965 -215.395 ;
        RECT 23.635 -217.085 23.965 -216.755 ;
        RECT 23.635 -218.445 23.965 -218.115 ;
        RECT 23.635 -219.805 23.965 -219.475 ;
        RECT 23.635 -221.165 23.965 -220.835 ;
        RECT 23.635 -222.525 23.965 -222.195 ;
        RECT 23.635 -223.885 23.965 -223.555 ;
        RECT 23.635 -225.245 23.965 -224.915 ;
        RECT 23.635 -226.605 23.965 -226.275 ;
        RECT 23.635 -227.965 23.965 -227.635 ;
        RECT 23.635 -229.325 23.965 -228.995 ;
        RECT 23.635 -230.685 23.965 -230.355 ;
        RECT 23.635 -232.045 23.965 -231.715 ;
        RECT 23.635 -233.405 23.965 -233.075 ;
        RECT 23.635 -234.765 23.965 -234.435 ;
        RECT 23.635 -236.125 23.965 -235.795 ;
        RECT 23.635 -237.485 23.965 -237.155 ;
        RECT 23.635 -238.845 23.965 -238.515 ;
        RECT 23.635 -241.09 23.965 -239.96 ;
        RECT 23.64 -241.205 23.96 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 244.04 25.325 245.17 ;
        RECT 24.995 242.595 25.325 242.925 ;
        RECT 24.995 241.235 25.325 241.565 ;
        RECT 24.995 239.875 25.325 240.205 ;
        RECT 24.995 238.515 25.325 238.845 ;
        RECT 24.995 237.155 25.325 237.485 ;
        RECT 25 237.155 25.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -127.325 25.325 -126.995 ;
        RECT 24.995 -128.685 25.325 -128.355 ;
        RECT 24.995 -130.045 25.325 -129.715 ;
        RECT 24.995 -131.405 25.325 -131.075 ;
        RECT 24.995 -132.765 25.325 -132.435 ;
        RECT 24.995 -134.125 25.325 -133.795 ;
        RECT 24.995 -135.485 25.325 -135.155 ;
        RECT 24.995 -136.845 25.325 -136.515 ;
        RECT 24.995 -138.205 25.325 -137.875 ;
        RECT 24.995 -139.565 25.325 -139.235 ;
        RECT 24.995 -140.925 25.325 -140.595 ;
        RECT 24.995 -142.285 25.325 -141.955 ;
        RECT 24.995 -143.645 25.325 -143.315 ;
        RECT 24.995 -145.005 25.325 -144.675 ;
        RECT 24.995 -146.365 25.325 -146.035 ;
        RECT 24.995 -147.725 25.325 -147.395 ;
        RECT 24.995 -149.085 25.325 -148.755 ;
        RECT 24.995 -150.445 25.325 -150.115 ;
        RECT 24.995 -151.805 25.325 -151.475 ;
        RECT 24.995 -153.165 25.325 -152.835 ;
        RECT 24.995 -154.525 25.325 -154.195 ;
        RECT 24.995 -155.885 25.325 -155.555 ;
        RECT 24.995 -157.245 25.325 -156.915 ;
        RECT 24.995 -158.605 25.325 -158.275 ;
        RECT 24.995 -159.965 25.325 -159.635 ;
        RECT 24.995 -161.325 25.325 -160.995 ;
        RECT 24.995 -162.685 25.325 -162.355 ;
        RECT 24.995 -164.045 25.325 -163.715 ;
        RECT 24.995 -165.405 25.325 -165.075 ;
        RECT 24.995 -166.765 25.325 -166.435 ;
        RECT 24.995 -168.125 25.325 -167.795 ;
        RECT 24.995 -169.485 25.325 -169.155 ;
        RECT 24.995 -170.845 25.325 -170.515 ;
        RECT 24.995 -172.205 25.325 -171.875 ;
        RECT 24.995 -173.565 25.325 -173.235 ;
        RECT 24.995 -174.925 25.325 -174.595 ;
        RECT 24.995 -176.285 25.325 -175.955 ;
        RECT 24.995 -177.645 25.325 -177.315 ;
        RECT 24.995 -179.005 25.325 -178.675 ;
        RECT 24.995 -180.365 25.325 -180.035 ;
        RECT 24.995 -181.725 25.325 -181.395 ;
        RECT 24.995 -183.085 25.325 -182.755 ;
        RECT 24.995 -184.445 25.325 -184.115 ;
        RECT 24.995 -185.805 25.325 -185.475 ;
        RECT 24.995 -187.165 25.325 -186.835 ;
        RECT 24.995 -188.525 25.325 -188.195 ;
        RECT 24.995 -189.885 25.325 -189.555 ;
        RECT 24.995 -191.245 25.325 -190.915 ;
        RECT 24.995 -192.605 25.325 -192.275 ;
        RECT 24.995 -193.965 25.325 -193.635 ;
        RECT 24.995 -195.325 25.325 -194.995 ;
        RECT 24.995 -196.685 25.325 -196.355 ;
        RECT 24.995 -198.045 25.325 -197.715 ;
        RECT 24.995 -199.405 25.325 -199.075 ;
        RECT 24.995 -200.765 25.325 -200.435 ;
        RECT 24.995 -202.125 25.325 -201.795 ;
        RECT 24.995 -203.485 25.325 -203.155 ;
        RECT 24.995 -204.845 25.325 -204.515 ;
        RECT 24.995 -206.205 25.325 -205.875 ;
        RECT 24.995 -207.565 25.325 -207.235 ;
        RECT 24.995 -208.925 25.325 -208.595 ;
        RECT 24.995 -210.285 25.325 -209.955 ;
        RECT 24.995 -211.645 25.325 -211.315 ;
        RECT 24.995 -213.005 25.325 -212.675 ;
        RECT 24.995 -214.365 25.325 -214.035 ;
        RECT 24.995 -215.725 25.325 -215.395 ;
        RECT 24.995 -217.085 25.325 -216.755 ;
        RECT 24.995 -218.445 25.325 -218.115 ;
        RECT 24.995 -219.805 25.325 -219.475 ;
        RECT 24.995 -221.165 25.325 -220.835 ;
        RECT 24.995 -222.525 25.325 -222.195 ;
        RECT 24.995 -223.885 25.325 -223.555 ;
        RECT 24.995 -225.245 25.325 -224.915 ;
        RECT 24.995 -226.605 25.325 -226.275 ;
        RECT 24.995 -227.965 25.325 -227.635 ;
        RECT 24.995 -229.325 25.325 -228.995 ;
        RECT 24.995 -230.685 25.325 -230.355 ;
        RECT 24.995 -232.045 25.325 -231.715 ;
        RECT 24.995 -233.405 25.325 -233.075 ;
        RECT 24.995 -234.765 25.325 -234.435 ;
        RECT 24.995 -236.125 25.325 -235.795 ;
        RECT 24.995 -237.485 25.325 -237.155 ;
        RECT 24.995 -238.845 25.325 -238.515 ;
        RECT 24.995 -241.09 25.325 -239.96 ;
        RECT 25 -241.205 25.32 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.11 -125.535 25.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 244.04 26.685 245.17 ;
        RECT 26.355 242.595 26.685 242.925 ;
        RECT 26.355 241.235 26.685 241.565 ;
        RECT 26.355 239.875 26.685 240.205 ;
        RECT 26.355 238.515 26.685 238.845 ;
        RECT 26.355 237.155 26.685 237.485 ;
        RECT 26.36 237.155 26.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -0.845 26.685 -0.515 ;
        RECT 26.355 -2.205 26.685 -1.875 ;
        RECT 26.355 -3.565 26.685 -3.235 ;
        RECT 26.36 -3.565 26.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 244.04 28.045 245.17 ;
        RECT 27.715 242.595 28.045 242.925 ;
        RECT 27.715 241.235 28.045 241.565 ;
        RECT 27.715 239.875 28.045 240.205 ;
        RECT 27.715 238.515 28.045 238.845 ;
        RECT 27.715 237.155 28.045 237.485 ;
        RECT 27.72 237.155 28.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 -0.845 28.045 -0.515 ;
        RECT 27.715 -2.205 28.045 -1.875 ;
        RECT 27.715 -3.565 28.045 -3.235 ;
        RECT 27.72 -3.565 28.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 244.04 29.405 245.17 ;
        RECT 29.075 242.595 29.405 242.925 ;
        RECT 29.075 241.235 29.405 241.565 ;
        RECT 29.075 239.875 29.405 240.205 ;
        RECT 29.075 238.515 29.405 238.845 ;
        RECT 29.075 237.155 29.405 237.485 ;
        RECT 29.08 237.155 29.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -0.845 29.405 -0.515 ;
        RECT 29.075 -2.205 29.405 -1.875 ;
        RECT 29.075 -3.565 29.405 -3.235 ;
        RECT 29.08 -3.565 29.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -123.245 29.405 -122.915 ;
        RECT 29.075 -124.605 29.405 -124.275 ;
        RECT 29.075 -125.965 29.405 -125.635 ;
        RECT 29.075 -127.325 29.405 -126.995 ;
        RECT 29.075 -128.685 29.405 -128.355 ;
        RECT 29.075 -130.045 29.405 -129.715 ;
        RECT 29.075 -131.405 29.405 -131.075 ;
        RECT 29.075 -132.765 29.405 -132.435 ;
        RECT 29.075 -134.125 29.405 -133.795 ;
        RECT 29.075 -135.485 29.405 -135.155 ;
        RECT 29.075 -136.845 29.405 -136.515 ;
        RECT 29.075 -138.205 29.405 -137.875 ;
        RECT 29.075 -139.565 29.405 -139.235 ;
        RECT 29.075 -140.925 29.405 -140.595 ;
        RECT 29.075 -142.285 29.405 -141.955 ;
        RECT 29.075 -143.645 29.405 -143.315 ;
        RECT 29.075 -145.005 29.405 -144.675 ;
        RECT 29.075 -146.365 29.405 -146.035 ;
        RECT 29.075 -147.725 29.405 -147.395 ;
        RECT 29.075 -149.085 29.405 -148.755 ;
        RECT 29.075 -150.445 29.405 -150.115 ;
        RECT 29.075 -151.805 29.405 -151.475 ;
        RECT 29.075 -153.165 29.405 -152.835 ;
        RECT 29.075 -154.525 29.405 -154.195 ;
        RECT 29.075 -155.885 29.405 -155.555 ;
        RECT 29.075 -157.245 29.405 -156.915 ;
        RECT 29.075 -158.605 29.405 -158.275 ;
        RECT 29.075 -159.965 29.405 -159.635 ;
        RECT 29.075 -161.325 29.405 -160.995 ;
        RECT 29.075 -162.685 29.405 -162.355 ;
        RECT 29.075 -164.045 29.405 -163.715 ;
        RECT 29.075 -165.405 29.405 -165.075 ;
        RECT 29.075 -166.765 29.405 -166.435 ;
        RECT 29.075 -168.125 29.405 -167.795 ;
        RECT 29.075 -169.485 29.405 -169.155 ;
        RECT 29.075 -170.845 29.405 -170.515 ;
        RECT 29.075 -172.205 29.405 -171.875 ;
        RECT 29.075 -173.565 29.405 -173.235 ;
        RECT 29.075 -174.925 29.405 -174.595 ;
        RECT 29.075 -176.285 29.405 -175.955 ;
        RECT 29.075 -177.645 29.405 -177.315 ;
        RECT 29.075 -179.005 29.405 -178.675 ;
        RECT 29.075 -180.365 29.405 -180.035 ;
        RECT 29.075 -181.725 29.405 -181.395 ;
        RECT 29.075 -183.085 29.405 -182.755 ;
        RECT 29.075 -184.445 29.405 -184.115 ;
        RECT 29.075 -185.805 29.405 -185.475 ;
        RECT 29.075 -187.165 29.405 -186.835 ;
        RECT 29.075 -188.525 29.405 -188.195 ;
        RECT 29.075 -189.885 29.405 -189.555 ;
        RECT 29.075 -191.245 29.405 -190.915 ;
        RECT 29.075 -192.605 29.405 -192.275 ;
        RECT 29.075 -193.965 29.405 -193.635 ;
        RECT 29.075 -195.325 29.405 -194.995 ;
        RECT 29.075 -196.685 29.405 -196.355 ;
        RECT 29.075 -198.045 29.405 -197.715 ;
        RECT 29.075 -199.405 29.405 -199.075 ;
        RECT 29.075 -200.765 29.405 -200.435 ;
        RECT 29.075 -202.125 29.405 -201.795 ;
        RECT 29.075 -203.485 29.405 -203.155 ;
        RECT 29.075 -204.845 29.405 -204.515 ;
        RECT 29.075 -206.205 29.405 -205.875 ;
        RECT 29.075 -207.565 29.405 -207.235 ;
        RECT 29.075 -208.925 29.405 -208.595 ;
        RECT 29.075 -210.285 29.405 -209.955 ;
        RECT 29.075 -211.645 29.405 -211.315 ;
        RECT 29.075 -213.005 29.405 -212.675 ;
        RECT 29.075 -214.365 29.405 -214.035 ;
        RECT 29.075 -215.725 29.405 -215.395 ;
        RECT 29.075 -217.085 29.405 -216.755 ;
        RECT 29.075 -218.445 29.405 -218.115 ;
        RECT 29.075 -219.805 29.405 -219.475 ;
        RECT 29.075 -221.165 29.405 -220.835 ;
        RECT 29.075 -222.525 29.405 -222.195 ;
        RECT 29.075 -223.885 29.405 -223.555 ;
        RECT 29.075 -225.245 29.405 -224.915 ;
        RECT 29.075 -226.605 29.405 -226.275 ;
        RECT 29.075 -227.965 29.405 -227.635 ;
        RECT 29.075 -229.325 29.405 -228.995 ;
        RECT 29.075 -230.685 29.405 -230.355 ;
        RECT 29.075 -232.045 29.405 -231.715 ;
        RECT 29.075 -233.405 29.405 -233.075 ;
        RECT 29.075 -234.765 29.405 -234.435 ;
        RECT 29.075 -236.125 29.405 -235.795 ;
        RECT 29.075 -237.485 29.405 -237.155 ;
        RECT 29.075 -238.845 29.405 -238.515 ;
        RECT 29.075 -241.09 29.405 -239.96 ;
        RECT 29.08 -241.205 29.4 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 244.04 30.765 245.17 ;
        RECT 30.435 242.595 30.765 242.925 ;
        RECT 30.435 241.235 30.765 241.565 ;
        RECT 30.435 239.875 30.765 240.205 ;
        RECT 30.435 238.515 30.765 238.845 ;
        RECT 30.435 237.155 30.765 237.485 ;
        RECT 30.44 237.155 30.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -0.845 30.765 -0.515 ;
        RECT 30.435 -2.205 30.765 -1.875 ;
        RECT 30.435 -3.565 30.765 -3.235 ;
        RECT 30.44 -3.565 30.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -123.245 30.765 -122.915 ;
        RECT 30.435 -124.605 30.765 -124.275 ;
        RECT 30.435 -125.965 30.765 -125.635 ;
        RECT 30.435 -127.325 30.765 -126.995 ;
        RECT 30.435 -128.685 30.765 -128.355 ;
        RECT 30.435 -130.045 30.765 -129.715 ;
        RECT 30.435 -131.405 30.765 -131.075 ;
        RECT 30.435 -132.765 30.765 -132.435 ;
        RECT 30.435 -134.125 30.765 -133.795 ;
        RECT 30.435 -135.485 30.765 -135.155 ;
        RECT 30.435 -136.845 30.765 -136.515 ;
        RECT 30.435 -138.205 30.765 -137.875 ;
        RECT 30.435 -139.565 30.765 -139.235 ;
        RECT 30.435 -140.925 30.765 -140.595 ;
        RECT 30.435 -142.285 30.765 -141.955 ;
        RECT 30.435 -143.645 30.765 -143.315 ;
        RECT 30.435 -145.005 30.765 -144.675 ;
        RECT 30.435 -146.365 30.765 -146.035 ;
        RECT 30.435 -147.725 30.765 -147.395 ;
        RECT 30.435 -149.085 30.765 -148.755 ;
        RECT 30.435 -150.445 30.765 -150.115 ;
        RECT 30.435 -151.805 30.765 -151.475 ;
        RECT 30.435 -153.165 30.765 -152.835 ;
        RECT 30.435 -154.525 30.765 -154.195 ;
        RECT 30.435 -155.885 30.765 -155.555 ;
        RECT 30.435 -157.245 30.765 -156.915 ;
        RECT 30.435 -158.605 30.765 -158.275 ;
        RECT 30.435 -159.965 30.765 -159.635 ;
        RECT 30.435 -161.325 30.765 -160.995 ;
        RECT 30.435 -162.685 30.765 -162.355 ;
        RECT 30.435 -164.045 30.765 -163.715 ;
        RECT 30.435 -165.405 30.765 -165.075 ;
        RECT 30.435 -166.765 30.765 -166.435 ;
        RECT 30.435 -168.125 30.765 -167.795 ;
        RECT 30.435 -169.485 30.765 -169.155 ;
        RECT 30.435 -170.845 30.765 -170.515 ;
        RECT 30.435 -172.205 30.765 -171.875 ;
        RECT 30.435 -173.565 30.765 -173.235 ;
        RECT 30.435 -174.925 30.765 -174.595 ;
        RECT 30.435 -176.285 30.765 -175.955 ;
        RECT 30.435 -177.645 30.765 -177.315 ;
        RECT 30.435 -179.005 30.765 -178.675 ;
        RECT 30.435 -180.365 30.765 -180.035 ;
        RECT 30.435 -181.725 30.765 -181.395 ;
        RECT 30.435 -183.085 30.765 -182.755 ;
        RECT 30.435 -184.445 30.765 -184.115 ;
        RECT 30.435 -185.805 30.765 -185.475 ;
        RECT 30.435 -187.165 30.765 -186.835 ;
        RECT 30.435 -188.525 30.765 -188.195 ;
        RECT 30.435 -189.885 30.765 -189.555 ;
        RECT 30.435 -191.245 30.765 -190.915 ;
        RECT 30.435 -192.605 30.765 -192.275 ;
        RECT 30.435 -193.965 30.765 -193.635 ;
        RECT 30.435 -195.325 30.765 -194.995 ;
        RECT 30.435 -196.685 30.765 -196.355 ;
        RECT 30.435 -198.045 30.765 -197.715 ;
        RECT 30.435 -199.405 30.765 -199.075 ;
        RECT 30.435 -200.765 30.765 -200.435 ;
        RECT 30.435 -202.125 30.765 -201.795 ;
        RECT 30.435 -203.485 30.765 -203.155 ;
        RECT 30.435 -204.845 30.765 -204.515 ;
        RECT 30.435 -206.205 30.765 -205.875 ;
        RECT 30.435 -207.565 30.765 -207.235 ;
        RECT 30.435 -208.925 30.765 -208.595 ;
        RECT 30.435 -210.285 30.765 -209.955 ;
        RECT 30.435 -211.645 30.765 -211.315 ;
        RECT 30.435 -213.005 30.765 -212.675 ;
        RECT 30.435 -214.365 30.765 -214.035 ;
        RECT 30.435 -215.725 30.765 -215.395 ;
        RECT 30.435 -217.085 30.765 -216.755 ;
        RECT 30.435 -218.445 30.765 -218.115 ;
        RECT 30.435 -219.805 30.765 -219.475 ;
        RECT 30.435 -221.165 30.765 -220.835 ;
        RECT 30.435 -222.525 30.765 -222.195 ;
        RECT 30.435 -223.885 30.765 -223.555 ;
        RECT 30.435 -225.245 30.765 -224.915 ;
        RECT 30.435 -226.605 30.765 -226.275 ;
        RECT 30.435 -227.965 30.765 -227.635 ;
        RECT 30.435 -229.325 30.765 -228.995 ;
        RECT 30.435 -230.685 30.765 -230.355 ;
        RECT 30.435 -232.045 30.765 -231.715 ;
        RECT 30.435 -233.405 30.765 -233.075 ;
        RECT 30.435 -234.765 30.765 -234.435 ;
        RECT 30.435 -236.125 30.765 -235.795 ;
        RECT 30.435 -237.485 30.765 -237.155 ;
        RECT 30.435 -238.845 30.765 -238.515 ;
        RECT 30.435 -241.09 30.765 -239.96 ;
        RECT 30.44 -241.205 30.76 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 244.04 32.125 245.17 ;
        RECT 31.795 242.595 32.125 242.925 ;
        RECT 31.795 241.235 32.125 241.565 ;
        RECT 31.795 239.875 32.125 240.205 ;
        RECT 31.795 238.515 32.125 238.845 ;
        RECT 31.795 237.155 32.125 237.485 ;
        RECT 31.8 237.155 32.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -0.845 32.125 -0.515 ;
        RECT 31.795 -2.205 32.125 -1.875 ;
        RECT 31.795 -3.565 32.125 -3.235 ;
        RECT 31.8 -3.565 32.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -123.245 32.125 -122.915 ;
        RECT 31.795 -124.605 32.125 -124.275 ;
        RECT 31.795 -125.965 32.125 -125.635 ;
        RECT 31.795 -127.325 32.125 -126.995 ;
        RECT 31.795 -128.685 32.125 -128.355 ;
        RECT 31.795 -130.045 32.125 -129.715 ;
        RECT 31.795 -131.405 32.125 -131.075 ;
        RECT 31.795 -132.765 32.125 -132.435 ;
        RECT 31.795 -134.125 32.125 -133.795 ;
        RECT 31.795 -135.485 32.125 -135.155 ;
        RECT 31.795 -136.845 32.125 -136.515 ;
        RECT 31.795 -138.205 32.125 -137.875 ;
        RECT 31.795 -139.565 32.125 -139.235 ;
        RECT 31.795 -140.925 32.125 -140.595 ;
        RECT 31.795 -142.285 32.125 -141.955 ;
        RECT 31.795 -143.645 32.125 -143.315 ;
        RECT 31.795 -145.005 32.125 -144.675 ;
        RECT 31.795 -146.365 32.125 -146.035 ;
        RECT 31.795 -147.725 32.125 -147.395 ;
        RECT 31.795 -149.085 32.125 -148.755 ;
        RECT 31.795 -150.445 32.125 -150.115 ;
        RECT 31.795 -151.805 32.125 -151.475 ;
        RECT 31.795 -153.165 32.125 -152.835 ;
        RECT 31.795 -154.525 32.125 -154.195 ;
        RECT 31.795 -155.885 32.125 -155.555 ;
        RECT 31.795 -157.245 32.125 -156.915 ;
        RECT 31.795 -158.605 32.125 -158.275 ;
        RECT 31.795 -159.965 32.125 -159.635 ;
        RECT 31.795 -161.325 32.125 -160.995 ;
        RECT 31.795 -162.685 32.125 -162.355 ;
        RECT 31.795 -164.045 32.125 -163.715 ;
        RECT 31.795 -165.405 32.125 -165.075 ;
        RECT 31.795 -166.765 32.125 -166.435 ;
        RECT 31.795 -168.125 32.125 -167.795 ;
        RECT 31.795 -169.485 32.125 -169.155 ;
        RECT 31.795 -170.845 32.125 -170.515 ;
        RECT 31.795 -172.205 32.125 -171.875 ;
        RECT 31.795 -173.565 32.125 -173.235 ;
        RECT 31.795 -174.925 32.125 -174.595 ;
        RECT 31.795 -176.285 32.125 -175.955 ;
        RECT 31.795 -177.645 32.125 -177.315 ;
        RECT 31.795 -179.005 32.125 -178.675 ;
        RECT 31.795 -180.365 32.125 -180.035 ;
        RECT 31.795 -181.725 32.125 -181.395 ;
        RECT 31.795 -183.085 32.125 -182.755 ;
        RECT 31.795 -184.445 32.125 -184.115 ;
        RECT 31.795 -185.805 32.125 -185.475 ;
        RECT 31.795 -187.165 32.125 -186.835 ;
        RECT 31.795 -188.525 32.125 -188.195 ;
        RECT 31.795 -189.885 32.125 -189.555 ;
        RECT 31.795 -191.245 32.125 -190.915 ;
        RECT 31.795 -192.605 32.125 -192.275 ;
        RECT 31.795 -193.965 32.125 -193.635 ;
        RECT 31.795 -195.325 32.125 -194.995 ;
        RECT 31.795 -196.685 32.125 -196.355 ;
        RECT 31.795 -198.045 32.125 -197.715 ;
        RECT 31.795 -199.405 32.125 -199.075 ;
        RECT 31.795 -200.765 32.125 -200.435 ;
        RECT 31.795 -202.125 32.125 -201.795 ;
        RECT 31.795 -203.485 32.125 -203.155 ;
        RECT 31.795 -204.845 32.125 -204.515 ;
        RECT 31.795 -206.205 32.125 -205.875 ;
        RECT 31.795 -207.565 32.125 -207.235 ;
        RECT 31.795 -208.925 32.125 -208.595 ;
        RECT 31.795 -210.285 32.125 -209.955 ;
        RECT 31.795 -211.645 32.125 -211.315 ;
        RECT 31.795 -213.005 32.125 -212.675 ;
        RECT 31.795 -214.365 32.125 -214.035 ;
        RECT 31.795 -215.725 32.125 -215.395 ;
        RECT 31.795 -217.085 32.125 -216.755 ;
        RECT 31.795 -218.445 32.125 -218.115 ;
        RECT 31.795 -219.805 32.125 -219.475 ;
        RECT 31.795 -221.165 32.125 -220.835 ;
        RECT 31.795 -222.525 32.125 -222.195 ;
        RECT 31.795 -223.885 32.125 -223.555 ;
        RECT 31.795 -225.245 32.125 -224.915 ;
        RECT 31.795 -226.605 32.125 -226.275 ;
        RECT 31.795 -227.965 32.125 -227.635 ;
        RECT 31.795 -229.325 32.125 -228.995 ;
        RECT 31.795 -230.685 32.125 -230.355 ;
        RECT 31.795 -232.045 32.125 -231.715 ;
        RECT 31.795 -233.405 32.125 -233.075 ;
        RECT 31.795 -234.765 32.125 -234.435 ;
        RECT 31.795 -236.125 32.125 -235.795 ;
        RECT 31.795 -237.485 32.125 -237.155 ;
        RECT 31.795 -238.845 32.125 -238.515 ;
        RECT 31.795 -241.09 32.125 -239.96 ;
        RECT 31.8 -241.205 32.12 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 244.04 33.485 245.17 ;
        RECT 33.155 242.595 33.485 242.925 ;
        RECT 33.155 241.235 33.485 241.565 ;
        RECT 33.155 239.875 33.485 240.205 ;
        RECT 33.155 238.515 33.485 238.845 ;
        RECT 33.155 237.155 33.485 237.485 ;
        RECT 33.16 237.155 33.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 -0.845 33.485 -0.515 ;
        RECT 33.155 -2.205 33.485 -1.875 ;
        RECT 33.155 -3.565 33.485 -3.235 ;
        RECT 33.16 -3.565 33.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 -123.245 33.485 -122.915 ;
        RECT 33.155 -124.605 33.485 -124.275 ;
        RECT 33.155 -125.965 33.485 -125.635 ;
        RECT 33.155 -127.325 33.485 -126.995 ;
        RECT 33.155 -128.685 33.485 -128.355 ;
        RECT 33.155 -130.045 33.485 -129.715 ;
        RECT 33.155 -131.405 33.485 -131.075 ;
        RECT 33.155 -132.765 33.485 -132.435 ;
        RECT 33.155 -134.125 33.485 -133.795 ;
        RECT 33.155 -135.485 33.485 -135.155 ;
        RECT 33.155 -136.845 33.485 -136.515 ;
        RECT 33.155 -138.205 33.485 -137.875 ;
        RECT 33.155 -139.565 33.485 -139.235 ;
        RECT 33.155 -140.925 33.485 -140.595 ;
        RECT 33.155 -142.285 33.485 -141.955 ;
        RECT 33.155 -143.645 33.485 -143.315 ;
        RECT 33.155 -145.005 33.485 -144.675 ;
        RECT 33.155 -146.365 33.485 -146.035 ;
        RECT 33.155 -147.725 33.485 -147.395 ;
        RECT 33.155 -149.085 33.485 -148.755 ;
        RECT 33.155 -150.445 33.485 -150.115 ;
        RECT 33.155 -151.805 33.485 -151.475 ;
        RECT 33.155 -153.165 33.485 -152.835 ;
        RECT 33.155 -154.525 33.485 -154.195 ;
        RECT 33.155 -155.885 33.485 -155.555 ;
        RECT 33.155 -157.245 33.485 -156.915 ;
        RECT 33.155 -158.605 33.485 -158.275 ;
        RECT 33.155 -159.965 33.485 -159.635 ;
        RECT 33.155 -161.325 33.485 -160.995 ;
        RECT 33.155 -162.685 33.485 -162.355 ;
        RECT 33.155 -164.045 33.485 -163.715 ;
        RECT 33.155 -165.405 33.485 -165.075 ;
        RECT 33.155 -166.765 33.485 -166.435 ;
        RECT 33.155 -168.125 33.485 -167.795 ;
        RECT 33.155 -169.485 33.485 -169.155 ;
        RECT 33.155 -170.845 33.485 -170.515 ;
        RECT 33.155 -172.205 33.485 -171.875 ;
        RECT 33.155 -173.565 33.485 -173.235 ;
        RECT 33.155 -174.925 33.485 -174.595 ;
        RECT 33.155 -176.285 33.485 -175.955 ;
        RECT 33.155 -177.645 33.485 -177.315 ;
        RECT 33.155 -179.005 33.485 -178.675 ;
        RECT 33.155 -180.365 33.485 -180.035 ;
        RECT 33.155 -181.725 33.485 -181.395 ;
        RECT 33.155 -183.085 33.485 -182.755 ;
        RECT 33.155 -184.445 33.485 -184.115 ;
        RECT 33.155 -185.805 33.485 -185.475 ;
        RECT 33.155 -187.165 33.485 -186.835 ;
        RECT 33.155 -188.525 33.485 -188.195 ;
        RECT 33.155 -189.885 33.485 -189.555 ;
        RECT 33.155 -191.245 33.485 -190.915 ;
        RECT 33.155 -192.605 33.485 -192.275 ;
        RECT 33.155 -193.965 33.485 -193.635 ;
        RECT 33.155 -195.325 33.485 -194.995 ;
        RECT 33.155 -196.685 33.485 -196.355 ;
        RECT 33.155 -198.045 33.485 -197.715 ;
        RECT 33.155 -199.405 33.485 -199.075 ;
        RECT 33.155 -200.765 33.485 -200.435 ;
        RECT 33.155 -202.125 33.485 -201.795 ;
        RECT 33.155 -203.485 33.485 -203.155 ;
        RECT 33.155 -204.845 33.485 -204.515 ;
        RECT 33.155 -206.205 33.485 -205.875 ;
        RECT 33.155 -207.565 33.485 -207.235 ;
        RECT 33.155 -208.925 33.485 -208.595 ;
        RECT 33.155 -210.285 33.485 -209.955 ;
        RECT 33.155 -211.645 33.485 -211.315 ;
        RECT 33.155 -213.005 33.485 -212.675 ;
        RECT 33.155 -214.365 33.485 -214.035 ;
        RECT 33.155 -215.725 33.485 -215.395 ;
        RECT 33.155 -217.085 33.485 -216.755 ;
        RECT 33.155 -218.445 33.485 -218.115 ;
        RECT 33.155 -219.805 33.485 -219.475 ;
        RECT 33.155 -221.165 33.485 -220.835 ;
        RECT 33.155 -222.525 33.485 -222.195 ;
        RECT 33.155 -223.885 33.485 -223.555 ;
        RECT 33.155 -225.245 33.485 -224.915 ;
        RECT 33.155 -226.605 33.485 -226.275 ;
        RECT 33.155 -227.965 33.485 -227.635 ;
        RECT 33.155 -229.325 33.485 -228.995 ;
        RECT 33.155 -230.685 33.485 -230.355 ;
        RECT 33.155 -232.045 33.485 -231.715 ;
        RECT 33.155 -233.405 33.485 -233.075 ;
        RECT 33.155 -234.765 33.485 -234.435 ;
        RECT 33.155 -236.125 33.485 -235.795 ;
        RECT 33.155 -237.485 33.485 -237.155 ;
        RECT 33.155 -238.845 33.485 -238.515 ;
        RECT 33.155 -241.09 33.485 -239.96 ;
        RECT 33.16 -241.205 33.48 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 244.04 34.845 245.17 ;
        RECT 34.515 242.595 34.845 242.925 ;
        RECT 34.515 241.235 34.845 241.565 ;
        RECT 34.515 239.875 34.845 240.205 ;
        RECT 34.515 238.515 34.845 238.845 ;
        RECT 34.515 237.155 34.845 237.485 ;
        RECT 34.52 237.155 34.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 -0.845 34.845 -0.515 ;
        RECT 34.515 -2.205 34.845 -1.875 ;
        RECT 34.515 -3.565 34.845 -3.235 ;
        RECT 34.52 -3.565 34.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 -123.245 34.845 -122.915 ;
        RECT 34.515 -124.605 34.845 -124.275 ;
        RECT 34.515 -125.965 34.845 -125.635 ;
        RECT 34.515 -127.325 34.845 -126.995 ;
        RECT 34.515 -128.685 34.845 -128.355 ;
        RECT 34.515 -130.045 34.845 -129.715 ;
        RECT 34.515 -131.405 34.845 -131.075 ;
        RECT 34.515 -132.765 34.845 -132.435 ;
        RECT 34.515 -134.125 34.845 -133.795 ;
        RECT 34.515 -135.485 34.845 -135.155 ;
        RECT 34.515 -136.845 34.845 -136.515 ;
        RECT 34.515 -138.205 34.845 -137.875 ;
        RECT 34.515 -139.565 34.845 -139.235 ;
        RECT 34.515 -140.925 34.845 -140.595 ;
        RECT 34.515 -142.285 34.845 -141.955 ;
        RECT 34.515 -143.645 34.845 -143.315 ;
        RECT 34.515 -145.005 34.845 -144.675 ;
        RECT 34.515 -146.365 34.845 -146.035 ;
        RECT 34.515 -147.725 34.845 -147.395 ;
        RECT 34.515 -149.085 34.845 -148.755 ;
        RECT 34.515 -150.445 34.845 -150.115 ;
        RECT 34.515 -151.805 34.845 -151.475 ;
        RECT 34.515 -153.165 34.845 -152.835 ;
        RECT 34.515 -154.525 34.845 -154.195 ;
        RECT 34.515 -155.885 34.845 -155.555 ;
        RECT 34.515 -157.245 34.845 -156.915 ;
        RECT 34.515 -158.605 34.845 -158.275 ;
        RECT 34.515 -159.965 34.845 -159.635 ;
        RECT 34.515 -161.325 34.845 -160.995 ;
        RECT 34.515 -162.685 34.845 -162.355 ;
        RECT 34.515 -164.045 34.845 -163.715 ;
        RECT 34.515 -165.405 34.845 -165.075 ;
        RECT 34.515 -166.765 34.845 -166.435 ;
        RECT 34.515 -168.125 34.845 -167.795 ;
        RECT 34.515 -169.485 34.845 -169.155 ;
        RECT 34.515 -170.845 34.845 -170.515 ;
        RECT 34.515 -172.205 34.845 -171.875 ;
        RECT 34.515 -173.565 34.845 -173.235 ;
        RECT 34.515 -174.925 34.845 -174.595 ;
        RECT 34.515 -176.285 34.845 -175.955 ;
        RECT 34.515 -177.645 34.845 -177.315 ;
        RECT 34.515 -179.005 34.845 -178.675 ;
        RECT 34.515 -180.365 34.845 -180.035 ;
        RECT 34.515 -181.725 34.845 -181.395 ;
        RECT 34.515 -183.085 34.845 -182.755 ;
        RECT 34.515 -184.445 34.845 -184.115 ;
        RECT 34.515 -185.805 34.845 -185.475 ;
        RECT 34.515 -187.165 34.845 -186.835 ;
        RECT 34.515 -188.525 34.845 -188.195 ;
        RECT 34.515 -189.885 34.845 -189.555 ;
        RECT 34.515 -191.245 34.845 -190.915 ;
        RECT 34.515 -192.605 34.845 -192.275 ;
        RECT 34.515 -193.965 34.845 -193.635 ;
        RECT 34.515 -195.325 34.845 -194.995 ;
        RECT 34.515 -196.685 34.845 -196.355 ;
        RECT 34.515 -198.045 34.845 -197.715 ;
        RECT 34.515 -199.405 34.845 -199.075 ;
        RECT 34.515 -200.765 34.845 -200.435 ;
        RECT 34.515 -202.125 34.845 -201.795 ;
        RECT 34.515 -203.485 34.845 -203.155 ;
        RECT 34.515 -204.845 34.845 -204.515 ;
        RECT 34.515 -206.205 34.845 -205.875 ;
        RECT 34.515 -207.565 34.845 -207.235 ;
        RECT 34.515 -208.925 34.845 -208.595 ;
        RECT 34.515 -210.285 34.845 -209.955 ;
        RECT 34.515 -211.645 34.845 -211.315 ;
        RECT 34.515 -213.005 34.845 -212.675 ;
        RECT 34.515 -214.365 34.845 -214.035 ;
        RECT 34.515 -215.725 34.845 -215.395 ;
        RECT 34.515 -217.085 34.845 -216.755 ;
        RECT 34.515 -218.445 34.845 -218.115 ;
        RECT 34.515 -219.805 34.845 -219.475 ;
        RECT 34.515 -221.165 34.845 -220.835 ;
        RECT 34.515 -222.525 34.845 -222.195 ;
        RECT 34.515 -223.885 34.845 -223.555 ;
        RECT 34.515 -225.245 34.845 -224.915 ;
        RECT 34.515 -226.605 34.845 -226.275 ;
        RECT 34.515 -227.965 34.845 -227.635 ;
        RECT 34.515 -229.325 34.845 -228.995 ;
        RECT 34.515 -230.685 34.845 -230.355 ;
        RECT 34.515 -232.045 34.845 -231.715 ;
        RECT 34.515 -233.405 34.845 -233.075 ;
        RECT 34.515 -234.765 34.845 -234.435 ;
        RECT 34.515 -236.125 34.845 -235.795 ;
        RECT 34.515 -237.485 34.845 -237.155 ;
        RECT 34.515 -238.845 34.845 -238.515 ;
        RECT 34.515 -241.09 34.845 -239.96 ;
        RECT 34.52 -241.205 34.84 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 244.04 36.205 245.17 ;
        RECT 35.875 242.595 36.205 242.925 ;
        RECT 35.875 241.235 36.205 241.565 ;
        RECT 35.875 239.875 36.205 240.205 ;
        RECT 35.875 238.515 36.205 238.845 ;
        RECT 35.875 237.155 36.205 237.485 ;
        RECT 35.88 237.155 36.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 -127.325 36.205 -126.995 ;
        RECT 35.875 -128.685 36.205 -128.355 ;
        RECT 35.875 -130.045 36.205 -129.715 ;
        RECT 35.875 -131.405 36.205 -131.075 ;
        RECT 35.875 -132.765 36.205 -132.435 ;
        RECT 35.875 -134.125 36.205 -133.795 ;
        RECT 35.875 -135.485 36.205 -135.155 ;
        RECT 35.875 -136.845 36.205 -136.515 ;
        RECT 35.875 -138.205 36.205 -137.875 ;
        RECT 35.875 -139.565 36.205 -139.235 ;
        RECT 35.875 -140.925 36.205 -140.595 ;
        RECT 35.875 -142.285 36.205 -141.955 ;
        RECT 35.875 -143.645 36.205 -143.315 ;
        RECT 35.875 -145.005 36.205 -144.675 ;
        RECT 35.875 -146.365 36.205 -146.035 ;
        RECT 35.875 -147.725 36.205 -147.395 ;
        RECT 35.875 -149.085 36.205 -148.755 ;
        RECT 35.875 -150.445 36.205 -150.115 ;
        RECT 35.875 -151.805 36.205 -151.475 ;
        RECT 35.875 -153.165 36.205 -152.835 ;
        RECT 35.875 -154.525 36.205 -154.195 ;
        RECT 35.875 -155.885 36.205 -155.555 ;
        RECT 35.875 -157.245 36.205 -156.915 ;
        RECT 35.875 -158.605 36.205 -158.275 ;
        RECT 35.875 -159.965 36.205 -159.635 ;
        RECT 35.875 -161.325 36.205 -160.995 ;
        RECT 35.875 -162.685 36.205 -162.355 ;
        RECT 35.875 -164.045 36.205 -163.715 ;
        RECT 35.875 -165.405 36.205 -165.075 ;
        RECT 35.875 -166.765 36.205 -166.435 ;
        RECT 35.875 -168.125 36.205 -167.795 ;
        RECT 35.875 -169.485 36.205 -169.155 ;
        RECT 35.875 -170.845 36.205 -170.515 ;
        RECT 35.875 -172.205 36.205 -171.875 ;
        RECT 35.875 -173.565 36.205 -173.235 ;
        RECT 35.875 -174.925 36.205 -174.595 ;
        RECT 35.875 -176.285 36.205 -175.955 ;
        RECT 35.875 -177.645 36.205 -177.315 ;
        RECT 35.875 -179.005 36.205 -178.675 ;
        RECT 35.875 -180.365 36.205 -180.035 ;
        RECT 35.875 -181.725 36.205 -181.395 ;
        RECT 35.875 -183.085 36.205 -182.755 ;
        RECT 35.875 -184.445 36.205 -184.115 ;
        RECT 35.875 -185.805 36.205 -185.475 ;
        RECT 35.875 -187.165 36.205 -186.835 ;
        RECT 35.875 -188.525 36.205 -188.195 ;
        RECT 35.875 -189.885 36.205 -189.555 ;
        RECT 35.875 -191.245 36.205 -190.915 ;
        RECT 35.875 -192.605 36.205 -192.275 ;
        RECT 35.875 -193.965 36.205 -193.635 ;
        RECT 35.875 -195.325 36.205 -194.995 ;
        RECT 35.875 -196.685 36.205 -196.355 ;
        RECT 35.875 -198.045 36.205 -197.715 ;
        RECT 35.875 -199.405 36.205 -199.075 ;
        RECT 35.875 -200.765 36.205 -200.435 ;
        RECT 35.875 -202.125 36.205 -201.795 ;
        RECT 35.875 -203.485 36.205 -203.155 ;
        RECT 35.875 -204.845 36.205 -204.515 ;
        RECT 35.875 -206.205 36.205 -205.875 ;
        RECT 35.875 -207.565 36.205 -207.235 ;
        RECT 35.875 -208.925 36.205 -208.595 ;
        RECT 35.875 -210.285 36.205 -209.955 ;
        RECT 35.875 -211.645 36.205 -211.315 ;
        RECT 35.875 -213.005 36.205 -212.675 ;
        RECT 35.875 -214.365 36.205 -214.035 ;
        RECT 35.875 -215.725 36.205 -215.395 ;
        RECT 35.875 -217.085 36.205 -216.755 ;
        RECT 35.875 -218.445 36.205 -218.115 ;
        RECT 35.875 -219.805 36.205 -219.475 ;
        RECT 35.875 -221.165 36.205 -220.835 ;
        RECT 35.875 -222.525 36.205 -222.195 ;
        RECT 35.875 -223.885 36.205 -223.555 ;
        RECT 35.875 -225.245 36.205 -224.915 ;
        RECT 35.875 -226.605 36.205 -226.275 ;
        RECT 35.875 -227.965 36.205 -227.635 ;
        RECT 35.875 -229.325 36.205 -228.995 ;
        RECT 35.875 -230.685 36.205 -230.355 ;
        RECT 35.875 -232.045 36.205 -231.715 ;
        RECT 35.875 -233.405 36.205 -233.075 ;
        RECT 35.875 -234.765 36.205 -234.435 ;
        RECT 35.875 -236.125 36.205 -235.795 ;
        RECT 35.875 -237.485 36.205 -237.155 ;
        RECT 35.875 -238.845 36.205 -238.515 ;
        RECT 35.875 -241.09 36.205 -239.96 ;
        RECT 35.88 -241.205 36.2 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.01 -125.535 36.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 244.04 37.565 245.17 ;
        RECT 37.235 242.595 37.565 242.925 ;
        RECT 37.235 241.235 37.565 241.565 ;
        RECT 37.235 239.875 37.565 240.205 ;
        RECT 37.235 238.515 37.565 238.845 ;
        RECT 37.235 237.155 37.565 237.485 ;
        RECT 37.24 237.155 37.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 -0.845 37.565 -0.515 ;
        RECT 37.235 -2.205 37.565 -1.875 ;
        RECT 37.235 -3.565 37.565 -3.235 ;
        RECT 37.24 -3.565 37.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 244.04 38.925 245.17 ;
        RECT 38.595 242.595 38.925 242.925 ;
        RECT 38.595 241.235 38.925 241.565 ;
        RECT 38.595 239.875 38.925 240.205 ;
        RECT 38.595 238.515 38.925 238.845 ;
        RECT 38.595 237.155 38.925 237.485 ;
        RECT 38.6 237.155 38.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 -0.845 38.925 -0.515 ;
        RECT 38.595 -2.205 38.925 -1.875 ;
        RECT 38.595 -3.565 38.925 -3.235 ;
        RECT 38.6 -3.565 38.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 244.04 40.285 245.17 ;
        RECT 39.955 242.595 40.285 242.925 ;
        RECT 39.955 241.235 40.285 241.565 ;
        RECT 39.955 239.875 40.285 240.205 ;
        RECT 39.955 238.515 40.285 238.845 ;
        RECT 39.955 237.155 40.285 237.485 ;
        RECT 39.96 237.155 40.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 -0.845 40.285 -0.515 ;
        RECT 39.955 -2.205 40.285 -1.875 ;
        RECT 39.955 -3.565 40.285 -3.235 ;
        RECT 39.96 -3.565 40.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 -139.565 40.285 -139.235 ;
        RECT 39.955 -140.925 40.285 -140.595 ;
        RECT 39.955 -142.285 40.285 -141.955 ;
        RECT 39.955 -143.645 40.285 -143.315 ;
        RECT 39.955 -145.005 40.285 -144.675 ;
        RECT 39.955 -146.365 40.285 -146.035 ;
        RECT 39.955 -147.725 40.285 -147.395 ;
        RECT 39.955 -149.085 40.285 -148.755 ;
        RECT 39.955 -150.445 40.285 -150.115 ;
        RECT 39.955 -151.805 40.285 -151.475 ;
        RECT 39.955 -153.165 40.285 -152.835 ;
        RECT 39.955 -154.525 40.285 -154.195 ;
        RECT 39.955 -155.885 40.285 -155.555 ;
        RECT 39.955 -157.245 40.285 -156.915 ;
        RECT 39.955 -158.605 40.285 -158.275 ;
        RECT 39.955 -159.965 40.285 -159.635 ;
        RECT 39.955 -161.325 40.285 -160.995 ;
        RECT 39.955 -162.685 40.285 -162.355 ;
        RECT 39.955 -164.045 40.285 -163.715 ;
        RECT 39.955 -165.405 40.285 -165.075 ;
        RECT 39.955 -166.765 40.285 -166.435 ;
        RECT 39.955 -168.125 40.285 -167.795 ;
        RECT 39.955 -169.485 40.285 -169.155 ;
        RECT 39.955 -170.845 40.285 -170.515 ;
        RECT 39.955 -172.205 40.285 -171.875 ;
        RECT 39.955 -173.565 40.285 -173.235 ;
        RECT 39.955 -174.925 40.285 -174.595 ;
        RECT 39.955 -176.285 40.285 -175.955 ;
        RECT 39.955 -177.645 40.285 -177.315 ;
        RECT 39.955 -179.005 40.285 -178.675 ;
        RECT 39.955 -180.365 40.285 -180.035 ;
        RECT 39.955 -181.725 40.285 -181.395 ;
        RECT 39.955 -183.085 40.285 -182.755 ;
        RECT 39.955 -184.445 40.285 -184.115 ;
        RECT 39.955 -185.805 40.285 -185.475 ;
        RECT 39.955 -187.165 40.285 -186.835 ;
        RECT 39.955 -188.525 40.285 -188.195 ;
        RECT 39.955 -189.885 40.285 -189.555 ;
        RECT 39.955 -191.245 40.285 -190.915 ;
        RECT 39.955 -192.605 40.285 -192.275 ;
        RECT 39.955 -193.965 40.285 -193.635 ;
        RECT 39.955 -195.325 40.285 -194.995 ;
        RECT 39.955 -196.685 40.285 -196.355 ;
        RECT 39.955 -198.045 40.285 -197.715 ;
        RECT 39.955 -199.405 40.285 -199.075 ;
        RECT 39.955 -200.765 40.285 -200.435 ;
        RECT 39.955 -202.125 40.285 -201.795 ;
        RECT 39.955 -203.485 40.285 -203.155 ;
        RECT 39.955 -204.845 40.285 -204.515 ;
        RECT 39.955 -206.205 40.285 -205.875 ;
        RECT 39.955 -207.565 40.285 -207.235 ;
        RECT 39.955 -208.925 40.285 -208.595 ;
        RECT 39.955 -210.285 40.285 -209.955 ;
        RECT 39.955 -211.645 40.285 -211.315 ;
        RECT 39.955 -213.005 40.285 -212.675 ;
        RECT 39.955 -214.365 40.285 -214.035 ;
        RECT 39.955 -215.725 40.285 -215.395 ;
        RECT 39.955 -217.085 40.285 -216.755 ;
        RECT 39.955 -218.445 40.285 -218.115 ;
        RECT 39.955 -219.805 40.285 -219.475 ;
        RECT 39.955 -221.165 40.285 -220.835 ;
        RECT 39.955 -222.525 40.285 -222.195 ;
        RECT 39.955 -223.885 40.285 -223.555 ;
        RECT 39.955 -225.245 40.285 -224.915 ;
        RECT 39.955 -226.605 40.285 -226.275 ;
        RECT 39.955 -227.965 40.285 -227.635 ;
        RECT 39.955 -229.325 40.285 -228.995 ;
        RECT 39.955 -230.685 40.285 -230.355 ;
        RECT 39.955 -232.045 40.285 -231.715 ;
        RECT 39.955 -233.405 40.285 -233.075 ;
        RECT 39.955 -234.765 40.285 -234.435 ;
        RECT 39.955 -236.125 40.285 -235.795 ;
        RECT 39.955 -237.485 40.285 -237.155 ;
        RECT 39.955 -238.845 40.285 -238.515 ;
        RECT 39.955 -241.09 40.285 -239.96 ;
        RECT 39.96 -241.205 40.28 -122.24 ;
        RECT 39.955 -123.245 40.285 -122.915 ;
        RECT 39.955 -124.605 40.285 -124.275 ;
        RECT 39.955 -125.965 40.285 -125.635 ;
        RECT 39.955 -127.325 40.285 -126.995 ;
        RECT 39.955 -128.685 40.285 -128.355 ;
        RECT 39.955 -130.045 40.285 -129.715 ;
        RECT 39.955 -131.405 40.285 -131.075 ;
        RECT 39.955 -132.765 40.285 -132.435 ;
        RECT 39.955 -134.125 40.285 -133.795 ;
        RECT 39.955 -135.485 40.285 -135.155 ;
        RECT 39.955 -136.845 40.285 -136.515 ;
        RECT 39.955 -138.205 40.285 -137.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.31 -125.535 3.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 244.04 4.925 245.17 ;
        RECT 4.595 242.595 4.925 242.925 ;
        RECT 4.595 241.235 4.925 241.565 ;
        RECT 4.595 239.875 4.925 240.205 ;
        RECT 4.595 238.515 4.925 238.845 ;
        RECT 4.595 237.155 4.925 237.485 ;
        RECT 4.6 237.155 4.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 -0.845 4.925 -0.515 ;
        RECT 4.595 -2.205 4.925 -1.875 ;
        RECT 4.595 -3.565 4.925 -3.235 ;
        RECT 4.6 -3.565 4.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 244.04 6.285 245.17 ;
        RECT 5.955 242.595 6.285 242.925 ;
        RECT 5.955 241.235 6.285 241.565 ;
        RECT 5.955 239.875 6.285 240.205 ;
        RECT 5.955 238.515 6.285 238.845 ;
        RECT 5.955 237.155 6.285 237.485 ;
        RECT 5.96 237.155 6.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 -0.845 6.285 -0.515 ;
        RECT 5.955 -2.205 6.285 -1.875 ;
        RECT 5.955 -3.565 6.285 -3.235 ;
        RECT 5.96 -3.565 6.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 244.04 7.645 245.17 ;
        RECT 7.315 242.595 7.645 242.925 ;
        RECT 7.315 241.235 7.645 241.565 ;
        RECT 7.315 239.875 7.645 240.205 ;
        RECT 7.315 238.515 7.645 238.845 ;
        RECT 7.315 237.155 7.645 237.485 ;
        RECT 7.32 237.155 7.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -0.845 7.645 -0.515 ;
        RECT 7.315 -2.205 7.645 -1.875 ;
        RECT 7.315 -3.565 7.645 -3.235 ;
        RECT 7.32 -3.565 7.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -123.245 7.645 -122.915 ;
        RECT 7.315 -124.605 7.645 -124.275 ;
        RECT 7.315 -125.965 7.645 -125.635 ;
        RECT 7.315 -127.325 7.645 -126.995 ;
        RECT 7.315 -128.685 7.645 -128.355 ;
        RECT 7.315 -130.045 7.645 -129.715 ;
        RECT 7.315 -131.405 7.645 -131.075 ;
        RECT 7.315 -132.765 7.645 -132.435 ;
        RECT 7.315 -134.125 7.645 -133.795 ;
        RECT 7.315 -135.485 7.645 -135.155 ;
        RECT 7.315 -136.845 7.645 -136.515 ;
        RECT 7.315 -138.205 7.645 -137.875 ;
        RECT 7.315 -139.565 7.645 -139.235 ;
        RECT 7.315 -140.925 7.645 -140.595 ;
        RECT 7.315 -142.285 7.645 -141.955 ;
        RECT 7.315 -143.645 7.645 -143.315 ;
        RECT 7.315 -145.005 7.645 -144.675 ;
        RECT 7.315 -146.365 7.645 -146.035 ;
        RECT 7.315 -147.725 7.645 -147.395 ;
        RECT 7.315 -149.085 7.645 -148.755 ;
        RECT 7.315 -150.445 7.645 -150.115 ;
        RECT 7.315 -151.805 7.645 -151.475 ;
        RECT 7.315 -153.165 7.645 -152.835 ;
        RECT 7.315 -154.525 7.645 -154.195 ;
        RECT 7.315 -155.885 7.645 -155.555 ;
        RECT 7.315 -157.245 7.645 -156.915 ;
        RECT 7.315 -158.605 7.645 -158.275 ;
        RECT 7.315 -159.965 7.645 -159.635 ;
        RECT 7.315 -161.325 7.645 -160.995 ;
        RECT 7.315 -162.685 7.645 -162.355 ;
        RECT 7.315 -164.045 7.645 -163.715 ;
        RECT 7.315 -165.405 7.645 -165.075 ;
        RECT 7.315 -166.765 7.645 -166.435 ;
        RECT 7.315 -168.125 7.645 -167.795 ;
        RECT 7.315 -169.485 7.645 -169.155 ;
        RECT 7.315 -170.845 7.645 -170.515 ;
        RECT 7.315 -172.205 7.645 -171.875 ;
        RECT 7.315 -173.565 7.645 -173.235 ;
        RECT 7.315 -174.925 7.645 -174.595 ;
        RECT 7.315 -176.285 7.645 -175.955 ;
        RECT 7.315 -177.645 7.645 -177.315 ;
        RECT 7.315 -179.005 7.645 -178.675 ;
        RECT 7.315 -180.365 7.645 -180.035 ;
        RECT 7.315 -181.725 7.645 -181.395 ;
        RECT 7.315 -183.085 7.645 -182.755 ;
        RECT 7.315 -184.445 7.645 -184.115 ;
        RECT 7.315 -185.805 7.645 -185.475 ;
        RECT 7.315 -187.165 7.645 -186.835 ;
        RECT 7.315 -188.525 7.645 -188.195 ;
        RECT 7.315 -189.885 7.645 -189.555 ;
        RECT 7.315 -191.245 7.645 -190.915 ;
        RECT 7.315 -192.605 7.645 -192.275 ;
        RECT 7.315 -193.965 7.645 -193.635 ;
        RECT 7.315 -195.325 7.645 -194.995 ;
        RECT 7.315 -196.685 7.645 -196.355 ;
        RECT 7.315 -198.045 7.645 -197.715 ;
        RECT 7.315 -199.405 7.645 -199.075 ;
        RECT 7.315 -200.765 7.645 -200.435 ;
        RECT 7.315 -202.125 7.645 -201.795 ;
        RECT 7.315 -203.485 7.645 -203.155 ;
        RECT 7.315 -204.845 7.645 -204.515 ;
        RECT 7.315 -206.205 7.645 -205.875 ;
        RECT 7.315 -207.565 7.645 -207.235 ;
        RECT 7.315 -208.925 7.645 -208.595 ;
        RECT 7.315 -210.285 7.645 -209.955 ;
        RECT 7.315 -211.645 7.645 -211.315 ;
        RECT 7.315 -213.005 7.645 -212.675 ;
        RECT 7.315 -214.365 7.645 -214.035 ;
        RECT 7.315 -215.725 7.645 -215.395 ;
        RECT 7.315 -217.085 7.645 -216.755 ;
        RECT 7.315 -218.445 7.645 -218.115 ;
        RECT 7.315 -219.805 7.645 -219.475 ;
        RECT 7.315 -221.165 7.645 -220.835 ;
        RECT 7.315 -222.525 7.645 -222.195 ;
        RECT 7.315 -223.885 7.645 -223.555 ;
        RECT 7.315 -225.245 7.645 -224.915 ;
        RECT 7.315 -226.605 7.645 -226.275 ;
        RECT 7.315 -227.965 7.645 -227.635 ;
        RECT 7.315 -229.325 7.645 -228.995 ;
        RECT 7.315 -230.685 7.645 -230.355 ;
        RECT 7.315 -232.045 7.645 -231.715 ;
        RECT 7.315 -233.405 7.645 -233.075 ;
        RECT 7.315 -234.765 7.645 -234.435 ;
        RECT 7.315 -236.125 7.645 -235.795 ;
        RECT 7.315 -237.485 7.645 -237.155 ;
        RECT 7.315 -238.845 7.645 -238.515 ;
        RECT 7.315 -241.09 7.645 -239.96 ;
        RECT 7.32 -241.205 7.64 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 244.04 9.005 245.17 ;
        RECT 8.675 242.595 9.005 242.925 ;
        RECT 8.675 241.235 9.005 241.565 ;
        RECT 8.675 239.875 9.005 240.205 ;
        RECT 8.675 238.515 9.005 238.845 ;
        RECT 8.675 237.155 9.005 237.485 ;
        RECT 8.68 237.155 9 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 -0.845 9.005 -0.515 ;
        RECT 8.675 -2.205 9.005 -1.875 ;
        RECT 8.675 -3.565 9.005 -3.235 ;
        RECT 8.68 -3.565 9 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 -123.245 9.005 -122.915 ;
        RECT 8.675 -124.605 9.005 -124.275 ;
        RECT 8.675 -125.965 9.005 -125.635 ;
        RECT 8.675 -127.325 9.005 -126.995 ;
        RECT 8.675 -128.685 9.005 -128.355 ;
        RECT 8.675 -130.045 9.005 -129.715 ;
        RECT 8.675 -131.405 9.005 -131.075 ;
        RECT 8.675 -132.765 9.005 -132.435 ;
        RECT 8.675 -134.125 9.005 -133.795 ;
        RECT 8.675 -135.485 9.005 -135.155 ;
        RECT 8.675 -136.845 9.005 -136.515 ;
        RECT 8.675 -138.205 9.005 -137.875 ;
        RECT 8.675 -139.565 9.005 -139.235 ;
        RECT 8.675 -140.925 9.005 -140.595 ;
        RECT 8.675 -142.285 9.005 -141.955 ;
        RECT 8.675 -143.645 9.005 -143.315 ;
        RECT 8.675 -145.005 9.005 -144.675 ;
        RECT 8.675 -146.365 9.005 -146.035 ;
        RECT 8.675 -147.725 9.005 -147.395 ;
        RECT 8.675 -149.085 9.005 -148.755 ;
        RECT 8.675 -150.445 9.005 -150.115 ;
        RECT 8.675 -151.805 9.005 -151.475 ;
        RECT 8.675 -153.165 9.005 -152.835 ;
        RECT 8.675 -154.525 9.005 -154.195 ;
        RECT 8.675 -155.885 9.005 -155.555 ;
        RECT 8.675 -157.245 9.005 -156.915 ;
        RECT 8.675 -158.605 9.005 -158.275 ;
        RECT 8.675 -159.965 9.005 -159.635 ;
        RECT 8.675 -161.325 9.005 -160.995 ;
        RECT 8.675 -162.685 9.005 -162.355 ;
        RECT 8.675 -164.045 9.005 -163.715 ;
        RECT 8.675 -165.405 9.005 -165.075 ;
        RECT 8.675 -166.765 9.005 -166.435 ;
        RECT 8.675 -168.125 9.005 -167.795 ;
        RECT 8.675 -169.485 9.005 -169.155 ;
        RECT 8.675 -170.845 9.005 -170.515 ;
        RECT 8.675 -172.205 9.005 -171.875 ;
        RECT 8.675 -173.565 9.005 -173.235 ;
        RECT 8.675 -174.925 9.005 -174.595 ;
        RECT 8.675 -176.285 9.005 -175.955 ;
        RECT 8.675 -177.645 9.005 -177.315 ;
        RECT 8.675 -179.005 9.005 -178.675 ;
        RECT 8.675 -180.365 9.005 -180.035 ;
        RECT 8.675 -181.725 9.005 -181.395 ;
        RECT 8.675 -183.085 9.005 -182.755 ;
        RECT 8.675 -184.445 9.005 -184.115 ;
        RECT 8.675 -185.805 9.005 -185.475 ;
        RECT 8.675 -187.165 9.005 -186.835 ;
        RECT 8.675 -188.525 9.005 -188.195 ;
        RECT 8.675 -189.885 9.005 -189.555 ;
        RECT 8.675 -191.245 9.005 -190.915 ;
        RECT 8.675 -192.605 9.005 -192.275 ;
        RECT 8.675 -193.965 9.005 -193.635 ;
        RECT 8.675 -195.325 9.005 -194.995 ;
        RECT 8.675 -196.685 9.005 -196.355 ;
        RECT 8.675 -198.045 9.005 -197.715 ;
        RECT 8.675 -199.405 9.005 -199.075 ;
        RECT 8.675 -200.765 9.005 -200.435 ;
        RECT 8.675 -202.125 9.005 -201.795 ;
        RECT 8.675 -203.485 9.005 -203.155 ;
        RECT 8.675 -204.845 9.005 -204.515 ;
        RECT 8.675 -206.205 9.005 -205.875 ;
        RECT 8.675 -207.565 9.005 -207.235 ;
        RECT 8.675 -208.925 9.005 -208.595 ;
        RECT 8.675 -210.285 9.005 -209.955 ;
        RECT 8.675 -211.645 9.005 -211.315 ;
        RECT 8.675 -213.005 9.005 -212.675 ;
        RECT 8.675 -214.365 9.005 -214.035 ;
        RECT 8.675 -215.725 9.005 -215.395 ;
        RECT 8.675 -217.085 9.005 -216.755 ;
        RECT 8.675 -218.445 9.005 -218.115 ;
        RECT 8.675 -219.805 9.005 -219.475 ;
        RECT 8.675 -221.165 9.005 -220.835 ;
        RECT 8.675 -222.525 9.005 -222.195 ;
        RECT 8.675 -223.885 9.005 -223.555 ;
        RECT 8.675 -225.245 9.005 -224.915 ;
        RECT 8.675 -226.605 9.005 -226.275 ;
        RECT 8.675 -227.965 9.005 -227.635 ;
        RECT 8.675 -229.325 9.005 -228.995 ;
        RECT 8.675 -230.685 9.005 -230.355 ;
        RECT 8.675 -232.045 9.005 -231.715 ;
        RECT 8.675 -233.405 9.005 -233.075 ;
        RECT 8.675 -234.765 9.005 -234.435 ;
        RECT 8.675 -236.125 9.005 -235.795 ;
        RECT 8.675 -237.485 9.005 -237.155 ;
        RECT 8.675 -238.845 9.005 -238.515 ;
        RECT 8.675 -241.09 9.005 -239.96 ;
        RECT 8.68 -241.205 9 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 244.04 10.365 245.17 ;
        RECT 10.035 242.595 10.365 242.925 ;
        RECT 10.035 241.235 10.365 241.565 ;
        RECT 10.035 239.875 10.365 240.205 ;
        RECT 10.035 238.515 10.365 238.845 ;
        RECT 10.035 237.155 10.365 237.485 ;
        RECT 10.04 237.155 10.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 -0.845 10.365 -0.515 ;
        RECT 10.035 -2.205 10.365 -1.875 ;
        RECT 10.035 -3.565 10.365 -3.235 ;
        RECT 10.04 -3.565 10.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 -123.245 10.365 -122.915 ;
        RECT 10.035 -124.605 10.365 -124.275 ;
        RECT 10.035 -125.965 10.365 -125.635 ;
        RECT 10.035 -127.325 10.365 -126.995 ;
        RECT 10.035 -128.685 10.365 -128.355 ;
        RECT 10.035 -130.045 10.365 -129.715 ;
        RECT 10.035 -131.405 10.365 -131.075 ;
        RECT 10.035 -132.765 10.365 -132.435 ;
        RECT 10.035 -134.125 10.365 -133.795 ;
        RECT 10.035 -135.485 10.365 -135.155 ;
        RECT 10.035 -136.845 10.365 -136.515 ;
        RECT 10.035 -138.205 10.365 -137.875 ;
        RECT 10.035 -139.565 10.365 -139.235 ;
        RECT 10.035 -140.925 10.365 -140.595 ;
        RECT 10.035 -142.285 10.365 -141.955 ;
        RECT 10.035 -143.645 10.365 -143.315 ;
        RECT 10.035 -145.005 10.365 -144.675 ;
        RECT 10.035 -146.365 10.365 -146.035 ;
        RECT 10.035 -147.725 10.365 -147.395 ;
        RECT 10.035 -149.085 10.365 -148.755 ;
        RECT 10.035 -150.445 10.365 -150.115 ;
        RECT 10.035 -151.805 10.365 -151.475 ;
        RECT 10.035 -153.165 10.365 -152.835 ;
        RECT 10.035 -154.525 10.365 -154.195 ;
        RECT 10.035 -155.885 10.365 -155.555 ;
        RECT 10.035 -157.245 10.365 -156.915 ;
        RECT 10.035 -158.605 10.365 -158.275 ;
        RECT 10.035 -159.965 10.365 -159.635 ;
        RECT 10.035 -161.325 10.365 -160.995 ;
        RECT 10.035 -162.685 10.365 -162.355 ;
        RECT 10.035 -164.045 10.365 -163.715 ;
        RECT 10.035 -165.405 10.365 -165.075 ;
        RECT 10.035 -166.765 10.365 -166.435 ;
        RECT 10.035 -168.125 10.365 -167.795 ;
        RECT 10.035 -169.485 10.365 -169.155 ;
        RECT 10.035 -170.845 10.365 -170.515 ;
        RECT 10.035 -172.205 10.365 -171.875 ;
        RECT 10.035 -173.565 10.365 -173.235 ;
        RECT 10.035 -174.925 10.365 -174.595 ;
        RECT 10.035 -176.285 10.365 -175.955 ;
        RECT 10.035 -177.645 10.365 -177.315 ;
        RECT 10.035 -179.005 10.365 -178.675 ;
        RECT 10.035 -180.365 10.365 -180.035 ;
        RECT 10.035 -181.725 10.365 -181.395 ;
        RECT 10.035 -183.085 10.365 -182.755 ;
        RECT 10.035 -184.445 10.365 -184.115 ;
        RECT 10.035 -185.805 10.365 -185.475 ;
        RECT 10.035 -187.165 10.365 -186.835 ;
        RECT 10.035 -188.525 10.365 -188.195 ;
        RECT 10.035 -189.885 10.365 -189.555 ;
        RECT 10.035 -191.245 10.365 -190.915 ;
        RECT 10.035 -192.605 10.365 -192.275 ;
        RECT 10.035 -193.965 10.365 -193.635 ;
        RECT 10.035 -195.325 10.365 -194.995 ;
        RECT 10.035 -196.685 10.365 -196.355 ;
        RECT 10.035 -198.045 10.365 -197.715 ;
        RECT 10.035 -199.405 10.365 -199.075 ;
        RECT 10.035 -200.765 10.365 -200.435 ;
        RECT 10.035 -202.125 10.365 -201.795 ;
        RECT 10.035 -203.485 10.365 -203.155 ;
        RECT 10.035 -204.845 10.365 -204.515 ;
        RECT 10.035 -206.205 10.365 -205.875 ;
        RECT 10.035 -207.565 10.365 -207.235 ;
        RECT 10.035 -208.925 10.365 -208.595 ;
        RECT 10.035 -210.285 10.365 -209.955 ;
        RECT 10.035 -211.645 10.365 -211.315 ;
        RECT 10.035 -213.005 10.365 -212.675 ;
        RECT 10.035 -214.365 10.365 -214.035 ;
        RECT 10.035 -215.725 10.365 -215.395 ;
        RECT 10.035 -217.085 10.365 -216.755 ;
        RECT 10.035 -218.445 10.365 -218.115 ;
        RECT 10.035 -219.805 10.365 -219.475 ;
        RECT 10.035 -221.165 10.365 -220.835 ;
        RECT 10.035 -222.525 10.365 -222.195 ;
        RECT 10.035 -223.885 10.365 -223.555 ;
        RECT 10.035 -225.245 10.365 -224.915 ;
        RECT 10.035 -226.605 10.365 -226.275 ;
        RECT 10.035 -227.965 10.365 -227.635 ;
        RECT 10.035 -229.325 10.365 -228.995 ;
        RECT 10.035 -230.685 10.365 -230.355 ;
        RECT 10.035 -232.045 10.365 -231.715 ;
        RECT 10.035 -233.405 10.365 -233.075 ;
        RECT 10.035 -234.765 10.365 -234.435 ;
        RECT 10.035 -236.125 10.365 -235.795 ;
        RECT 10.035 -237.485 10.365 -237.155 ;
        RECT 10.035 -238.845 10.365 -238.515 ;
        RECT 10.035 -241.09 10.365 -239.96 ;
        RECT 10.04 -241.205 10.36 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 244.04 11.725 245.17 ;
        RECT 11.395 242.595 11.725 242.925 ;
        RECT 11.395 241.235 11.725 241.565 ;
        RECT 11.395 239.875 11.725 240.205 ;
        RECT 11.395 238.515 11.725 238.845 ;
        RECT 11.395 237.155 11.725 237.485 ;
        RECT 11.4 237.155 11.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 -0.845 11.725 -0.515 ;
        RECT 11.395 -2.205 11.725 -1.875 ;
        RECT 11.395 -3.565 11.725 -3.235 ;
        RECT 11.4 -3.565 11.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 -123.245 11.725 -122.915 ;
        RECT 11.395 -124.605 11.725 -124.275 ;
        RECT 11.395 -125.965 11.725 -125.635 ;
        RECT 11.395 -127.325 11.725 -126.995 ;
        RECT 11.395 -128.685 11.725 -128.355 ;
        RECT 11.395 -130.045 11.725 -129.715 ;
        RECT 11.395 -131.405 11.725 -131.075 ;
        RECT 11.395 -132.765 11.725 -132.435 ;
        RECT 11.395 -134.125 11.725 -133.795 ;
        RECT 11.395 -135.485 11.725 -135.155 ;
        RECT 11.395 -136.845 11.725 -136.515 ;
        RECT 11.395 -138.205 11.725 -137.875 ;
        RECT 11.395 -139.565 11.725 -139.235 ;
        RECT 11.395 -140.925 11.725 -140.595 ;
        RECT 11.395 -142.285 11.725 -141.955 ;
        RECT 11.395 -143.645 11.725 -143.315 ;
        RECT 11.395 -145.005 11.725 -144.675 ;
        RECT 11.395 -146.365 11.725 -146.035 ;
        RECT 11.395 -147.725 11.725 -147.395 ;
        RECT 11.395 -149.085 11.725 -148.755 ;
        RECT 11.395 -150.445 11.725 -150.115 ;
        RECT 11.395 -151.805 11.725 -151.475 ;
        RECT 11.395 -153.165 11.725 -152.835 ;
        RECT 11.395 -154.525 11.725 -154.195 ;
        RECT 11.395 -155.885 11.725 -155.555 ;
        RECT 11.395 -157.245 11.725 -156.915 ;
        RECT 11.395 -158.605 11.725 -158.275 ;
        RECT 11.395 -159.965 11.725 -159.635 ;
        RECT 11.395 -161.325 11.725 -160.995 ;
        RECT 11.395 -162.685 11.725 -162.355 ;
        RECT 11.395 -164.045 11.725 -163.715 ;
        RECT 11.395 -165.405 11.725 -165.075 ;
        RECT 11.395 -166.765 11.725 -166.435 ;
        RECT 11.395 -168.125 11.725 -167.795 ;
        RECT 11.395 -169.485 11.725 -169.155 ;
        RECT 11.395 -170.845 11.725 -170.515 ;
        RECT 11.395 -172.205 11.725 -171.875 ;
        RECT 11.395 -173.565 11.725 -173.235 ;
        RECT 11.395 -174.925 11.725 -174.595 ;
        RECT 11.395 -176.285 11.725 -175.955 ;
        RECT 11.395 -177.645 11.725 -177.315 ;
        RECT 11.395 -179.005 11.725 -178.675 ;
        RECT 11.395 -180.365 11.725 -180.035 ;
        RECT 11.395 -181.725 11.725 -181.395 ;
        RECT 11.395 -183.085 11.725 -182.755 ;
        RECT 11.395 -184.445 11.725 -184.115 ;
        RECT 11.395 -185.805 11.725 -185.475 ;
        RECT 11.395 -187.165 11.725 -186.835 ;
        RECT 11.395 -188.525 11.725 -188.195 ;
        RECT 11.395 -189.885 11.725 -189.555 ;
        RECT 11.395 -191.245 11.725 -190.915 ;
        RECT 11.395 -192.605 11.725 -192.275 ;
        RECT 11.395 -193.965 11.725 -193.635 ;
        RECT 11.395 -195.325 11.725 -194.995 ;
        RECT 11.395 -196.685 11.725 -196.355 ;
        RECT 11.395 -198.045 11.725 -197.715 ;
        RECT 11.395 -199.405 11.725 -199.075 ;
        RECT 11.395 -200.765 11.725 -200.435 ;
        RECT 11.395 -202.125 11.725 -201.795 ;
        RECT 11.395 -203.485 11.725 -203.155 ;
        RECT 11.395 -204.845 11.725 -204.515 ;
        RECT 11.395 -206.205 11.725 -205.875 ;
        RECT 11.395 -207.565 11.725 -207.235 ;
        RECT 11.395 -208.925 11.725 -208.595 ;
        RECT 11.395 -210.285 11.725 -209.955 ;
        RECT 11.395 -211.645 11.725 -211.315 ;
        RECT 11.395 -213.005 11.725 -212.675 ;
        RECT 11.395 -214.365 11.725 -214.035 ;
        RECT 11.395 -215.725 11.725 -215.395 ;
        RECT 11.395 -217.085 11.725 -216.755 ;
        RECT 11.395 -218.445 11.725 -218.115 ;
        RECT 11.395 -219.805 11.725 -219.475 ;
        RECT 11.395 -221.165 11.725 -220.835 ;
        RECT 11.395 -222.525 11.725 -222.195 ;
        RECT 11.395 -223.885 11.725 -223.555 ;
        RECT 11.395 -225.245 11.725 -224.915 ;
        RECT 11.395 -226.605 11.725 -226.275 ;
        RECT 11.395 -227.965 11.725 -227.635 ;
        RECT 11.395 -229.325 11.725 -228.995 ;
        RECT 11.395 -230.685 11.725 -230.355 ;
        RECT 11.395 -232.045 11.725 -231.715 ;
        RECT 11.395 -233.405 11.725 -233.075 ;
        RECT 11.395 -234.765 11.725 -234.435 ;
        RECT 11.395 -236.125 11.725 -235.795 ;
        RECT 11.395 -237.485 11.725 -237.155 ;
        RECT 11.395 -238.845 11.725 -238.515 ;
        RECT 11.395 -241.09 11.725 -239.96 ;
        RECT 11.4 -241.205 11.72 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 244.04 13.085 245.17 ;
        RECT 12.755 242.595 13.085 242.925 ;
        RECT 12.755 241.235 13.085 241.565 ;
        RECT 12.755 239.875 13.085 240.205 ;
        RECT 12.755 238.515 13.085 238.845 ;
        RECT 12.755 237.155 13.085 237.485 ;
        RECT 12.76 237.155 13.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -0.845 13.085 -0.515 ;
        RECT 12.755 -2.205 13.085 -1.875 ;
        RECT 12.755 -3.565 13.085 -3.235 ;
        RECT 12.76 -3.565 13.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -123.245 13.085 -122.915 ;
        RECT 12.755 -124.605 13.085 -124.275 ;
        RECT 12.755 -125.965 13.085 -125.635 ;
        RECT 12.755 -127.325 13.085 -126.995 ;
        RECT 12.755 -128.685 13.085 -128.355 ;
        RECT 12.755 -130.045 13.085 -129.715 ;
        RECT 12.755 -131.405 13.085 -131.075 ;
        RECT 12.755 -132.765 13.085 -132.435 ;
        RECT 12.755 -134.125 13.085 -133.795 ;
        RECT 12.755 -135.485 13.085 -135.155 ;
        RECT 12.755 -136.845 13.085 -136.515 ;
        RECT 12.755 -138.205 13.085 -137.875 ;
        RECT 12.755 -139.565 13.085 -139.235 ;
        RECT 12.755 -140.925 13.085 -140.595 ;
        RECT 12.755 -142.285 13.085 -141.955 ;
        RECT 12.755 -143.645 13.085 -143.315 ;
        RECT 12.755 -145.005 13.085 -144.675 ;
        RECT 12.755 -146.365 13.085 -146.035 ;
        RECT 12.755 -147.725 13.085 -147.395 ;
        RECT 12.755 -149.085 13.085 -148.755 ;
        RECT 12.755 -150.445 13.085 -150.115 ;
        RECT 12.755 -151.805 13.085 -151.475 ;
        RECT 12.755 -153.165 13.085 -152.835 ;
        RECT 12.755 -154.525 13.085 -154.195 ;
        RECT 12.755 -155.885 13.085 -155.555 ;
        RECT 12.755 -157.245 13.085 -156.915 ;
        RECT 12.755 -158.605 13.085 -158.275 ;
        RECT 12.755 -159.965 13.085 -159.635 ;
        RECT 12.755 -161.325 13.085 -160.995 ;
        RECT 12.755 -162.685 13.085 -162.355 ;
        RECT 12.755 -164.045 13.085 -163.715 ;
        RECT 12.755 -165.405 13.085 -165.075 ;
        RECT 12.755 -166.765 13.085 -166.435 ;
        RECT 12.755 -168.125 13.085 -167.795 ;
        RECT 12.755 -169.485 13.085 -169.155 ;
        RECT 12.755 -170.845 13.085 -170.515 ;
        RECT 12.755 -172.205 13.085 -171.875 ;
        RECT 12.755 -173.565 13.085 -173.235 ;
        RECT 12.755 -174.925 13.085 -174.595 ;
        RECT 12.755 -176.285 13.085 -175.955 ;
        RECT 12.755 -177.645 13.085 -177.315 ;
        RECT 12.755 -179.005 13.085 -178.675 ;
        RECT 12.755 -180.365 13.085 -180.035 ;
        RECT 12.755 -181.725 13.085 -181.395 ;
        RECT 12.755 -183.085 13.085 -182.755 ;
        RECT 12.755 -184.445 13.085 -184.115 ;
        RECT 12.755 -185.805 13.085 -185.475 ;
        RECT 12.755 -187.165 13.085 -186.835 ;
        RECT 12.755 -188.525 13.085 -188.195 ;
        RECT 12.755 -189.885 13.085 -189.555 ;
        RECT 12.755 -191.245 13.085 -190.915 ;
        RECT 12.755 -192.605 13.085 -192.275 ;
        RECT 12.755 -193.965 13.085 -193.635 ;
        RECT 12.755 -195.325 13.085 -194.995 ;
        RECT 12.755 -196.685 13.085 -196.355 ;
        RECT 12.755 -198.045 13.085 -197.715 ;
        RECT 12.755 -199.405 13.085 -199.075 ;
        RECT 12.755 -200.765 13.085 -200.435 ;
        RECT 12.755 -202.125 13.085 -201.795 ;
        RECT 12.755 -203.485 13.085 -203.155 ;
        RECT 12.755 -204.845 13.085 -204.515 ;
        RECT 12.755 -206.205 13.085 -205.875 ;
        RECT 12.755 -207.565 13.085 -207.235 ;
        RECT 12.755 -208.925 13.085 -208.595 ;
        RECT 12.755 -210.285 13.085 -209.955 ;
        RECT 12.755 -211.645 13.085 -211.315 ;
        RECT 12.755 -213.005 13.085 -212.675 ;
        RECT 12.755 -214.365 13.085 -214.035 ;
        RECT 12.755 -215.725 13.085 -215.395 ;
        RECT 12.755 -217.085 13.085 -216.755 ;
        RECT 12.755 -218.445 13.085 -218.115 ;
        RECT 12.755 -219.805 13.085 -219.475 ;
        RECT 12.755 -221.165 13.085 -220.835 ;
        RECT 12.755 -222.525 13.085 -222.195 ;
        RECT 12.755 -223.885 13.085 -223.555 ;
        RECT 12.755 -225.245 13.085 -224.915 ;
        RECT 12.755 -226.605 13.085 -226.275 ;
        RECT 12.755 -227.965 13.085 -227.635 ;
        RECT 12.755 -229.325 13.085 -228.995 ;
        RECT 12.755 -230.685 13.085 -230.355 ;
        RECT 12.755 -232.045 13.085 -231.715 ;
        RECT 12.755 -233.405 13.085 -233.075 ;
        RECT 12.755 -234.765 13.085 -234.435 ;
        RECT 12.755 -236.125 13.085 -235.795 ;
        RECT 12.755 -237.485 13.085 -237.155 ;
        RECT 12.755 -238.845 13.085 -238.515 ;
        RECT 12.755 -241.09 13.085 -239.96 ;
        RECT 12.76 -241.205 13.08 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 244.04 14.445 245.17 ;
        RECT 14.115 242.595 14.445 242.925 ;
        RECT 14.115 241.235 14.445 241.565 ;
        RECT 14.115 239.875 14.445 240.205 ;
        RECT 14.115 238.515 14.445 238.845 ;
        RECT 14.115 237.155 14.445 237.485 ;
        RECT 14.12 237.155 14.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -127.325 14.445 -126.995 ;
        RECT 14.115 -128.685 14.445 -128.355 ;
        RECT 14.115 -130.045 14.445 -129.715 ;
        RECT 14.115 -131.405 14.445 -131.075 ;
        RECT 14.115 -132.765 14.445 -132.435 ;
        RECT 14.115 -134.125 14.445 -133.795 ;
        RECT 14.115 -135.485 14.445 -135.155 ;
        RECT 14.115 -136.845 14.445 -136.515 ;
        RECT 14.115 -138.205 14.445 -137.875 ;
        RECT 14.115 -139.565 14.445 -139.235 ;
        RECT 14.115 -140.925 14.445 -140.595 ;
        RECT 14.115 -142.285 14.445 -141.955 ;
        RECT 14.115 -143.645 14.445 -143.315 ;
        RECT 14.115 -145.005 14.445 -144.675 ;
        RECT 14.115 -146.365 14.445 -146.035 ;
        RECT 14.115 -147.725 14.445 -147.395 ;
        RECT 14.115 -149.085 14.445 -148.755 ;
        RECT 14.115 -150.445 14.445 -150.115 ;
        RECT 14.115 -151.805 14.445 -151.475 ;
        RECT 14.115 -153.165 14.445 -152.835 ;
        RECT 14.115 -154.525 14.445 -154.195 ;
        RECT 14.115 -155.885 14.445 -155.555 ;
        RECT 14.115 -157.245 14.445 -156.915 ;
        RECT 14.115 -158.605 14.445 -158.275 ;
        RECT 14.115 -159.965 14.445 -159.635 ;
        RECT 14.115 -161.325 14.445 -160.995 ;
        RECT 14.115 -162.685 14.445 -162.355 ;
        RECT 14.115 -164.045 14.445 -163.715 ;
        RECT 14.115 -165.405 14.445 -165.075 ;
        RECT 14.115 -166.765 14.445 -166.435 ;
        RECT 14.115 -168.125 14.445 -167.795 ;
        RECT 14.115 -169.485 14.445 -169.155 ;
        RECT 14.115 -170.845 14.445 -170.515 ;
        RECT 14.115 -172.205 14.445 -171.875 ;
        RECT 14.115 -173.565 14.445 -173.235 ;
        RECT 14.115 -174.925 14.445 -174.595 ;
        RECT 14.115 -176.285 14.445 -175.955 ;
        RECT 14.115 -177.645 14.445 -177.315 ;
        RECT 14.115 -179.005 14.445 -178.675 ;
        RECT 14.115 -180.365 14.445 -180.035 ;
        RECT 14.115 -181.725 14.445 -181.395 ;
        RECT 14.115 -183.085 14.445 -182.755 ;
        RECT 14.115 -184.445 14.445 -184.115 ;
        RECT 14.115 -185.805 14.445 -185.475 ;
        RECT 14.115 -187.165 14.445 -186.835 ;
        RECT 14.115 -188.525 14.445 -188.195 ;
        RECT 14.115 -189.885 14.445 -189.555 ;
        RECT 14.115 -191.245 14.445 -190.915 ;
        RECT 14.115 -192.605 14.445 -192.275 ;
        RECT 14.115 -193.965 14.445 -193.635 ;
        RECT 14.115 -195.325 14.445 -194.995 ;
        RECT 14.115 -196.685 14.445 -196.355 ;
        RECT 14.115 -198.045 14.445 -197.715 ;
        RECT 14.115 -199.405 14.445 -199.075 ;
        RECT 14.115 -200.765 14.445 -200.435 ;
        RECT 14.115 -202.125 14.445 -201.795 ;
        RECT 14.115 -203.485 14.445 -203.155 ;
        RECT 14.115 -204.845 14.445 -204.515 ;
        RECT 14.115 -206.205 14.445 -205.875 ;
        RECT 14.115 -207.565 14.445 -207.235 ;
        RECT 14.115 -208.925 14.445 -208.595 ;
        RECT 14.115 -210.285 14.445 -209.955 ;
        RECT 14.115 -211.645 14.445 -211.315 ;
        RECT 14.115 -213.005 14.445 -212.675 ;
        RECT 14.115 -214.365 14.445 -214.035 ;
        RECT 14.115 -215.725 14.445 -215.395 ;
        RECT 14.115 -217.085 14.445 -216.755 ;
        RECT 14.115 -218.445 14.445 -218.115 ;
        RECT 14.115 -219.805 14.445 -219.475 ;
        RECT 14.115 -221.165 14.445 -220.835 ;
        RECT 14.115 -222.525 14.445 -222.195 ;
        RECT 14.115 -223.885 14.445 -223.555 ;
        RECT 14.115 -225.245 14.445 -224.915 ;
        RECT 14.115 -226.605 14.445 -226.275 ;
        RECT 14.115 -227.965 14.445 -227.635 ;
        RECT 14.115 -229.325 14.445 -228.995 ;
        RECT 14.115 -230.685 14.445 -230.355 ;
        RECT 14.115 -232.045 14.445 -231.715 ;
        RECT 14.115 -233.405 14.445 -233.075 ;
        RECT 14.115 -234.765 14.445 -234.435 ;
        RECT 14.115 -236.125 14.445 -235.795 ;
        RECT 14.115 -237.485 14.445 -237.155 ;
        RECT 14.115 -238.845 14.445 -238.515 ;
        RECT 14.115 -241.09 14.445 -239.96 ;
        RECT 14.12 -241.205 14.44 -126.32 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.21 -125.535 14.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 244.04 15.805 245.17 ;
        RECT 15.475 242.595 15.805 242.925 ;
        RECT 15.475 241.235 15.805 241.565 ;
        RECT 15.475 239.875 15.805 240.205 ;
        RECT 15.475 238.515 15.805 238.845 ;
        RECT 15.475 237.155 15.805 237.485 ;
        RECT 15.48 237.155 15.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 -0.845 15.805 -0.515 ;
        RECT 15.475 -2.205 15.805 -1.875 ;
        RECT 15.475 -3.565 15.805 -3.235 ;
        RECT 15.48 -3.565 15.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 244.04 17.165 245.17 ;
        RECT 16.835 242.595 17.165 242.925 ;
        RECT 16.835 241.235 17.165 241.565 ;
        RECT 16.835 239.875 17.165 240.205 ;
        RECT 16.835 238.515 17.165 238.845 ;
        RECT 16.835 237.155 17.165 237.485 ;
        RECT 16.84 237.155 17.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 -0.845 17.165 -0.515 ;
        RECT 16.835 -2.205 17.165 -1.875 ;
        RECT 16.835 -3.565 17.165 -3.235 ;
        RECT 16.84 -3.565 17.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 244.04 18.525 245.17 ;
        RECT 18.195 242.595 18.525 242.925 ;
        RECT 18.195 241.235 18.525 241.565 ;
        RECT 18.195 239.875 18.525 240.205 ;
        RECT 18.195 238.515 18.525 238.845 ;
        RECT 18.195 237.155 18.525 237.485 ;
        RECT 18.2 237.155 18.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 -0.845 18.525 -0.515 ;
        RECT 18.195 -2.205 18.525 -1.875 ;
        RECT 18.195 -3.565 18.525 -3.235 ;
        RECT 18.2 -3.565 18.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 -123.245 18.525 -122.915 ;
        RECT 18.195 -124.605 18.525 -124.275 ;
        RECT 18.195 -125.965 18.525 -125.635 ;
        RECT 18.195 -127.325 18.525 -126.995 ;
        RECT 18.195 -128.685 18.525 -128.355 ;
        RECT 18.195 -130.045 18.525 -129.715 ;
        RECT 18.195 -131.405 18.525 -131.075 ;
        RECT 18.195 -132.765 18.525 -132.435 ;
        RECT 18.195 -134.125 18.525 -133.795 ;
        RECT 18.195 -135.485 18.525 -135.155 ;
        RECT 18.195 -136.845 18.525 -136.515 ;
        RECT 18.195 -138.205 18.525 -137.875 ;
        RECT 18.195 -139.565 18.525 -139.235 ;
        RECT 18.195 -140.925 18.525 -140.595 ;
        RECT 18.195 -142.285 18.525 -141.955 ;
        RECT 18.195 -143.645 18.525 -143.315 ;
        RECT 18.195 -145.005 18.525 -144.675 ;
        RECT 18.195 -146.365 18.525 -146.035 ;
        RECT 18.195 -147.725 18.525 -147.395 ;
        RECT 18.195 -149.085 18.525 -148.755 ;
        RECT 18.195 -150.445 18.525 -150.115 ;
        RECT 18.195 -151.805 18.525 -151.475 ;
        RECT 18.195 -153.165 18.525 -152.835 ;
        RECT 18.195 -154.525 18.525 -154.195 ;
        RECT 18.195 -155.885 18.525 -155.555 ;
        RECT 18.195 -157.245 18.525 -156.915 ;
        RECT 18.195 -158.605 18.525 -158.275 ;
        RECT 18.195 -159.965 18.525 -159.635 ;
        RECT 18.195 -161.325 18.525 -160.995 ;
        RECT 18.195 -162.685 18.525 -162.355 ;
        RECT 18.195 -164.045 18.525 -163.715 ;
        RECT 18.195 -165.405 18.525 -165.075 ;
        RECT 18.195 -166.765 18.525 -166.435 ;
        RECT 18.195 -168.125 18.525 -167.795 ;
        RECT 18.195 -169.485 18.525 -169.155 ;
        RECT 18.195 -170.845 18.525 -170.515 ;
        RECT 18.195 -172.205 18.525 -171.875 ;
        RECT 18.195 -173.565 18.525 -173.235 ;
        RECT 18.195 -174.925 18.525 -174.595 ;
        RECT 18.195 -176.285 18.525 -175.955 ;
        RECT 18.195 -177.645 18.525 -177.315 ;
        RECT 18.195 -179.005 18.525 -178.675 ;
        RECT 18.195 -180.365 18.525 -180.035 ;
        RECT 18.195 -181.725 18.525 -181.395 ;
        RECT 18.195 -183.085 18.525 -182.755 ;
        RECT 18.195 -184.445 18.525 -184.115 ;
        RECT 18.195 -185.805 18.525 -185.475 ;
        RECT 18.195 -187.165 18.525 -186.835 ;
        RECT 18.195 -188.525 18.525 -188.195 ;
        RECT 18.195 -189.885 18.525 -189.555 ;
        RECT 18.195 -191.245 18.525 -190.915 ;
        RECT 18.195 -192.605 18.525 -192.275 ;
        RECT 18.195 -193.965 18.525 -193.635 ;
        RECT 18.195 -195.325 18.525 -194.995 ;
        RECT 18.195 -196.685 18.525 -196.355 ;
        RECT 18.195 -198.045 18.525 -197.715 ;
        RECT 18.195 -199.405 18.525 -199.075 ;
        RECT 18.195 -200.765 18.525 -200.435 ;
        RECT 18.195 -202.125 18.525 -201.795 ;
        RECT 18.195 -203.485 18.525 -203.155 ;
        RECT 18.195 -204.845 18.525 -204.515 ;
        RECT 18.195 -206.205 18.525 -205.875 ;
        RECT 18.195 -207.565 18.525 -207.235 ;
        RECT 18.195 -208.925 18.525 -208.595 ;
        RECT 18.195 -210.285 18.525 -209.955 ;
        RECT 18.195 -211.645 18.525 -211.315 ;
        RECT 18.195 -213.005 18.525 -212.675 ;
        RECT 18.195 -214.365 18.525 -214.035 ;
        RECT 18.195 -215.725 18.525 -215.395 ;
        RECT 18.195 -217.085 18.525 -216.755 ;
        RECT 18.195 -218.445 18.525 -218.115 ;
        RECT 18.195 -219.805 18.525 -219.475 ;
        RECT 18.195 -221.165 18.525 -220.835 ;
        RECT 18.195 -222.525 18.525 -222.195 ;
        RECT 18.195 -223.885 18.525 -223.555 ;
        RECT 18.195 -225.245 18.525 -224.915 ;
        RECT 18.195 -226.605 18.525 -226.275 ;
        RECT 18.195 -227.965 18.525 -227.635 ;
        RECT 18.195 -229.325 18.525 -228.995 ;
        RECT 18.195 -230.685 18.525 -230.355 ;
        RECT 18.195 -232.045 18.525 -231.715 ;
        RECT 18.195 -233.405 18.525 -233.075 ;
        RECT 18.195 -234.765 18.525 -234.435 ;
        RECT 18.195 -236.125 18.525 -235.795 ;
        RECT 18.195 -237.485 18.525 -237.155 ;
        RECT 18.195 -238.845 18.525 -238.515 ;
        RECT 18.195 -241.09 18.525 -239.96 ;
        RECT 18.2 -241.205 18.52 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 244.04 19.885 245.17 ;
        RECT 19.555 242.595 19.885 242.925 ;
        RECT 19.555 241.235 19.885 241.565 ;
        RECT 19.555 239.875 19.885 240.205 ;
        RECT 19.555 238.515 19.885 238.845 ;
        RECT 19.555 237.155 19.885 237.485 ;
        RECT 19.56 237.155 19.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -0.845 19.885 -0.515 ;
        RECT 19.555 -2.205 19.885 -1.875 ;
        RECT 19.555 -3.565 19.885 -3.235 ;
        RECT 19.56 -3.565 19.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -123.245 19.885 -122.915 ;
        RECT 19.555 -124.605 19.885 -124.275 ;
        RECT 19.555 -125.965 19.885 -125.635 ;
        RECT 19.555 -127.325 19.885 -126.995 ;
        RECT 19.555 -128.685 19.885 -128.355 ;
        RECT 19.555 -130.045 19.885 -129.715 ;
        RECT 19.555 -131.405 19.885 -131.075 ;
        RECT 19.555 -132.765 19.885 -132.435 ;
        RECT 19.555 -134.125 19.885 -133.795 ;
        RECT 19.555 -135.485 19.885 -135.155 ;
        RECT 19.555 -136.845 19.885 -136.515 ;
        RECT 19.555 -138.205 19.885 -137.875 ;
        RECT 19.555 -139.565 19.885 -139.235 ;
        RECT 19.555 -140.925 19.885 -140.595 ;
        RECT 19.555 -142.285 19.885 -141.955 ;
        RECT 19.555 -143.645 19.885 -143.315 ;
        RECT 19.555 -145.005 19.885 -144.675 ;
        RECT 19.555 -146.365 19.885 -146.035 ;
        RECT 19.555 -147.725 19.885 -147.395 ;
        RECT 19.555 -149.085 19.885 -148.755 ;
        RECT 19.555 -150.445 19.885 -150.115 ;
        RECT 19.555 -151.805 19.885 -151.475 ;
        RECT 19.555 -153.165 19.885 -152.835 ;
        RECT 19.555 -154.525 19.885 -154.195 ;
        RECT 19.555 -155.885 19.885 -155.555 ;
        RECT 19.555 -157.245 19.885 -156.915 ;
        RECT 19.555 -158.605 19.885 -158.275 ;
        RECT 19.555 -159.965 19.885 -159.635 ;
        RECT 19.555 -161.325 19.885 -160.995 ;
        RECT 19.555 -162.685 19.885 -162.355 ;
        RECT 19.555 -164.045 19.885 -163.715 ;
        RECT 19.555 -165.405 19.885 -165.075 ;
        RECT 19.555 -166.765 19.885 -166.435 ;
        RECT 19.555 -168.125 19.885 -167.795 ;
        RECT 19.555 -169.485 19.885 -169.155 ;
        RECT 19.555 -170.845 19.885 -170.515 ;
        RECT 19.555 -172.205 19.885 -171.875 ;
        RECT 19.555 -173.565 19.885 -173.235 ;
        RECT 19.555 -174.925 19.885 -174.595 ;
        RECT 19.555 -176.285 19.885 -175.955 ;
        RECT 19.555 -177.645 19.885 -177.315 ;
        RECT 19.555 -179.005 19.885 -178.675 ;
        RECT 19.555 -180.365 19.885 -180.035 ;
        RECT 19.555 -181.725 19.885 -181.395 ;
        RECT 19.555 -183.085 19.885 -182.755 ;
        RECT 19.555 -184.445 19.885 -184.115 ;
        RECT 19.555 -185.805 19.885 -185.475 ;
        RECT 19.555 -187.165 19.885 -186.835 ;
        RECT 19.555 -188.525 19.885 -188.195 ;
        RECT 19.555 -189.885 19.885 -189.555 ;
        RECT 19.555 -191.245 19.885 -190.915 ;
        RECT 19.555 -192.605 19.885 -192.275 ;
        RECT 19.555 -193.965 19.885 -193.635 ;
        RECT 19.555 -195.325 19.885 -194.995 ;
        RECT 19.555 -196.685 19.885 -196.355 ;
        RECT 19.555 -198.045 19.885 -197.715 ;
        RECT 19.555 -199.405 19.885 -199.075 ;
        RECT 19.555 -200.765 19.885 -200.435 ;
        RECT 19.555 -202.125 19.885 -201.795 ;
        RECT 19.555 -203.485 19.885 -203.155 ;
        RECT 19.555 -204.845 19.885 -204.515 ;
        RECT 19.555 -206.205 19.885 -205.875 ;
        RECT 19.555 -207.565 19.885 -207.235 ;
        RECT 19.555 -208.925 19.885 -208.595 ;
        RECT 19.555 -210.285 19.885 -209.955 ;
        RECT 19.555 -211.645 19.885 -211.315 ;
        RECT 19.555 -213.005 19.885 -212.675 ;
        RECT 19.555 -214.365 19.885 -214.035 ;
        RECT 19.555 -215.725 19.885 -215.395 ;
        RECT 19.555 -217.085 19.885 -216.755 ;
        RECT 19.555 -218.445 19.885 -218.115 ;
        RECT 19.555 -219.805 19.885 -219.475 ;
        RECT 19.555 -221.165 19.885 -220.835 ;
        RECT 19.555 -222.525 19.885 -222.195 ;
        RECT 19.555 -223.885 19.885 -223.555 ;
        RECT 19.555 -225.245 19.885 -224.915 ;
        RECT 19.555 -226.605 19.885 -226.275 ;
        RECT 19.555 -227.965 19.885 -227.635 ;
        RECT 19.555 -229.325 19.885 -228.995 ;
        RECT 19.555 -230.685 19.885 -230.355 ;
        RECT 19.555 -232.045 19.885 -231.715 ;
        RECT 19.555 -233.405 19.885 -233.075 ;
        RECT 19.555 -234.765 19.885 -234.435 ;
        RECT 19.555 -236.125 19.885 -235.795 ;
        RECT 19.555 -237.485 19.885 -237.155 ;
        RECT 19.555 -238.845 19.885 -238.515 ;
        RECT 19.555 -241.09 19.885 -239.96 ;
        RECT 19.56 -241.205 19.88 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 244.04 21.245 245.17 ;
        RECT 20.915 242.595 21.245 242.925 ;
        RECT 20.915 241.235 21.245 241.565 ;
        RECT 20.915 239.875 21.245 240.205 ;
        RECT 20.915 238.515 21.245 238.845 ;
        RECT 20.915 237.155 21.245 237.485 ;
        RECT 20.92 237.155 21.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 -0.845 21.245 -0.515 ;
        RECT 20.915 -2.205 21.245 -1.875 ;
        RECT 20.915 -3.565 21.245 -3.235 ;
        RECT 20.92 -3.565 21.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 -123.245 21.245 -122.915 ;
        RECT 20.915 -124.605 21.245 -124.275 ;
        RECT 20.915 -125.965 21.245 -125.635 ;
        RECT 20.915 -127.325 21.245 -126.995 ;
        RECT 20.915 -128.685 21.245 -128.355 ;
        RECT 20.915 -130.045 21.245 -129.715 ;
        RECT 20.915 -131.405 21.245 -131.075 ;
        RECT 20.915 -132.765 21.245 -132.435 ;
        RECT 20.915 -134.125 21.245 -133.795 ;
        RECT 20.915 -135.485 21.245 -135.155 ;
        RECT 20.915 -136.845 21.245 -136.515 ;
        RECT 20.915 -138.205 21.245 -137.875 ;
        RECT 20.915 -139.565 21.245 -139.235 ;
        RECT 20.915 -140.925 21.245 -140.595 ;
        RECT 20.915 -142.285 21.245 -141.955 ;
        RECT 20.915 -143.645 21.245 -143.315 ;
        RECT 20.915 -145.005 21.245 -144.675 ;
        RECT 20.915 -146.365 21.245 -146.035 ;
        RECT 20.915 -147.725 21.245 -147.395 ;
        RECT 20.915 -149.085 21.245 -148.755 ;
        RECT 20.915 -150.445 21.245 -150.115 ;
        RECT 20.915 -151.805 21.245 -151.475 ;
        RECT 20.915 -153.165 21.245 -152.835 ;
        RECT 20.915 -154.525 21.245 -154.195 ;
        RECT 20.915 -155.885 21.245 -155.555 ;
        RECT 20.915 -157.245 21.245 -156.915 ;
        RECT 20.915 -158.605 21.245 -158.275 ;
        RECT 20.915 -159.965 21.245 -159.635 ;
        RECT 20.915 -161.325 21.245 -160.995 ;
        RECT 20.915 -162.685 21.245 -162.355 ;
        RECT 20.915 -164.045 21.245 -163.715 ;
        RECT 20.915 -165.405 21.245 -165.075 ;
        RECT 20.915 -166.765 21.245 -166.435 ;
        RECT 20.915 -168.125 21.245 -167.795 ;
        RECT 20.915 -169.485 21.245 -169.155 ;
        RECT 20.915 -170.845 21.245 -170.515 ;
        RECT 20.915 -172.205 21.245 -171.875 ;
        RECT 20.915 -173.565 21.245 -173.235 ;
        RECT 20.915 -174.925 21.245 -174.595 ;
        RECT 20.915 -176.285 21.245 -175.955 ;
        RECT 20.915 -177.645 21.245 -177.315 ;
        RECT 20.915 -179.005 21.245 -178.675 ;
        RECT 20.915 -180.365 21.245 -180.035 ;
        RECT 20.915 -181.725 21.245 -181.395 ;
        RECT 20.915 -183.085 21.245 -182.755 ;
        RECT 20.915 -184.445 21.245 -184.115 ;
        RECT 20.915 -185.805 21.245 -185.475 ;
        RECT 20.915 -187.165 21.245 -186.835 ;
        RECT 20.915 -188.525 21.245 -188.195 ;
        RECT 20.915 -189.885 21.245 -189.555 ;
        RECT 20.915 -191.245 21.245 -190.915 ;
        RECT 20.915 -192.605 21.245 -192.275 ;
        RECT 20.915 -193.965 21.245 -193.635 ;
        RECT 20.915 -195.325 21.245 -194.995 ;
        RECT 20.915 -196.685 21.245 -196.355 ;
        RECT 20.915 -198.045 21.245 -197.715 ;
        RECT 20.915 -199.405 21.245 -199.075 ;
        RECT 20.915 -200.765 21.245 -200.435 ;
        RECT 20.915 -202.125 21.245 -201.795 ;
        RECT 20.915 -203.485 21.245 -203.155 ;
        RECT 20.915 -204.845 21.245 -204.515 ;
        RECT 20.915 -206.205 21.245 -205.875 ;
        RECT 20.915 -207.565 21.245 -207.235 ;
        RECT 20.915 -208.925 21.245 -208.595 ;
        RECT 20.915 -210.285 21.245 -209.955 ;
        RECT 20.915 -211.645 21.245 -211.315 ;
        RECT 20.915 -213.005 21.245 -212.675 ;
        RECT 20.915 -214.365 21.245 -214.035 ;
        RECT 20.915 -215.725 21.245 -215.395 ;
        RECT 20.915 -217.085 21.245 -216.755 ;
        RECT 20.915 -218.445 21.245 -218.115 ;
        RECT 20.915 -219.805 21.245 -219.475 ;
        RECT 20.915 -221.165 21.245 -220.835 ;
        RECT 20.915 -222.525 21.245 -222.195 ;
        RECT 20.915 -223.885 21.245 -223.555 ;
        RECT 20.915 -225.245 21.245 -224.915 ;
        RECT 20.915 -226.605 21.245 -226.275 ;
        RECT 20.915 -227.965 21.245 -227.635 ;
        RECT 20.915 -229.325 21.245 -228.995 ;
        RECT 20.915 -230.685 21.245 -230.355 ;
        RECT 20.915 -232.045 21.245 -231.715 ;
        RECT 20.915 -233.405 21.245 -233.075 ;
        RECT 20.915 -234.765 21.245 -234.435 ;
        RECT 20.915 -236.125 21.245 -235.795 ;
        RECT 20.915 -237.485 21.245 -237.155 ;
        RECT 20.915 -238.845 21.245 -238.515 ;
        RECT 20.915 -241.09 21.245 -239.96 ;
        RECT 20.92 -241.205 21.24 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 244.04 22.605 245.17 ;
        RECT 22.275 242.595 22.605 242.925 ;
        RECT 22.275 241.235 22.605 241.565 ;
        RECT 22.275 239.875 22.605 240.205 ;
        RECT 22.275 238.515 22.605 238.845 ;
        RECT 22.275 237.155 22.605 237.485 ;
        RECT 22.28 237.155 22.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 -2.205 22.605 -1.875 ;
        RECT 22.275 -3.565 22.605 -3.235 ;
        RECT 22.28 -3.565 22.6 -0.515 ;
        RECT 22.275 -0.845 22.605 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.565 -140.925 -3.235 -140.595 ;
        RECT -3.565 -142.285 -3.235 -141.955 ;
        RECT -3.565 -143.645 -3.235 -143.315 ;
        RECT -3.565 -145.005 -3.235 -144.675 ;
        RECT -3.565 -146.365 -3.235 -146.035 ;
        RECT -3.565 -147.725 -3.235 -147.395 ;
        RECT -3.565 -149.085 -3.235 -148.755 ;
        RECT -3.565 -150.445 -3.235 -150.115 ;
        RECT -3.565 -151.805 -3.235 -151.475 ;
        RECT -3.565 -153.165 -3.235 -152.835 ;
        RECT -3.565 -154.525 -3.235 -154.195 ;
        RECT -3.565 -155.885 -3.235 -155.555 ;
        RECT -3.565 -157.245 -3.235 -156.915 ;
        RECT -3.565 -158.605 -3.235 -158.275 ;
        RECT -3.565 -159.965 -3.235 -159.635 ;
        RECT -3.565 -161.325 -3.235 -160.995 ;
        RECT -3.565 -162.685 -3.235 -162.355 ;
        RECT -3.565 -164.045 -3.235 -163.715 ;
        RECT -3.565 -165.405 -3.235 -165.075 ;
        RECT -3.565 -166.765 -3.235 -166.435 ;
        RECT -3.565 -168.125 -3.235 -167.795 ;
        RECT -3.565 -169.485 -3.235 -169.155 ;
        RECT -3.565 -170.845 -3.235 -170.515 ;
        RECT -3.565 -172.205 -3.235 -171.875 ;
        RECT -3.565 -173.565 -3.235 -173.235 ;
        RECT -3.565 -174.925 -3.235 -174.595 ;
        RECT -3.565 -176.285 -3.235 -175.955 ;
        RECT -3.565 -177.645 -3.235 -177.315 ;
        RECT -3.565 -179.005 -3.235 -178.675 ;
        RECT -3.565 -180.365 -3.235 -180.035 ;
        RECT -3.565 -181.725 -3.235 -181.395 ;
        RECT -3.565 -183.085 -3.235 -182.755 ;
        RECT -3.565 -184.445 -3.235 -184.115 ;
        RECT -3.565 -185.805 -3.235 -185.475 ;
        RECT -3.565 -187.165 -3.235 -186.835 ;
        RECT -3.565 -188.525 -3.235 -188.195 ;
        RECT -3.565 -189.885 -3.235 -189.555 ;
        RECT -3.565 -191.245 -3.235 -190.915 ;
        RECT -3.565 -192.605 -3.235 -192.275 ;
        RECT -3.565 -193.965 -3.235 -193.635 ;
        RECT -3.565 -195.325 -3.235 -194.995 ;
        RECT -3.565 -196.685 -3.235 -196.355 ;
        RECT -3.565 -198.045 -3.235 -197.715 ;
        RECT -3.565 -199.405 -3.235 -199.075 ;
        RECT -3.565 -200.765 -3.235 -200.435 ;
        RECT -3.565 -202.125 -3.235 -201.795 ;
        RECT -3.565 -203.485 -3.235 -203.155 ;
        RECT -3.565 -204.845 -3.235 -204.515 ;
        RECT -3.565 -206.205 -3.235 -205.875 ;
        RECT -3.565 -207.565 -3.235 -207.235 ;
        RECT -3.565 -208.925 -3.235 -208.595 ;
        RECT -3.565 -210.285 -3.235 -209.955 ;
        RECT -3.565 -211.645 -3.235 -211.315 ;
        RECT -3.565 -213.005 -3.235 -212.675 ;
        RECT -3.565 -214.365 -3.235 -214.035 ;
        RECT -3.565 -215.725 -3.235 -215.395 ;
        RECT -3.565 -217.085 -3.235 -216.755 ;
        RECT -3.565 -218.445 -3.235 -218.115 ;
        RECT -3.565 -219.805 -3.235 -219.475 ;
        RECT -3.565 -221.165 -3.235 -220.835 ;
        RECT -3.565 -222.525 -3.235 -222.195 ;
        RECT -3.565 -223.885 -3.235 -223.555 ;
        RECT -3.565 -225.245 -3.235 -224.915 ;
        RECT -3.565 -226.605 -3.235 -226.275 ;
        RECT -3.565 -227.965 -3.235 -227.635 ;
        RECT -3.565 -229.325 -3.235 -228.995 ;
        RECT -3.565 -230.685 -3.235 -230.355 ;
        RECT -3.565 -232.045 -3.235 -231.715 ;
        RECT -3.565 -233.405 -3.235 -233.075 ;
        RECT -3.565 -234.765 -3.235 -234.435 ;
        RECT -3.565 -236.125 -3.235 -235.795 ;
        RECT -3.565 -237.485 -3.235 -237.155 ;
        RECT -3.565 -238.845 -3.235 -238.515 ;
        RECT -3.565 -241.09 -3.235 -239.96 ;
        RECT -3.56 -241.205 -3.24 -139.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 244.04 -1.875 245.17 ;
        RECT -2.205 242.595 -1.875 242.925 ;
        RECT -2.205 241.235 -1.875 241.565 ;
        RECT -2.205 239.875 -1.875 240.205 ;
        RECT -2.205 238.515 -1.875 238.845 ;
        RECT -2.205 237.155 -1.875 237.485 ;
        RECT -2.205 235.975 -1.875 236.305 ;
        RECT -2.205 233.925 -1.875 234.255 ;
        RECT -2.205 231.995 -1.875 232.325 ;
        RECT -2.205 230.155 -1.875 230.485 ;
        RECT -2.205 228.665 -1.875 228.995 ;
        RECT -2.205 226.995 -1.875 227.325 ;
        RECT -2.205 225.505 -1.875 225.835 ;
        RECT -2.205 223.835 -1.875 224.165 ;
        RECT -2.205 222.345 -1.875 222.675 ;
        RECT -2.205 220.675 -1.875 221.005 ;
        RECT -2.205 219.185 -1.875 219.515 ;
        RECT -2.205 217.775 -1.875 218.105 ;
        RECT -2.205 215.935 -1.875 216.265 ;
        RECT -2.205 214.445 -1.875 214.775 ;
        RECT -2.205 212.775 -1.875 213.105 ;
        RECT -2.205 211.285 -1.875 211.615 ;
        RECT -2.205 209.615 -1.875 209.945 ;
        RECT -2.205 208.125 -1.875 208.455 ;
        RECT -2.205 206.455 -1.875 206.785 ;
        RECT -2.205 204.965 -1.875 205.295 ;
        RECT -2.205 203.555 -1.875 203.885 ;
        RECT -2.205 201.715 -1.875 202.045 ;
        RECT -2.205 200.225 -1.875 200.555 ;
        RECT -2.205 198.555 -1.875 198.885 ;
        RECT -2.205 197.065 -1.875 197.395 ;
        RECT -2.205 195.395 -1.875 195.725 ;
        RECT -2.205 193.905 -1.875 194.235 ;
        RECT -2.205 192.235 -1.875 192.565 ;
        RECT -2.205 190.745 -1.875 191.075 ;
        RECT -2.205 189.335 -1.875 189.665 ;
        RECT -2.205 187.495 -1.875 187.825 ;
        RECT -2.205 186.005 -1.875 186.335 ;
        RECT -2.205 184.335 -1.875 184.665 ;
        RECT -2.205 182.845 -1.875 183.175 ;
        RECT -2.205 181.175 -1.875 181.505 ;
        RECT -2.205 179.685 -1.875 180.015 ;
        RECT -2.205 178.015 -1.875 178.345 ;
        RECT -2.205 176.525 -1.875 176.855 ;
        RECT -2.205 175.115 -1.875 175.445 ;
        RECT -2.205 173.275 -1.875 173.605 ;
        RECT -2.205 171.785 -1.875 172.115 ;
        RECT -2.205 170.115 -1.875 170.445 ;
        RECT -2.205 168.625 -1.875 168.955 ;
        RECT -2.205 166.955 -1.875 167.285 ;
        RECT -2.205 165.465 -1.875 165.795 ;
        RECT -2.205 163.795 -1.875 164.125 ;
        RECT -2.205 162.305 -1.875 162.635 ;
        RECT -2.205 160.895 -1.875 161.225 ;
        RECT -2.205 159.055 -1.875 159.385 ;
        RECT -2.205 157.565 -1.875 157.895 ;
        RECT -2.205 155.895 -1.875 156.225 ;
        RECT -2.205 154.405 -1.875 154.735 ;
        RECT -2.205 152.735 -1.875 153.065 ;
        RECT -2.205 151.245 -1.875 151.575 ;
        RECT -2.205 149.575 -1.875 149.905 ;
        RECT -2.205 148.085 -1.875 148.415 ;
        RECT -2.205 146.675 -1.875 147.005 ;
        RECT -2.205 144.835 -1.875 145.165 ;
        RECT -2.205 143.345 -1.875 143.675 ;
        RECT -2.205 141.675 -1.875 142.005 ;
        RECT -2.205 140.185 -1.875 140.515 ;
        RECT -2.205 138.515 -1.875 138.845 ;
        RECT -2.205 137.025 -1.875 137.355 ;
        RECT -2.205 135.355 -1.875 135.685 ;
        RECT -2.205 133.865 -1.875 134.195 ;
        RECT -2.205 132.455 -1.875 132.785 ;
        RECT -2.205 130.615 -1.875 130.945 ;
        RECT -2.205 129.125 -1.875 129.455 ;
        RECT -2.205 127.455 -1.875 127.785 ;
        RECT -2.205 125.965 -1.875 126.295 ;
        RECT -2.205 124.295 -1.875 124.625 ;
        RECT -2.205 122.805 -1.875 123.135 ;
        RECT -2.205 121.135 -1.875 121.465 ;
        RECT -2.205 119.645 -1.875 119.975 ;
        RECT -2.205 118.235 -1.875 118.565 ;
        RECT -2.205 116.395 -1.875 116.725 ;
        RECT -2.205 114.905 -1.875 115.235 ;
        RECT -2.205 113.235 -1.875 113.565 ;
        RECT -2.205 111.745 -1.875 112.075 ;
        RECT -2.205 110.075 -1.875 110.405 ;
        RECT -2.205 108.585 -1.875 108.915 ;
        RECT -2.205 106.915 -1.875 107.245 ;
        RECT -2.205 105.425 -1.875 105.755 ;
        RECT -2.205 104.015 -1.875 104.345 ;
        RECT -2.205 102.175 -1.875 102.505 ;
        RECT -2.205 100.685 -1.875 101.015 ;
        RECT -2.205 99.015 -1.875 99.345 ;
        RECT -2.205 97.525 -1.875 97.855 ;
        RECT -2.205 95.855 -1.875 96.185 ;
        RECT -2.205 94.365 -1.875 94.695 ;
        RECT -2.205 92.695 -1.875 93.025 ;
        RECT -2.205 91.205 -1.875 91.535 ;
        RECT -2.205 89.795 -1.875 90.125 ;
        RECT -2.205 87.955 -1.875 88.285 ;
        RECT -2.205 86.465 -1.875 86.795 ;
        RECT -2.205 84.795 -1.875 85.125 ;
        RECT -2.205 83.305 -1.875 83.635 ;
        RECT -2.205 81.635 -1.875 81.965 ;
        RECT -2.205 80.145 -1.875 80.475 ;
        RECT -2.205 78.475 -1.875 78.805 ;
        RECT -2.205 76.985 -1.875 77.315 ;
        RECT -2.205 75.575 -1.875 75.905 ;
        RECT -2.205 73.735 -1.875 74.065 ;
        RECT -2.205 72.245 -1.875 72.575 ;
        RECT -2.205 70.575 -1.875 70.905 ;
        RECT -2.205 69.085 -1.875 69.415 ;
        RECT -2.205 67.415 -1.875 67.745 ;
        RECT -2.205 65.925 -1.875 66.255 ;
        RECT -2.205 64.255 -1.875 64.585 ;
        RECT -2.205 62.765 -1.875 63.095 ;
        RECT -2.205 61.355 -1.875 61.685 ;
        RECT -2.205 59.515 -1.875 59.845 ;
        RECT -2.205 58.025 -1.875 58.355 ;
        RECT -2.205 56.355 -1.875 56.685 ;
        RECT -2.205 54.865 -1.875 55.195 ;
        RECT -2.205 53.195 -1.875 53.525 ;
        RECT -2.205 51.705 -1.875 52.035 ;
        RECT -2.205 50.035 -1.875 50.365 ;
        RECT -2.205 48.545 -1.875 48.875 ;
        RECT -2.205 47.135 -1.875 47.465 ;
        RECT -2.205 45.295 -1.875 45.625 ;
        RECT -2.205 43.805 -1.875 44.135 ;
        RECT -2.205 42.135 -1.875 42.465 ;
        RECT -2.205 40.645 -1.875 40.975 ;
        RECT -2.205 38.975 -1.875 39.305 ;
        RECT -2.205 37.485 -1.875 37.815 ;
        RECT -2.205 35.815 -1.875 36.145 ;
        RECT -2.205 34.325 -1.875 34.655 ;
        RECT -2.205 32.915 -1.875 33.245 ;
        RECT -2.205 31.075 -1.875 31.405 ;
        RECT -2.205 29.585 -1.875 29.915 ;
        RECT -2.205 27.915 -1.875 28.245 ;
        RECT -2.205 26.425 -1.875 26.755 ;
        RECT -2.205 24.755 -1.875 25.085 ;
        RECT -2.205 23.265 -1.875 23.595 ;
        RECT -2.205 21.595 -1.875 21.925 ;
        RECT -2.205 20.105 -1.875 20.435 ;
        RECT -2.205 18.695 -1.875 19.025 ;
        RECT -2.205 16.855 -1.875 17.185 ;
        RECT -2.205 15.365 -1.875 15.695 ;
        RECT -2.205 13.695 -1.875 14.025 ;
        RECT -2.205 12.205 -1.875 12.535 ;
        RECT -2.205 10.535 -1.875 10.865 ;
        RECT -2.205 9.045 -1.875 9.375 ;
        RECT -2.205 7.375 -1.875 7.705 ;
        RECT -2.205 5.885 -1.875 6.215 ;
        RECT -2.205 4.475 -1.875 4.805 ;
        RECT -2.205 2.115 -1.875 2.445 ;
        RECT -2.205 0.06 -1.875 0.39 ;
        RECT -2.205 -0.845 -1.875 -0.515 ;
        RECT -2.205 -2.205 -1.875 -1.875 ;
        RECT -2.205 -3.565 -1.875 -3.235 ;
        RECT -2.205 -4.925 -1.875 -4.595 ;
        RECT -2.205 -6.285 -1.875 -5.955 ;
        RECT -2.205 -7.645 -1.875 -7.315 ;
        RECT -2.205 -9.005 -1.875 -8.675 ;
        RECT -2.205 -10.365 -1.875 -10.035 ;
        RECT -2.205 -11.725 -1.875 -11.395 ;
        RECT -2.205 -13.085 -1.875 -12.755 ;
        RECT -2.205 -14.445 -1.875 -14.115 ;
        RECT -2.205 -15.805 -1.875 -15.475 ;
        RECT -2.205 -17.165 -1.875 -16.835 ;
        RECT -2.205 -18.525 -1.875 -18.195 ;
        RECT -2.205 -19.885 -1.875 -19.555 ;
        RECT -2.2 -23.28 -1.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 -138.205 -1.875 -137.875 ;
        RECT -2.205 -139.565 -1.875 -139.235 ;
        RECT -2.205 -140.925 -1.875 -140.595 ;
        RECT -2.205 -142.285 -1.875 -141.955 ;
        RECT -2.205 -143.645 -1.875 -143.315 ;
        RECT -2.205 -145.005 -1.875 -144.675 ;
        RECT -2.205 -146.365 -1.875 -146.035 ;
        RECT -2.205 -147.725 -1.875 -147.395 ;
        RECT -2.205 -149.085 -1.875 -148.755 ;
        RECT -2.205 -150.445 -1.875 -150.115 ;
        RECT -2.205 -151.805 -1.875 -151.475 ;
        RECT -2.205 -153.165 -1.875 -152.835 ;
        RECT -2.205 -154.525 -1.875 -154.195 ;
        RECT -2.205 -155.885 -1.875 -155.555 ;
        RECT -2.205 -157.245 -1.875 -156.915 ;
        RECT -2.205 -158.605 -1.875 -158.275 ;
        RECT -2.205 -159.965 -1.875 -159.635 ;
        RECT -2.205 -161.325 -1.875 -160.995 ;
        RECT -2.205 -162.685 -1.875 -162.355 ;
        RECT -2.205 -164.045 -1.875 -163.715 ;
        RECT -2.205 -165.405 -1.875 -165.075 ;
        RECT -2.205 -166.765 -1.875 -166.435 ;
        RECT -2.205 -168.125 -1.875 -167.795 ;
        RECT -2.205 -169.485 -1.875 -169.155 ;
        RECT -2.205 -170.845 -1.875 -170.515 ;
        RECT -2.205 -172.205 -1.875 -171.875 ;
        RECT -2.205 -173.565 -1.875 -173.235 ;
        RECT -2.205 -174.925 -1.875 -174.595 ;
        RECT -2.205 -176.285 -1.875 -175.955 ;
        RECT -2.205 -177.645 -1.875 -177.315 ;
        RECT -2.205 -179.005 -1.875 -178.675 ;
        RECT -2.205 -180.365 -1.875 -180.035 ;
        RECT -2.205 -181.725 -1.875 -181.395 ;
        RECT -2.205 -183.085 -1.875 -182.755 ;
        RECT -2.205 -184.445 -1.875 -184.115 ;
        RECT -2.205 -185.805 -1.875 -185.475 ;
        RECT -2.205 -187.165 -1.875 -186.835 ;
        RECT -2.205 -188.525 -1.875 -188.195 ;
        RECT -2.205 -189.885 -1.875 -189.555 ;
        RECT -2.205 -191.245 -1.875 -190.915 ;
        RECT -2.205 -192.605 -1.875 -192.275 ;
        RECT -2.205 -193.965 -1.875 -193.635 ;
        RECT -2.205 -195.325 -1.875 -194.995 ;
        RECT -2.205 -196.685 -1.875 -196.355 ;
        RECT -2.205 -198.045 -1.875 -197.715 ;
        RECT -2.205 -199.405 -1.875 -199.075 ;
        RECT -2.205 -200.765 -1.875 -200.435 ;
        RECT -2.205 -202.125 -1.875 -201.795 ;
        RECT -2.205 -203.485 -1.875 -203.155 ;
        RECT -2.205 -204.845 -1.875 -204.515 ;
        RECT -2.205 -206.205 -1.875 -205.875 ;
        RECT -2.205 -207.565 -1.875 -207.235 ;
        RECT -2.205 -208.925 -1.875 -208.595 ;
        RECT -2.205 -210.285 -1.875 -209.955 ;
        RECT -2.205 -211.645 -1.875 -211.315 ;
        RECT -2.205 -213.005 -1.875 -212.675 ;
        RECT -2.205 -214.365 -1.875 -214.035 ;
        RECT -2.205 -215.725 -1.875 -215.395 ;
        RECT -2.205 -217.085 -1.875 -216.755 ;
        RECT -2.205 -218.445 -1.875 -218.115 ;
        RECT -2.205 -219.805 -1.875 -219.475 ;
        RECT -2.205 -221.165 -1.875 -220.835 ;
        RECT -2.205 -222.525 -1.875 -222.195 ;
        RECT -2.205 -223.885 -1.875 -223.555 ;
        RECT -2.205 -225.245 -1.875 -224.915 ;
        RECT -2.205 -226.605 -1.875 -226.275 ;
        RECT -2.205 -227.965 -1.875 -227.635 ;
        RECT -2.205 -229.325 -1.875 -228.995 ;
        RECT -2.205 -230.685 -1.875 -230.355 ;
        RECT -2.205 -232.045 -1.875 -231.715 ;
        RECT -2.205 -233.405 -1.875 -233.075 ;
        RECT -2.205 -234.765 -1.875 -234.435 ;
        RECT -2.205 -236.125 -1.875 -235.795 ;
        RECT -2.205 -237.485 -1.875 -237.155 ;
        RECT -2.205 -238.845 -1.875 -238.515 ;
        RECT -2.205 -241.09 -1.875 -239.96 ;
        RECT -2.2 -241.205 -1.88 -136.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 244.04 -0.515 245.17 ;
        RECT -0.845 242.595 -0.515 242.925 ;
        RECT -0.845 241.235 -0.515 241.565 ;
        RECT -0.845 239.875 -0.515 240.205 ;
        RECT -0.845 238.515 -0.515 238.845 ;
        RECT -0.845 237.155 -0.515 237.485 ;
        RECT -0.845 235.975 -0.515 236.305 ;
        RECT -0.845 233.925 -0.515 234.255 ;
        RECT -0.845 231.995 -0.515 232.325 ;
        RECT -0.845 230.155 -0.515 230.485 ;
        RECT -0.845 228.665 -0.515 228.995 ;
        RECT -0.845 226.995 -0.515 227.325 ;
        RECT -0.845 225.505 -0.515 225.835 ;
        RECT -0.845 223.835 -0.515 224.165 ;
        RECT -0.845 222.345 -0.515 222.675 ;
        RECT -0.845 220.675 -0.515 221.005 ;
        RECT -0.845 219.185 -0.515 219.515 ;
        RECT -0.845 217.775 -0.515 218.105 ;
        RECT -0.845 215.935 -0.515 216.265 ;
        RECT -0.845 214.445 -0.515 214.775 ;
        RECT -0.845 212.775 -0.515 213.105 ;
        RECT -0.845 211.285 -0.515 211.615 ;
        RECT -0.845 209.615 -0.515 209.945 ;
        RECT -0.845 208.125 -0.515 208.455 ;
        RECT -0.845 206.455 -0.515 206.785 ;
        RECT -0.845 204.965 -0.515 205.295 ;
        RECT -0.845 203.555 -0.515 203.885 ;
        RECT -0.845 201.715 -0.515 202.045 ;
        RECT -0.845 200.225 -0.515 200.555 ;
        RECT -0.845 198.555 -0.515 198.885 ;
        RECT -0.845 197.065 -0.515 197.395 ;
        RECT -0.845 195.395 -0.515 195.725 ;
        RECT -0.845 193.905 -0.515 194.235 ;
        RECT -0.845 192.235 -0.515 192.565 ;
        RECT -0.845 190.745 -0.515 191.075 ;
        RECT -0.845 189.335 -0.515 189.665 ;
        RECT -0.845 187.495 -0.515 187.825 ;
        RECT -0.845 186.005 -0.515 186.335 ;
        RECT -0.845 184.335 -0.515 184.665 ;
        RECT -0.845 182.845 -0.515 183.175 ;
        RECT -0.845 181.175 -0.515 181.505 ;
        RECT -0.845 179.685 -0.515 180.015 ;
        RECT -0.845 178.015 -0.515 178.345 ;
        RECT -0.845 176.525 -0.515 176.855 ;
        RECT -0.845 175.115 -0.515 175.445 ;
        RECT -0.845 173.275 -0.515 173.605 ;
        RECT -0.845 171.785 -0.515 172.115 ;
        RECT -0.845 170.115 -0.515 170.445 ;
        RECT -0.845 168.625 -0.515 168.955 ;
        RECT -0.845 166.955 -0.515 167.285 ;
        RECT -0.845 165.465 -0.515 165.795 ;
        RECT -0.845 163.795 -0.515 164.125 ;
        RECT -0.845 162.305 -0.515 162.635 ;
        RECT -0.845 160.895 -0.515 161.225 ;
        RECT -0.845 159.055 -0.515 159.385 ;
        RECT -0.845 157.565 -0.515 157.895 ;
        RECT -0.845 155.895 -0.515 156.225 ;
        RECT -0.845 154.405 -0.515 154.735 ;
        RECT -0.845 152.735 -0.515 153.065 ;
        RECT -0.845 151.245 -0.515 151.575 ;
        RECT -0.845 149.575 -0.515 149.905 ;
        RECT -0.845 148.085 -0.515 148.415 ;
        RECT -0.845 146.675 -0.515 147.005 ;
        RECT -0.845 144.835 -0.515 145.165 ;
        RECT -0.845 143.345 -0.515 143.675 ;
        RECT -0.845 141.675 -0.515 142.005 ;
        RECT -0.845 140.185 -0.515 140.515 ;
        RECT -0.845 138.515 -0.515 138.845 ;
        RECT -0.845 137.025 -0.515 137.355 ;
        RECT -0.845 135.355 -0.515 135.685 ;
        RECT -0.845 133.865 -0.515 134.195 ;
        RECT -0.845 132.455 -0.515 132.785 ;
        RECT -0.845 130.615 -0.515 130.945 ;
        RECT -0.845 129.125 -0.515 129.455 ;
        RECT -0.845 127.455 -0.515 127.785 ;
        RECT -0.845 125.965 -0.515 126.295 ;
        RECT -0.845 124.295 -0.515 124.625 ;
        RECT -0.845 122.805 -0.515 123.135 ;
        RECT -0.845 121.135 -0.515 121.465 ;
        RECT -0.845 119.645 -0.515 119.975 ;
        RECT -0.845 118.235 -0.515 118.565 ;
        RECT -0.845 116.395 -0.515 116.725 ;
        RECT -0.845 114.905 -0.515 115.235 ;
        RECT -0.845 113.235 -0.515 113.565 ;
        RECT -0.845 111.745 -0.515 112.075 ;
        RECT -0.845 110.075 -0.515 110.405 ;
        RECT -0.845 108.585 -0.515 108.915 ;
        RECT -0.845 106.915 -0.515 107.245 ;
        RECT -0.845 105.425 -0.515 105.755 ;
        RECT -0.845 104.015 -0.515 104.345 ;
        RECT -0.845 102.175 -0.515 102.505 ;
        RECT -0.845 100.685 -0.515 101.015 ;
        RECT -0.845 99.015 -0.515 99.345 ;
        RECT -0.845 97.525 -0.515 97.855 ;
        RECT -0.845 95.855 -0.515 96.185 ;
        RECT -0.845 94.365 -0.515 94.695 ;
        RECT -0.845 92.695 -0.515 93.025 ;
        RECT -0.845 91.205 -0.515 91.535 ;
        RECT -0.845 89.795 -0.515 90.125 ;
        RECT -0.845 87.955 -0.515 88.285 ;
        RECT -0.845 86.465 -0.515 86.795 ;
        RECT -0.845 84.795 -0.515 85.125 ;
        RECT -0.845 83.305 -0.515 83.635 ;
        RECT -0.845 81.635 -0.515 81.965 ;
        RECT -0.845 80.145 -0.515 80.475 ;
        RECT -0.845 78.475 -0.515 78.805 ;
        RECT -0.845 76.985 -0.515 77.315 ;
        RECT -0.845 75.575 -0.515 75.905 ;
        RECT -0.845 73.735 -0.515 74.065 ;
        RECT -0.845 72.245 -0.515 72.575 ;
        RECT -0.845 70.575 -0.515 70.905 ;
        RECT -0.845 69.085 -0.515 69.415 ;
        RECT -0.845 67.415 -0.515 67.745 ;
        RECT -0.845 65.925 -0.515 66.255 ;
        RECT -0.845 64.255 -0.515 64.585 ;
        RECT -0.845 62.765 -0.515 63.095 ;
        RECT -0.845 61.355 -0.515 61.685 ;
        RECT -0.845 59.515 -0.515 59.845 ;
        RECT -0.845 58.025 -0.515 58.355 ;
        RECT -0.845 56.355 -0.515 56.685 ;
        RECT -0.845 54.865 -0.515 55.195 ;
        RECT -0.845 53.195 -0.515 53.525 ;
        RECT -0.845 51.705 -0.515 52.035 ;
        RECT -0.845 50.035 -0.515 50.365 ;
        RECT -0.845 48.545 -0.515 48.875 ;
        RECT -0.845 47.135 -0.515 47.465 ;
        RECT -0.845 45.295 -0.515 45.625 ;
        RECT -0.845 43.805 -0.515 44.135 ;
        RECT -0.845 42.135 -0.515 42.465 ;
        RECT -0.845 40.645 -0.515 40.975 ;
        RECT -0.845 38.975 -0.515 39.305 ;
        RECT -0.845 37.485 -0.515 37.815 ;
        RECT -0.845 35.815 -0.515 36.145 ;
        RECT -0.845 34.325 -0.515 34.655 ;
        RECT -0.845 32.915 -0.515 33.245 ;
        RECT -0.845 31.075 -0.515 31.405 ;
        RECT -0.845 29.585 -0.515 29.915 ;
        RECT -0.845 27.915 -0.515 28.245 ;
        RECT -0.845 26.425 -0.515 26.755 ;
        RECT -0.845 24.755 -0.515 25.085 ;
        RECT -0.845 23.265 -0.515 23.595 ;
        RECT -0.845 21.595 -0.515 21.925 ;
        RECT -0.845 20.105 -0.515 20.435 ;
        RECT -0.845 18.695 -0.515 19.025 ;
        RECT -0.845 16.855 -0.515 17.185 ;
        RECT -0.845 15.365 -0.515 15.695 ;
        RECT -0.845 13.695 -0.515 14.025 ;
        RECT -0.845 12.205 -0.515 12.535 ;
        RECT -0.845 10.535 -0.515 10.865 ;
        RECT -0.845 9.045 -0.515 9.375 ;
        RECT -0.845 7.375 -0.515 7.705 ;
        RECT -0.845 5.885 -0.515 6.215 ;
        RECT -0.845 4.475 -0.515 4.805 ;
        RECT -0.845 2.115 -0.515 2.445 ;
        RECT -0.845 0.06 -0.515 0.39 ;
        RECT -0.845 -0.845 -0.515 -0.515 ;
        RECT -0.845 -2.205 -0.515 -1.875 ;
        RECT -0.845 -3.565 -0.515 -3.235 ;
        RECT -0.845 -4.925 -0.515 -4.595 ;
        RECT -0.845 -6.285 -0.515 -5.955 ;
        RECT -0.845 -7.645 -0.515 -7.315 ;
        RECT -0.845 -9.005 -0.515 -8.675 ;
        RECT -0.845 -10.365 -0.515 -10.035 ;
        RECT -0.845 -13.085 -0.515 -12.755 ;
        RECT -0.845 -14.445 -0.515 -14.115 ;
        RECT -0.845 -15.805 -0.515 -15.475 ;
        RECT -0.845 -17.165 -0.515 -16.835 ;
        RECT -0.845 -18.525 -0.515 -18.195 ;
        RECT -0.845 -26.685 -0.515 -26.355 ;
        RECT -0.845 -28.045 -0.515 -27.715 ;
        RECT -0.845 -29.405 -0.515 -29.075 ;
        RECT -0.845 -30.765 -0.515 -30.435 ;
        RECT -0.845 -32.125 -0.515 -31.795 ;
        RECT -0.845 -33.485 -0.515 -33.155 ;
        RECT -0.845 -34.845 -0.515 -34.515 ;
        RECT -0.845 -36.205 -0.515 -35.875 ;
        RECT -0.845 -37.565 -0.515 -37.235 ;
        RECT -0.845 -38.925 -0.515 -38.595 ;
        RECT -0.845 -40.285 -0.515 -39.955 ;
        RECT -0.845 -41.645 -0.515 -41.315 ;
        RECT -0.845 -43.005 -0.515 -42.675 ;
        RECT -0.845 -44.365 -0.515 -44.035 ;
        RECT -0.845 -45.725 -0.515 -45.395 ;
        RECT -0.845 -47.085 -0.515 -46.755 ;
        RECT -0.845 -48.445 -0.515 -48.115 ;
        RECT -0.845 -49.805 -0.515 -49.475 ;
        RECT -0.845 -51.165 -0.515 -50.835 ;
        RECT -0.845 -52.525 -0.515 -52.195 ;
        RECT -0.845 -53.885 -0.515 -53.555 ;
        RECT -0.845 -55.245 -0.515 -54.915 ;
        RECT -0.845 -56.605 -0.515 -56.275 ;
        RECT -0.845 -57.965 -0.515 -57.635 ;
        RECT -0.845 -59.325 -0.515 -58.995 ;
        RECT -0.845 -60.685 -0.515 -60.355 ;
        RECT -0.845 -62.045 -0.515 -61.715 ;
        RECT -0.845 -68.845 -0.515 -68.515 ;
        RECT -0.845 -70.205 -0.515 -69.875 ;
        RECT -0.845 -72.925 -0.515 -72.595 ;
        RECT -0.845 -74.285 -0.515 -73.955 ;
        RECT -0.845 -75.645 -0.515 -75.315 ;
        RECT -0.845 -77.005 -0.515 -76.675 ;
        RECT -0.845 -78.365 -0.515 -78.035 ;
        RECT -0.845 -79.725 -0.515 -79.395 ;
        RECT -0.845 -81.085 -0.515 -80.755 ;
        RECT -0.845 -82.445 -0.515 -82.115 ;
        RECT -0.845 -83.805 -0.515 -83.475 ;
        RECT -0.845 -85.165 -0.515 -84.835 ;
        RECT -0.845 -86.525 -0.515 -86.195 ;
        RECT -0.845 -87.885 -0.515 -87.555 ;
        RECT -0.845 -89.245 -0.515 -88.915 ;
        RECT -0.845 -90.605 -0.515 -90.275 ;
        RECT -0.845 -91.965 -0.515 -91.635 ;
        RECT -0.845 -93.325 -0.515 -92.995 ;
        RECT -0.845 -94.685 -0.515 -94.355 ;
        RECT -0.845 -96.045 -0.515 -95.715 ;
        RECT -0.845 -97.405 -0.515 -97.075 ;
        RECT -0.845 -98.765 -0.515 -98.435 ;
        RECT -0.845 -100.125 -0.515 -99.795 ;
        RECT -0.845 -101.485 -0.515 -101.155 ;
        RECT -0.845 -102.845 -0.515 -102.515 ;
        RECT -0.845 -104.205 -0.515 -103.875 ;
        RECT -0.845 -105.565 -0.515 -105.235 ;
        RECT -0.845 -106.925 -0.515 -106.595 ;
        RECT -0.845 -108.285 -0.515 -107.955 ;
        RECT -0.845 -109.645 -0.515 -109.315 ;
        RECT -0.845 -111.005 -0.515 -110.675 ;
        RECT -0.845 -112.365 -0.515 -112.035 ;
        RECT -0.845 -113.725 -0.515 -113.395 ;
        RECT -0.845 -115.085 -0.515 -114.755 ;
        RECT -0.845 -116.445 -0.515 -116.115 ;
        RECT -0.845 -119.165 -0.515 -118.835 ;
        RECT -0.845 -120.525 -0.515 -120.195 ;
        RECT -0.845 -121.885 -0.515 -121.555 ;
        RECT -0.845 -123.245 -0.515 -122.915 ;
        RECT -0.845 -124.605 -0.515 -124.275 ;
        RECT -0.845 -125.965 -0.515 -125.635 ;
        RECT -0.845 -127.325 -0.515 -126.995 ;
        RECT -0.845 -128.685 -0.515 -128.355 ;
        RECT -0.845 -130.045 -0.515 -129.715 ;
        RECT -0.845 -131.405 -0.515 -131.075 ;
        RECT -0.845 -132.765 -0.515 -132.435 ;
        RECT -0.845 -134.125 -0.515 -133.795 ;
        RECT -0.845 -135.485 -0.515 -135.155 ;
        RECT -0.845 -136.845 -0.515 -136.515 ;
        RECT -0.845 -138.205 -0.515 -137.875 ;
        RECT -0.845 -139.565 -0.515 -139.235 ;
        RECT -0.845 -140.925 -0.515 -140.595 ;
        RECT -0.845 -142.285 -0.515 -141.955 ;
        RECT -0.845 -143.645 -0.515 -143.315 ;
        RECT -0.845 -145.005 -0.515 -144.675 ;
        RECT -0.845 -146.365 -0.515 -146.035 ;
        RECT -0.845 -147.725 -0.515 -147.395 ;
        RECT -0.845 -149.085 -0.515 -148.755 ;
        RECT -0.845 -150.445 -0.515 -150.115 ;
        RECT -0.845 -151.805 -0.515 -151.475 ;
        RECT -0.845 -153.165 -0.515 -152.835 ;
        RECT -0.845 -154.525 -0.515 -154.195 ;
        RECT -0.845 -155.885 -0.515 -155.555 ;
        RECT -0.845 -157.245 -0.515 -156.915 ;
        RECT -0.845 -158.605 -0.515 -158.275 ;
        RECT -0.845 -159.965 -0.515 -159.635 ;
        RECT -0.845 -161.325 -0.515 -160.995 ;
        RECT -0.845 -162.685 -0.515 -162.355 ;
        RECT -0.845 -164.045 -0.515 -163.715 ;
        RECT -0.845 -165.405 -0.515 -165.075 ;
        RECT -0.845 -166.765 -0.515 -166.435 ;
        RECT -0.845 -168.125 -0.515 -167.795 ;
        RECT -0.845 -169.485 -0.515 -169.155 ;
        RECT -0.845 -170.845 -0.515 -170.515 ;
        RECT -0.845 -172.205 -0.515 -171.875 ;
        RECT -0.845 -173.565 -0.515 -173.235 ;
        RECT -0.845 -174.925 -0.515 -174.595 ;
        RECT -0.845 -176.285 -0.515 -175.955 ;
        RECT -0.845 -177.645 -0.515 -177.315 ;
        RECT -0.845 -179.005 -0.515 -178.675 ;
        RECT -0.845 -180.365 -0.515 -180.035 ;
        RECT -0.845 -181.725 -0.515 -181.395 ;
        RECT -0.845 -183.085 -0.515 -182.755 ;
        RECT -0.845 -184.445 -0.515 -184.115 ;
        RECT -0.845 -185.805 -0.515 -185.475 ;
        RECT -0.845 -187.165 -0.515 -186.835 ;
        RECT -0.845 -188.525 -0.515 -188.195 ;
        RECT -0.845 -189.885 -0.515 -189.555 ;
        RECT -0.845 -191.245 -0.515 -190.915 ;
        RECT -0.845 -192.605 -0.515 -192.275 ;
        RECT -0.845 -193.965 -0.515 -193.635 ;
        RECT -0.845 -195.325 -0.515 -194.995 ;
        RECT -0.845 -196.685 -0.515 -196.355 ;
        RECT -0.845 -198.045 -0.515 -197.715 ;
        RECT -0.845 -199.405 -0.515 -199.075 ;
        RECT -0.845 -200.765 -0.515 -200.435 ;
        RECT -0.845 -202.125 -0.515 -201.795 ;
        RECT -0.845 -203.485 -0.515 -203.155 ;
        RECT -0.845 -204.845 -0.515 -204.515 ;
        RECT -0.845 -206.205 -0.515 -205.875 ;
        RECT -0.845 -207.565 -0.515 -207.235 ;
        RECT -0.845 -208.925 -0.515 -208.595 ;
        RECT -0.845 -210.285 -0.515 -209.955 ;
        RECT -0.845 -211.645 -0.515 -211.315 ;
        RECT -0.845 -213.005 -0.515 -212.675 ;
        RECT -0.845 -214.365 -0.515 -214.035 ;
        RECT -0.845 -215.725 -0.515 -215.395 ;
        RECT -0.845 -217.085 -0.515 -216.755 ;
        RECT -0.845 -218.445 -0.515 -218.115 ;
        RECT -0.845 -219.805 -0.515 -219.475 ;
        RECT -0.845 -221.165 -0.515 -220.835 ;
        RECT -0.845 -222.525 -0.515 -222.195 ;
        RECT -0.845 -223.885 -0.515 -223.555 ;
        RECT -0.845 -225.245 -0.515 -224.915 ;
        RECT -0.845 -226.605 -0.515 -226.275 ;
        RECT -0.845 -227.965 -0.515 -227.635 ;
        RECT -0.845 -229.325 -0.515 -228.995 ;
        RECT -0.845 -230.685 -0.515 -230.355 ;
        RECT -0.845 -232.045 -0.515 -231.715 ;
        RECT -0.845 -233.405 -0.515 -233.075 ;
        RECT -0.845 -234.765 -0.515 -234.435 ;
        RECT -0.845 -236.125 -0.515 -235.795 ;
        RECT -0.845 -237.485 -0.515 -237.155 ;
        RECT -0.845 -238.845 -0.515 -238.515 ;
        RECT -0.845 -241.09 -0.515 -239.96 ;
        RECT -0.84 -241.205 -0.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 244.04 0.845 245.17 ;
        RECT 0.515 242.595 0.845 242.925 ;
        RECT 0.515 241.235 0.845 241.565 ;
        RECT 0.515 239.875 0.845 240.205 ;
        RECT 0.515 238.515 0.845 238.845 ;
        RECT 0.515 237.155 0.845 237.485 ;
        RECT 0.52 237.155 0.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -0.845 0.845 -0.515 ;
        RECT 0.515 -2.205 0.845 -1.875 ;
        RECT 0.515 -3.565 0.845 -3.235 ;
        RECT 0.52 -3.565 0.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -123.245 0.845 -122.915 ;
        RECT 0.515 -124.605 0.845 -124.275 ;
        RECT 0.515 -125.965 0.845 -125.635 ;
        RECT 0.515 -127.325 0.845 -126.995 ;
        RECT 0.515 -128.685 0.845 -128.355 ;
        RECT 0.515 -130.045 0.845 -129.715 ;
        RECT 0.515 -131.405 0.845 -131.075 ;
        RECT 0.515 -132.765 0.845 -132.435 ;
        RECT 0.515 -134.125 0.845 -133.795 ;
        RECT 0.515 -135.485 0.845 -135.155 ;
        RECT 0.515 -136.845 0.845 -136.515 ;
        RECT 0.515 -138.205 0.845 -137.875 ;
        RECT 0.515 -139.565 0.845 -139.235 ;
        RECT 0.515 -140.925 0.845 -140.595 ;
        RECT 0.515 -142.285 0.845 -141.955 ;
        RECT 0.515 -143.645 0.845 -143.315 ;
        RECT 0.515 -145.005 0.845 -144.675 ;
        RECT 0.515 -146.365 0.845 -146.035 ;
        RECT 0.515 -147.725 0.845 -147.395 ;
        RECT 0.515 -149.085 0.845 -148.755 ;
        RECT 0.515 -150.445 0.845 -150.115 ;
        RECT 0.515 -151.805 0.845 -151.475 ;
        RECT 0.515 -153.165 0.845 -152.835 ;
        RECT 0.515 -154.525 0.845 -154.195 ;
        RECT 0.515 -155.885 0.845 -155.555 ;
        RECT 0.515 -157.245 0.845 -156.915 ;
        RECT 0.515 -158.605 0.845 -158.275 ;
        RECT 0.515 -159.965 0.845 -159.635 ;
        RECT 0.515 -161.325 0.845 -160.995 ;
        RECT 0.515 -162.685 0.845 -162.355 ;
        RECT 0.515 -164.045 0.845 -163.715 ;
        RECT 0.515 -165.405 0.845 -165.075 ;
        RECT 0.515 -166.765 0.845 -166.435 ;
        RECT 0.515 -168.125 0.845 -167.795 ;
        RECT 0.515 -169.485 0.845 -169.155 ;
        RECT 0.515 -170.845 0.845 -170.515 ;
        RECT 0.515 -172.205 0.845 -171.875 ;
        RECT 0.515 -173.565 0.845 -173.235 ;
        RECT 0.515 -174.925 0.845 -174.595 ;
        RECT 0.515 -176.285 0.845 -175.955 ;
        RECT 0.515 -177.645 0.845 -177.315 ;
        RECT 0.515 -179.005 0.845 -178.675 ;
        RECT 0.515 -180.365 0.845 -180.035 ;
        RECT 0.515 -181.725 0.845 -181.395 ;
        RECT 0.515 -183.085 0.845 -182.755 ;
        RECT 0.515 -184.445 0.845 -184.115 ;
        RECT 0.515 -185.805 0.845 -185.475 ;
        RECT 0.515 -187.165 0.845 -186.835 ;
        RECT 0.515 -188.525 0.845 -188.195 ;
        RECT 0.515 -189.885 0.845 -189.555 ;
        RECT 0.515 -191.245 0.845 -190.915 ;
        RECT 0.515 -192.605 0.845 -192.275 ;
        RECT 0.515 -193.965 0.845 -193.635 ;
        RECT 0.515 -195.325 0.845 -194.995 ;
        RECT 0.515 -196.685 0.845 -196.355 ;
        RECT 0.515 -198.045 0.845 -197.715 ;
        RECT 0.515 -199.405 0.845 -199.075 ;
        RECT 0.515 -200.765 0.845 -200.435 ;
        RECT 0.515 -202.125 0.845 -201.795 ;
        RECT 0.515 -203.485 0.845 -203.155 ;
        RECT 0.515 -204.845 0.845 -204.515 ;
        RECT 0.515 -206.205 0.845 -205.875 ;
        RECT 0.515 -207.565 0.845 -207.235 ;
        RECT 0.515 -208.925 0.845 -208.595 ;
        RECT 0.515 -210.285 0.845 -209.955 ;
        RECT 0.515 -211.645 0.845 -211.315 ;
        RECT 0.515 -213.005 0.845 -212.675 ;
        RECT 0.515 -214.365 0.845 -214.035 ;
        RECT 0.515 -215.725 0.845 -215.395 ;
        RECT 0.515 -217.085 0.845 -216.755 ;
        RECT 0.515 -218.445 0.845 -218.115 ;
        RECT 0.515 -219.805 0.845 -219.475 ;
        RECT 0.515 -221.165 0.845 -220.835 ;
        RECT 0.515 -222.525 0.845 -222.195 ;
        RECT 0.515 -223.885 0.845 -223.555 ;
        RECT 0.515 -225.245 0.845 -224.915 ;
        RECT 0.515 -226.605 0.845 -226.275 ;
        RECT 0.515 -227.965 0.845 -227.635 ;
        RECT 0.515 -229.325 0.845 -228.995 ;
        RECT 0.515 -230.685 0.845 -230.355 ;
        RECT 0.515 -232.045 0.845 -231.715 ;
        RECT 0.515 -233.405 0.845 -233.075 ;
        RECT 0.515 -234.765 0.845 -234.435 ;
        RECT 0.515 -236.125 0.845 -235.795 ;
        RECT 0.515 -237.485 0.845 -237.155 ;
        RECT 0.515 -238.845 0.845 -238.515 ;
        RECT 0.515 -241.09 0.845 -239.96 ;
        RECT 0.52 -241.205 0.84 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 244.04 2.205 245.17 ;
        RECT 1.875 242.595 2.205 242.925 ;
        RECT 1.875 241.235 2.205 241.565 ;
        RECT 1.875 239.875 2.205 240.205 ;
        RECT 1.875 238.515 2.205 238.845 ;
        RECT 1.875 237.155 2.205 237.485 ;
        RECT 1.88 237.155 2.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -0.845 2.205 -0.515 ;
        RECT 1.875 -2.205 2.205 -1.875 ;
        RECT 1.875 -3.565 2.205 -3.235 ;
        RECT 1.88 -3.565 2.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -123.245 2.205 -122.915 ;
        RECT 1.875 -124.605 2.205 -124.275 ;
        RECT 1.875 -125.965 2.205 -125.635 ;
        RECT 1.875 -127.325 2.205 -126.995 ;
        RECT 1.875 -128.685 2.205 -128.355 ;
        RECT 1.875 -130.045 2.205 -129.715 ;
        RECT 1.875 -131.405 2.205 -131.075 ;
        RECT 1.875 -132.765 2.205 -132.435 ;
        RECT 1.875 -134.125 2.205 -133.795 ;
        RECT 1.875 -135.485 2.205 -135.155 ;
        RECT 1.875 -136.845 2.205 -136.515 ;
        RECT 1.875 -138.205 2.205 -137.875 ;
        RECT 1.875 -139.565 2.205 -139.235 ;
        RECT 1.875 -140.925 2.205 -140.595 ;
        RECT 1.875 -142.285 2.205 -141.955 ;
        RECT 1.875 -143.645 2.205 -143.315 ;
        RECT 1.875 -145.005 2.205 -144.675 ;
        RECT 1.875 -146.365 2.205 -146.035 ;
        RECT 1.875 -147.725 2.205 -147.395 ;
        RECT 1.875 -149.085 2.205 -148.755 ;
        RECT 1.875 -150.445 2.205 -150.115 ;
        RECT 1.875 -151.805 2.205 -151.475 ;
        RECT 1.875 -153.165 2.205 -152.835 ;
        RECT 1.875 -154.525 2.205 -154.195 ;
        RECT 1.875 -155.885 2.205 -155.555 ;
        RECT 1.875 -157.245 2.205 -156.915 ;
        RECT 1.875 -158.605 2.205 -158.275 ;
        RECT 1.875 -159.965 2.205 -159.635 ;
        RECT 1.875 -161.325 2.205 -160.995 ;
        RECT 1.875 -162.685 2.205 -162.355 ;
        RECT 1.875 -164.045 2.205 -163.715 ;
        RECT 1.875 -165.405 2.205 -165.075 ;
        RECT 1.875 -166.765 2.205 -166.435 ;
        RECT 1.875 -168.125 2.205 -167.795 ;
        RECT 1.875 -169.485 2.205 -169.155 ;
        RECT 1.875 -170.845 2.205 -170.515 ;
        RECT 1.875 -172.205 2.205 -171.875 ;
        RECT 1.875 -173.565 2.205 -173.235 ;
        RECT 1.875 -174.925 2.205 -174.595 ;
        RECT 1.875 -176.285 2.205 -175.955 ;
        RECT 1.875 -177.645 2.205 -177.315 ;
        RECT 1.875 -179.005 2.205 -178.675 ;
        RECT 1.875 -180.365 2.205 -180.035 ;
        RECT 1.875 -181.725 2.205 -181.395 ;
        RECT 1.875 -183.085 2.205 -182.755 ;
        RECT 1.875 -184.445 2.205 -184.115 ;
        RECT 1.875 -185.805 2.205 -185.475 ;
        RECT 1.875 -187.165 2.205 -186.835 ;
        RECT 1.875 -188.525 2.205 -188.195 ;
        RECT 1.875 -189.885 2.205 -189.555 ;
        RECT 1.875 -191.245 2.205 -190.915 ;
        RECT 1.875 -192.605 2.205 -192.275 ;
        RECT 1.875 -193.965 2.205 -193.635 ;
        RECT 1.875 -195.325 2.205 -194.995 ;
        RECT 1.875 -196.685 2.205 -196.355 ;
        RECT 1.875 -198.045 2.205 -197.715 ;
        RECT 1.875 -199.405 2.205 -199.075 ;
        RECT 1.875 -200.765 2.205 -200.435 ;
        RECT 1.875 -202.125 2.205 -201.795 ;
        RECT 1.875 -203.485 2.205 -203.155 ;
        RECT 1.875 -204.845 2.205 -204.515 ;
        RECT 1.875 -206.205 2.205 -205.875 ;
        RECT 1.875 -207.565 2.205 -207.235 ;
        RECT 1.875 -208.925 2.205 -208.595 ;
        RECT 1.875 -210.285 2.205 -209.955 ;
        RECT 1.875 -211.645 2.205 -211.315 ;
        RECT 1.875 -213.005 2.205 -212.675 ;
        RECT 1.875 -214.365 2.205 -214.035 ;
        RECT 1.875 -215.725 2.205 -215.395 ;
        RECT 1.875 -217.085 2.205 -216.755 ;
        RECT 1.875 -218.445 2.205 -218.115 ;
        RECT 1.875 -219.805 2.205 -219.475 ;
        RECT 1.875 -221.165 2.205 -220.835 ;
        RECT 1.875 -222.525 2.205 -222.195 ;
        RECT 1.875 -223.885 2.205 -223.555 ;
        RECT 1.875 -225.245 2.205 -224.915 ;
        RECT 1.875 -226.605 2.205 -226.275 ;
        RECT 1.875 -227.965 2.205 -227.635 ;
        RECT 1.875 -229.325 2.205 -228.995 ;
        RECT 1.875 -230.685 2.205 -230.355 ;
        RECT 1.875 -232.045 2.205 -231.715 ;
        RECT 1.875 -233.405 2.205 -233.075 ;
        RECT 1.875 -234.765 2.205 -234.435 ;
        RECT 1.875 -236.125 2.205 -235.795 ;
        RECT 1.875 -237.485 2.205 -237.155 ;
        RECT 1.875 -238.845 2.205 -238.515 ;
        RECT 1.875 -241.09 2.205 -239.96 ;
        RECT 1.88 -241.205 2.2 -122.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 244.04 3.565 245.17 ;
        RECT 3.235 242.595 3.565 242.925 ;
        RECT 3.235 241.235 3.565 241.565 ;
        RECT 3.235 239.875 3.565 240.205 ;
        RECT 3.235 238.515 3.565 238.845 ;
        RECT 3.235 237.155 3.565 237.485 ;
        RECT 3.24 237.155 3.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 -208.925 3.565 -208.595 ;
        RECT 3.235 -210.285 3.565 -209.955 ;
        RECT 3.235 -211.645 3.565 -211.315 ;
        RECT 3.235 -213.005 3.565 -212.675 ;
        RECT 3.235 -214.365 3.565 -214.035 ;
        RECT 3.235 -215.725 3.565 -215.395 ;
        RECT 3.235 -217.085 3.565 -216.755 ;
        RECT 3.235 -218.445 3.565 -218.115 ;
        RECT 3.235 -219.805 3.565 -219.475 ;
        RECT 3.235 -221.165 3.565 -220.835 ;
        RECT 3.235 -222.525 3.565 -222.195 ;
        RECT 3.235 -223.885 3.565 -223.555 ;
        RECT 3.235 -225.245 3.565 -224.915 ;
        RECT 3.235 -226.605 3.565 -226.275 ;
        RECT 3.235 -227.965 3.565 -227.635 ;
        RECT 3.235 -229.325 3.565 -228.995 ;
        RECT 3.235 -230.685 3.565 -230.355 ;
        RECT 3.235 -232.045 3.565 -231.715 ;
        RECT 3.235 -233.405 3.565 -233.075 ;
        RECT 3.235 -234.765 3.565 -234.435 ;
        RECT 3.235 -236.125 3.565 -235.795 ;
        RECT 3.235 -237.485 3.565 -237.155 ;
        RECT 3.235 -238.845 3.565 -238.515 ;
        RECT 3.235 -241.09 3.565 -239.96 ;
        RECT 3.24 -241.205 3.56 -126.32 ;
        RECT 3.235 -127.325 3.565 -126.995 ;
        RECT 3.235 -128.685 3.565 -128.355 ;
        RECT 3.235 -130.045 3.565 -129.715 ;
        RECT 3.235 -131.405 3.565 -131.075 ;
        RECT 3.235 -132.765 3.565 -132.435 ;
        RECT 3.235 -134.125 3.565 -133.795 ;
        RECT 3.235 -135.485 3.565 -135.155 ;
        RECT 3.235 -136.845 3.565 -136.515 ;
        RECT 3.235 -138.205 3.565 -137.875 ;
        RECT 3.235 -139.565 3.565 -139.235 ;
        RECT 3.235 -140.925 3.565 -140.595 ;
        RECT 3.235 -142.285 3.565 -141.955 ;
        RECT 3.235 -143.645 3.565 -143.315 ;
        RECT 3.235 -145.005 3.565 -144.675 ;
        RECT 3.235 -146.365 3.565 -146.035 ;
        RECT 3.235 -147.725 3.565 -147.395 ;
        RECT 3.235 -149.085 3.565 -148.755 ;
        RECT 3.235 -150.445 3.565 -150.115 ;
        RECT 3.235 -151.805 3.565 -151.475 ;
        RECT 3.235 -153.165 3.565 -152.835 ;
        RECT 3.235 -154.525 3.565 -154.195 ;
        RECT 3.235 -155.885 3.565 -155.555 ;
        RECT 3.235 -157.245 3.565 -156.915 ;
        RECT 3.235 -158.605 3.565 -158.275 ;
        RECT 3.235 -159.965 3.565 -159.635 ;
        RECT 3.235 -161.325 3.565 -160.995 ;
        RECT 3.235 -162.685 3.565 -162.355 ;
        RECT 3.235 -164.045 3.565 -163.715 ;
        RECT 3.235 -165.405 3.565 -165.075 ;
        RECT 3.235 -166.765 3.565 -166.435 ;
        RECT 3.235 -168.125 3.565 -167.795 ;
        RECT 3.235 -169.485 3.565 -169.155 ;
        RECT 3.235 -170.845 3.565 -170.515 ;
        RECT 3.235 -172.205 3.565 -171.875 ;
        RECT 3.235 -173.565 3.565 -173.235 ;
        RECT 3.235 -174.925 3.565 -174.595 ;
        RECT 3.235 -176.285 3.565 -175.955 ;
        RECT 3.235 -177.645 3.565 -177.315 ;
        RECT 3.235 -179.005 3.565 -178.675 ;
        RECT 3.235 -180.365 3.565 -180.035 ;
        RECT 3.235 -181.725 3.565 -181.395 ;
        RECT 3.235 -183.085 3.565 -182.755 ;
        RECT 3.235 -184.445 3.565 -184.115 ;
        RECT 3.235 -185.805 3.565 -185.475 ;
        RECT 3.235 -187.165 3.565 -186.835 ;
        RECT 3.235 -188.525 3.565 -188.195 ;
        RECT 3.235 -189.885 3.565 -189.555 ;
        RECT 3.235 -191.245 3.565 -190.915 ;
        RECT 3.235 -192.605 3.565 -192.275 ;
        RECT 3.235 -193.965 3.565 -193.635 ;
        RECT 3.235 -195.325 3.565 -194.995 ;
        RECT 3.235 -196.685 3.565 -196.355 ;
        RECT 3.235 -198.045 3.565 -197.715 ;
        RECT 3.235 -199.405 3.565 -199.075 ;
        RECT 3.235 -200.765 3.565 -200.435 ;
        RECT 3.235 -202.125 3.565 -201.795 ;
        RECT 3.235 -203.485 3.565 -203.155 ;
        RECT 3.235 -204.845 3.565 -204.515 ;
        RECT 3.235 -206.205 3.565 -205.875 ;
        RECT 3.235 -207.565 3.565 -207.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.645 244.04 -7.315 245.17 ;
        RECT -7.645 242.595 -7.315 242.925 ;
        RECT -7.645 241.235 -7.315 241.565 ;
        RECT -7.645 239.875 -7.315 240.205 ;
        RECT -7.645 238.515 -7.315 238.845 ;
        RECT -7.645 237.155 -7.315 237.485 ;
        RECT -7.645 235.795 -7.315 236.125 ;
        RECT -7.645 234.435 -7.315 234.765 ;
        RECT -7.645 233.075 -7.315 233.405 ;
        RECT -7.645 231.715 -7.315 232.045 ;
        RECT -7.645 227.635 -7.315 227.965 ;
        RECT -7.645 224.915 -7.315 225.245 ;
        RECT -7.645 218.115 -7.315 218.445 ;
        RECT -7.645 216.755 -7.315 217.085 ;
        RECT -7.645 207.235 -7.315 207.565 ;
        RECT -7.645 204.515 -7.315 204.845 ;
        RECT -7.645 203.155 -7.315 203.485 ;
        RECT -7.645 199.075 -7.315 199.405 ;
        RECT -7.645 196.355 -7.315 196.685 ;
        RECT -7.645 189.555 -7.315 189.885 ;
        RECT -7.645 188.195 -7.315 188.525 ;
        RECT -7.645 185.475 -7.315 185.805 ;
        RECT -7.645 178.675 -7.315 179.005 ;
        RECT -7.645 175.955 -7.315 176.285 ;
        RECT -7.645 174.595 -7.315 174.925 ;
        RECT -7.645 167.795 -7.315 168.125 ;
        RECT -7.645 160.995 -7.315 161.325 ;
        RECT -7.645 159.635 -7.315 159.965 ;
        RECT -7.645 156.915 -7.315 157.245 ;
        RECT -7.645 150.115 -7.315 150.445 ;
        RECT -7.645 147.395 -7.315 147.725 ;
        RECT -7.645 146.035 -7.315 146.365 ;
        RECT -7.645 139.235 -7.315 139.565 ;
        RECT -7.645 136.515 -7.315 136.845 ;
        RECT -7.645 132.435 -7.315 132.765 ;
        RECT -7.645 131.075 -7.315 131.405 ;
        RECT -7.645 128.355 -7.315 128.685 ;
        RECT -7.645 118.835 -7.315 119.165 ;
        RECT -7.645 117.475 -7.315 117.805 ;
        RECT -7.645 110.675 -7.315 111.005 ;
        RECT -7.645 107.955 -7.315 108.285 ;
        RECT -7.645 103.875 -7.315 104.205 ;
        RECT -7.645 99.795 -7.315 100.125 ;
        RECT -7.645 97.075 -7.315 97.405 ;
        RECT -7.645 90.275 -7.315 90.605 ;
        RECT -7.645 88.915 -7.315 89.245 ;
        RECT -7.645 82.115 -7.315 82.445 ;
        RECT -7.645 79.395 -7.315 79.725 ;
        RECT -7.645 75.315 -7.315 75.645 ;
        RECT -7.645 71.235 -7.315 71.565 ;
        RECT -7.645 68.515 -7.315 68.845 ;
        RECT -7.645 61.715 -7.315 62.045 ;
        RECT -7.645 60.355 -7.315 60.685 ;
        RECT -7.645 50.835 -7.315 51.165 ;
        RECT -7.645 46.755 -7.315 47.085 ;
        RECT -7.645 42.675 -7.315 43.005 ;
        RECT -7.645 39.955 -7.315 40.285 ;
        RECT -7.645 33.155 -7.315 33.485 ;
        RECT -7.645 31.795 -7.315 32.125 ;
        RECT -7.645 29.075 -7.315 29.405 ;
        RECT -7.645 22.275 -7.315 22.605 ;
        RECT -7.645 19.555 -7.315 19.885 ;
        RECT -7.645 18.195 -7.315 18.525 ;
        RECT -7.645 11.395 -7.315 11.725 ;
        RECT -7.645 4.595 -7.315 4.925 ;
        RECT -7.645 3.235 -7.315 3.565 ;
        RECT -7.645 1.875 -7.315 2.205 ;
        RECT -7.645 0.515 -7.315 0.845 ;
        RECT -7.645 -0.845 -7.315 -0.515 ;
        RECT -7.645 -2.205 -7.315 -1.875 ;
        RECT -7.645 -3.565 -7.315 -3.235 ;
        RECT -7.645 -4.925 -7.315 -4.595 ;
        RECT -7.645 -6.285 -7.315 -5.955 ;
        RECT -7.645 -7.645 -7.315 -7.315 ;
        RECT -7.645 -9.005 -7.315 -8.675 ;
        RECT -7.645 -10.365 -7.315 -10.035 ;
        RECT -7.645 -11.725 -7.315 -11.395 ;
        RECT -7.645 -13.085 -7.315 -12.755 ;
        RECT -7.645 -14.445 -7.315 -14.115 ;
        RECT -7.645 -15.805 -7.315 -15.475 ;
        RECT -7.645 -17.165 -7.315 -16.835 ;
        RECT -7.645 -18.525 -7.315 -18.195 ;
        RECT -7.645 -19.885 -7.315 -19.555 ;
        RECT -7.645 -21.245 -7.315 -20.915 ;
        RECT -7.645 -22.605 -7.315 -22.275 ;
        RECT -7.645 -23.965 -7.315 -23.635 ;
        RECT -7.645 -25.325 -7.315 -24.995 ;
        RECT -7.645 -26.685 -7.315 -26.355 ;
        RECT -7.645 -28.045 -7.315 -27.715 ;
        RECT -7.645 -29.405 -7.315 -29.075 ;
        RECT -7.645 -30.765 -7.315 -30.435 ;
        RECT -7.645 -32.125 -7.315 -31.795 ;
        RECT -7.645 -33.485 -7.315 -33.155 ;
        RECT -7.645 -34.845 -7.315 -34.515 ;
        RECT -7.645 -36.205 -7.315 -35.875 ;
        RECT -7.645 -37.565 -7.315 -37.235 ;
        RECT -7.645 -38.925 -7.315 -38.595 ;
        RECT -7.645 -40.285 -7.315 -39.955 ;
        RECT -7.645 -41.645 -7.315 -41.315 ;
        RECT -7.645 -43.005 -7.315 -42.675 ;
        RECT -7.645 -44.365 -7.315 -44.035 ;
        RECT -7.645 -45.725 -7.315 -45.395 ;
        RECT -7.645 -47.085 -7.315 -46.755 ;
        RECT -7.645 -48.445 -7.315 -48.115 ;
        RECT -7.645 -49.805 -7.315 -49.475 ;
        RECT -7.645 -51.165 -7.315 -50.835 ;
        RECT -7.645 -52.525 -7.315 -52.195 ;
        RECT -7.645 -53.885 -7.315 -53.555 ;
        RECT -7.645 -55.245 -7.315 -54.915 ;
        RECT -7.645 -56.605 -7.315 -56.275 ;
        RECT -7.645 -57.965 -7.315 -57.635 ;
        RECT -7.645 -59.325 -7.315 -58.995 ;
        RECT -7.645 -60.685 -7.315 -60.355 ;
        RECT -7.645 -62.045 -7.315 -61.715 ;
        RECT -7.645 -68.845 -7.315 -68.515 ;
        RECT -7.645 -70.205 -7.315 -69.875 ;
        RECT -7.645 -72.925 -7.315 -72.595 ;
        RECT -7.645 -74.285 -7.315 -73.955 ;
        RECT -7.645 -75.645 -7.315 -75.315 ;
        RECT -7.645 -77.005 -7.315 -76.675 ;
        RECT -7.645 -78.365 -7.315 -78.035 ;
        RECT -7.645 -79.725 -7.315 -79.395 ;
        RECT -7.645 -81.085 -7.315 -80.755 ;
        RECT -7.645 -82.445 -7.315 -82.115 ;
        RECT -7.645 -83.805 -7.315 -83.475 ;
        RECT -7.645 -85.165 -7.315 -84.835 ;
        RECT -7.645 -86.525 -7.315 -86.195 ;
        RECT -7.645 -87.885 -7.315 -87.555 ;
        RECT -7.645 -89.245 -7.315 -88.915 ;
        RECT -7.645 -90.605 -7.315 -90.275 ;
        RECT -7.645 -91.965 -7.315 -91.635 ;
        RECT -7.645 -93.325 -7.315 -92.995 ;
        RECT -7.645 -94.685 -7.315 -94.355 ;
        RECT -7.645 -96.045 -7.315 -95.715 ;
        RECT -7.645 -97.405 -7.315 -97.075 ;
        RECT -7.645 -98.765 -7.315 -98.435 ;
        RECT -7.645 -100.125 -7.315 -99.795 ;
        RECT -7.645 -101.485 -7.315 -101.155 ;
        RECT -7.645 -102.845 -7.315 -102.515 ;
        RECT -7.645 -104.205 -7.315 -103.875 ;
        RECT -7.645 -105.565 -7.315 -105.235 ;
        RECT -7.645 -106.925 -7.315 -106.595 ;
        RECT -7.645 -108.285 -7.315 -107.955 ;
        RECT -7.645 -109.645 -7.315 -109.315 ;
        RECT -7.645 -111.005 -7.315 -110.675 ;
        RECT -7.645 -112.365 -7.315 -112.035 ;
        RECT -7.645 -113.725 -7.315 -113.395 ;
        RECT -7.645 -115.085 -7.315 -114.755 ;
        RECT -7.645 -116.445 -7.315 -116.115 ;
        RECT -7.645 -119.165 -7.315 -118.835 ;
        RECT -7.645 -120.525 -7.315 -120.195 ;
        RECT -7.645 -121.885 -7.315 -121.555 ;
        RECT -7.645 -123.245 -7.315 -122.915 ;
        RECT -7.645 -124.605 -7.315 -124.275 ;
        RECT -7.645 -125.965 -7.315 -125.635 ;
        RECT -7.645 -127.325 -7.315 -126.995 ;
        RECT -7.645 -128.685 -7.315 -128.355 ;
        RECT -7.645 -130.045 -7.315 -129.715 ;
        RECT -7.645 -131.405 -7.315 -131.075 ;
        RECT -7.645 -132.765 -7.315 -132.435 ;
        RECT -7.645 -134.125 -7.315 -133.795 ;
        RECT -7.645 -140.925 -7.315 -140.595 ;
        RECT -7.645 -142.285 -7.315 -141.955 ;
        RECT -7.645 -143.645 -7.315 -143.315 ;
        RECT -7.645 -145.005 -7.315 -144.675 ;
        RECT -7.645 -146.365 -7.315 -146.035 ;
        RECT -7.645 -147.725 -7.315 -147.395 ;
        RECT -7.645 -149.085 -7.315 -148.755 ;
        RECT -7.645 -150.445 -7.315 -150.115 ;
        RECT -7.645 -151.805 -7.315 -151.475 ;
        RECT -7.645 -153.165 -7.315 -152.835 ;
        RECT -7.645 -154.525 -7.315 -154.195 ;
        RECT -7.645 -155.885 -7.315 -155.555 ;
        RECT -7.645 -157.245 -7.315 -156.915 ;
        RECT -7.645 -158.605 -7.315 -158.275 ;
        RECT -7.645 -159.965 -7.315 -159.635 ;
        RECT -7.645 -161.325 -7.315 -160.995 ;
        RECT -7.645 -162.685 -7.315 -162.355 ;
        RECT -7.645 -164.045 -7.315 -163.715 ;
        RECT -7.645 -165.405 -7.315 -165.075 ;
        RECT -7.645 -166.765 -7.315 -166.435 ;
        RECT -7.645 -168.125 -7.315 -167.795 ;
        RECT -7.645 -169.485 -7.315 -169.155 ;
        RECT -7.645 -170.845 -7.315 -170.515 ;
        RECT -7.645 -172.205 -7.315 -171.875 ;
        RECT -7.645 -173.565 -7.315 -173.235 ;
        RECT -7.645 -174.925 -7.315 -174.595 ;
        RECT -7.645 -176.285 -7.315 -175.955 ;
        RECT -7.645 -177.645 -7.315 -177.315 ;
        RECT -7.645 -179.005 -7.315 -178.675 ;
        RECT -7.645 -180.365 -7.315 -180.035 ;
        RECT -7.645 -181.725 -7.315 -181.395 ;
        RECT -7.645 -183.085 -7.315 -182.755 ;
        RECT -7.645 -184.445 -7.315 -184.115 ;
        RECT -7.645 -185.805 -7.315 -185.475 ;
        RECT -7.645 -187.165 -7.315 -186.835 ;
        RECT -7.645 -188.525 -7.315 -188.195 ;
        RECT -7.645 -189.885 -7.315 -189.555 ;
        RECT -7.645 -191.245 -7.315 -190.915 ;
        RECT -7.645 -192.605 -7.315 -192.275 ;
        RECT -7.645 -193.965 -7.315 -193.635 ;
        RECT -7.645 -195.325 -7.315 -194.995 ;
        RECT -7.645 -196.685 -7.315 -196.355 ;
        RECT -7.645 -198.045 -7.315 -197.715 ;
        RECT -7.645 -199.405 -7.315 -199.075 ;
        RECT -7.645 -200.765 -7.315 -200.435 ;
        RECT -7.645 -202.125 -7.315 -201.795 ;
        RECT -7.645 -203.485 -7.315 -203.155 ;
        RECT -7.645 -204.845 -7.315 -204.515 ;
        RECT -7.645 -206.205 -7.315 -205.875 ;
        RECT -7.645 -207.565 -7.315 -207.235 ;
        RECT -7.645 -208.925 -7.315 -208.595 ;
        RECT -7.645 -210.285 -7.315 -209.955 ;
        RECT -7.645 -211.645 -7.315 -211.315 ;
        RECT -7.645 -213.005 -7.315 -212.675 ;
        RECT -7.645 -214.365 -7.315 -214.035 ;
        RECT -7.645 -215.725 -7.315 -215.395 ;
        RECT -7.645 -217.085 -7.315 -216.755 ;
        RECT -7.645 -218.445 -7.315 -218.115 ;
        RECT -7.645 -219.805 -7.315 -219.475 ;
        RECT -7.645 -221.165 -7.315 -220.835 ;
        RECT -7.645 -222.525 -7.315 -222.195 ;
        RECT -7.645 -223.885 -7.315 -223.555 ;
        RECT -7.645 -225.245 -7.315 -224.915 ;
        RECT -7.645 -226.605 -7.315 -226.275 ;
        RECT -7.645 -227.965 -7.315 -227.635 ;
        RECT -7.645 -229.325 -7.315 -228.995 ;
        RECT -7.645 -230.685 -7.315 -230.355 ;
        RECT -7.645 -232.045 -7.315 -231.715 ;
        RECT -7.645 -233.405 -7.315 -233.075 ;
        RECT -7.645 -234.765 -7.315 -234.435 ;
        RECT -7.645 -236.125 -7.315 -235.795 ;
        RECT -7.645 -237.485 -7.315 -237.155 ;
        RECT -7.645 -238.845 -7.315 -238.515 ;
        RECT -7.645 -241.09 -7.315 -239.96 ;
        RECT -7.64 -241.205 -7.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.285 244.04 -5.955 245.17 ;
        RECT -6.285 242.595 -5.955 242.925 ;
        RECT -6.285 241.235 -5.955 241.565 ;
        RECT -6.285 239.875 -5.955 240.205 ;
        RECT -6.285 238.515 -5.955 238.845 ;
        RECT -6.285 237.155 -5.955 237.485 ;
        RECT -6.285 -0.845 -5.955 -0.515 ;
        RECT -6.285 -2.205 -5.955 -1.875 ;
        RECT -6.285 -3.565 -5.955 -3.235 ;
        RECT -6.285 -4.925 -5.955 -4.595 ;
        RECT -6.285 -6.285 -5.955 -5.955 ;
        RECT -6.285 -7.645 -5.955 -7.315 ;
        RECT -6.285 -9.005 -5.955 -8.675 ;
        RECT -6.285 -10.365 -5.955 -10.035 ;
        RECT -6.285 -11.725 -5.955 -11.395 ;
        RECT -6.285 -13.085 -5.955 -12.755 ;
        RECT -6.285 -14.445 -5.955 -14.115 ;
        RECT -6.285 -15.805 -5.955 -15.475 ;
        RECT -6.285 -17.165 -5.955 -16.835 ;
        RECT -6.285 -18.525 -5.955 -18.195 ;
        RECT -6.285 -19.885 -5.955 -19.555 ;
        RECT -6.285 -21.245 -5.955 -20.915 ;
        RECT -6.285 -22.605 -5.955 -22.275 ;
        RECT -6.285 -23.965 -5.955 -23.635 ;
        RECT -6.285 -25.325 -5.955 -24.995 ;
        RECT -6.285 -26.685 -5.955 -26.355 ;
        RECT -6.285 -28.045 -5.955 -27.715 ;
        RECT -6.285 -29.405 -5.955 -29.075 ;
        RECT -6.285 -30.765 -5.955 -30.435 ;
        RECT -6.285 -32.125 -5.955 -31.795 ;
        RECT -6.285 -33.485 -5.955 -33.155 ;
        RECT -6.285 -34.845 -5.955 -34.515 ;
        RECT -6.285 -36.205 -5.955 -35.875 ;
        RECT -6.285 -37.565 -5.955 -37.235 ;
        RECT -6.285 -38.925 -5.955 -38.595 ;
        RECT -6.285 -40.285 -5.955 -39.955 ;
        RECT -6.285 -41.645 -5.955 -41.315 ;
        RECT -6.285 -43.005 -5.955 -42.675 ;
        RECT -6.285 -44.365 -5.955 -44.035 ;
        RECT -6.285 -45.725 -5.955 -45.395 ;
        RECT -6.285 -47.085 -5.955 -46.755 ;
        RECT -6.285 -48.445 -5.955 -48.115 ;
        RECT -6.285 -49.805 -5.955 -49.475 ;
        RECT -6.285 -51.165 -5.955 -50.835 ;
        RECT -6.285 -52.525 -5.955 -52.195 ;
        RECT -6.285 -53.885 -5.955 -53.555 ;
        RECT -6.285 -55.245 -5.955 -54.915 ;
        RECT -6.285 -56.605 -5.955 -56.275 ;
        RECT -6.285 -57.965 -5.955 -57.635 ;
        RECT -6.285 -59.325 -5.955 -58.995 ;
        RECT -6.285 -60.685 -5.955 -60.355 ;
        RECT -6.285 -62.045 -5.955 -61.715 ;
        RECT -6.285 -68.845 -5.955 -68.515 ;
        RECT -6.285 -70.205 -5.955 -69.875 ;
        RECT -6.285 -72.925 -5.955 -72.595 ;
        RECT -6.285 -74.285 -5.955 -73.955 ;
        RECT -6.285 -75.645 -5.955 -75.315 ;
        RECT -6.285 -77.005 -5.955 -76.675 ;
        RECT -6.285 -78.365 -5.955 -78.035 ;
        RECT -6.285 -79.725 -5.955 -79.395 ;
        RECT -6.285 -81.085 -5.955 -80.755 ;
        RECT -6.285 -82.445 -5.955 -82.115 ;
        RECT -6.285 -83.805 -5.955 -83.475 ;
        RECT -6.285 -85.165 -5.955 -84.835 ;
        RECT -6.285 -86.525 -5.955 -86.195 ;
        RECT -6.285 -87.885 -5.955 -87.555 ;
        RECT -6.285 -89.245 -5.955 -88.915 ;
        RECT -6.285 -90.605 -5.955 -90.275 ;
        RECT -6.285 -91.965 -5.955 -91.635 ;
        RECT -6.285 -93.325 -5.955 -92.995 ;
        RECT -6.285 -94.685 -5.955 -94.355 ;
        RECT -6.285 -96.045 -5.955 -95.715 ;
        RECT -6.285 -97.405 -5.955 -97.075 ;
        RECT -6.285 -98.765 -5.955 -98.435 ;
        RECT -6.285 -100.125 -5.955 -99.795 ;
        RECT -6.285 -101.485 -5.955 -101.155 ;
        RECT -6.285 -102.845 -5.955 -102.515 ;
        RECT -6.285 -104.205 -5.955 -103.875 ;
        RECT -6.285 -105.565 -5.955 -105.235 ;
        RECT -6.285 -106.925 -5.955 -106.595 ;
        RECT -6.285 -108.285 -5.955 -107.955 ;
        RECT -6.285 -109.645 -5.955 -109.315 ;
        RECT -6.285 -111.005 -5.955 -110.675 ;
        RECT -6.285 -112.365 -5.955 -112.035 ;
        RECT -6.285 -113.725 -5.955 -113.395 ;
        RECT -6.285 -115.085 -5.955 -114.755 ;
        RECT -6.285 -116.445 -5.955 -116.115 ;
        RECT -6.285 -119.165 -5.955 -118.835 ;
        RECT -6.285 -120.525 -5.955 -120.195 ;
        RECT -6.285 -121.885 -5.955 -121.555 ;
        RECT -6.285 -123.245 -5.955 -122.915 ;
        RECT -6.285 -124.605 -5.955 -124.275 ;
        RECT -6.285 -125.965 -5.955 -125.635 ;
        RECT -6.285 -127.325 -5.955 -126.995 ;
        RECT -6.285 -128.685 -5.955 -128.355 ;
        RECT -6.285 -130.045 -5.955 -129.715 ;
        RECT -6.285 -131.405 -5.955 -131.075 ;
        RECT -6.285 -132.765 -5.955 -132.435 ;
        RECT -6.285 -134.125 -5.955 -133.795 ;
        RECT -6.285 -140.925 -5.955 -140.595 ;
        RECT -6.285 -142.285 -5.955 -141.955 ;
        RECT -6.285 -143.645 -5.955 -143.315 ;
        RECT -6.285 -145.005 -5.955 -144.675 ;
        RECT -6.285 -146.365 -5.955 -146.035 ;
        RECT -6.285 -147.725 -5.955 -147.395 ;
        RECT -6.285 -149.085 -5.955 -148.755 ;
        RECT -6.285 -150.445 -5.955 -150.115 ;
        RECT -6.285 -151.805 -5.955 -151.475 ;
        RECT -6.285 -153.165 -5.955 -152.835 ;
        RECT -6.285 -154.525 -5.955 -154.195 ;
        RECT -6.285 -155.885 -5.955 -155.555 ;
        RECT -6.285 -157.245 -5.955 -156.915 ;
        RECT -6.285 -158.605 -5.955 -158.275 ;
        RECT -6.285 -159.965 -5.955 -159.635 ;
        RECT -6.285 -161.325 -5.955 -160.995 ;
        RECT -6.285 -162.685 -5.955 -162.355 ;
        RECT -6.285 -164.045 -5.955 -163.715 ;
        RECT -6.285 -165.405 -5.955 -165.075 ;
        RECT -6.285 -166.765 -5.955 -166.435 ;
        RECT -6.285 -168.125 -5.955 -167.795 ;
        RECT -6.285 -169.485 -5.955 -169.155 ;
        RECT -6.285 -170.845 -5.955 -170.515 ;
        RECT -6.285 -172.205 -5.955 -171.875 ;
        RECT -6.285 -173.565 -5.955 -173.235 ;
        RECT -6.285 -174.925 -5.955 -174.595 ;
        RECT -6.285 -176.285 -5.955 -175.955 ;
        RECT -6.285 -177.645 -5.955 -177.315 ;
        RECT -6.285 -179.005 -5.955 -178.675 ;
        RECT -6.285 -180.365 -5.955 -180.035 ;
        RECT -6.285 -181.725 -5.955 -181.395 ;
        RECT -6.285 -183.085 -5.955 -182.755 ;
        RECT -6.285 -184.445 -5.955 -184.115 ;
        RECT -6.285 -185.805 -5.955 -185.475 ;
        RECT -6.285 -187.165 -5.955 -186.835 ;
        RECT -6.285 -188.525 -5.955 -188.195 ;
        RECT -6.285 -189.885 -5.955 -189.555 ;
        RECT -6.285 -191.245 -5.955 -190.915 ;
        RECT -6.285 -192.605 -5.955 -192.275 ;
        RECT -6.285 -193.965 -5.955 -193.635 ;
        RECT -6.285 -195.325 -5.955 -194.995 ;
        RECT -6.285 -196.685 -5.955 -196.355 ;
        RECT -6.285 -198.045 -5.955 -197.715 ;
        RECT -6.285 -199.405 -5.955 -199.075 ;
        RECT -6.285 -200.765 -5.955 -200.435 ;
        RECT -6.285 -202.125 -5.955 -201.795 ;
        RECT -6.285 -203.485 -5.955 -203.155 ;
        RECT -6.285 -204.845 -5.955 -204.515 ;
        RECT -6.285 -206.205 -5.955 -205.875 ;
        RECT -6.285 -207.565 -5.955 -207.235 ;
        RECT -6.285 -208.925 -5.955 -208.595 ;
        RECT -6.285 -210.285 -5.955 -209.955 ;
        RECT -6.285 -211.645 -5.955 -211.315 ;
        RECT -6.285 -213.005 -5.955 -212.675 ;
        RECT -6.285 -214.365 -5.955 -214.035 ;
        RECT -6.285 -215.725 -5.955 -215.395 ;
        RECT -6.285 -217.085 -5.955 -216.755 ;
        RECT -6.285 -218.445 -5.955 -218.115 ;
        RECT -6.285 -219.805 -5.955 -219.475 ;
        RECT -6.285 -221.165 -5.955 -220.835 ;
        RECT -6.285 -222.525 -5.955 -222.195 ;
        RECT -6.285 -223.885 -5.955 -223.555 ;
        RECT -6.285 -225.245 -5.955 -224.915 ;
        RECT -6.285 -226.605 -5.955 -226.275 ;
        RECT -6.285 -227.965 -5.955 -227.635 ;
        RECT -6.285 -229.325 -5.955 -228.995 ;
        RECT -6.285 -230.685 -5.955 -230.355 ;
        RECT -6.285 -232.045 -5.955 -231.715 ;
        RECT -6.285 -233.405 -5.955 -233.075 ;
        RECT -6.285 -234.765 -5.955 -234.435 ;
        RECT -6.285 -236.125 -5.955 -235.795 ;
        RECT -6.285 -237.485 -5.955 -237.155 ;
        RECT -6.285 -238.845 -5.955 -238.515 ;
        RECT -6.285 -241.09 -5.955 -239.96 ;
        RECT -6.28 -241.205 -5.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.925 244.04 -4.595 245.17 ;
        RECT -4.925 242.595 -4.595 242.925 ;
        RECT -4.925 241.235 -4.595 241.565 ;
        RECT -4.925 239.875 -4.595 240.205 ;
        RECT -4.925 238.515 -4.595 238.845 ;
        RECT -4.925 237.155 -4.595 237.485 ;
        RECT -4.925 235.975 -4.595 236.305 ;
        RECT -4.925 233.925 -4.595 234.255 ;
        RECT -4.925 231.995 -4.595 232.325 ;
        RECT -4.925 230.155 -4.595 230.485 ;
        RECT -4.925 228.665 -4.595 228.995 ;
        RECT -4.925 226.995 -4.595 227.325 ;
        RECT -4.925 225.505 -4.595 225.835 ;
        RECT -4.925 223.835 -4.595 224.165 ;
        RECT -4.925 222.345 -4.595 222.675 ;
        RECT -4.925 220.675 -4.595 221.005 ;
        RECT -4.925 219.185 -4.595 219.515 ;
        RECT -4.925 217.775 -4.595 218.105 ;
        RECT -4.925 215.935 -4.595 216.265 ;
        RECT -4.925 214.445 -4.595 214.775 ;
        RECT -4.925 212.775 -4.595 213.105 ;
        RECT -4.925 211.285 -4.595 211.615 ;
        RECT -4.925 209.615 -4.595 209.945 ;
        RECT -4.925 208.125 -4.595 208.455 ;
        RECT -4.925 206.455 -4.595 206.785 ;
        RECT -4.925 204.965 -4.595 205.295 ;
        RECT -4.925 203.555 -4.595 203.885 ;
        RECT -4.925 201.715 -4.595 202.045 ;
        RECT -4.925 200.225 -4.595 200.555 ;
        RECT -4.925 198.555 -4.595 198.885 ;
        RECT -4.925 197.065 -4.595 197.395 ;
        RECT -4.925 195.395 -4.595 195.725 ;
        RECT -4.925 193.905 -4.595 194.235 ;
        RECT -4.925 192.235 -4.595 192.565 ;
        RECT -4.925 190.745 -4.595 191.075 ;
        RECT -4.925 189.335 -4.595 189.665 ;
        RECT -4.925 187.495 -4.595 187.825 ;
        RECT -4.925 186.005 -4.595 186.335 ;
        RECT -4.925 184.335 -4.595 184.665 ;
        RECT -4.925 182.845 -4.595 183.175 ;
        RECT -4.925 181.175 -4.595 181.505 ;
        RECT -4.925 179.685 -4.595 180.015 ;
        RECT -4.925 178.015 -4.595 178.345 ;
        RECT -4.925 176.525 -4.595 176.855 ;
        RECT -4.925 175.115 -4.595 175.445 ;
        RECT -4.925 173.275 -4.595 173.605 ;
        RECT -4.925 171.785 -4.595 172.115 ;
        RECT -4.925 170.115 -4.595 170.445 ;
        RECT -4.925 168.625 -4.595 168.955 ;
        RECT -4.925 166.955 -4.595 167.285 ;
        RECT -4.925 165.465 -4.595 165.795 ;
        RECT -4.925 163.795 -4.595 164.125 ;
        RECT -4.925 162.305 -4.595 162.635 ;
        RECT -4.925 160.895 -4.595 161.225 ;
        RECT -4.925 159.055 -4.595 159.385 ;
        RECT -4.925 157.565 -4.595 157.895 ;
        RECT -4.925 155.895 -4.595 156.225 ;
        RECT -4.925 154.405 -4.595 154.735 ;
        RECT -4.925 152.735 -4.595 153.065 ;
        RECT -4.925 151.245 -4.595 151.575 ;
        RECT -4.925 149.575 -4.595 149.905 ;
        RECT -4.925 148.085 -4.595 148.415 ;
        RECT -4.925 146.675 -4.595 147.005 ;
        RECT -4.925 144.835 -4.595 145.165 ;
        RECT -4.925 143.345 -4.595 143.675 ;
        RECT -4.925 141.675 -4.595 142.005 ;
        RECT -4.925 140.185 -4.595 140.515 ;
        RECT -4.925 138.515 -4.595 138.845 ;
        RECT -4.925 137.025 -4.595 137.355 ;
        RECT -4.925 135.355 -4.595 135.685 ;
        RECT -4.925 133.865 -4.595 134.195 ;
        RECT -4.925 132.455 -4.595 132.785 ;
        RECT -4.925 130.615 -4.595 130.945 ;
        RECT -4.925 129.125 -4.595 129.455 ;
        RECT -4.925 127.455 -4.595 127.785 ;
        RECT -4.925 125.965 -4.595 126.295 ;
        RECT -4.925 124.295 -4.595 124.625 ;
        RECT -4.925 122.805 -4.595 123.135 ;
        RECT -4.925 121.135 -4.595 121.465 ;
        RECT -4.925 119.645 -4.595 119.975 ;
        RECT -4.925 118.235 -4.595 118.565 ;
        RECT -4.925 116.395 -4.595 116.725 ;
        RECT -4.925 114.905 -4.595 115.235 ;
        RECT -4.925 113.235 -4.595 113.565 ;
        RECT -4.925 111.745 -4.595 112.075 ;
        RECT -4.925 110.075 -4.595 110.405 ;
        RECT -4.925 108.585 -4.595 108.915 ;
        RECT -4.925 106.915 -4.595 107.245 ;
        RECT -4.925 105.425 -4.595 105.755 ;
        RECT -4.925 104.015 -4.595 104.345 ;
        RECT -4.925 102.175 -4.595 102.505 ;
        RECT -4.925 100.685 -4.595 101.015 ;
        RECT -4.925 99.015 -4.595 99.345 ;
        RECT -4.925 97.525 -4.595 97.855 ;
        RECT -4.925 95.855 -4.595 96.185 ;
        RECT -4.925 94.365 -4.595 94.695 ;
        RECT -4.925 92.695 -4.595 93.025 ;
        RECT -4.925 91.205 -4.595 91.535 ;
        RECT -4.925 89.795 -4.595 90.125 ;
        RECT -4.925 87.955 -4.595 88.285 ;
        RECT -4.925 86.465 -4.595 86.795 ;
        RECT -4.925 84.795 -4.595 85.125 ;
        RECT -4.925 83.305 -4.595 83.635 ;
        RECT -4.925 81.635 -4.595 81.965 ;
        RECT -4.925 80.145 -4.595 80.475 ;
        RECT -4.925 78.475 -4.595 78.805 ;
        RECT -4.925 76.985 -4.595 77.315 ;
        RECT -4.925 75.575 -4.595 75.905 ;
        RECT -4.925 73.735 -4.595 74.065 ;
        RECT -4.925 72.245 -4.595 72.575 ;
        RECT -4.925 70.575 -4.595 70.905 ;
        RECT -4.925 69.085 -4.595 69.415 ;
        RECT -4.925 67.415 -4.595 67.745 ;
        RECT -4.925 65.925 -4.595 66.255 ;
        RECT -4.925 64.255 -4.595 64.585 ;
        RECT -4.925 62.765 -4.595 63.095 ;
        RECT -4.925 61.355 -4.595 61.685 ;
        RECT -4.925 59.515 -4.595 59.845 ;
        RECT -4.925 58.025 -4.595 58.355 ;
        RECT -4.925 56.355 -4.595 56.685 ;
        RECT -4.925 54.865 -4.595 55.195 ;
        RECT -4.925 53.195 -4.595 53.525 ;
        RECT -4.925 51.705 -4.595 52.035 ;
        RECT -4.925 50.035 -4.595 50.365 ;
        RECT -4.925 48.545 -4.595 48.875 ;
        RECT -4.925 47.135 -4.595 47.465 ;
        RECT -4.925 45.295 -4.595 45.625 ;
        RECT -4.925 43.805 -4.595 44.135 ;
        RECT -4.925 42.135 -4.595 42.465 ;
        RECT -4.925 40.645 -4.595 40.975 ;
        RECT -4.925 38.975 -4.595 39.305 ;
        RECT -4.925 37.485 -4.595 37.815 ;
        RECT -4.925 35.815 -4.595 36.145 ;
        RECT -4.925 34.325 -4.595 34.655 ;
        RECT -4.925 32.915 -4.595 33.245 ;
        RECT -4.925 31.075 -4.595 31.405 ;
        RECT -4.925 29.585 -4.595 29.915 ;
        RECT -4.925 27.915 -4.595 28.245 ;
        RECT -4.925 26.425 -4.595 26.755 ;
        RECT -4.925 24.755 -4.595 25.085 ;
        RECT -4.925 23.265 -4.595 23.595 ;
        RECT -4.925 21.595 -4.595 21.925 ;
        RECT -4.925 20.105 -4.595 20.435 ;
        RECT -4.925 18.695 -4.595 19.025 ;
        RECT -4.925 16.855 -4.595 17.185 ;
        RECT -4.925 15.365 -4.595 15.695 ;
        RECT -4.925 13.695 -4.595 14.025 ;
        RECT -4.925 12.205 -4.595 12.535 ;
        RECT -4.925 10.535 -4.595 10.865 ;
        RECT -4.925 9.045 -4.595 9.375 ;
        RECT -4.925 7.375 -4.595 7.705 ;
        RECT -4.925 5.885 -4.595 6.215 ;
        RECT -4.925 4.475 -4.595 4.805 ;
        RECT -4.925 2.115 -4.595 2.445 ;
        RECT -4.925 0.06 -4.595 0.39 ;
        RECT -4.925 -0.845 -4.595 -0.515 ;
        RECT -4.925 -2.205 -4.595 -1.875 ;
        RECT -4.925 -3.565 -4.595 -3.235 ;
        RECT -4.925 -4.925 -4.595 -4.595 ;
        RECT -4.925 -6.285 -4.595 -5.955 ;
        RECT -4.925 -7.645 -4.595 -7.315 ;
        RECT -4.925 -9.005 -4.595 -8.675 ;
        RECT -4.925 -10.365 -4.595 -10.035 ;
        RECT -4.925 -11.725 -4.595 -11.395 ;
        RECT -4.925 -13.085 -4.595 -12.755 ;
        RECT -4.925 -14.445 -4.595 -14.115 ;
        RECT -4.925 -15.805 -4.595 -15.475 ;
        RECT -4.925 -17.165 -4.595 -16.835 ;
        RECT -4.925 -18.525 -4.595 -18.195 ;
        RECT -4.925 -19.885 -4.595 -19.555 ;
        RECT -4.925 -21.245 -4.595 -20.915 ;
        RECT -4.925 -22.605 -4.595 -22.275 ;
        RECT -4.925 -23.965 -4.595 -23.635 ;
        RECT -4.925 -25.325 -4.595 -24.995 ;
        RECT -4.925 -26.685 -4.595 -26.355 ;
        RECT -4.925 -28.045 -4.595 -27.715 ;
        RECT -4.925 -29.405 -4.595 -29.075 ;
        RECT -4.925 -30.765 -4.595 -30.435 ;
        RECT -4.925 -32.125 -4.595 -31.795 ;
        RECT -4.925 -33.485 -4.595 -33.155 ;
        RECT -4.925 -34.845 -4.595 -34.515 ;
        RECT -4.925 -36.205 -4.595 -35.875 ;
        RECT -4.925 -37.565 -4.595 -37.235 ;
        RECT -4.925 -38.925 -4.595 -38.595 ;
        RECT -4.925 -40.285 -4.595 -39.955 ;
        RECT -4.925 -41.645 -4.595 -41.315 ;
        RECT -4.925 -43.005 -4.595 -42.675 ;
        RECT -4.925 -44.365 -4.595 -44.035 ;
        RECT -4.925 -45.725 -4.595 -45.395 ;
        RECT -4.925 -47.085 -4.595 -46.755 ;
        RECT -4.925 -48.445 -4.595 -48.115 ;
        RECT -4.925 -49.805 -4.595 -49.475 ;
        RECT -4.925 -51.165 -4.595 -50.835 ;
        RECT -4.925 -52.525 -4.595 -52.195 ;
        RECT -4.925 -53.885 -4.595 -53.555 ;
        RECT -4.925 -55.245 -4.595 -54.915 ;
        RECT -4.925 -56.605 -4.595 -56.275 ;
        RECT -4.925 -57.965 -4.595 -57.635 ;
        RECT -4.925 -59.325 -4.595 -58.995 ;
        RECT -4.925 -60.685 -4.595 -60.355 ;
        RECT -4.925 -62.045 -4.595 -61.715 ;
        RECT -4.925 -68.845 -4.595 -68.515 ;
        RECT -4.925 -70.205 -4.595 -69.875 ;
        RECT -4.925 -72.925 -4.595 -72.595 ;
        RECT -4.925 -74.285 -4.595 -73.955 ;
        RECT -4.925 -75.645 -4.595 -75.315 ;
        RECT -4.925 -77.005 -4.595 -76.675 ;
        RECT -4.925 -78.365 -4.595 -78.035 ;
        RECT -4.925 -79.725 -4.595 -79.395 ;
        RECT -4.925 -81.085 -4.595 -80.755 ;
        RECT -4.925 -82.445 -4.595 -82.115 ;
        RECT -4.925 -83.805 -4.595 -83.475 ;
        RECT -4.925 -85.165 -4.595 -84.835 ;
        RECT -4.925 -86.525 -4.595 -86.195 ;
        RECT -4.925 -87.885 -4.595 -87.555 ;
        RECT -4.925 -89.245 -4.595 -88.915 ;
        RECT -4.925 -90.605 -4.595 -90.275 ;
        RECT -4.925 -91.965 -4.595 -91.635 ;
        RECT -4.925 -93.325 -4.595 -92.995 ;
        RECT -4.925 -94.685 -4.595 -94.355 ;
        RECT -4.925 -96.045 -4.595 -95.715 ;
        RECT -4.925 -97.405 -4.595 -97.075 ;
        RECT -4.925 -98.765 -4.595 -98.435 ;
        RECT -4.925 -100.125 -4.595 -99.795 ;
        RECT -4.925 -101.485 -4.595 -101.155 ;
        RECT -4.925 -102.845 -4.595 -102.515 ;
        RECT -4.925 -104.205 -4.595 -103.875 ;
        RECT -4.925 -105.565 -4.595 -105.235 ;
        RECT -4.925 -106.925 -4.595 -106.595 ;
        RECT -4.925 -108.285 -4.595 -107.955 ;
        RECT -4.925 -109.645 -4.595 -109.315 ;
        RECT -4.925 -111.005 -4.595 -110.675 ;
        RECT -4.925 -112.365 -4.595 -112.035 ;
        RECT -4.925 -113.725 -4.595 -113.395 ;
        RECT -4.925 -115.085 -4.595 -114.755 ;
        RECT -4.925 -116.445 -4.595 -116.115 ;
        RECT -4.925 -119.165 -4.595 -118.835 ;
        RECT -4.925 -120.525 -4.595 -120.195 ;
        RECT -4.925 -121.885 -4.595 -121.555 ;
        RECT -4.925 -123.245 -4.595 -122.915 ;
        RECT -4.925 -124.605 -4.595 -124.275 ;
        RECT -4.925 -125.965 -4.595 -125.635 ;
        RECT -4.925 -127.325 -4.595 -126.995 ;
        RECT -4.925 -128.685 -4.595 -128.355 ;
        RECT -4.925 -130.045 -4.595 -129.715 ;
        RECT -4.925 -131.405 -4.595 -131.075 ;
        RECT -4.925 -132.765 -4.595 -132.435 ;
        RECT -4.925 -134.125 -4.595 -133.795 ;
        RECT -4.925 -140.925 -4.595 -140.595 ;
        RECT -4.925 -142.285 -4.595 -141.955 ;
        RECT -4.925 -143.645 -4.595 -143.315 ;
        RECT -4.925 -145.005 -4.595 -144.675 ;
        RECT -4.925 -146.365 -4.595 -146.035 ;
        RECT -4.925 -147.725 -4.595 -147.395 ;
        RECT -4.925 -149.085 -4.595 -148.755 ;
        RECT -4.925 -150.445 -4.595 -150.115 ;
        RECT -4.925 -151.805 -4.595 -151.475 ;
        RECT -4.925 -153.165 -4.595 -152.835 ;
        RECT -4.925 -154.525 -4.595 -154.195 ;
        RECT -4.925 -155.885 -4.595 -155.555 ;
        RECT -4.925 -157.245 -4.595 -156.915 ;
        RECT -4.925 -158.605 -4.595 -158.275 ;
        RECT -4.925 -159.965 -4.595 -159.635 ;
        RECT -4.925 -161.325 -4.595 -160.995 ;
        RECT -4.925 -162.685 -4.595 -162.355 ;
        RECT -4.925 -164.045 -4.595 -163.715 ;
        RECT -4.925 -165.405 -4.595 -165.075 ;
        RECT -4.925 -166.765 -4.595 -166.435 ;
        RECT -4.925 -168.125 -4.595 -167.795 ;
        RECT -4.925 -169.485 -4.595 -169.155 ;
        RECT -4.925 -170.845 -4.595 -170.515 ;
        RECT -4.925 -172.205 -4.595 -171.875 ;
        RECT -4.925 -173.565 -4.595 -173.235 ;
        RECT -4.925 -174.925 -4.595 -174.595 ;
        RECT -4.925 -176.285 -4.595 -175.955 ;
        RECT -4.925 -177.645 -4.595 -177.315 ;
        RECT -4.925 -179.005 -4.595 -178.675 ;
        RECT -4.925 -180.365 -4.595 -180.035 ;
        RECT -4.925 -181.725 -4.595 -181.395 ;
        RECT -4.925 -183.085 -4.595 -182.755 ;
        RECT -4.925 -184.445 -4.595 -184.115 ;
        RECT -4.925 -185.805 -4.595 -185.475 ;
        RECT -4.925 -187.165 -4.595 -186.835 ;
        RECT -4.925 -188.525 -4.595 -188.195 ;
        RECT -4.925 -189.885 -4.595 -189.555 ;
        RECT -4.925 -191.245 -4.595 -190.915 ;
        RECT -4.925 -192.605 -4.595 -192.275 ;
        RECT -4.925 -193.965 -4.595 -193.635 ;
        RECT -4.925 -195.325 -4.595 -194.995 ;
        RECT -4.925 -196.685 -4.595 -196.355 ;
        RECT -4.925 -198.045 -4.595 -197.715 ;
        RECT -4.925 -199.405 -4.595 -199.075 ;
        RECT -4.925 -200.765 -4.595 -200.435 ;
        RECT -4.925 -202.125 -4.595 -201.795 ;
        RECT -4.925 -203.485 -4.595 -203.155 ;
        RECT -4.925 -204.845 -4.595 -204.515 ;
        RECT -4.925 -206.205 -4.595 -205.875 ;
        RECT -4.925 -207.565 -4.595 -207.235 ;
        RECT -4.925 -208.925 -4.595 -208.595 ;
        RECT -4.925 -210.285 -4.595 -209.955 ;
        RECT -4.925 -211.645 -4.595 -211.315 ;
        RECT -4.925 -213.005 -4.595 -212.675 ;
        RECT -4.925 -214.365 -4.595 -214.035 ;
        RECT -4.925 -215.725 -4.595 -215.395 ;
        RECT -4.925 -217.085 -4.595 -216.755 ;
        RECT -4.925 -218.445 -4.595 -218.115 ;
        RECT -4.925 -219.805 -4.595 -219.475 ;
        RECT -4.925 -221.165 -4.595 -220.835 ;
        RECT -4.925 -222.525 -4.595 -222.195 ;
        RECT -4.925 -223.885 -4.595 -223.555 ;
        RECT -4.925 -225.245 -4.595 -224.915 ;
        RECT -4.925 -226.605 -4.595 -226.275 ;
        RECT -4.925 -227.965 -4.595 -227.635 ;
        RECT -4.925 -229.325 -4.595 -228.995 ;
        RECT -4.925 -230.685 -4.595 -230.355 ;
        RECT -4.925 -232.045 -4.595 -231.715 ;
        RECT -4.925 -233.405 -4.595 -233.075 ;
        RECT -4.925 -234.765 -4.595 -234.435 ;
        RECT -4.925 -236.125 -4.595 -235.795 ;
        RECT -4.925 -237.485 -4.595 -237.155 ;
        RECT -4.925 -238.845 -4.595 -238.515 ;
        RECT -4.925 -241.09 -4.595 -239.96 ;
        RECT -4.92 -241.205 -4.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.565 45.295 -3.235 45.625 ;
        RECT -3.565 43.805 -3.235 44.135 ;
        RECT -3.565 42.135 -3.235 42.465 ;
        RECT -3.565 40.645 -3.235 40.975 ;
        RECT -3.565 38.975 -3.235 39.305 ;
        RECT -3.565 37.485 -3.235 37.815 ;
        RECT -3.565 35.815 -3.235 36.145 ;
        RECT -3.565 34.325 -3.235 34.655 ;
        RECT -3.565 32.915 -3.235 33.245 ;
        RECT -3.565 31.075 -3.235 31.405 ;
        RECT -3.565 29.585 -3.235 29.915 ;
        RECT -3.565 27.915 -3.235 28.245 ;
        RECT -3.565 26.425 -3.235 26.755 ;
        RECT -3.565 24.755 -3.235 25.085 ;
        RECT -3.565 23.265 -3.235 23.595 ;
        RECT -3.565 21.595 -3.235 21.925 ;
        RECT -3.565 20.105 -3.235 20.435 ;
        RECT -3.565 18.695 -3.235 19.025 ;
        RECT -3.565 16.855 -3.235 17.185 ;
        RECT -3.565 15.365 -3.235 15.695 ;
        RECT -3.565 13.695 -3.235 14.025 ;
        RECT -3.565 12.205 -3.235 12.535 ;
        RECT -3.565 10.535 -3.235 10.865 ;
        RECT -3.565 9.045 -3.235 9.375 ;
        RECT -3.565 7.375 -3.235 7.705 ;
        RECT -3.565 5.885 -3.235 6.215 ;
        RECT -3.565 4.475 -3.235 4.805 ;
        RECT -3.565 2.115 -3.235 2.445 ;
        RECT -3.565 0.06 -3.235 0.39 ;
        RECT -3.565 -0.845 -3.235 -0.515 ;
        RECT -3.565 -2.205 -3.235 -1.875 ;
        RECT -3.565 -3.565 -3.235 -3.235 ;
        RECT -3.565 -4.925 -3.235 -4.595 ;
        RECT -3.565 -6.285 -3.235 -5.955 ;
        RECT -3.565 -7.645 -3.235 -7.315 ;
        RECT -3.565 -9.005 -3.235 -8.675 ;
        RECT -3.565 -10.365 -3.235 -10.035 ;
        RECT -3.565 -11.725 -3.235 -11.395 ;
        RECT -3.565 -13.085 -3.235 -12.755 ;
        RECT -3.565 -14.445 -3.235 -14.115 ;
        RECT -3.565 -15.805 -3.235 -15.475 ;
        RECT -3.565 -17.165 -3.235 -16.835 ;
        RECT -3.565 -18.525 -3.235 -18.195 ;
        RECT -3.565 -19.885 -3.235 -19.555 ;
        RECT -3.56 -20.56 -3.24 245.285 ;
        RECT -3.565 244.04 -3.235 245.17 ;
        RECT -3.565 242.595 -3.235 242.925 ;
        RECT -3.565 241.235 -3.235 241.565 ;
        RECT -3.565 239.875 -3.235 240.205 ;
        RECT -3.565 238.515 -3.235 238.845 ;
        RECT -3.565 237.155 -3.235 237.485 ;
        RECT -3.565 235.975 -3.235 236.305 ;
        RECT -3.565 233.925 -3.235 234.255 ;
        RECT -3.565 231.995 -3.235 232.325 ;
        RECT -3.565 230.155 -3.235 230.485 ;
        RECT -3.565 228.665 -3.235 228.995 ;
        RECT -3.565 226.995 -3.235 227.325 ;
        RECT -3.565 225.505 -3.235 225.835 ;
        RECT -3.565 223.835 -3.235 224.165 ;
        RECT -3.565 222.345 -3.235 222.675 ;
        RECT -3.565 220.675 -3.235 221.005 ;
        RECT -3.565 219.185 -3.235 219.515 ;
        RECT -3.565 217.775 -3.235 218.105 ;
        RECT -3.565 215.935 -3.235 216.265 ;
        RECT -3.565 214.445 -3.235 214.775 ;
        RECT -3.565 212.775 -3.235 213.105 ;
        RECT -3.565 211.285 -3.235 211.615 ;
        RECT -3.565 209.615 -3.235 209.945 ;
        RECT -3.565 208.125 -3.235 208.455 ;
        RECT -3.565 206.455 -3.235 206.785 ;
        RECT -3.565 204.965 -3.235 205.295 ;
        RECT -3.565 203.555 -3.235 203.885 ;
        RECT -3.565 201.715 -3.235 202.045 ;
        RECT -3.565 200.225 -3.235 200.555 ;
        RECT -3.565 198.555 -3.235 198.885 ;
        RECT -3.565 197.065 -3.235 197.395 ;
        RECT -3.565 195.395 -3.235 195.725 ;
        RECT -3.565 193.905 -3.235 194.235 ;
        RECT -3.565 192.235 -3.235 192.565 ;
        RECT -3.565 190.745 -3.235 191.075 ;
        RECT -3.565 189.335 -3.235 189.665 ;
        RECT -3.565 187.495 -3.235 187.825 ;
        RECT -3.565 186.005 -3.235 186.335 ;
        RECT -3.565 184.335 -3.235 184.665 ;
        RECT -3.565 182.845 -3.235 183.175 ;
        RECT -3.565 181.175 -3.235 181.505 ;
        RECT -3.565 179.685 -3.235 180.015 ;
        RECT -3.565 178.015 -3.235 178.345 ;
        RECT -3.565 176.525 -3.235 176.855 ;
        RECT -3.565 175.115 -3.235 175.445 ;
        RECT -3.565 173.275 -3.235 173.605 ;
        RECT -3.565 171.785 -3.235 172.115 ;
        RECT -3.565 170.115 -3.235 170.445 ;
        RECT -3.565 168.625 -3.235 168.955 ;
        RECT -3.565 166.955 -3.235 167.285 ;
        RECT -3.565 165.465 -3.235 165.795 ;
        RECT -3.565 163.795 -3.235 164.125 ;
        RECT -3.565 162.305 -3.235 162.635 ;
        RECT -3.565 160.895 -3.235 161.225 ;
        RECT -3.565 159.055 -3.235 159.385 ;
        RECT -3.565 157.565 -3.235 157.895 ;
        RECT -3.565 155.895 -3.235 156.225 ;
        RECT -3.565 154.405 -3.235 154.735 ;
        RECT -3.565 152.735 -3.235 153.065 ;
        RECT -3.565 151.245 -3.235 151.575 ;
        RECT -3.565 149.575 -3.235 149.905 ;
        RECT -3.565 148.085 -3.235 148.415 ;
        RECT -3.565 146.675 -3.235 147.005 ;
        RECT -3.565 144.835 -3.235 145.165 ;
        RECT -3.565 143.345 -3.235 143.675 ;
        RECT -3.565 141.675 -3.235 142.005 ;
        RECT -3.565 140.185 -3.235 140.515 ;
        RECT -3.565 138.515 -3.235 138.845 ;
        RECT -3.565 137.025 -3.235 137.355 ;
        RECT -3.565 135.355 -3.235 135.685 ;
        RECT -3.565 133.865 -3.235 134.195 ;
        RECT -3.565 132.455 -3.235 132.785 ;
        RECT -3.565 130.615 -3.235 130.945 ;
        RECT -3.565 129.125 -3.235 129.455 ;
        RECT -3.565 127.455 -3.235 127.785 ;
        RECT -3.565 125.965 -3.235 126.295 ;
        RECT -3.565 124.295 -3.235 124.625 ;
        RECT -3.565 122.805 -3.235 123.135 ;
        RECT -3.565 121.135 -3.235 121.465 ;
        RECT -3.565 119.645 -3.235 119.975 ;
        RECT -3.565 118.235 -3.235 118.565 ;
        RECT -3.565 116.395 -3.235 116.725 ;
        RECT -3.565 114.905 -3.235 115.235 ;
        RECT -3.565 113.235 -3.235 113.565 ;
        RECT -3.565 111.745 -3.235 112.075 ;
        RECT -3.565 110.075 -3.235 110.405 ;
        RECT -3.565 108.585 -3.235 108.915 ;
        RECT -3.565 106.915 -3.235 107.245 ;
        RECT -3.565 105.425 -3.235 105.755 ;
        RECT -3.565 104.015 -3.235 104.345 ;
        RECT -3.565 102.175 -3.235 102.505 ;
        RECT -3.565 100.685 -3.235 101.015 ;
        RECT -3.565 99.015 -3.235 99.345 ;
        RECT -3.565 97.525 -3.235 97.855 ;
        RECT -3.565 95.855 -3.235 96.185 ;
        RECT -3.565 94.365 -3.235 94.695 ;
        RECT -3.565 92.695 -3.235 93.025 ;
        RECT -3.565 91.205 -3.235 91.535 ;
        RECT -3.565 89.795 -3.235 90.125 ;
        RECT -3.565 87.955 -3.235 88.285 ;
        RECT -3.565 86.465 -3.235 86.795 ;
        RECT -3.565 84.795 -3.235 85.125 ;
        RECT -3.565 83.305 -3.235 83.635 ;
        RECT -3.565 81.635 -3.235 81.965 ;
        RECT -3.565 80.145 -3.235 80.475 ;
        RECT -3.565 78.475 -3.235 78.805 ;
        RECT -3.565 76.985 -3.235 77.315 ;
        RECT -3.565 75.575 -3.235 75.905 ;
        RECT -3.565 73.735 -3.235 74.065 ;
        RECT -3.565 72.245 -3.235 72.575 ;
        RECT -3.565 70.575 -3.235 70.905 ;
        RECT -3.565 69.085 -3.235 69.415 ;
        RECT -3.565 67.415 -3.235 67.745 ;
        RECT -3.565 65.925 -3.235 66.255 ;
        RECT -3.565 64.255 -3.235 64.585 ;
        RECT -3.565 62.765 -3.235 63.095 ;
        RECT -3.565 61.355 -3.235 61.685 ;
        RECT -3.565 59.515 -3.235 59.845 ;
        RECT -3.565 58.025 -3.235 58.355 ;
        RECT -3.565 56.355 -3.235 56.685 ;
        RECT -3.565 54.865 -3.235 55.195 ;
        RECT -3.565 53.195 -3.235 53.525 ;
        RECT -3.565 51.705 -3.235 52.035 ;
        RECT -3.565 50.035 -3.235 50.365 ;
        RECT -3.565 48.545 -3.235 48.875 ;
        RECT -3.565 47.135 -3.235 47.465 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 244.04 -12.755 245.17 ;
        RECT -13.085 242.595 -12.755 242.925 ;
        RECT -13.085 241.235 -12.755 241.565 ;
        RECT -13.085 239.875 -12.755 240.205 ;
        RECT -13.085 238.515 -12.755 238.845 ;
        RECT -13.085 237.155 -12.755 237.485 ;
        RECT -13.085 235.795 -12.755 236.125 ;
        RECT -13.085 234.435 -12.755 234.765 ;
        RECT -13.085 233.075 -12.755 233.405 ;
        RECT -13.085 231.715 -12.755 232.045 ;
        RECT -13.085 230.355 -12.755 230.685 ;
        RECT -13.085 228.995 -12.755 229.325 ;
        RECT -13.085 227.635 -12.755 227.965 ;
        RECT -13.085 226.275 -12.755 226.605 ;
        RECT -13.085 224.915 -12.755 225.245 ;
        RECT -13.085 223.555 -12.755 223.885 ;
        RECT -13.085 222.195 -12.755 222.525 ;
        RECT -13.085 220.835 -12.755 221.165 ;
        RECT -13.085 219.475 -12.755 219.805 ;
        RECT -13.085 218.115 -12.755 218.445 ;
        RECT -13.085 216.755 -12.755 217.085 ;
        RECT -13.085 215.395 -12.755 215.725 ;
        RECT -13.085 214.035 -12.755 214.365 ;
        RECT -13.085 212.675 -12.755 213.005 ;
        RECT -13.085 211.315 -12.755 211.645 ;
        RECT -13.085 209.955 -12.755 210.285 ;
        RECT -13.085 208.595 -12.755 208.925 ;
        RECT -13.085 207.235 -12.755 207.565 ;
        RECT -13.085 205.875 -12.755 206.205 ;
        RECT -13.085 204.515 -12.755 204.845 ;
        RECT -13.085 203.155 -12.755 203.485 ;
        RECT -13.085 201.795 -12.755 202.125 ;
        RECT -13.085 200.435 -12.755 200.765 ;
        RECT -13.085 199.075 -12.755 199.405 ;
        RECT -13.085 197.715 -12.755 198.045 ;
        RECT -13.085 196.355 -12.755 196.685 ;
        RECT -13.085 194.995 -12.755 195.325 ;
        RECT -13.085 193.635 -12.755 193.965 ;
        RECT -13.085 192.275 -12.755 192.605 ;
        RECT -13.085 190.915 -12.755 191.245 ;
        RECT -13.085 189.555 -12.755 189.885 ;
        RECT -13.085 188.195 -12.755 188.525 ;
        RECT -13.085 186.835 -12.755 187.165 ;
        RECT -13.085 185.475 -12.755 185.805 ;
        RECT -13.085 184.115 -12.755 184.445 ;
        RECT -13.085 182.755 -12.755 183.085 ;
        RECT -13.085 181.395 -12.755 181.725 ;
        RECT -13.085 180.035 -12.755 180.365 ;
        RECT -13.085 178.675 -12.755 179.005 ;
        RECT -13.085 177.315 -12.755 177.645 ;
        RECT -13.085 175.955 -12.755 176.285 ;
        RECT -13.085 174.595 -12.755 174.925 ;
        RECT -13.085 173.235 -12.755 173.565 ;
        RECT -13.085 171.875 -12.755 172.205 ;
        RECT -13.085 170.515 -12.755 170.845 ;
        RECT -13.085 169.155 -12.755 169.485 ;
        RECT -13.085 167.795 -12.755 168.125 ;
        RECT -13.085 166.435 -12.755 166.765 ;
        RECT -13.085 165.075 -12.755 165.405 ;
        RECT -13.085 163.715 -12.755 164.045 ;
        RECT -13.085 162.355 -12.755 162.685 ;
        RECT -13.085 160.995 -12.755 161.325 ;
        RECT -13.085 159.635 -12.755 159.965 ;
        RECT -13.085 158.275 -12.755 158.605 ;
        RECT -13.085 156.915 -12.755 157.245 ;
        RECT -13.085 155.555 -12.755 155.885 ;
        RECT -13.085 154.195 -12.755 154.525 ;
        RECT -13.085 152.835 -12.755 153.165 ;
        RECT -13.085 151.475 -12.755 151.805 ;
        RECT -13.085 150.115 -12.755 150.445 ;
        RECT -13.085 148.755 -12.755 149.085 ;
        RECT -13.085 147.395 -12.755 147.725 ;
        RECT -13.085 146.035 -12.755 146.365 ;
        RECT -13.085 144.675 -12.755 145.005 ;
        RECT -13.085 143.315 -12.755 143.645 ;
        RECT -13.085 141.955 -12.755 142.285 ;
        RECT -13.085 140.595 -12.755 140.925 ;
        RECT -13.085 139.235 -12.755 139.565 ;
        RECT -13.085 137.875 -12.755 138.205 ;
        RECT -13.085 136.515 -12.755 136.845 ;
        RECT -13.085 135.155 -12.755 135.485 ;
        RECT -13.085 133.795 -12.755 134.125 ;
        RECT -13.085 132.435 -12.755 132.765 ;
        RECT -13.085 131.075 -12.755 131.405 ;
        RECT -13.085 129.715 -12.755 130.045 ;
        RECT -13.085 128.355 -12.755 128.685 ;
        RECT -13.085 126.995 -12.755 127.325 ;
        RECT -13.085 125.635 -12.755 125.965 ;
        RECT -13.085 124.275 -12.755 124.605 ;
        RECT -13.085 122.915 -12.755 123.245 ;
        RECT -13.085 121.555 -12.755 121.885 ;
        RECT -13.085 120.195 -12.755 120.525 ;
        RECT -13.085 118.835 -12.755 119.165 ;
        RECT -13.085 117.475 -12.755 117.805 ;
        RECT -13.085 116.115 -12.755 116.445 ;
        RECT -13.085 114.755 -12.755 115.085 ;
        RECT -13.085 113.395 -12.755 113.725 ;
        RECT -13.085 112.035 -12.755 112.365 ;
        RECT -13.085 110.675 -12.755 111.005 ;
        RECT -13.085 109.315 -12.755 109.645 ;
        RECT -13.085 107.955 -12.755 108.285 ;
        RECT -13.085 106.595 -12.755 106.925 ;
        RECT -13.085 105.235 -12.755 105.565 ;
        RECT -13.085 103.875 -12.755 104.205 ;
        RECT -13.085 102.515 -12.755 102.845 ;
        RECT -13.085 101.155 -12.755 101.485 ;
        RECT -13.085 99.795 -12.755 100.125 ;
        RECT -13.085 98.435 -12.755 98.765 ;
        RECT -13.085 97.075 -12.755 97.405 ;
        RECT -13.085 95.715 -12.755 96.045 ;
        RECT -13.085 94.355 -12.755 94.685 ;
        RECT -13.085 92.995 -12.755 93.325 ;
        RECT -13.085 91.635 -12.755 91.965 ;
        RECT -13.085 90.275 -12.755 90.605 ;
        RECT -13.085 88.915 -12.755 89.245 ;
        RECT -13.085 87.555 -12.755 87.885 ;
        RECT -13.085 86.195 -12.755 86.525 ;
        RECT -13.085 84.835 -12.755 85.165 ;
        RECT -13.085 83.475 -12.755 83.805 ;
        RECT -13.085 82.115 -12.755 82.445 ;
        RECT -13.085 80.755 -12.755 81.085 ;
        RECT -13.085 79.395 -12.755 79.725 ;
        RECT -13.085 78.035 -12.755 78.365 ;
        RECT -13.085 76.675 -12.755 77.005 ;
        RECT -13.085 75.315 -12.755 75.645 ;
        RECT -13.085 73.955 -12.755 74.285 ;
        RECT -13.085 72.595 -12.755 72.925 ;
        RECT -13.085 71.235 -12.755 71.565 ;
        RECT -13.085 69.875 -12.755 70.205 ;
        RECT -13.085 68.515 -12.755 68.845 ;
        RECT -13.085 67.155 -12.755 67.485 ;
        RECT -13.085 65.795 -12.755 66.125 ;
        RECT -13.085 64.435 -12.755 64.765 ;
        RECT -13.085 63.075 -12.755 63.405 ;
        RECT -13.085 61.715 -12.755 62.045 ;
        RECT -13.085 60.355 -12.755 60.685 ;
        RECT -13.085 58.995 -12.755 59.325 ;
        RECT -13.085 57.635 -12.755 57.965 ;
        RECT -13.085 56.275 -12.755 56.605 ;
        RECT -13.085 54.915 -12.755 55.245 ;
        RECT -13.085 53.555 -12.755 53.885 ;
        RECT -13.085 52.195 -12.755 52.525 ;
        RECT -13.085 50.835 -12.755 51.165 ;
        RECT -13.085 49.475 -12.755 49.805 ;
        RECT -13.085 48.115 -12.755 48.445 ;
        RECT -13.085 46.755 -12.755 47.085 ;
        RECT -13.085 45.395 -12.755 45.725 ;
        RECT -13.085 44.035 -12.755 44.365 ;
        RECT -13.085 42.675 -12.755 43.005 ;
        RECT -13.085 41.315 -12.755 41.645 ;
        RECT -13.085 39.955 -12.755 40.285 ;
        RECT -13.085 38.595 -12.755 38.925 ;
        RECT -13.085 37.235 -12.755 37.565 ;
        RECT -13.085 35.875 -12.755 36.205 ;
        RECT -13.085 34.515 -12.755 34.845 ;
        RECT -13.085 33.155 -12.755 33.485 ;
        RECT -13.085 31.795 -12.755 32.125 ;
        RECT -13.085 30.435 -12.755 30.765 ;
        RECT -13.085 29.075 -12.755 29.405 ;
        RECT -13.085 27.715 -12.755 28.045 ;
        RECT -13.085 26.355 -12.755 26.685 ;
        RECT -13.085 24.995 -12.755 25.325 ;
        RECT -13.085 23.635 -12.755 23.965 ;
        RECT -13.085 22.275 -12.755 22.605 ;
        RECT -13.085 20.915 -12.755 21.245 ;
        RECT -13.085 19.555 -12.755 19.885 ;
        RECT -13.085 18.195 -12.755 18.525 ;
        RECT -13.085 16.835 -12.755 17.165 ;
        RECT -13.085 15.475 -12.755 15.805 ;
        RECT -13.085 14.115 -12.755 14.445 ;
        RECT -13.085 12.755 -12.755 13.085 ;
        RECT -13.085 11.395 -12.755 11.725 ;
        RECT -13.085 10.035 -12.755 10.365 ;
        RECT -13.085 8.675 -12.755 9.005 ;
        RECT -13.085 7.315 -12.755 7.645 ;
        RECT -13.085 5.955 -12.755 6.285 ;
        RECT -13.085 4.595 -12.755 4.925 ;
        RECT -13.085 3.235 -12.755 3.565 ;
        RECT -13.085 1.875 -12.755 2.205 ;
        RECT -13.085 0.515 -12.755 0.845 ;
        RECT -13.085 -2.205 -12.755 -1.875 ;
        RECT -13.085 -3.565 -12.755 -3.235 ;
        RECT -13.085 -4.925 -12.755 -4.595 ;
        RECT -13.085 -6.285 -12.755 -5.955 ;
        RECT -13.085 -7.645 -12.755 -7.315 ;
        RECT -13.085 -10.365 -12.755 -10.035 ;
        RECT -13.085 -11.725 -12.755 -11.395 ;
        RECT -13.085 -13.7 -12.755 -13.37 ;
        RECT -13.085 -14.445 -12.755 -14.115 ;
        RECT -13.085 -15.805 -12.755 -15.475 ;
        RECT -13.085 -18.79 -12.755 -18.46 ;
        RECT -13.085 -19.885 -12.755 -19.555 ;
        RECT -13.085 -23.965 -12.755 -23.635 ;
        RECT -13.085 -25.325 -12.755 -24.995 ;
        RECT -13.085 -26.685 -12.755 -26.355 ;
        RECT -13.085 -28.045 -12.755 -27.715 ;
        RECT -13.085 -29.405 -12.755 -29.075 ;
        RECT -13.085 -32.125 -12.755 -31.795 ;
        RECT -13.085 -33.485 -12.755 -33.155 ;
        RECT -13.085 -34.88 -12.755 -34.55 ;
        RECT -13.085 -36.205 -12.755 -35.875 ;
        RECT -13.085 -38.925 -12.755 -38.595 ;
        RECT -13.085 -39.97 -12.755 -39.64 ;
        RECT -13.085 -47.085 -12.755 -46.755 ;
        RECT -13.085 -48.445 -12.755 -48.115 ;
        RECT -13.085 -49.805 -12.755 -49.475 ;
        RECT -13.085 -51.165 -12.755 -50.835 ;
        RECT -13.085 -52.525 -12.755 -52.195 ;
        RECT -13.085 -53.885 -12.755 -53.555 ;
        RECT -13.085 -55.245 -12.755 -54.915 ;
        RECT -13.085 -56.605 -12.755 -56.275 ;
        RECT -13.085 -57.965 -12.755 -57.635 ;
        RECT -13.085 -59.325 -12.755 -58.995 ;
        RECT -13.085 -60.685 -12.755 -60.355 ;
        RECT -13.085 -62.045 -12.755 -61.715 ;
        RECT -13.085 -68.845 -12.755 -68.515 ;
        RECT -13.085 -72.925 -12.755 -72.595 ;
        RECT -13.085 -74.285 -12.755 -73.955 ;
        RECT -13.085 -75.645 -12.755 -75.315 ;
        RECT -13.085 -77.005 -12.755 -76.675 ;
        RECT -13.085 -78.365 -12.755 -78.035 ;
        RECT -13.085 -80.31 -12.755 -79.98 ;
        RECT -13.085 -81.085 -12.755 -80.755 ;
        RECT -13.085 -82.445 -12.755 -82.115 ;
        RECT -13.085 -83.805 -12.755 -83.475 ;
        RECT -13.085 -85.165 -12.755 -84.835 ;
        RECT -13.085 -86.525 -12.755 -86.195 ;
        RECT -13.085 -87.885 -12.755 -87.555 ;
        RECT -13.085 -90.605 -12.755 -90.275 ;
        RECT -13.085 -91.965 -12.755 -91.635 ;
        RECT -13.085 -93.325 -12.755 -92.995 ;
        RECT -13.085 -94.685 -12.755 -94.355 ;
        RECT -13.085 -96.045 -12.755 -95.715 ;
        RECT -13.085 -97.405 -12.755 -97.075 ;
        RECT -13.085 -98.85 -12.755 -98.52 ;
        RECT -13.085 -100.125 -12.755 -99.795 ;
        RECT -13.085 -101.485 -12.755 -101.155 ;
        RECT -13.085 -102.845 -12.755 -102.515 ;
        RECT -13.085 -105.565 -12.755 -105.235 ;
        RECT -13.085 -106.925 -12.755 -106.595 ;
        RECT -13.085 -108.285 -12.755 -107.955 ;
        RECT -13.085 -109.645 -12.755 -109.315 ;
        RECT -13.085 -111.005 -12.755 -110.675 ;
        RECT -13.085 -112.365 -12.755 -112.035 ;
        RECT -13.085 -113.725 -12.755 -113.395 ;
        RECT -13.085 -116.445 -12.755 -116.115 ;
        RECT -13.08 -117.12 -12.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 -217.085 -12.755 -216.755 ;
        RECT -13.085 -218.445 -12.755 -218.115 ;
        RECT -13.085 -219.805 -12.755 -219.475 ;
        RECT -13.085 -221.165 -12.755 -220.835 ;
        RECT -13.085 -222.525 -12.755 -222.195 ;
        RECT -13.085 -223.885 -12.755 -223.555 ;
        RECT -13.085 -227.965 -12.755 -227.635 ;
        RECT -13.085 -230.685 -12.755 -230.355 ;
        RECT -13.085 -232.045 -12.755 -231.715 ;
        RECT -13.085 -233.225 -12.755 -232.895 ;
        RECT -13.085 -234.765 -12.755 -234.435 ;
        RECT -13.085 -236.125 -12.755 -235.795 ;
        RECT -13.085 -237.485 -12.755 -237.155 ;
        RECT -13.085 -238.845 -12.755 -238.515 ;
        RECT -13.085 -241.09 -12.755 -239.96 ;
        RECT -13.08 -241.205 -12.76 -216.755 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.725 244.04 -11.395 245.17 ;
        RECT -11.725 242.595 -11.395 242.925 ;
        RECT -11.725 241.235 -11.395 241.565 ;
        RECT -11.725 239.875 -11.395 240.205 ;
        RECT -11.725 238.515 -11.395 238.845 ;
        RECT -11.725 237.155 -11.395 237.485 ;
        RECT -11.725 235.795 -11.395 236.125 ;
        RECT -11.725 234.435 -11.395 234.765 ;
        RECT -11.725 233.075 -11.395 233.405 ;
        RECT -11.725 231.715 -11.395 232.045 ;
        RECT -11.725 230.355 -11.395 230.685 ;
        RECT -11.725 228.995 -11.395 229.325 ;
        RECT -11.725 227.635 -11.395 227.965 ;
        RECT -11.725 226.275 -11.395 226.605 ;
        RECT -11.725 224.915 -11.395 225.245 ;
        RECT -11.725 223.555 -11.395 223.885 ;
        RECT -11.725 222.195 -11.395 222.525 ;
        RECT -11.725 220.835 -11.395 221.165 ;
        RECT -11.725 219.475 -11.395 219.805 ;
        RECT -11.725 218.115 -11.395 218.445 ;
        RECT -11.725 216.755 -11.395 217.085 ;
        RECT -11.725 215.395 -11.395 215.725 ;
        RECT -11.725 214.035 -11.395 214.365 ;
        RECT -11.725 212.675 -11.395 213.005 ;
        RECT -11.725 211.315 -11.395 211.645 ;
        RECT -11.725 209.955 -11.395 210.285 ;
        RECT -11.725 208.595 -11.395 208.925 ;
        RECT -11.725 207.235 -11.395 207.565 ;
        RECT -11.725 205.875 -11.395 206.205 ;
        RECT -11.725 204.515 -11.395 204.845 ;
        RECT -11.725 203.155 -11.395 203.485 ;
        RECT -11.725 201.795 -11.395 202.125 ;
        RECT -11.725 200.435 -11.395 200.765 ;
        RECT -11.725 199.075 -11.395 199.405 ;
        RECT -11.725 197.715 -11.395 198.045 ;
        RECT -11.725 196.355 -11.395 196.685 ;
        RECT -11.725 194.995 -11.395 195.325 ;
        RECT -11.725 193.635 -11.395 193.965 ;
        RECT -11.725 192.275 -11.395 192.605 ;
        RECT -11.725 190.915 -11.395 191.245 ;
        RECT -11.725 189.555 -11.395 189.885 ;
        RECT -11.725 188.195 -11.395 188.525 ;
        RECT -11.725 186.835 -11.395 187.165 ;
        RECT -11.725 185.475 -11.395 185.805 ;
        RECT -11.725 184.115 -11.395 184.445 ;
        RECT -11.725 182.755 -11.395 183.085 ;
        RECT -11.725 181.395 -11.395 181.725 ;
        RECT -11.725 180.035 -11.395 180.365 ;
        RECT -11.725 178.675 -11.395 179.005 ;
        RECT -11.725 177.315 -11.395 177.645 ;
        RECT -11.725 175.955 -11.395 176.285 ;
        RECT -11.725 174.595 -11.395 174.925 ;
        RECT -11.725 173.235 -11.395 173.565 ;
        RECT -11.725 171.875 -11.395 172.205 ;
        RECT -11.725 170.515 -11.395 170.845 ;
        RECT -11.725 169.155 -11.395 169.485 ;
        RECT -11.725 167.795 -11.395 168.125 ;
        RECT -11.725 166.435 -11.395 166.765 ;
        RECT -11.725 165.075 -11.395 165.405 ;
        RECT -11.725 163.715 -11.395 164.045 ;
        RECT -11.725 162.355 -11.395 162.685 ;
        RECT -11.725 160.995 -11.395 161.325 ;
        RECT -11.725 159.635 -11.395 159.965 ;
        RECT -11.725 158.275 -11.395 158.605 ;
        RECT -11.725 156.915 -11.395 157.245 ;
        RECT -11.725 155.555 -11.395 155.885 ;
        RECT -11.725 154.195 -11.395 154.525 ;
        RECT -11.725 152.835 -11.395 153.165 ;
        RECT -11.725 151.475 -11.395 151.805 ;
        RECT -11.725 150.115 -11.395 150.445 ;
        RECT -11.725 148.755 -11.395 149.085 ;
        RECT -11.725 147.395 -11.395 147.725 ;
        RECT -11.725 146.035 -11.395 146.365 ;
        RECT -11.725 144.675 -11.395 145.005 ;
        RECT -11.725 143.315 -11.395 143.645 ;
        RECT -11.725 141.955 -11.395 142.285 ;
        RECT -11.725 140.595 -11.395 140.925 ;
        RECT -11.725 139.235 -11.395 139.565 ;
        RECT -11.725 137.875 -11.395 138.205 ;
        RECT -11.725 136.515 -11.395 136.845 ;
        RECT -11.725 135.155 -11.395 135.485 ;
        RECT -11.725 133.795 -11.395 134.125 ;
        RECT -11.725 132.435 -11.395 132.765 ;
        RECT -11.725 131.075 -11.395 131.405 ;
        RECT -11.725 129.715 -11.395 130.045 ;
        RECT -11.725 128.355 -11.395 128.685 ;
        RECT -11.725 126.995 -11.395 127.325 ;
        RECT -11.725 125.635 -11.395 125.965 ;
        RECT -11.725 124.275 -11.395 124.605 ;
        RECT -11.725 122.915 -11.395 123.245 ;
        RECT -11.725 121.555 -11.395 121.885 ;
        RECT -11.725 120.195 -11.395 120.525 ;
        RECT -11.725 118.835 -11.395 119.165 ;
        RECT -11.725 117.475 -11.395 117.805 ;
        RECT -11.725 116.115 -11.395 116.445 ;
        RECT -11.725 114.755 -11.395 115.085 ;
        RECT -11.725 113.395 -11.395 113.725 ;
        RECT -11.725 112.035 -11.395 112.365 ;
        RECT -11.725 110.675 -11.395 111.005 ;
        RECT -11.725 109.315 -11.395 109.645 ;
        RECT -11.725 107.955 -11.395 108.285 ;
        RECT -11.725 106.595 -11.395 106.925 ;
        RECT -11.725 105.235 -11.395 105.565 ;
        RECT -11.725 103.875 -11.395 104.205 ;
        RECT -11.725 102.515 -11.395 102.845 ;
        RECT -11.725 101.155 -11.395 101.485 ;
        RECT -11.725 99.795 -11.395 100.125 ;
        RECT -11.725 98.435 -11.395 98.765 ;
        RECT -11.725 97.075 -11.395 97.405 ;
        RECT -11.725 95.715 -11.395 96.045 ;
        RECT -11.725 94.355 -11.395 94.685 ;
        RECT -11.725 92.995 -11.395 93.325 ;
        RECT -11.725 91.635 -11.395 91.965 ;
        RECT -11.725 90.275 -11.395 90.605 ;
        RECT -11.725 88.915 -11.395 89.245 ;
        RECT -11.725 87.555 -11.395 87.885 ;
        RECT -11.725 86.195 -11.395 86.525 ;
        RECT -11.725 84.835 -11.395 85.165 ;
        RECT -11.725 83.475 -11.395 83.805 ;
        RECT -11.725 82.115 -11.395 82.445 ;
        RECT -11.725 80.755 -11.395 81.085 ;
        RECT -11.725 79.395 -11.395 79.725 ;
        RECT -11.725 78.035 -11.395 78.365 ;
        RECT -11.725 76.675 -11.395 77.005 ;
        RECT -11.725 75.315 -11.395 75.645 ;
        RECT -11.725 73.955 -11.395 74.285 ;
        RECT -11.725 72.595 -11.395 72.925 ;
        RECT -11.725 71.235 -11.395 71.565 ;
        RECT -11.725 69.875 -11.395 70.205 ;
        RECT -11.725 68.515 -11.395 68.845 ;
        RECT -11.725 67.155 -11.395 67.485 ;
        RECT -11.725 65.795 -11.395 66.125 ;
        RECT -11.725 64.435 -11.395 64.765 ;
        RECT -11.725 63.075 -11.395 63.405 ;
        RECT -11.725 61.715 -11.395 62.045 ;
        RECT -11.725 60.355 -11.395 60.685 ;
        RECT -11.725 58.995 -11.395 59.325 ;
        RECT -11.725 57.635 -11.395 57.965 ;
        RECT -11.725 56.275 -11.395 56.605 ;
        RECT -11.725 54.915 -11.395 55.245 ;
        RECT -11.725 53.555 -11.395 53.885 ;
        RECT -11.725 52.195 -11.395 52.525 ;
        RECT -11.725 50.835 -11.395 51.165 ;
        RECT -11.725 49.475 -11.395 49.805 ;
        RECT -11.725 48.115 -11.395 48.445 ;
        RECT -11.725 46.755 -11.395 47.085 ;
        RECT -11.725 45.395 -11.395 45.725 ;
        RECT -11.725 44.035 -11.395 44.365 ;
        RECT -11.725 42.675 -11.395 43.005 ;
        RECT -11.725 41.315 -11.395 41.645 ;
        RECT -11.725 39.955 -11.395 40.285 ;
        RECT -11.725 38.595 -11.395 38.925 ;
        RECT -11.725 37.235 -11.395 37.565 ;
        RECT -11.725 35.875 -11.395 36.205 ;
        RECT -11.725 34.515 -11.395 34.845 ;
        RECT -11.725 33.155 -11.395 33.485 ;
        RECT -11.725 31.795 -11.395 32.125 ;
        RECT -11.725 30.435 -11.395 30.765 ;
        RECT -11.725 29.075 -11.395 29.405 ;
        RECT -11.725 27.715 -11.395 28.045 ;
        RECT -11.725 26.355 -11.395 26.685 ;
        RECT -11.725 24.995 -11.395 25.325 ;
        RECT -11.725 23.635 -11.395 23.965 ;
        RECT -11.725 22.275 -11.395 22.605 ;
        RECT -11.725 20.915 -11.395 21.245 ;
        RECT -11.725 19.555 -11.395 19.885 ;
        RECT -11.725 18.195 -11.395 18.525 ;
        RECT -11.725 16.835 -11.395 17.165 ;
        RECT -11.725 15.475 -11.395 15.805 ;
        RECT -11.725 14.115 -11.395 14.445 ;
        RECT -11.725 12.755 -11.395 13.085 ;
        RECT -11.725 11.395 -11.395 11.725 ;
        RECT -11.725 10.035 -11.395 10.365 ;
        RECT -11.725 8.675 -11.395 9.005 ;
        RECT -11.725 7.315 -11.395 7.645 ;
        RECT -11.725 5.955 -11.395 6.285 ;
        RECT -11.725 4.595 -11.395 4.925 ;
        RECT -11.725 3.235 -11.395 3.565 ;
        RECT -11.725 1.875 -11.395 2.205 ;
        RECT -11.725 0.515 -11.395 0.845 ;
        RECT -11.725 -0.845 -11.395 -0.515 ;
        RECT -11.725 -2.205 -11.395 -1.875 ;
        RECT -11.725 -3.565 -11.395 -3.235 ;
        RECT -11.725 -4.925 -11.395 -4.595 ;
        RECT -11.725 -6.285 -11.395 -5.955 ;
        RECT -11.725 -7.645 -11.395 -7.315 ;
        RECT -11.725 -10.365 -11.395 -10.035 ;
        RECT -11.725 -11.725 -11.395 -11.395 ;
        RECT -11.725 -13.7 -11.395 -13.37 ;
        RECT -11.725 -14.445 -11.395 -14.115 ;
        RECT -11.725 -15.805 -11.395 -15.475 ;
        RECT -11.725 -18.79 -11.395 -18.46 ;
        RECT -11.725 -19.885 -11.395 -19.555 ;
        RECT -11.725 -23.965 -11.395 -23.635 ;
        RECT -11.725 -25.325 -11.395 -24.995 ;
        RECT -11.725 -26.685 -11.395 -26.355 ;
        RECT -11.725 -28.045 -11.395 -27.715 ;
        RECT -11.725 -29.405 -11.395 -29.075 ;
        RECT -11.725 -32.125 -11.395 -31.795 ;
        RECT -11.725 -33.485 -11.395 -33.155 ;
        RECT -11.725 -34.88 -11.395 -34.55 ;
        RECT -11.725 -36.205 -11.395 -35.875 ;
        RECT -11.725 -38.925 -11.395 -38.595 ;
        RECT -11.725 -39.97 -11.395 -39.64 ;
        RECT -11.725 -47.085 -11.395 -46.755 ;
        RECT -11.725 -48.445 -11.395 -48.115 ;
        RECT -11.725 -49.805 -11.395 -49.475 ;
        RECT -11.725 -51.165 -11.395 -50.835 ;
        RECT -11.725 -52.525 -11.395 -52.195 ;
        RECT -11.725 -53.885 -11.395 -53.555 ;
        RECT -11.725 -55.245 -11.395 -54.915 ;
        RECT -11.725 -56.605 -11.395 -56.275 ;
        RECT -11.725 -57.965 -11.395 -57.635 ;
        RECT -11.725 -59.325 -11.395 -58.995 ;
        RECT -11.725 -60.685 -11.395 -60.355 ;
        RECT -11.725 -62.045 -11.395 -61.715 ;
        RECT -11.725 -68.845 -11.395 -68.515 ;
        RECT -11.725 -72.925 -11.395 -72.595 ;
        RECT -11.725 -74.285 -11.395 -73.955 ;
        RECT -11.725 -75.645 -11.395 -75.315 ;
        RECT -11.725 -77.005 -11.395 -76.675 ;
        RECT -11.725 -78.365 -11.395 -78.035 ;
        RECT -11.725 -80.31 -11.395 -79.98 ;
        RECT -11.725 -81.085 -11.395 -80.755 ;
        RECT -11.725 -82.445 -11.395 -82.115 ;
        RECT -11.725 -83.805 -11.395 -83.475 ;
        RECT -11.725 -85.165 -11.395 -84.835 ;
        RECT -11.725 -86.525 -11.395 -86.195 ;
        RECT -11.725 -87.885 -11.395 -87.555 ;
        RECT -11.725 -90.605 -11.395 -90.275 ;
        RECT -11.725 -91.965 -11.395 -91.635 ;
        RECT -11.725 -93.325 -11.395 -92.995 ;
        RECT -11.725 -94.685 -11.395 -94.355 ;
        RECT -11.725 -96.045 -11.395 -95.715 ;
        RECT -11.725 -97.405 -11.395 -97.075 ;
        RECT -11.725 -98.85 -11.395 -98.52 ;
        RECT -11.725 -100.125 -11.395 -99.795 ;
        RECT -11.725 -101.485 -11.395 -101.155 ;
        RECT -11.725 -102.845 -11.395 -102.515 ;
        RECT -11.725 -105.565 -11.395 -105.235 ;
        RECT -11.725 -106.925 -11.395 -106.595 ;
        RECT -11.725 -108.285 -11.395 -107.955 ;
        RECT -11.725 -109.645 -11.395 -109.315 ;
        RECT -11.725 -111.005 -11.395 -110.675 ;
        RECT -11.725 -112.365 -11.395 -112.035 ;
        RECT -11.725 -113.725 -11.395 -113.395 ;
        RECT -11.725 -116.445 -11.395 -116.115 ;
        RECT -11.725 -119.165 -11.395 -118.835 ;
        RECT -11.725 -120.525 -11.395 -120.195 ;
        RECT -11.725 -121.885 -11.395 -121.555 ;
        RECT -11.725 -123.245 -11.395 -122.915 ;
        RECT -11.725 -124.49 -11.395 -124.16 ;
        RECT -11.725 -125.965 -11.395 -125.635 ;
        RECT -11.725 -127.325 -11.395 -126.995 ;
        RECT -11.725 -128.685 -11.395 -128.355 ;
        RECT -11.725 -130.045 -11.395 -129.715 ;
        RECT -11.725 -131.405 -11.395 -131.075 ;
        RECT -11.725 -132.765 -11.395 -132.435 ;
        RECT -11.725 -140.925 -11.395 -140.595 ;
        RECT -11.725 -142.285 -11.395 -141.955 ;
        RECT -11.725 -143.03 -11.395 -142.7 ;
        RECT -11.725 -145.005 -11.395 -144.675 ;
        RECT -11.725 -146.365 -11.395 -146.035 ;
        RECT -11.725 -147.725 -11.395 -147.395 ;
        RECT -11.725 -153.165 -11.395 -152.835 ;
        RECT -11.725 -154.525 -11.395 -154.195 ;
        RECT -11.725 -155.885 -11.395 -155.555 ;
        RECT -11.725 -157.245 -11.395 -156.915 ;
        RECT -11.725 -158.605 -11.395 -158.275 ;
        RECT -11.725 -159.965 -11.395 -159.635 ;
        RECT -11.725 -161.325 -11.395 -160.995 ;
        RECT -11.725 -164.045 -11.395 -163.715 ;
        RECT -11.725 -168.125 -11.395 -167.795 ;
        RECT -11.725 -172.205 -11.395 -171.875 ;
        RECT -11.725 -173.565 -11.395 -173.235 ;
        RECT -11.725 -174.925 -11.395 -174.595 ;
        RECT -11.725 -176.285 -11.395 -175.955 ;
        RECT -11.725 -177.645 -11.395 -177.315 ;
        RECT -11.725 -179.005 -11.395 -178.675 ;
        RECT -11.725 -180.365 -11.395 -180.035 ;
        RECT -11.725 -181.725 -11.395 -181.395 ;
        RECT -11.725 -183.085 -11.395 -182.755 ;
        RECT -11.725 -184.445 -11.395 -184.115 ;
        RECT -11.725 -185.805 -11.395 -185.475 ;
        RECT -11.725 -188.525 -11.395 -188.195 ;
        RECT -11.725 -189.885 -11.395 -189.555 ;
        RECT -11.725 -191.245 -11.395 -190.915 ;
        RECT -11.725 -192.605 -11.395 -192.275 ;
        RECT -11.725 -193.965 -11.395 -193.635 ;
        RECT -11.725 -195.325 -11.395 -194.995 ;
        RECT -11.725 -196.685 -11.395 -196.355 ;
        RECT -11.725 -198.045 -11.395 -197.715 ;
        RECT -11.725 -199.405 -11.395 -199.075 ;
        RECT -11.725 -203.485 -11.395 -203.155 ;
        RECT -11.725 -204.845 -11.395 -204.515 ;
        RECT -11.725 -206.205 -11.395 -205.875 ;
        RECT -11.725 -207.565 -11.395 -207.235 ;
        RECT -11.725 -208.925 -11.395 -208.595 ;
        RECT -11.725 -210.285 -11.395 -209.955 ;
        RECT -11.725 -211.645 -11.395 -211.315 ;
        RECT -11.725 -213.005 -11.395 -212.675 ;
        RECT -11.725 -214.365 -11.395 -214.035 ;
        RECT -11.725 -215.725 -11.395 -215.395 ;
        RECT -11.725 -217.085 -11.395 -216.755 ;
        RECT -11.725 -218.445 -11.395 -218.115 ;
        RECT -11.725 -219.805 -11.395 -219.475 ;
        RECT -11.725 -221.165 -11.395 -220.835 ;
        RECT -11.725 -222.525 -11.395 -222.195 ;
        RECT -11.725 -223.885 -11.395 -223.555 ;
        RECT -11.725 -227.965 -11.395 -227.635 ;
        RECT -11.725 -232.045 -11.395 -231.715 ;
        RECT -11.725 -233.225 -11.395 -232.895 ;
        RECT -11.725 -234.765 -11.395 -234.435 ;
        RECT -11.725 -236.125 -11.395 -235.795 ;
        RECT -11.725 -237.485 -11.395 -237.155 ;
        RECT -11.725 -238.845 -11.395 -238.515 ;
        RECT -11.725 -241.09 -11.395 -239.96 ;
        RECT -11.72 -241.205 -11.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 244.04 -10.035 245.17 ;
        RECT -10.365 242.595 -10.035 242.925 ;
        RECT -10.365 241.235 -10.035 241.565 ;
        RECT -10.365 239.875 -10.035 240.205 ;
        RECT -10.365 238.515 -10.035 238.845 ;
        RECT -10.365 237.155 -10.035 237.485 ;
        RECT -10.365 235.795 -10.035 236.125 ;
        RECT -10.365 234.435 -10.035 234.765 ;
        RECT -10.365 233.075 -10.035 233.405 ;
        RECT -10.365 231.715 -10.035 232.045 ;
        RECT -10.365 227.635 -10.035 227.965 ;
        RECT -10.365 224.915 -10.035 225.245 ;
        RECT -10.365 218.115 -10.035 218.445 ;
        RECT -10.365 216.755 -10.035 217.085 ;
        RECT -10.365 207.235 -10.035 207.565 ;
        RECT -10.365 204.515 -10.035 204.845 ;
        RECT -10.365 203.155 -10.035 203.485 ;
        RECT -10.365 199.075 -10.035 199.405 ;
        RECT -10.365 196.355 -10.035 196.685 ;
        RECT -10.365 189.555 -10.035 189.885 ;
        RECT -10.365 188.195 -10.035 188.525 ;
        RECT -10.365 185.475 -10.035 185.805 ;
        RECT -10.365 178.675 -10.035 179.005 ;
        RECT -10.365 175.955 -10.035 176.285 ;
        RECT -10.365 174.595 -10.035 174.925 ;
        RECT -10.365 167.795 -10.035 168.125 ;
        RECT -10.365 160.995 -10.035 161.325 ;
        RECT -10.365 159.635 -10.035 159.965 ;
        RECT -10.365 156.915 -10.035 157.245 ;
        RECT -10.365 150.115 -10.035 150.445 ;
        RECT -10.365 147.395 -10.035 147.725 ;
        RECT -10.365 146.035 -10.035 146.365 ;
        RECT -10.365 139.235 -10.035 139.565 ;
        RECT -10.365 136.515 -10.035 136.845 ;
        RECT -10.365 132.435 -10.035 132.765 ;
        RECT -10.365 131.075 -10.035 131.405 ;
        RECT -10.365 128.355 -10.035 128.685 ;
        RECT -10.365 118.835 -10.035 119.165 ;
        RECT -10.365 117.475 -10.035 117.805 ;
        RECT -10.365 110.675 -10.035 111.005 ;
        RECT -10.365 107.955 -10.035 108.285 ;
        RECT -10.365 103.875 -10.035 104.205 ;
        RECT -10.365 99.795 -10.035 100.125 ;
        RECT -10.365 97.075 -10.035 97.405 ;
        RECT -10.365 90.275 -10.035 90.605 ;
        RECT -10.365 88.915 -10.035 89.245 ;
        RECT -10.365 82.115 -10.035 82.445 ;
        RECT -10.365 79.395 -10.035 79.725 ;
        RECT -10.365 75.315 -10.035 75.645 ;
        RECT -10.365 71.235 -10.035 71.565 ;
        RECT -10.365 68.515 -10.035 68.845 ;
        RECT -10.365 61.715 -10.035 62.045 ;
        RECT -10.365 60.355 -10.035 60.685 ;
        RECT -10.365 50.835 -10.035 51.165 ;
        RECT -10.365 46.755 -10.035 47.085 ;
        RECT -10.365 42.675 -10.035 43.005 ;
        RECT -10.365 39.955 -10.035 40.285 ;
        RECT -10.365 33.155 -10.035 33.485 ;
        RECT -10.365 31.795 -10.035 32.125 ;
        RECT -10.365 29.075 -10.035 29.405 ;
        RECT -10.365 22.275 -10.035 22.605 ;
        RECT -10.365 19.555 -10.035 19.885 ;
        RECT -10.365 18.195 -10.035 18.525 ;
        RECT -10.365 11.395 -10.035 11.725 ;
        RECT -10.365 4.595 -10.035 4.925 ;
        RECT -10.365 3.235 -10.035 3.565 ;
        RECT -10.365 1.875 -10.035 2.205 ;
        RECT -10.365 0.515 -10.035 0.845 ;
        RECT -10.365 -0.845 -10.035 -0.515 ;
        RECT -10.365 -2.205 -10.035 -1.875 ;
        RECT -10.365 -3.565 -10.035 -3.235 ;
        RECT -10.365 -4.925 -10.035 -4.595 ;
        RECT -10.365 -6.285 -10.035 -5.955 ;
        RECT -10.365 -7.645 -10.035 -7.315 ;
        RECT -10.365 -10.365 -10.035 -10.035 ;
        RECT -10.365 -11.725 -10.035 -11.395 ;
        RECT -10.365 -14.445 -10.035 -14.115 ;
        RECT -10.365 -15.805 -10.035 -15.475 ;
        RECT -10.365 -19.885 -10.035 -19.555 ;
        RECT -10.365 -23.965 -10.035 -23.635 ;
        RECT -10.365 -25.325 -10.035 -24.995 ;
        RECT -10.365 -26.685 -10.035 -26.355 ;
        RECT -10.365 -28.045 -10.035 -27.715 ;
        RECT -10.365 -29.405 -10.035 -29.075 ;
        RECT -10.365 -32.125 -10.035 -31.795 ;
        RECT -10.365 -33.485 -10.035 -33.155 ;
        RECT -10.365 -36.205 -10.035 -35.875 ;
        RECT -10.365 -38.925 -10.035 -38.595 ;
        RECT -10.365 -47.085 -10.035 -46.755 ;
        RECT -10.365 -48.445 -10.035 -48.115 ;
        RECT -10.365 -49.805 -10.035 -49.475 ;
        RECT -10.365 -51.165 -10.035 -50.835 ;
        RECT -10.365 -52.525 -10.035 -52.195 ;
        RECT -10.365 -53.885 -10.035 -53.555 ;
        RECT -10.365 -55.245 -10.035 -54.915 ;
        RECT -10.365 -56.605 -10.035 -56.275 ;
        RECT -10.365 -57.965 -10.035 -57.635 ;
        RECT -10.365 -59.325 -10.035 -58.995 ;
        RECT -10.365 -60.685 -10.035 -60.355 ;
        RECT -10.365 -62.045 -10.035 -61.715 ;
        RECT -10.365 -68.845 -10.035 -68.515 ;
        RECT -10.365 -72.925 -10.035 -72.595 ;
        RECT -10.365 -74.285 -10.035 -73.955 ;
        RECT -10.365 -75.645 -10.035 -75.315 ;
        RECT -10.365 -77.005 -10.035 -76.675 ;
        RECT -10.365 -78.365 -10.035 -78.035 ;
        RECT -10.365 -81.085 -10.035 -80.755 ;
        RECT -10.365 -82.445 -10.035 -82.115 ;
        RECT -10.365 -83.805 -10.035 -83.475 ;
        RECT -10.365 -85.165 -10.035 -84.835 ;
        RECT -10.365 -86.525 -10.035 -86.195 ;
        RECT -10.365 -87.885 -10.035 -87.555 ;
        RECT -10.365 -90.605 -10.035 -90.275 ;
        RECT -10.365 -91.965 -10.035 -91.635 ;
        RECT -10.365 -93.325 -10.035 -92.995 ;
        RECT -10.365 -94.685 -10.035 -94.355 ;
        RECT -10.365 -96.045 -10.035 -95.715 ;
        RECT -10.365 -97.405 -10.035 -97.075 ;
        RECT -10.365 -100.125 -10.035 -99.795 ;
        RECT -10.365 -101.485 -10.035 -101.155 ;
        RECT -10.365 -102.845 -10.035 -102.515 ;
        RECT -10.365 -105.565 -10.035 -105.235 ;
        RECT -10.365 -106.925 -10.035 -106.595 ;
        RECT -10.365 -108.285 -10.035 -107.955 ;
        RECT -10.365 -109.645 -10.035 -109.315 ;
        RECT -10.365 -111.005 -10.035 -110.675 ;
        RECT -10.365 -112.365 -10.035 -112.035 ;
        RECT -10.365 -113.725 -10.035 -113.395 ;
        RECT -10.365 -116.445 -10.035 -116.115 ;
        RECT -10.365 -119.165 -10.035 -118.835 ;
        RECT -10.365 -120.525 -10.035 -120.195 ;
        RECT -10.365 -121.885 -10.035 -121.555 ;
        RECT -10.365 -123.245 -10.035 -122.915 ;
        RECT -10.365 -125.965 -10.035 -125.635 ;
        RECT -10.365 -127.325 -10.035 -126.995 ;
        RECT -10.365 -128.685 -10.035 -128.355 ;
        RECT -10.365 -130.045 -10.035 -129.715 ;
        RECT -10.365 -131.405 -10.035 -131.075 ;
        RECT -10.365 -132.765 -10.035 -132.435 ;
        RECT -10.365 -140.925 -10.035 -140.595 ;
        RECT -10.365 -142.285 -10.035 -141.955 ;
        RECT -10.365 -145.005 -10.035 -144.675 ;
        RECT -10.365 -146.365 -10.035 -146.035 ;
        RECT -10.365 -147.725 -10.035 -147.395 ;
        RECT -10.365 -153.165 -10.035 -152.835 ;
        RECT -10.365 -154.525 -10.035 -154.195 ;
        RECT -10.365 -155.885 -10.035 -155.555 ;
        RECT -10.365 -157.245 -10.035 -156.915 ;
        RECT -10.365 -158.605 -10.035 -158.275 ;
        RECT -10.365 -159.965 -10.035 -159.635 ;
        RECT -10.365 -161.325 -10.035 -160.995 ;
        RECT -10.365 -164.045 -10.035 -163.715 ;
        RECT -10.365 -165.405 -10.035 -165.075 ;
        RECT -10.365 -166.765 -10.035 -166.435 ;
        RECT -10.365 -168.125 -10.035 -167.795 ;
        RECT -10.365 -170.845 -10.035 -170.515 ;
        RECT -10.365 -172.205 -10.035 -171.875 ;
        RECT -10.365 -173.565 -10.035 -173.235 ;
        RECT -10.365 -174.925 -10.035 -174.595 ;
        RECT -10.365 -176.285 -10.035 -175.955 ;
        RECT -10.365 -177.645 -10.035 -177.315 ;
        RECT -10.365 -179.005 -10.035 -178.675 ;
        RECT -10.365 -180.365 -10.035 -180.035 ;
        RECT -10.365 -181.725 -10.035 -181.395 ;
        RECT -10.365 -183.085 -10.035 -182.755 ;
        RECT -10.365 -184.445 -10.035 -184.115 ;
        RECT -10.365 -185.805 -10.035 -185.475 ;
        RECT -10.365 -187.165 -10.035 -186.835 ;
        RECT -10.365 -188.525 -10.035 -188.195 ;
        RECT -10.365 -189.885 -10.035 -189.555 ;
        RECT -10.365 -191.245 -10.035 -190.915 ;
        RECT -10.365 -192.605 -10.035 -192.275 ;
        RECT -10.365 -193.965 -10.035 -193.635 ;
        RECT -10.365 -195.325 -10.035 -194.995 ;
        RECT -10.365 -196.685 -10.035 -196.355 ;
        RECT -10.365 -198.045 -10.035 -197.715 ;
        RECT -10.365 -199.405 -10.035 -199.075 ;
        RECT -10.365 -203.485 -10.035 -203.155 ;
        RECT -10.365 -204.845 -10.035 -204.515 ;
        RECT -10.365 -206.205 -10.035 -205.875 ;
        RECT -10.365 -207.565 -10.035 -207.235 ;
        RECT -10.365 -208.925 -10.035 -208.595 ;
        RECT -10.365 -210.285 -10.035 -209.955 ;
        RECT -10.365 -211.645 -10.035 -211.315 ;
        RECT -10.365 -213.005 -10.035 -212.675 ;
        RECT -10.365 -214.365 -10.035 -214.035 ;
        RECT -10.365 -215.725 -10.035 -215.395 ;
        RECT -10.365 -217.085 -10.035 -216.755 ;
        RECT -10.365 -218.445 -10.035 -218.115 ;
        RECT -10.365 -219.805 -10.035 -219.475 ;
        RECT -10.365 -221.165 -10.035 -220.835 ;
        RECT -10.365 -222.525 -10.035 -222.195 ;
        RECT -10.365 -223.885 -10.035 -223.555 ;
        RECT -10.365 -225.245 -10.035 -224.915 ;
        RECT -10.365 -227.965 -10.035 -227.635 ;
        RECT -10.365 -232.045 -10.035 -231.715 ;
        RECT -10.365 -234.765 -10.035 -234.435 ;
        RECT -10.365 -236.125 -10.035 -235.795 ;
        RECT -10.365 -237.485 -10.035 -237.155 ;
        RECT -10.365 -238.845 -10.035 -238.515 ;
        RECT -10.365 -241.09 -10.035 -239.96 ;
        RECT -10.36 -241.205 -10.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 -223.885 -8.675 -223.555 ;
        RECT -9.005 -225.245 -8.675 -224.915 ;
        RECT -9.005 -226.605 -8.675 -226.275 ;
        RECT -9.005 -227.965 -8.675 -227.635 ;
        RECT -9.005 -229.325 -8.675 -228.995 ;
        RECT -9.005 -230.685 -8.675 -230.355 ;
        RECT -9.005 -232.045 -8.675 -231.715 ;
        RECT -9.005 -233.405 -8.675 -233.075 ;
        RECT -9.005 -234.765 -8.675 -234.435 ;
        RECT -9.005 -236.125 -8.675 -235.795 ;
        RECT -9.005 -237.485 -8.675 -237.155 ;
        RECT -9.005 -238.845 -8.675 -238.515 ;
        RECT -9.005 -241.09 -8.675 -239.96 ;
        RECT -9 -241.205 -8.68 245.285 ;
        RECT -9.005 244.04 -8.675 245.17 ;
        RECT -9.005 242.595 -8.675 242.925 ;
        RECT -9.005 241.235 -8.675 241.565 ;
        RECT -9.005 239.875 -8.675 240.205 ;
        RECT -9.005 238.515 -8.675 238.845 ;
        RECT -9.005 237.155 -8.675 237.485 ;
        RECT -9.005 235.795 -8.675 236.125 ;
        RECT -9.005 234.435 -8.675 234.765 ;
        RECT -9.005 233.075 -8.675 233.405 ;
        RECT -9.005 231.715 -8.675 232.045 ;
        RECT -9.005 227.635 -8.675 227.965 ;
        RECT -9.005 224.915 -8.675 225.245 ;
        RECT -9.005 218.115 -8.675 218.445 ;
        RECT -9.005 216.755 -8.675 217.085 ;
        RECT -9.005 207.235 -8.675 207.565 ;
        RECT -9.005 204.515 -8.675 204.845 ;
        RECT -9.005 203.155 -8.675 203.485 ;
        RECT -9.005 199.075 -8.675 199.405 ;
        RECT -9.005 196.355 -8.675 196.685 ;
        RECT -9.005 189.555 -8.675 189.885 ;
        RECT -9.005 188.195 -8.675 188.525 ;
        RECT -9.005 185.475 -8.675 185.805 ;
        RECT -9.005 178.675 -8.675 179.005 ;
        RECT -9.005 175.955 -8.675 176.285 ;
        RECT -9.005 174.595 -8.675 174.925 ;
        RECT -9.005 167.795 -8.675 168.125 ;
        RECT -9.005 160.995 -8.675 161.325 ;
        RECT -9.005 159.635 -8.675 159.965 ;
        RECT -9.005 156.915 -8.675 157.245 ;
        RECT -9.005 150.115 -8.675 150.445 ;
        RECT -9.005 147.395 -8.675 147.725 ;
        RECT -9.005 146.035 -8.675 146.365 ;
        RECT -9.005 139.235 -8.675 139.565 ;
        RECT -9.005 136.515 -8.675 136.845 ;
        RECT -9.005 132.435 -8.675 132.765 ;
        RECT -9.005 131.075 -8.675 131.405 ;
        RECT -9.005 128.355 -8.675 128.685 ;
        RECT -9.005 118.835 -8.675 119.165 ;
        RECT -9.005 117.475 -8.675 117.805 ;
        RECT -9.005 110.675 -8.675 111.005 ;
        RECT -9.005 107.955 -8.675 108.285 ;
        RECT -9.005 103.875 -8.675 104.205 ;
        RECT -9.005 99.795 -8.675 100.125 ;
        RECT -9.005 97.075 -8.675 97.405 ;
        RECT -9.005 90.275 -8.675 90.605 ;
        RECT -9.005 88.915 -8.675 89.245 ;
        RECT -9.005 82.115 -8.675 82.445 ;
        RECT -9.005 79.395 -8.675 79.725 ;
        RECT -9.005 75.315 -8.675 75.645 ;
        RECT -9.005 71.235 -8.675 71.565 ;
        RECT -9.005 68.515 -8.675 68.845 ;
        RECT -9.005 61.715 -8.675 62.045 ;
        RECT -9.005 60.355 -8.675 60.685 ;
        RECT -9.005 50.835 -8.675 51.165 ;
        RECT -9.005 46.755 -8.675 47.085 ;
        RECT -9.005 42.675 -8.675 43.005 ;
        RECT -9.005 39.955 -8.675 40.285 ;
        RECT -9.005 33.155 -8.675 33.485 ;
        RECT -9.005 31.795 -8.675 32.125 ;
        RECT -9.005 29.075 -8.675 29.405 ;
        RECT -9.005 22.275 -8.675 22.605 ;
        RECT -9.005 19.555 -8.675 19.885 ;
        RECT -9.005 18.195 -8.675 18.525 ;
        RECT -9.005 11.395 -8.675 11.725 ;
        RECT -9.005 4.595 -8.675 4.925 ;
        RECT -9.005 3.235 -8.675 3.565 ;
        RECT -9.005 1.875 -8.675 2.205 ;
        RECT -9.005 0.515 -8.675 0.845 ;
        RECT -9.005 -0.845 -8.675 -0.515 ;
        RECT -9.005 -2.205 -8.675 -1.875 ;
        RECT -9.005 -3.565 -8.675 -3.235 ;
        RECT -9.005 -4.925 -8.675 -4.595 ;
        RECT -9.005 -6.285 -8.675 -5.955 ;
        RECT -9.005 -7.645 -8.675 -7.315 ;
        RECT -9.005 -9.005 -8.675 -8.675 ;
        RECT -9.005 -10.365 -8.675 -10.035 ;
        RECT -9.005 -11.725 -8.675 -11.395 ;
        RECT -9.005 -13.085 -8.675 -12.755 ;
        RECT -9.005 -14.445 -8.675 -14.115 ;
        RECT -9.005 -15.805 -8.675 -15.475 ;
        RECT -9.005 -17.165 -8.675 -16.835 ;
        RECT -9.005 -18.525 -8.675 -18.195 ;
        RECT -9.005 -19.885 -8.675 -19.555 ;
        RECT -9.005 -21.245 -8.675 -20.915 ;
        RECT -9.005 -22.605 -8.675 -22.275 ;
        RECT -9.005 -23.965 -8.675 -23.635 ;
        RECT -9.005 -25.325 -8.675 -24.995 ;
        RECT -9.005 -26.685 -8.675 -26.355 ;
        RECT -9.005 -28.045 -8.675 -27.715 ;
        RECT -9.005 -29.405 -8.675 -29.075 ;
        RECT -9.005 -30.765 -8.675 -30.435 ;
        RECT -9.005 -32.125 -8.675 -31.795 ;
        RECT -9.005 -33.485 -8.675 -33.155 ;
        RECT -9.005 -34.845 -8.675 -34.515 ;
        RECT -9.005 -36.205 -8.675 -35.875 ;
        RECT -9.005 -37.565 -8.675 -37.235 ;
        RECT -9.005 -38.925 -8.675 -38.595 ;
        RECT -9.005 -40.285 -8.675 -39.955 ;
        RECT -9.005 -41.645 -8.675 -41.315 ;
        RECT -9.005 -43.005 -8.675 -42.675 ;
        RECT -9.005 -44.365 -8.675 -44.035 ;
        RECT -9.005 -45.725 -8.675 -45.395 ;
        RECT -9.005 -47.085 -8.675 -46.755 ;
        RECT -9.005 -48.445 -8.675 -48.115 ;
        RECT -9.005 -49.805 -8.675 -49.475 ;
        RECT -9.005 -51.165 -8.675 -50.835 ;
        RECT -9.005 -52.525 -8.675 -52.195 ;
        RECT -9.005 -53.885 -8.675 -53.555 ;
        RECT -9.005 -55.245 -8.675 -54.915 ;
        RECT -9.005 -56.605 -8.675 -56.275 ;
        RECT -9.005 -57.965 -8.675 -57.635 ;
        RECT -9.005 -59.325 -8.675 -58.995 ;
        RECT -9.005 -60.685 -8.675 -60.355 ;
        RECT -9.005 -62.045 -8.675 -61.715 ;
        RECT -9.005 -68.845 -8.675 -68.515 ;
        RECT -9.005 -70.205 -8.675 -69.875 ;
        RECT -9.005 -72.925 -8.675 -72.595 ;
        RECT -9.005 -74.285 -8.675 -73.955 ;
        RECT -9.005 -75.645 -8.675 -75.315 ;
        RECT -9.005 -77.005 -8.675 -76.675 ;
        RECT -9.005 -78.365 -8.675 -78.035 ;
        RECT -9.005 -79.725 -8.675 -79.395 ;
        RECT -9.005 -81.085 -8.675 -80.755 ;
        RECT -9.005 -82.445 -8.675 -82.115 ;
        RECT -9.005 -83.805 -8.675 -83.475 ;
        RECT -9.005 -85.165 -8.675 -84.835 ;
        RECT -9.005 -86.525 -8.675 -86.195 ;
        RECT -9.005 -87.885 -8.675 -87.555 ;
        RECT -9.005 -89.245 -8.675 -88.915 ;
        RECT -9.005 -90.605 -8.675 -90.275 ;
        RECT -9.005 -91.965 -8.675 -91.635 ;
        RECT -9.005 -93.325 -8.675 -92.995 ;
        RECT -9.005 -94.685 -8.675 -94.355 ;
        RECT -9.005 -96.045 -8.675 -95.715 ;
        RECT -9.005 -97.405 -8.675 -97.075 ;
        RECT -9.005 -98.765 -8.675 -98.435 ;
        RECT -9.005 -100.125 -8.675 -99.795 ;
        RECT -9.005 -101.485 -8.675 -101.155 ;
        RECT -9.005 -102.845 -8.675 -102.515 ;
        RECT -9.005 -104.205 -8.675 -103.875 ;
        RECT -9.005 -105.565 -8.675 -105.235 ;
        RECT -9.005 -106.925 -8.675 -106.595 ;
        RECT -9.005 -108.285 -8.675 -107.955 ;
        RECT -9.005 -109.645 -8.675 -109.315 ;
        RECT -9.005 -111.005 -8.675 -110.675 ;
        RECT -9.005 -112.365 -8.675 -112.035 ;
        RECT -9.005 -113.725 -8.675 -113.395 ;
        RECT -9.005 -115.085 -8.675 -114.755 ;
        RECT -9.005 -116.445 -8.675 -116.115 ;
        RECT -9.005 -119.165 -8.675 -118.835 ;
        RECT -9.005 -120.525 -8.675 -120.195 ;
        RECT -9.005 -121.885 -8.675 -121.555 ;
        RECT -9.005 -123.245 -8.675 -122.915 ;
        RECT -9.005 -124.605 -8.675 -124.275 ;
        RECT -9.005 -125.965 -8.675 -125.635 ;
        RECT -9.005 -127.325 -8.675 -126.995 ;
        RECT -9.005 -128.685 -8.675 -128.355 ;
        RECT -9.005 -130.045 -8.675 -129.715 ;
        RECT -9.005 -131.405 -8.675 -131.075 ;
        RECT -9.005 -132.765 -8.675 -132.435 ;
        RECT -9.005 -134.125 -8.675 -133.795 ;
        RECT -9.005 -140.925 -8.675 -140.595 ;
        RECT -9.005 -142.285 -8.675 -141.955 ;
        RECT -9.005 -143.645 -8.675 -143.315 ;
        RECT -9.005 -145.005 -8.675 -144.675 ;
        RECT -9.005 -146.365 -8.675 -146.035 ;
        RECT -9.005 -147.725 -8.675 -147.395 ;
        RECT -9.005 -149.085 -8.675 -148.755 ;
        RECT -9.005 -150.445 -8.675 -150.115 ;
        RECT -9.005 -151.805 -8.675 -151.475 ;
        RECT -9.005 -153.165 -8.675 -152.835 ;
        RECT -9.005 -154.525 -8.675 -154.195 ;
        RECT -9.005 -155.885 -8.675 -155.555 ;
        RECT -9.005 -157.245 -8.675 -156.915 ;
        RECT -9.005 -158.605 -8.675 -158.275 ;
        RECT -9.005 -159.965 -8.675 -159.635 ;
        RECT -9.005 -161.325 -8.675 -160.995 ;
        RECT -9.005 -162.685 -8.675 -162.355 ;
        RECT -9.005 -164.045 -8.675 -163.715 ;
        RECT -9.005 -165.405 -8.675 -165.075 ;
        RECT -9.005 -166.765 -8.675 -166.435 ;
        RECT -9.005 -168.125 -8.675 -167.795 ;
        RECT -9.005 -169.485 -8.675 -169.155 ;
        RECT -9.005 -170.845 -8.675 -170.515 ;
        RECT -9.005 -172.205 -8.675 -171.875 ;
        RECT -9.005 -173.565 -8.675 -173.235 ;
        RECT -9.005 -174.925 -8.675 -174.595 ;
        RECT -9.005 -176.285 -8.675 -175.955 ;
        RECT -9.005 -177.645 -8.675 -177.315 ;
        RECT -9.005 -179.005 -8.675 -178.675 ;
        RECT -9.005 -180.365 -8.675 -180.035 ;
        RECT -9.005 -181.725 -8.675 -181.395 ;
        RECT -9.005 -183.085 -8.675 -182.755 ;
        RECT -9.005 -184.445 -8.675 -184.115 ;
        RECT -9.005 -185.805 -8.675 -185.475 ;
        RECT -9.005 -187.165 -8.675 -186.835 ;
        RECT -9.005 -188.525 -8.675 -188.195 ;
        RECT -9.005 -189.885 -8.675 -189.555 ;
        RECT -9.005 -191.245 -8.675 -190.915 ;
        RECT -9.005 -192.605 -8.675 -192.275 ;
        RECT -9.005 -193.965 -8.675 -193.635 ;
        RECT -9.005 -195.325 -8.675 -194.995 ;
        RECT -9.005 -196.685 -8.675 -196.355 ;
        RECT -9.005 -198.045 -8.675 -197.715 ;
        RECT -9.005 -199.405 -8.675 -199.075 ;
        RECT -9.005 -200.765 -8.675 -200.435 ;
        RECT -9.005 -202.125 -8.675 -201.795 ;
        RECT -9.005 -203.485 -8.675 -203.155 ;
        RECT -9.005 -204.845 -8.675 -204.515 ;
        RECT -9.005 -206.205 -8.675 -205.875 ;
        RECT -9.005 -207.565 -8.675 -207.235 ;
        RECT -9.005 -208.925 -8.675 -208.595 ;
        RECT -9.005 -210.285 -8.675 -209.955 ;
        RECT -9.005 -211.645 -8.675 -211.315 ;
        RECT -9.005 -213.005 -8.675 -212.675 ;
        RECT -9.005 -214.365 -8.675 -214.035 ;
        RECT -9.005 -215.725 -8.675 -215.395 ;
        RECT -9.005 -217.085 -8.675 -216.755 ;
        RECT -9.005 -218.445 -8.675 -218.115 ;
        RECT -9.005 -219.805 -8.675 -219.475 ;
        RECT -9.005 -221.165 -8.675 -220.835 ;
        RECT -9.005 -222.525 -8.675 -222.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -128.685 -19.555 -128.355 ;
        RECT -19.885 -130.045 -19.555 -129.715 ;
        RECT -19.885 -131.405 -19.555 -131.075 ;
        RECT -19.885 -132.765 -19.555 -132.435 ;
        RECT -19.885 -138.205 -19.555 -137.875 ;
        RECT -19.885 -139.565 -19.555 -139.235 ;
        RECT -19.885 -140.925 -19.555 -140.595 ;
        RECT -19.885 -142.285 -19.555 -141.955 ;
        RECT -19.885 -143.03 -19.555 -142.7 ;
        RECT -19.885 -145.005 -19.555 -144.675 ;
        RECT -19.885 -146.365 -19.555 -146.035 ;
        RECT -19.885 -147.725 -19.555 -147.395 ;
        RECT -19.88 -148.4 -19.56 -127 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -230.685 -19.555 -230.355 ;
        RECT -19.885 -232.045 -19.555 -231.715 ;
        RECT -19.885 -233.225 -19.555 -232.895 ;
        RECT -19.885 -234.765 -19.555 -234.435 ;
        RECT -19.885 -236.125 -19.555 -235.795 ;
        RECT -19.885 -237.485 -19.555 -237.155 ;
        RECT -19.885 -238.845 -19.555 -238.515 ;
        RECT -19.885 -241.09 -19.555 -239.96 ;
        RECT -19.88 -241.205 -19.56 -227.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 244.04 -18.195 245.17 ;
        RECT -18.525 242.595 -18.195 242.925 ;
        RECT -18.525 241.235 -18.195 241.565 ;
        RECT -18.525 239.875 -18.195 240.205 ;
        RECT -18.525 238.515 -18.195 238.845 ;
        RECT -18.525 237.155 -18.195 237.485 ;
        RECT -18.525 235.795 -18.195 236.125 ;
        RECT -18.525 234.435 -18.195 234.765 ;
        RECT -18.525 233.075 -18.195 233.405 ;
        RECT -18.525 231.715 -18.195 232.045 ;
        RECT -18.525 230.355 -18.195 230.685 ;
        RECT -18.525 228.995 -18.195 229.325 ;
        RECT -18.525 227.635 -18.195 227.965 ;
        RECT -18.525 226.275 -18.195 226.605 ;
        RECT -18.525 224.915 -18.195 225.245 ;
        RECT -18.525 223.555 -18.195 223.885 ;
        RECT -18.525 222.195 -18.195 222.525 ;
        RECT -18.525 220.835 -18.195 221.165 ;
        RECT -18.525 219.475 -18.195 219.805 ;
        RECT -18.525 218.115 -18.195 218.445 ;
        RECT -18.525 216.755 -18.195 217.085 ;
        RECT -18.525 215.395 -18.195 215.725 ;
        RECT -18.525 214.035 -18.195 214.365 ;
        RECT -18.525 212.675 -18.195 213.005 ;
        RECT -18.525 211.315 -18.195 211.645 ;
        RECT -18.525 209.955 -18.195 210.285 ;
        RECT -18.525 208.595 -18.195 208.925 ;
        RECT -18.525 207.235 -18.195 207.565 ;
        RECT -18.525 205.875 -18.195 206.205 ;
        RECT -18.525 204.515 -18.195 204.845 ;
        RECT -18.525 203.155 -18.195 203.485 ;
        RECT -18.525 201.795 -18.195 202.125 ;
        RECT -18.525 200.435 -18.195 200.765 ;
        RECT -18.525 199.075 -18.195 199.405 ;
        RECT -18.525 197.715 -18.195 198.045 ;
        RECT -18.525 196.355 -18.195 196.685 ;
        RECT -18.525 194.995 -18.195 195.325 ;
        RECT -18.525 193.635 -18.195 193.965 ;
        RECT -18.525 192.275 -18.195 192.605 ;
        RECT -18.525 190.915 -18.195 191.245 ;
        RECT -18.525 189.555 -18.195 189.885 ;
        RECT -18.525 188.195 -18.195 188.525 ;
        RECT -18.525 186.835 -18.195 187.165 ;
        RECT -18.525 185.475 -18.195 185.805 ;
        RECT -18.525 184.115 -18.195 184.445 ;
        RECT -18.525 182.755 -18.195 183.085 ;
        RECT -18.525 181.395 -18.195 181.725 ;
        RECT -18.525 180.035 -18.195 180.365 ;
        RECT -18.525 178.675 -18.195 179.005 ;
        RECT -18.525 177.315 -18.195 177.645 ;
        RECT -18.525 175.955 -18.195 176.285 ;
        RECT -18.525 174.595 -18.195 174.925 ;
        RECT -18.525 173.235 -18.195 173.565 ;
        RECT -18.525 171.875 -18.195 172.205 ;
        RECT -18.525 170.515 -18.195 170.845 ;
        RECT -18.525 169.155 -18.195 169.485 ;
        RECT -18.525 167.795 -18.195 168.125 ;
        RECT -18.525 166.435 -18.195 166.765 ;
        RECT -18.525 165.075 -18.195 165.405 ;
        RECT -18.525 163.715 -18.195 164.045 ;
        RECT -18.525 162.355 -18.195 162.685 ;
        RECT -18.525 160.995 -18.195 161.325 ;
        RECT -18.525 159.635 -18.195 159.965 ;
        RECT -18.525 158.275 -18.195 158.605 ;
        RECT -18.525 156.915 -18.195 157.245 ;
        RECT -18.525 155.555 -18.195 155.885 ;
        RECT -18.525 154.195 -18.195 154.525 ;
        RECT -18.525 152.835 -18.195 153.165 ;
        RECT -18.525 151.475 -18.195 151.805 ;
        RECT -18.525 150.115 -18.195 150.445 ;
        RECT -18.525 148.755 -18.195 149.085 ;
        RECT -18.525 147.395 -18.195 147.725 ;
        RECT -18.525 146.035 -18.195 146.365 ;
        RECT -18.525 144.675 -18.195 145.005 ;
        RECT -18.525 143.315 -18.195 143.645 ;
        RECT -18.525 141.955 -18.195 142.285 ;
        RECT -18.525 140.595 -18.195 140.925 ;
        RECT -18.525 139.235 -18.195 139.565 ;
        RECT -18.525 137.875 -18.195 138.205 ;
        RECT -18.525 136.515 -18.195 136.845 ;
        RECT -18.525 135.155 -18.195 135.485 ;
        RECT -18.525 133.795 -18.195 134.125 ;
        RECT -18.525 132.435 -18.195 132.765 ;
        RECT -18.525 131.075 -18.195 131.405 ;
        RECT -18.525 129.715 -18.195 130.045 ;
        RECT -18.525 128.355 -18.195 128.685 ;
        RECT -18.525 126.995 -18.195 127.325 ;
        RECT -18.525 125.635 -18.195 125.965 ;
        RECT -18.525 124.275 -18.195 124.605 ;
        RECT -18.525 122.915 -18.195 123.245 ;
        RECT -18.525 121.555 -18.195 121.885 ;
        RECT -18.525 120.195 -18.195 120.525 ;
        RECT -18.525 118.835 -18.195 119.165 ;
        RECT -18.525 117.475 -18.195 117.805 ;
        RECT -18.525 116.115 -18.195 116.445 ;
        RECT -18.525 114.755 -18.195 115.085 ;
        RECT -18.525 113.395 -18.195 113.725 ;
        RECT -18.525 112.035 -18.195 112.365 ;
        RECT -18.525 110.675 -18.195 111.005 ;
        RECT -18.525 109.315 -18.195 109.645 ;
        RECT -18.525 107.955 -18.195 108.285 ;
        RECT -18.525 106.595 -18.195 106.925 ;
        RECT -18.525 105.235 -18.195 105.565 ;
        RECT -18.525 103.875 -18.195 104.205 ;
        RECT -18.525 102.515 -18.195 102.845 ;
        RECT -18.525 101.155 -18.195 101.485 ;
        RECT -18.525 99.795 -18.195 100.125 ;
        RECT -18.525 98.435 -18.195 98.765 ;
        RECT -18.525 97.075 -18.195 97.405 ;
        RECT -18.525 95.715 -18.195 96.045 ;
        RECT -18.525 94.355 -18.195 94.685 ;
        RECT -18.525 92.995 -18.195 93.325 ;
        RECT -18.525 91.635 -18.195 91.965 ;
        RECT -18.525 90.275 -18.195 90.605 ;
        RECT -18.525 88.915 -18.195 89.245 ;
        RECT -18.525 87.555 -18.195 87.885 ;
        RECT -18.525 86.195 -18.195 86.525 ;
        RECT -18.525 84.835 -18.195 85.165 ;
        RECT -18.525 83.475 -18.195 83.805 ;
        RECT -18.525 82.115 -18.195 82.445 ;
        RECT -18.525 80.755 -18.195 81.085 ;
        RECT -18.525 79.395 -18.195 79.725 ;
        RECT -18.525 78.035 -18.195 78.365 ;
        RECT -18.525 76.675 -18.195 77.005 ;
        RECT -18.525 75.315 -18.195 75.645 ;
        RECT -18.525 73.955 -18.195 74.285 ;
        RECT -18.525 72.595 -18.195 72.925 ;
        RECT -18.525 71.235 -18.195 71.565 ;
        RECT -18.525 69.875 -18.195 70.205 ;
        RECT -18.525 68.515 -18.195 68.845 ;
        RECT -18.525 67.155 -18.195 67.485 ;
        RECT -18.525 65.795 -18.195 66.125 ;
        RECT -18.525 64.435 -18.195 64.765 ;
        RECT -18.525 63.075 -18.195 63.405 ;
        RECT -18.525 61.715 -18.195 62.045 ;
        RECT -18.525 60.355 -18.195 60.685 ;
        RECT -18.525 58.995 -18.195 59.325 ;
        RECT -18.525 57.635 -18.195 57.965 ;
        RECT -18.525 56.275 -18.195 56.605 ;
        RECT -18.525 54.915 -18.195 55.245 ;
        RECT -18.525 53.555 -18.195 53.885 ;
        RECT -18.525 52.195 -18.195 52.525 ;
        RECT -18.525 50.835 -18.195 51.165 ;
        RECT -18.525 49.475 -18.195 49.805 ;
        RECT -18.525 48.115 -18.195 48.445 ;
        RECT -18.525 46.755 -18.195 47.085 ;
        RECT -18.525 45.395 -18.195 45.725 ;
        RECT -18.525 44.035 -18.195 44.365 ;
        RECT -18.525 42.675 -18.195 43.005 ;
        RECT -18.525 41.315 -18.195 41.645 ;
        RECT -18.525 39.955 -18.195 40.285 ;
        RECT -18.525 38.595 -18.195 38.925 ;
        RECT -18.525 37.235 -18.195 37.565 ;
        RECT -18.525 35.875 -18.195 36.205 ;
        RECT -18.525 34.515 -18.195 34.845 ;
        RECT -18.525 33.155 -18.195 33.485 ;
        RECT -18.525 31.795 -18.195 32.125 ;
        RECT -18.525 30.435 -18.195 30.765 ;
        RECT -18.525 29.075 -18.195 29.405 ;
        RECT -18.525 27.715 -18.195 28.045 ;
        RECT -18.525 26.355 -18.195 26.685 ;
        RECT -18.525 24.995 -18.195 25.325 ;
        RECT -18.525 23.635 -18.195 23.965 ;
        RECT -18.525 22.275 -18.195 22.605 ;
        RECT -18.525 20.915 -18.195 21.245 ;
        RECT -18.525 19.555 -18.195 19.885 ;
        RECT -18.525 18.195 -18.195 18.525 ;
        RECT -18.525 16.835 -18.195 17.165 ;
        RECT -18.525 15.475 -18.195 15.805 ;
        RECT -18.525 14.115 -18.195 14.445 ;
        RECT -18.525 12.755 -18.195 13.085 ;
        RECT -18.525 11.395 -18.195 11.725 ;
        RECT -18.525 10.035 -18.195 10.365 ;
        RECT -18.525 8.675 -18.195 9.005 ;
        RECT -18.525 7.315 -18.195 7.645 ;
        RECT -18.525 5.955 -18.195 6.285 ;
        RECT -18.525 4.595 -18.195 4.925 ;
        RECT -18.525 3.235 -18.195 3.565 ;
        RECT -18.525 1.875 -18.195 2.205 ;
        RECT -18.525 0.515 -18.195 0.845 ;
        RECT -18.525 -2.205 -18.195 -1.875 ;
        RECT -18.525 -3.565 -18.195 -3.235 ;
        RECT -18.525 -7.645 -18.195 -7.315 ;
        RECT -18.525 -10.365 -18.195 -10.035 ;
        RECT -18.525 -11.725 -18.195 -11.395 ;
        RECT -18.525 -13.7 -18.195 -13.37 ;
        RECT -18.525 -14.445 -18.195 -14.115 ;
        RECT -18.525 -15.805 -18.195 -15.475 ;
        RECT -18.525 -18.79 -18.195 -18.46 ;
        RECT -18.525 -19.885 -18.195 -19.555 ;
        RECT -18.52 -19.885 -18.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -128.685 -18.195 -128.355 ;
        RECT -18.525 -130.045 -18.195 -129.715 ;
        RECT -18.525 -131.405 -18.195 -131.075 ;
        RECT -18.525 -132.765 -18.195 -132.435 ;
        RECT -18.525 -138.205 -18.195 -137.875 ;
        RECT -18.525 -139.565 -18.195 -139.235 ;
        RECT -18.525 -140.925 -18.195 -140.595 ;
        RECT -18.525 -142.285 -18.195 -141.955 ;
        RECT -18.525 -143.03 -18.195 -142.7 ;
        RECT -18.525 -145.005 -18.195 -144.675 ;
        RECT -18.525 -146.365 -18.195 -146.035 ;
        RECT -18.525 -147.725 -18.195 -147.395 ;
        RECT -18.52 -147.725 -18.2 -128.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -230.685 -18.195 -230.355 ;
        RECT -18.525 -232.045 -18.195 -231.715 ;
        RECT -18.525 -233.225 -18.195 -232.895 ;
        RECT -18.525 -234.765 -18.195 -234.435 ;
        RECT -18.525 -236.125 -18.195 -235.795 ;
        RECT -18.525 -237.485 -18.195 -237.155 ;
        RECT -18.525 -238.845 -18.195 -238.515 ;
        RECT -18.525 -241.09 -18.195 -239.96 ;
        RECT -18.52 -241.205 -18.2 -229 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 244.04 -16.835 245.17 ;
        RECT -17.165 242.595 -16.835 242.925 ;
        RECT -17.165 241.235 -16.835 241.565 ;
        RECT -17.165 239.875 -16.835 240.205 ;
        RECT -17.165 238.515 -16.835 238.845 ;
        RECT -17.165 237.155 -16.835 237.485 ;
        RECT -17.165 235.795 -16.835 236.125 ;
        RECT -17.165 234.435 -16.835 234.765 ;
        RECT -17.165 233.075 -16.835 233.405 ;
        RECT -17.165 231.715 -16.835 232.045 ;
        RECT -17.165 230.355 -16.835 230.685 ;
        RECT -17.165 228.995 -16.835 229.325 ;
        RECT -17.165 227.635 -16.835 227.965 ;
        RECT -17.165 226.275 -16.835 226.605 ;
        RECT -17.165 224.915 -16.835 225.245 ;
        RECT -17.165 223.555 -16.835 223.885 ;
        RECT -17.165 222.195 -16.835 222.525 ;
        RECT -17.165 220.835 -16.835 221.165 ;
        RECT -17.165 219.475 -16.835 219.805 ;
        RECT -17.165 218.115 -16.835 218.445 ;
        RECT -17.165 216.755 -16.835 217.085 ;
        RECT -17.165 215.395 -16.835 215.725 ;
        RECT -17.165 214.035 -16.835 214.365 ;
        RECT -17.165 212.675 -16.835 213.005 ;
        RECT -17.165 211.315 -16.835 211.645 ;
        RECT -17.165 209.955 -16.835 210.285 ;
        RECT -17.165 208.595 -16.835 208.925 ;
        RECT -17.165 207.235 -16.835 207.565 ;
        RECT -17.165 205.875 -16.835 206.205 ;
        RECT -17.165 204.515 -16.835 204.845 ;
        RECT -17.165 203.155 -16.835 203.485 ;
        RECT -17.165 201.795 -16.835 202.125 ;
        RECT -17.165 200.435 -16.835 200.765 ;
        RECT -17.165 199.075 -16.835 199.405 ;
        RECT -17.165 197.715 -16.835 198.045 ;
        RECT -17.165 196.355 -16.835 196.685 ;
        RECT -17.165 194.995 -16.835 195.325 ;
        RECT -17.165 193.635 -16.835 193.965 ;
        RECT -17.165 192.275 -16.835 192.605 ;
        RECT -17.165 190.915 -16.835 191.245 ;
        RECT -17.165 189.555 -16.835 189.885 ;
        RECT -17.165 188.195 -16.835 188.525 ;
        RECT -17.165 186.835 -16.835 187.165 ;
        RECT -17.165 185.475 -16.835 185.805 ;
        RECT -17.165 184.115 -16.835 184.445 ;
        RECT -17.165 182.755 -16.835 183.085 ;
        RECT -17.165 181.395 -16.835 181.725 ;
        RECT -17.165 180.035 -16.835 180.365 ;
        RECT -17.165 178.675 -16.835 179.005 ;
        RECT -17.165 177.315 -16.835 177.645 ;
        RECT -17.165 175.955 -16.835 176.285 ;
        RECT -17.165 174.595 -16.835 174.925 ;
        RECT -17.165 173.235 -16.835 173.565 ;
        RECT -17.165 171.875 -16.835 172.205 ;
        RECT -17.165 170.515 -16.835 170.845 ;
        RECT -17.165 169.155 -16.835 169.485 ;
        RECT -17.165 167.795 -16.835 168.125 ;
        RECT -17.165 166.435 -16.835 166.765 ;
        RECT -17.165 165.075 -16.835 165.405 ;
        RECT -17.165 163.715 -16.835 164.045 ;
        RECT -17.165 162.355 -16.835 162.685 ;
        RECT -17.165 160.995 -16.835 161.325 ;
        RECT -17.165 159.635 -16.835 159.965 ;
        RECT -17.165 158.275 -16.835 158.605 ;
        RECT -17.165 156.915 -16.835 157.245 ;
        RECT -17.165 155.555 -16.835 155.885 ;
        RECT -17.165 154.195 -16.835 154.525 ;
        RECT -17.165 152.835 -16.835 153.165 ;
        RECT -17.165 151.475 -16.835 151.805 ;
        RECT -17.165 150.115 -16.835 150.445 ;
        RECT -17.165 148.755 -16.835 149.085 ;
        RECT -17.165 147.395 -16.835 147.725 ;
        RECT -17.165 146.035 -16.835 146.365 ;
        RECT -17.165 144.675 -16.835 145.005 ;
        RECT -17.165 143.315 -16.835 143.645 ;
        RECT -17.165 141.955 -16.835 142.285 ;
        RECT -17.165 140.595 -16.835 140.925 ;
        RECT -17.165 139.235 -16.835 139.565 ;
        RECT -17.165 137.875 -16.835 138.205 ;
        RECT -17.165 136.515 -16.835 136.845 ;
        RECT -17.165 135.155 -16.835 135.485 ;
        RECT -17.165 133.795 -16.835 134.125 ;
        RECT -17.165 132.435 -16.835 132.765 ;
        RECT -17.165 131.075 -16.835 131.405 ;
        RECT -17.165 129.715 -16.835 130.045 ;
        RECT -17.165 128.355 -16.835 128.685 ;
        RECT -17.165 126.995 -16.835 127.325 ;
        RECT -17.165 125.635 -16.835 125.965 ;
        RECT -17.165 124.275 -16.835 124.605 ;
        RECT -17.165 122.915 -16.835 123.245 ;
        RECT -17.165 121.555 -16.835 121.885 ;
        RECT -17.165 120.195 -16.835 120.525 ;
        RECT -17.165 118.835 -16.835 119.165 ;
        RECT -17.165 117.475 -16.835 117.805 ;
        RECT -17.165 116.115 -16.835 116.445 ;
        RECT -17.165 114.755 -16.835 115.085 ;
        RECT -17.165 113.395 -16.835 113.725 ;
        RECT -17.165 112.035 -16.835 112.365 ;
        RECT -17.165 110.675 -16.835 111.005 ;
        RECT -17.165 109.315 -16.835 109.645 ;
        RECT -17.165 107.955 -16.835 108.285 ;
        RECT -17.165 106.595 -16.835 106.925 ;
        RECT -17.165 105.235 -16.835 105.565 ;
        RECT -17.165 103.875 -16.835 104.205 ;
        RECT -17.165 102.515 -16.835 102.845 ;
        RECT -17.165 101.155 -16.835 101.485 ;
        RECT -17.165 99.795 -16.835 100.125 ;
        RECT -17.165 98.435 -16.835 98.765 ;
        RECT -17.165 97.075 -16.835 97.405 ;
        RECT -17.165 95.715 -16.835 96.045 ;
        RECT -17.165 94.355 -16.835 94.685 ;
        RECT -17.165 92.995 -16.835 93.325 ;
        RECT -17.165 91.635 -16.835 91.965 ;
        RECT -17.165 90.275 -16.835 90.605 ;
        RECT -17.165 88.915 -16.835 89.245 ;
        RECT -17.165 87.555 -16.835 87.885 ;
        RECT -17.165 86.195 -16.835 86.525 ;
        RECT -17.165 84.835 -16.835 85.165 ;
        RECT -17.165 83.475 -16.835 83.805 ;
        RECT -17.165 82.115 -16.835 82.445 ;
        RECT -17.165 80.755 -16.835 81.085 ;
        RECT -17.165 79.395 -16.835 79.725 ;
        RECT -17.165 78.035 -16.835 78.365 ;
        RECT -17.165 76.675 -16.835 77.005 ;
        RECT -17.165 75.315 -16.835 75.645 ;
        RECT -17.165 73.955 -16.835 74.285 ;
        RECT -17.165 72.595 -16.835 72.925 ;
        RECT -17.165 71.235 -16.835 71.565 ;
        RECT -17.165 69.875 -16.835 70.205 ;
        RECT -17.165 68.515 -16.835 68.845 ;
        RECT -17.165 67.155 -16.835 67.485 ;
        RECT -17.165 65.795 -16.835 66.125 ;
        RECT -17.165 64.435 -16.835 64.765 ;
        RECT -17.165 63.075 -16.835 63.405 ;
        RECT -17.165 61.715 -16.835 62.045 ;
        RECT -17.165 60.355 -16.835 60.685 ;
        RECT -17.165 58.995 -16.835 59.325 ;
        RECT -17.165 57.635 -16.835 57.965 ;
        RECT -17.165 56.275 -16.835 56.605 ;
        RECT -17.165 54.915 -16.835 55.245 ;
        RECT -17.165 53.555 -16.835 53.885 ;
        RECT -17.165 52.195 -16.835 52.525 ;
        RECT -17.165 50.835 -16.835 51.165 ;
        RECT -17.165 49.475 -16.835 49.805 ;
        RECT -17.165 48.115 -16.835 48.445 ;
        RECT -17.165 46.755 -16.835 47.085 ;
        RECT -17.165 45.395 -16.835 45.725 ;
        RECT -17.165 44.035 -16.835 44.365 ;
        RECT -17.165 42.675 -16.835 43.005 ;
        RECT -17.165 41.315 -16.835 41.645 ;
        RECT -17.165 39.955 -16.835 40.285 ;
        RECT -17.165 38.595 -16.835 38.925 ;
        RECT -17.165 37.235 -16.835 37.565 ;
        RECT -17.165 35.875 -16.835 36.205 ;
        RECT -17.165 34.515 -16.835 34.845 ;
        RECT -17.165 33.155 -16.835 33.485 ;
        RECT -17.165 31.795 -16.835 32.125 ;
        RECT -17.165 30.435 -16.835 30.765 ;
        RECT -17.165 29.075 -16.835 29.405 ;
        RECT -17.165 27.715 -16.835 28.045 ;
        RECT -17.165 26.355 -16.835 26.685 ;
        RECT -17.165 24.995 -16.835 25.325 ;
        RECT -17.165 23.635 -16.835 23.965 ;
        RECT -17.165 22.275 -16.835 22.605 ;
        RECT -17.165 20.915 -16.835 21.245 ;
        RECT -17.165 19.555 -16.835 19.885 ;
        RECT -17.165 18.195 -16.835 18.525 ;
        RECT -17.165 16.835 -16.835 17.165 ;
        RECT -17.165 15.475 -16.835 15.805 ;
        RECT -17.165 14.115 -16.835 14.445 ;
        RECT -17.165 12.755 -16.835 13.085 ;
        RECT -17.165 11.395 -16.835 11.725 ;
        RECT -17.165 10.035 -16.835 10.365 ;
        RECT -17.165 8.675 -16.835 9.005 ;
        RECT -17.165 7.315 -16.835 7.645 ;
        RECT -17.165 5.955 -16.835 6.285 ;
        RECT -17.165 4.595 -16.835 4.925 ;
        RECT -17.165 3.235 -16.835 3.565 ;
        RECT -17.165 1.875 -16.835 2.205 ;
        RECT -17.165 0.515 -16.835 0.845 ;
        RECT -17.165 -2.205 -16.835 -1.875 ;
        RECT -17.165 -3.565 -16.835 -3.235 ;
        RECT -17.165 -4.925 -16.835 -4.595 ;
        RECT -17.165 -7.645 -16.835 -7.315 ;
        RECT -17.165 -10.365 -16.835 -10.035 ;
        RECT -17.165 -11.725 -16.835 -11.395 ;
        RECT -17.165 -13.7 -16.835 -13.37 ;
        RECT -17.165 -14.445 -16.835 -14.115 ;
        RECT -17.165 -15.805 -16.835 -15.475 ;
        RECT -17.165 -18.79 -16.835 -18.46 ;
        RECT -17.165 -19.885 -16.835 -19.555 ;
        RECT -17.165 -23.965 -16.835 -23.635 ;
        RECT -17.165 -25.325 -16.835 -24.995 ;
        RECT -17.165 -26.685 -16.835 -26.355 ;
        RECT -17.165 -29.405 -16.835 -29.075 ;
        RECT -17.165 -32.125 -16.835 -31.795 ;
        RECT -17.165 -33.485 -16.835 -33.155 ;
        RECT -17.165 -34.88 -16.835 -34.55 ;
        RECT -17.165 -36.205 -16.835 -35.875 ;
        RECT -17.165 -38.925 -16.835 -38.595 ;
        RECT -17.165 -39.97 -16.835 -39.64 ;
        RECT -17.165 -47.085 -16.835 -46.755 ;
        RECT -17.165 -48.445 -16.835 -48.115 ;
        RECT -17.165 -49.805 -16.835 -49.475 ;
        RECT -17.165 -51.165 -16.835 -50.835 ;
        RECT -17.165 -52.525 -16.835 -52.195 ;
        RECT -17.165 -53.885 -16.835 -53.555 ;
        RECT -17.165 -55.245 -16.835 -54.915 ;
        RECT -17.165 -56.605 -16.835 -56.275 ;
        RECT -17.165 -57.965 -16.835 -57.635 ;
        RECT -17.165 -59.325 -16.835 -58.995 ;
        RECT -17.165 -60.685 -16.835 -60.355 ;
        RECT -17.165 -62.045 -16.835 -61.715 ;
        RECT -17.165 -63.405 -16.835 -63.075 ;
        RECT -17.165 -68.845 -16.835 -68.515 ;
        RECT -17.165 -71.565 -16.835 -71.235 ;
        RECT -17.165 -72.925 -16.835 -72.595 ;
        RECT -17.165 -74.285 -16.835 -73.955 ;
        RECT -17.165 -75.645 -16.835 -75.315 ;
        RECT -17.165 -77.005 -16.835 -76.675 ;
        RECT -17.165 -78.365 -16.835 -78.035 ;
        RECT -17.165 -80.31 -16.835 -79.98 ;
        RECT -17.165 -81.085 -16.835 -80.755 ;
        RECT -17.165 -82.445 -16.835 -82.115 ;
        RECT -17.165 -83.805 -16.835 -83.475 ;
        RECT -17.165 -85.165 -16.835 -84.835 ;
        RECT -17.165 -86.525 -16.835 -86.195 ;
        RECT -17.165 -87.885 -16.835 -87.555 ;
        RECT -17.165 -90.605 -16.835 -90.275 ;
        RECT -17.165 -91.965 -16.835 -91.635 ;
        RECT -17.165 -93.325 -16.835 -92.995 ;
        RECT -17.165 -94.685 -16.835 -94.355 ;
        RECT -17.165 -96.045 -16.835 -95.715 ;
        RECT -17.165 -97.405 -16.835 -97.075 ;
        RECT -17.165 -98.85 -16.835 -98.52 ;
        RECT -17.165 -100.125 -16.835 -99.795 ;
        RECT -17.165 -101.485 -16.835 -101.155 ;
        RECT -17.165 -102.845 -16.835 -102.515 ;
        RECT -17.165 -105.565 -16.835 -105.235 ;
        RECT -17.165 -106.925 -16.835 -106.595 ;
        RECT -17.165 -108.285 -16.835 -107.955 ;
        RECT -17.165 -109.645 -16.835 -109.315 ;
        RECT -17.165 -111.005 -16.835 -110.675 ;
        RECT -17.165 -112.365 -16.835 -112.035 ;
        RECT -17.165 -113.725 -16.835 -113.395 ;
        RECT -17.165 -116.445 -16.835 -116.115 ;
        RECT -17.165 -117.805 -16.835 -117.475 ;
        RECT -17.165 -119.165 -16.835 -118.835 ;
        RECT -17.165 -120.525 -16.835 -120.195 ;
        RECT -17.165 -121.885 -16.835 -121.555 ;
        RECT -17.165 -123.245 -16.835 -122.915 ;
        RECT -17.165 -124.49 -16.835 -124.16 ;
        RECT -17.165 -125.965 -16.835 -125.635 ;
        RECT -17.165 -127.325 -16.835 -126.995 ;
        RECT -17.165 -128.685 -16.835 -128.355 ;
        RECT -17.165 -130.045 -16.835 -129.715 ;
        RECT -17.165 -131.405 -16.835 -131.075 ;
        RECT -17.165 -132.765 -16.835 -132.435 ;
        RECT -17.165 -139.565 -16.835 -139.235 ;
        RECT -17.165 -140.925 -16.835 -140.595 ;
        RECT -17.165 -142.285 -16.835 -141.955 ;
        RECT -17.165 -143.03 -16.835 -142.7 ;
        RECT -17.165 -145.005 -16.835 -144.675 ;
        RECT -17.165 -146.365 -16.835 -146.035 ;
        RECT -17.165 -147.725 -16.835 -147.395 ;
        RECT -17.165 -153.165 -16.835 -152.835 ;
        RECT -17.165 -154.525 -16.835 -154.195 ;
        RECT -17.165 -155.885 -16.835 -155.555 ;
        RECT -17.165 -157.245 -16.835 -156.915 ;
        RECT -17.165 -164.045 -16.835 -163.715 ;
        RECT -17.165 -168.125 -16.835 -167.795 ;
        RECT -17.165 -169.485 -16.835 -169.155 ;
        RECT -17.165 -170.845 -16.835 -170.515 ;
        RECT -17.165 -172.205 -16.835 -171.875 ;
        RECT -17.165 -174.925 -16.835 -174.595 ;
        RECT -17.165 -176.285 -16.835 -175.955 ;
        RECT -17.165 -177.645 -16.835 -177.315 ;
        RECT -17.165 -179.005 -16.835 -178.675 ;
        RECT -17.165 -180.365 -16.835 -180.035 ;
        RECT -17.165 -181.725 -16.835 -181.395 ;
        RECT -17.165 -183.085 -16.835 -182.755 ;
        RECT -17.165 -192.605 -16.835 -192.275 ;
        RECT -17.165 -195.325 -16.835 -194.995 ;
        RECT -17.165 -198.045 -16.835 -197.715 ;
        RECT -17.165 -202.125 -16.835 -201.795 ;
        RECT -17.165 -203.485 -16.835 -203.155 ;
        RECT -17.165 -208.925 -16.835 -208.595 ;
        RECT -17.165 -210.285 -16.835 -209.955 ;
        RECT -17.165 -214.365 -16.835 -214.035 ;
        RECT -17.165 -215.725 -16.835 -215.395 ;
        RECT -17.165 -217.085 -16.835 -216.755 ;
        RECT -17.165 -218.445 -16.835 -218.115 ;
        RECT -17.165 -219.805 -16.835 -219.475 ;
        RECT -17.165 -221.165 -16.835 -220.835 ;
        RECT -17.165 -222.525 -16.835 -222.195 ;
        RECT -17.165 -223.885 -16.835 -223.555 ;
        RECT -17.16 -224.56 -16.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -232.045 -16.835 -231.715 ;
        RECT -17.165 -233.225 -16.835 -232.895 ;
        RECT -17.165 -234.765 -16.835 -234.435 ;
        RECT -17.165 -236.125 -16.835 -235.795 ;
        RECT -17.165 -237.485 -16.835 -237.155 ;
        RECT -17.165 -238.845 -16.835 -238.515 ;
        RECT -17.165 -241.09 -16.835 -239.96 ;
        RECT -17.16 -241.205 -16.84 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 244.04 -15.475 245.17 ;
        RECT -15.805 242.595 -15.475 242.925 ;
        RECT -15.805 241.235 -15.475 241.565 ;
        RECT -15.805 239.875 -15.475 240.205 ;
        RECT -15.805 238.515 -15.475 238.845 ;
        RECT -15.805 237.155 -15.475 237.485 ;
        RECT -15.805 235.795 -15.475 236.125 ;
        RECT -15.805 234.435 -15.475 234.765 ;
        RECT -15.805 233.075 -15.475 233.405 ;
        RECT -15.805 231.715 -15.475 232.045 ;
        RECT -15.805 230.355 -15.475 230.685 ;
        RECT -15.805 228.995 -15.475 229.325 ;
        RECT -15.805 227.635 -15.475 227.965 ;
        RECT -15.805 226.275 -15.475 226.605 ;
        RECT -15.805 224.915 -15.475 225.245 ;
        RECT -15.805 223.555 -15.475 223.885 ;
        RECT -15.805 222.195 -15.475 222.525 ;
        RECT -15.805 220.835 -15.475 221.165 ;
        RECT -15.805 219.475 -15.475 219.805 ;
        RECT -15.805 218.115 -15.475 218.445 ;
        RECT -15.805 216.755 -15.475 217.085 ;
        RECT -15.805 215.395 -15.475 215.725 ;
        RECT -15.805 214.035 -15.475 214.365 ;
        RECT -15.805 212.675 -15.475 213.005 ;
        RECT -15.805 211.315 -15.475 211.645 ;
        RECT -15.805 209.955 -15.475 210.285 ;
        RECT -15.805 208.595 -15.475 208.925 ;
        RECT -15.805 207.235 -15.475 207.565 ;
        RECT -15.805 205.875 -15.475 206.205 ;
        RECT -15.805 204.515 -15.475 204.845 ;
        RECT -15.805 203.155 -15.475 203.485 ;
        RECT -15.805 201.795 -15.475 202.125 ;
        RECT -15.805 200.435 -15.475 200.765 ;
        RECT -15.805 199.075 -15.475 199.405 ;
        RECT -15.805 197.715 -15.475 198.045 ;
        RECT -15.805 196.355 -15.475 196.685 ;
        RECT -15.805 194.995 -15.475 195.325 ;
        RECT -15.805 193.635 -15.475 193.965 ;
        RECT -15.805 192.275 -15.475 192.605 ;
        RECT -15.805 190.915 -15.475 191.245 ;
        RECT -15.805 189.555 -15.475 189.885 ;
        RECT -15.805 188.195 -15.475 188.525 ;
        RECT -15.805 186.835 -15.475 187.165 ;
        RECT -15.805 185.475 -15.475 185.805 ;
        RECT -15.805 184.115 -15.475 184.445 ;
        RECT -15.805 182.755 -15.475 183.085 ;
        RECT -15.805 181.395 -15.475 181.725 ;
        RECT -15.805 180.035 -15.475 180.365 ;
        RECT -15.805 178.675 -15.475 179.005 ;
        RECT -15.805 177.315 -15.475 177.645 ;
        RECT -15.805 175.955 -15.475 176.285 ;
        RECT -15.805 174.595 -15.475 174.925 ;
        RECT -15.805 173.235 -15.475 173.565 ;
        RECT -15.805 171.875 -15.475 172.205 ;
        RECT -15.805 170.515 -15.475 170.845 ;
        RECT -15.805 169.155 -15.475 169.485 ;
        RECT -15.805 167.795 -15.475 168.125 ;
        RECT -15.805 166.435 -15.475 166.765 ;
        RECT -15.805 165.075 -15.475 165.405 ;
        RECT -15.805 163.715 -15.475 164.045 ;
        RECT -15.805 162.355 -15.475 162.685 ;
        RECT -15.805 160.995 -15.475 161.325 ;
        RECT -15.805 159.635 -15.475 159.965 ;
        RECT -15.805 158.275 -15.475 158.605 ;
        RECT -15.805 156.915 -15.475 157.245 ;
        RECT -15.805 155.555 -15.475 155.885 ;
        RECT -15.805 154.195 -15.475 154.525 ;
        RECT -15.805 152.835 -15.475 153.165 ;
        RECT -15.805 151.475 -15.475 151.805 ;
        RECT -15.805 150.115 -15.475 150.445 ;
        RECT -15.805 148.755 -15.475 149.085 ;
        RECT -15.805 147.395 -15.475 147.725 ;
        RECT -15.805 146.035 -15.475 146.365 ;
        RECT -15.805 144.675 -15.475 145.005 ;
        RECT -15.805 143.315 -15.475 143.645 ;
        RECT -15.805 141.955 -15.475 142.285 ;
        RECT -15.805 140.595 -15.475 140.925 ;
        RECT -15.805 139.235 -15.475 139.565 ;
        RECT -15.805 137.875 -15.475 138.205 ;
        RECT -15.805 136.515 -15.475 136.845 ;
        RECT -15.805 135.155 -15.475 135.485 ;
        RECT -15.805 133.795 -15.475 134.125 ;
        RECT -15.805 132.435 -15.475 132.765 ;
        RECT -15.805 131.075 -15.475 131.405 ;
        RECT -15.805 129.715 -15.475 130.045 ;
        RECT -15.805 128.355 -15.475 128.685 ;
        RECT -15.805 126.995 -15.475 127.325 ;
        RECT -15.805 125.635 -15.475 125.965 ;
        RECT -15.805 124.275 -15.475 124.605 ;
        RECT -15.805 122.915 -15.475 123.245 ;
        RECT -15.805 121.555 -15.475 121.885 ;
        RECT -15.805 120.195 -15.475 120.525 ;
        RECT -15.805 118.835 -15.475 119.165 ;
        RECT -15.805 117.475 -15.475 117.805 ;
        RECT -15.805 116.115 -15.475 116.445 ;
        RECT -15.805 114.755 -15.475 115.085 ;
        RECT -15.805 113.395 -15.475 113.725 ;
        RECT -15.805 112.035 -15.475 112.365 ;
        RECT -15.805 110.675 -15.475 111.005 ;
        RECT -15.805 109.315 -15.475 109.645 ;
        RECT -15.805 107.955 -15.475 108.285 ;
        RECT -15.805 106.595 -15.475 106.925 ;
        RECT -15.805 105.235 -15.475 105.565 ;
        RECT -15.805 103.875 -15.475 104.205 ;
        RECT -15.805 102.515 -15.475 102.845 ;
        RECT -15.805 101.155 -15.475 101.485 ;
        RECT -15.805 99.795 -15.475 100.125 ;
        RECT -15.805 98.435 -15.475 98.765 ;
        RECT -15.805 97.075 -15.475 97.405 ;
        RECT -15.805 95.715 -15.475 96.045 ;
        RECT -15.805 94.355 -15.475 94.685 ;
        RECT -15.805 92.995 -15.475 93.325 ;
        RECT -15.805 91.635 -15.475 91.965 ;
        RECT -15.805 90.275 -15.475 90.605 ;
        RECT -15.805 88.915 -15.475 89.245 ;
        RECT -15.805 87.555 -15.475 87.885 ;
        RECT -15.805 86.195 -15.475 86.525 ;
        RECT -15.805 84.835 -15.475 85.165 ;
        RECT -15.805 83.475 -15.475 83.805 ;
        RECT -15.805 82.115 -15.475 82.445 ;
        RECT -15.805 80.755 -15.475 81.085 ;
        RECT -15.805 79.395 -15.475 79.725 ;
        RECT -15.805 78.035 -15.475 78.365 ;
        RECT -15.805 76.675 -15.475 77.005 ;
        RECT -15.805 75.315 -15.475 75.645 ;
        RECT -15.805 73.955 -15.475 74.285 ;
        RECT -15.805 72.595 -15.475 72.925 ;
        RECT -15.805 71.235 -15.475 71.565 ;
        RECT -15.805 69.875 -15.475 70.205 ;
        RECT -15.805 68.515 -15.475 68.845 ;
        RECT -15.805 67.155 -15.475 67.485 ;
        RECT -15.805 65.795 -15.475 66.125 ;
        RECT -15.805 64.435 -15.475 64.765 ;
        RECT -15.805 63.075 -15.475 63.405 ;
        RECT -15.805 61.715 -15.475 62.045 ;
        RECT -15.805 60.355 -15.475 60.685 ;
        RECT -15.805 58.995 -15.475 59.325 ;
        RECT -15.805 57.635 -15.475 57.965 ;
        RECT -15.805 56.275 -15.475 56.605 ;
        RECT -15.805 54.915 -15.475 55.245 ;
        RECT -15.805 53.555 -15.475 53.885 ;
        RECT -15.805 52.195 -15.475 52.525 ;
        RECT -15.805 50.835 -15.475 51.165 ;
        RECT -15.805 49.475 -15.475 49.805 ;
        RECT -15.805 48.115 -15.475 48.445 ;
        RECT -15.805 46.755 -15.475 47.085 ;
        RECT -15.805 45.395 -15.475 45.725 ;
        RECT -15.805 44.035 -15.475 44.365 ;
        RECT -15.805 42.675 -15.475 43.005 ;
        RECT -15.805 41.315 -15.475 41.645 ;
        RECT -15.805 39.955 -15.475 40.285 ;
        RECT -15.805 38.595 -15.475 38.925 ;
        RECT -15.805 37.235 -15.475 37.565 ;
        RECT -15.805 35.875 -15.475 36.205 ;
        RECT -15.805 34.515 -15.475 34.845 ;
        RECT -15.805 33.155 -15.475 33.485 ;
        RECT -15.805 31.795 -15.475 32.125 ;
        RECT -15.805 30.435 -15.475 30.765 ;
        RECT -15.805 29.075 -15.475 29.405 ;
        RECT -15.805 27.715 -15.475 28.045 ;
        RECT -15.805 26.355 -15.475 26.685 ;
        RECT -15.805 24.995 -15.475 25.325 ;
        RECT -15.805 23.635 -15.475 23.965 ;
        RECT -15.805 22.275 -15.475 22.605 ;
        RECT -15.805 20.915 -15.475 21.245 ;
        RECT -15.805 19.555 -15.475 19.885 ;
        RECT -15.805 18.195 -15.475 18.525 ;
        RECT -15.805 16.835 -15.475 17.165 ;
        RECT -15.805 15.475 -15.475 15.805 ;
        RECT -15.805 14.115 -15.475 14.445 ;
        RECT -15.805 12.755 -15.475 13.085 ;
        RECT -15.805 11.395 -15.475 11.725 ;
        RECT -15.805 10.035 -15.475 10.365 ;
        RECT -15.805 8.675 -15.475 9.005 ;
        RECT -15.805 7.315 -15.475 7.645 ;
        RECT -15.805 5.955 -15.475 6.285 ;
        RECT -15.805 4.595 -15.475 4.925 ;
        RECT -15.805 3.235 -15.475 3.565 ;
        RECT -15.805 1.875 -15.475 2.205 ;
        RECT -15.805 0.515 -15.475 0.845 ;
        RECT -15.805 -2.205 -15.475 -1.875 ;
        RECT -15.805 -3.565 -15.475 -3.235 ;
        RECT -15.805 -4.925 -15.475 -4.595 ;
        RECT -15.805 -7.645 -15.475 -7.315 ;
        RECT -15.805 -10.365 -15.475 -10.035 ;
        RECT -15.805 -11.725 -15.475 -11.395 ;
        RECT -15.805 -13.7 -15.475 -13.37 ;
        RECT -15.805 -14.445 -15.475 -14.115 ;
        RECT -15.805 -15.805 -15.475 -15.475 ;
        RECT -15.805 -18.79 -15.475 -18.46 ;
        RECT -15.805 -19.885 -15.475 -19.555 ;
        RECT -15.805 -23.965 -15.475 -23.635 ;
        RECT -15.805 -25.325 -15.475 -24.995 ;
        RECT -15.805 -26.685 -15.475 -26.355 ;
        RECT -15.805 -29.405 -15.475 -29.075 ;
        RECT -15.805 -32.125 -15.475 -31.795 ;
        RECT -15.805 -33.485 -15.475 -33.155 ;
        RECT -15.805 -34.88 -15.475 -34.55 ;
        RECT -15.805 -36.205 -15.475 -35.875 ;
        RECT -15.805 -38.925 -15.475 -38.595 ;
        RECT -15.805 -39.97 -15.475 -39.64 ;
        RECT -15.805 -47.085 -15.475 -46.755 ;
        RECT -15.805 -48.445 -15.475 -48.115 ;
        RECT -15.805 -49.805 -15.475 -49.475 ;
        RECT -15.805 -51.165 -15.475 -50.835 ;
        RECT -15.805 -52.525 -15.475 -52.195 ;
        RECT -15.805 -53.885 -15.475 -53.555 ;
        RECT -15.805 -55.245 -15.475 -54.915 ;
        RECT -15.805 -56.605 -15.475 -56.275 ;
        RECT -15.805 -57.965 -15.475 -57.635 ;
        RECT -15.805 -59.325 -15.475 -58.995 ;
        RECT -15.805 -60.685 -15.475 -60.355 ;
        RECT -15.805 -62.045 -15.475 -61.715 ;
        RECT -15.805 -63.405 -15.475 -63.075 ;
        RECT -15.805 -68.845 -15.475 -68.515 ;
        RECT -15.805 -72.925 -15.475 -72.595 ;
        RECT -15.805 -74.285 -15.475 -73.955 ;
        RECT -15.805 -75.645 -15.475 -75.315 ;
        RECT -15.805 -77.005 -15.475 -76.675 ;
        RECT -15.805 -78.365 -15.475 -78.035 ;
        RECT -15.805 -80.31 -15.475 -79.98 ;
        RECT -15.805 -81.085 -15.475 -80.755 ;
        RECT -15.805 -82.445 -15.475 -82.115 ;
        RECT -15.805 -83.805 -15.475 -83.475 ;
        RECT -15.805 -85.165 -15.475 -84.835 ;
        RECT -15.805 -86.525 -15.475 -86.195 ;
        RECT -15.805 -87.885 -15.475 -87.555 ;
        RECT -15.805 -90.605 -15.475 -90.275 ;
        RECT -15.805 -91.965 -15.475 -91.635 ;
        RECT -15.805 -93.325 -15.475 -92.995 ;
        RECT -15.805 -94.685 -15.475 -94.355 ;
        RECT -15.805 -96.045 -15.475 -95.715 ;
        RECT -15.805 -97.405 -15.475 -97.075 ;
        RECT -15.805 -98.85 -15.475 -98.52 ;
        RECT -15.805 -100.125 -15.475 -99.795 ;
        RECT -15.805 -101.485 -15.475 -101.155 ;
        RECT -15.805 -102.845 -15.475 -102.515 ;
        RECT -15.805 -105.565 -15.475 -105.235 ;
        RECT -15.805 -106.925 -15.475 -106.595 ;
        RECT -15.805 -108.285 -15.475 -107.955 ;
        RECT -15.805 -109.645 -15.475 -109.315 ;
        RECT -15.805 -111.005 -15.475 -110.675 ;
        RECT -15.805 -112.365 -15.475 -112.035 ;
        RECT -15.805 -113.725 -15.475 -113.395 ;
        RECT -15.805 -116.445 -15.475 -116.115 ;
        RECT -15.805 -117.805 -15.475 -117.475 ;
        RECT -15.805 -119.165 -15.475 -118.835 ;
        RECT -15.805 -120.525 -15.475 -120.195 ;
        RECT -15.805 -121.885 -15.475 -121.555 ;
        RECT -15.805 -123.245 -15.475 -122.915 ;
        RECT -15.805 -124.49 -15.475 -124.16 ;
        RECT -15.805 -125.965 -15.475 -125.635 ;
        RECT -15.805 -127.325 -15.475 -126.995 ;
        RECT -15.805 -128.685 -15.475 -128.355 ;
        RECT -15.805 -130.045 -15.475 -129.715 ;
        RECT -15.805 -131.405 -15.475 -131.075 ;
        RECT -15.805 -132.765 -15.475 -132.435 ;
        RECT -15.805 -139.565 -15.475 -139.235 ;
        RECT -15.805 -140.925 -15.475 -140.595 ;
        RECT -15.805 -142.285 -15.475 -141.955 ;
        RECT -15.805 -143.03 -15.475 -142.7 ;
        RECT -15.805 -145.005 -15.475 -144.675 ;
        RECT -15.805 -146.365 -15.475 -146.035 ;
        RECT -15.805 -147.725 -15.475 -147.395 ;
        RECT -15.805 -153.165 -15.475 -152.835 ;
        RECT -15.805 -154.525 -15.475 -154.195 ;
        RECT -15.805 -155.885 -15.475 -155.555 ;
        RECT -15.805 -157.245 -15.475 -156.915 ;
        RECT -15.805 -161.325 -15.475 -160.995 ;
        RECT -15.805 -164.045 -15.475 -163.715 ;
        RECT -15.805 -168.125 -15.475 -167.795 ;
        RECT -15.805 -169.485 -15.475 -169.155 ;
        RECT -15.805 -170.845 -15.475 -170.515 ;
        RECT -15.805 -172.205 -15.475 -171.875 ;
        RECT -15.805 -174.925 -15.475 -174.595 ;
        RECT -15.805 -176.285 -15.475 -175.955 ;
        RECT -15.805 -177.645 -15.475 -177.315 ;
        RECT -15.805 -179.005 -15.475 -178.675 ;
        RECT -15.805 -180.365 -15.475 -180.035 ;
        RECT -15.805 -181.725 -15.475 -181.395 ;
        RECT -15.805 -183.085 -15.475 -182.755 ;
        RECT -15.805 -195.325 -15.475 -194.995 ;
        RECT -15.805 -198.045 -15.475 -197.715 ;
        RECT -15.805 -203.485 -15.475 -203.155 ;
        RECT -15.805 -214.365 -15.475 -214.035 ;
        RECT -15.805 -215.725 -15.475 -215.395 ;
        RECT -15.805 -217.085 -15.475 -216.755 ;
        RECT -15.805 -218.445 -15.475 -218.115 ;
        RECT -15.805 -219.805 -15.475 -219.475 ;
        RECT -15.805 -221.165 -15.475 -220.835 ;
        RECT -15.805 -222.525 -15.475 -222.195 ;
        RECT -15.805 -223.885 -15.475 -223.555 ;
        RECT -15.805 -225.245 -15.475 -224.915 ;
        RECT -15.805 -227.965 -15.475 -227.635 ;
        RECT -15.8 -229.32 -15.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -49.805 -14.115 -49.475 ;
        RECT -14.445 -51.165 -14.115 -50.835 ;
        RECT -14.445 -52.525 -14.115 -52.195 ;
        RECT -14.445 -53.885 -14.115 -53.555 ;
        RECT -14.445 -55.245 -14.115 -54.915 ;
        RECT -14.445 -56.605 -14.115 -56.275 ;
        RECT -14.445 -57.965 -14.115 -57.635 ;
        RECT -14.445 -59.325 -14.115 -58.995 ;
        RECT -14.445 -60.685 -14.115 -60.355 ;
        RECT -14.445 -62.045 -14.115 -61.715 ;
        RECT -14.445 -63.405 -14.115 -63.075 ;
        RECT -14.445 -68.845 -14.115 -68.515 ;
        RECT -14.445 -72.925 -14.115 -72.595 ;
        RECT -14.445 -74.285 -14.115 -73.955 ;
        RECT -14.445 -75.645 -14.115 -75.315 ;
        RECT -14.445 -77.005 -14.115 -76.675 ;
        RECT -14.445 -78.365 -14.115 -78.035 ;
        RECT -14.445 -80.31 -14.115 -79.98 ;
        RECT -14.445 -81.085 -14.115 -80.755 ;
        RECT -14.445 -82.445 -14.115 -82.115 ;
        RECT -14.445 -83.805 -14.115 -83.475 ;
        RECT -14.445 -85.165 -14.115 -84.835 ;
        RECT -14.445 -86.525 -14.115 -86.195 ;
        RECT -14.445 -87.885 -14.115 -87.555 ;
        RECT -14.445 -90.605 -14.115 -90.275 ;
        RECT -14.445 -91.965 -14.115 -91.635 ;
        RECT -14.445 -93.325 -14.115 -92.995 ;
        RECT -14.445 -94.685 -14.115 -94.355 ;
        RECT -14.445 -96.045 -14.115 -95.715 ;
        RECT -14.445 -97.405 -14.115 -97.075 ;
        RECT -14.445 -98.85 -14.115 -98.52 ;
        RECT -14.445 -100.125 -14.115 -99.795 ;
        RECT -14.445 -101.485 -14.115 -101.155 ;
        RECT -14.445 -102.845 -14.115 -102.515 ;
        RECT -14.445 -105.565 -14.115 -105.235 ;
        RECT -14.445 -106.925 -14.115 -106.595 ;
        RECT -14.445 -108.285 -14.115 -107.955 ;
        RECT -14.445 -109.645 -14.115 -109.315 ;
        RECT -14.445 -111.005 -14.115 -110.675 ;
        RECT -14.445 -112.365 -14.115 -112.035 ;
        RECT -14.445 -113.725 -14.115 -113.395 ;
        RECT -14.445 -116.445 -14.115 -116.115 ;
        RECT -14.445 -117.805 -14.115 -117.475 ;
        RECT -14.445 -119.165 -14.115 -118.835 ;
        RECT -14.445 -120.525 -14.115 -120.195 ;
        RECT -14.445 -121.885 -14.115 -121.555 ;
        RECT -14.445 -123.245 -14.115 -122.915 ;
        RECT -14.445 -124.49 -14.115 -124.16 ;
        RECT -14.445 -125.965 -14.115 -125.635 ;
        RECT -14.445 -127.325 -14.115 -126.995 ;
        RECT -14.445 -128.685 -14.115 -128.355 ;
        RECT -14.445 -130.045 -14.115 -129.715 ;
        RECT -14.445 -131.405 -14.115 -131.075 ;
        RECT -14.445 -132.765 -14.115 -132.435 ;
        RECT -14.445 -139.565 -14.115 -139.235 ;
        RECT -14.445 -140.925 -14.115 -140.595 ;
        RECT -14.445 -142.285 -14.115 -141.955 ;
        RECT -14.445 -143.03 -14.115 -142.7 ;
        RECT -14.445 -145.005 -14.115 -144.675 ;
        RECT -14.445 -146.365 -14.115 -146.035 ;
        RECT -14.445 -147.725 -14.115 -147.395 ;
        RECT -14.445 -153.165 -14.115 -152.835 ;
        RECT -14.445 -154.525 -14.115 -154.195 ;
        RECT -14.445 -155.885 -14.115 -155.555 ;
        RECT -14.445 -157.245 -14.115 -156.915 ;
        RECT -14.445 -159.965 -14.115 -159.635 ;
        RECT -14.445 -161.325 -14.115 -160.995 ;
        RECT -14.445 -164.045 -14.115 -163.715 ;
        RECT -14.445 -168.125 -14.115 -167.795 ;
        RECT -14.445 -169.485 -14.115 -169.155 ;
        RECT -14.445 -170.845 -14.115 -170.515 ;
        RECT -14.445 -172.205 -14.115 -171.875 ;
        RECT -14.445 -174.925 -14.115 -174.595 ;
        RECT -14.445 -176.285 -14.115 -175.955 ;
        RECT -14.445 -177.645 -14.115 -177.315 ;
        RECT -14.445 -179.005 -14.115 -178.675 ;
        RECT -14.445 -180.365 -14.115 -180.035 ;
        RECT -14.445 -181.725 -14.115 -181.395 ;
        RECT -14.445 -183.085 -14.115 -182.755 ;
        RECT -14.445 -185.805 -14.115 -185.475 ;
        RECT -14.445 -188.525 -14.115 -188.195 ;
        RECT -14.445 -189.885 -14.115 -189.555 ;
        RECT -14.445 -191.245 -14.115 -190.915 ;
        RECT -14.445 -193.965 -14.115 -193.635 ;
        RECT -14.445 -195.325 -14.115 -194.995 ;
        RECT -14.445 -196.685 -14.115 -196.355 ;
        RECT -14.445 -198.045 -14.115 -197.715 ;
        RECT -14.445 -199.405 -14.115 -199.075 ;
        RECT -14.445 -203.485 -14.115 -203.155 ;
        RECT -14.445 -204.845 -14.115 -204.515 ;
        RECT -14.445 -207.565 -14.115 -207.235 ;
        RECT -14.445 -211.645 -14.115 -211.315 ;
        RECT -14.445 -214.365 -14.115 -214.035 ;
        RECT -14.445 -215.725 -14.115 -215.395 ;
        RECT -14.445 -217.085 -14.115 -216.755 ;
        RECT -14.445 -218.445 -14.115 -218.115 ;
        RECT -14.445 -219.805 -14.115 -219.475 ;
        RECT -14.445 -221.165 -14.115 -220.835 ;
        RECT -14.445 -222.525 -14.115 -222.195 ;
        RECT -14.445 -223.885 -14.115 -223.555 ;
        RECT -14.445 -225.245 -14.115 -224.915 ;
        RECT -14.445 -227.965 -14.115 -227.635 ;
        RECT -14.445 -230.685 -14.115 -230.355 ;
        RECT -14.445 -232.045 -14.115 -231.715 ;
        RECT -14.445 -233.225 -14.115 -232.895 ;
        RECT -14.445 -234.765 -14.115 -234.435 ;
        RECT -14.445 -236.125 -14.115 -235.795 ;
        RECT -14.445 -237.485 -14.115 -237.155 ;
        RECT -14.445 -238.845 -14.115 -238.515 ;
        RECT -14.445 -241.09 -14.115 -239.96 ;
        RECT -14.44 -241.205 -14.12 245.285 ;
        RECT -14.445 244.04 -14.115 245.17 ;
        RECT -14.445 242.595 -14.115 242.925 ;
        RECT -14.445 241.235 -14.115 241.565 ;
        RECT -14.445 239.875 -14.115 240.205 ;
        RECT -14.445 238.515 -14.115 238.845 ;
        RECT -14.445 237.155 -14.115 237.485 ;
        RECT -14.445 235.795 -14.115 236.125 ;
        RECT -14.445 234.435 -14.115 234.765 ;
        RECT -14.445 233.075 -14.115 233.405 ;
        RECT -14.445 231.715 -14.115 232.045 ;
        RECT -14.445 230.355 -14.115 230.685 ;
        RECT -14.445 228.995 -14.115 229.325 ;
        RECT -14.445 227.635 -14.115 227.965 ;
        RECT -14.445 226.275 -14.115 226.605 ;
        RECT -14.445 224.915 -14.115 225.245 ;
        RECT -14.445 223.555 -14.115 223.885 ;
        RECT -14.445 222.195 -14.115 222.525 ;
        RECT -14.445 220.835 -14.115 221.165 ;
        RECT -14.445 219.475 -14.115 219.805 ;
        RECT -14.445 218.115 -14.115 218.445 ;
        RECT -14.445 216.755 -14.115 217.085 ;
        RECT -14.445 215.395 -14.115 215.725 ;
        RECT -14.445 214.035 -14.115 214.365 ;
        RECT -14.445 212.675 -14.115 213.005 ;
        RECT -14.445 211.315 -14.115 211.645 ;
        RECT -14.445 209.955 -14.115 210.285 ;
        RECT -14.445 208.595 -14.115 208.925 ;
        RECT -14.445 207.235 -14.115 207.565 ;
        RECT -14.445 205.875 -14.115 206.205 ;
        RECT -14.445 204.515 -14.115 204.845 ;
        RECT -14.445 203.155 -14.115 203.485 ;
        RECT -14.445 201.795 -14.115 202.125 ;
        RECT -14.445 200.435 -14.115 200.765 ;
        RECT -14.445 199.075 -14.115 199.405 ;
        RECT -14.445 197.715 -14.115 198.045 ;
        RECT -14.445 196.355 -14.115 196.685 ;
        RECT -14.445 194.995 -14.115 195.325 ;
        RECT -14.445 193.635 -14.115 193.965 ;
        RECT -14.445 192.275 -14.115 192.605 ;
        RECT -14.445 190.915 -14.115 191.245 ;
        RECT -14.445 189.555 -14.115 189.885 ;
        RECT -14.445 188.195 -14.115 188.525 ;
        RECT -14.445 186.835 -14.115 187.165 ;
        RECT -14.445 185.475 -14.115 185.805 ;
        RECT -14.445 184.115 -14.115 184.445 ;
        RECT -14.445 182.755 -14.115 183.085 ;
        RECT -14.445 181.395 -14.115 181.725 ;
        RECT -14.445 180.035 -14.115 180.365 ;
        RECT -14.445 178.675 -14.115 179.005 ;
        RECT -14.445 177.315 -14.115 177.645 ;
        RECT -14.445 175.955 -14.115 176.285 ;
        RECT -14.445 174.595 -14.115 174.925 ;
        RECT -14.445 173.235 -14.115 173.565 ;
        RECT -14.445 171.875 -14.115 172.205 ;
        RECT -14.445 170.515 -14.115 170.845 ;
        RECT -14.445 169.155 -14.115 169.485 ;
        RECT -14.445 167.795 -14.115 168.125 ;
        RECT -14.445 166.435 -14.115 166.765 ;
        RECT -14.445 165.075 -14.115 165.405 ;
        RECT -14.445 163.715 -14.115 164.045 ;
        RECT -14.445 162.355 -14.115 162.685 ;
        RECT -14.445 160.995 -14.115 161.325 ;
        RECT -14.445 159.635 -14.115 159.965 ;
        RECT -14.445 158.275 -14.115 158.605 ;
        RECT -14.445 156.915 -14.115 157.245 ;
        RECT -14.445 155.555 -14.115 155.885 ;
        RECT -14.445 154.195 -14.115 154.525 ;
        RECT -14.445 152.835 -14.115 153.165 ;
        RECT -14.445 151.475 -14.115 151.805 ;
        RECT -14.445 150.115 -14.115 150.445 ;
        RECT -14.445 148.755 -14.115 149.085 ;
        RECT -14.445 147.395 -14.115 147.725 ;
        RECT -14.445 146.035 -14.115 146.365 ;
        RECT -14.445 144.675 -14.115 145.005 ;
        RECT -14.445 143.315 -14.115 143.645 ;
        RECT -14.445 141.955 -14.115 142.285 ;
        RECT -14.445 140.595 -14.115 140.925 ;
        RECT -14.445 139.235 -14.115 139.565 ;
        RECT -14.445 137.875 -14.115 138.205 ;
        RECT -14.445 136.515 -14.115 136.845 ;
        RECT -14.445 135.155 -14.115 135.485 ;
        RECT -14.445 133.795 -14.115 134.125 ;
        RECT -14.445 132.435 -14.115 132.765 ;
        RECT -14.445 131.075 -14.115 131.405 ;
        RECT -14.445 129.715 -14.115 130.045 ;
        RECT -14.445 128.355 -14.115 128.685 ;
        RECT -14.445 126.995 -14.115 127.325 ;
        RECT -14.445 125.635 -14.115 125.965 ;
        RECT -14.445 124.275 -14.115 124.605 ;
        RECT -14.445 122.915 -14.115 123.245 ;
        RECT -14.445 121.555 -14.115 121.885 ;
        RECT -14.445 120.195 -14.115 120.525 ;
        RECT -14.445 118.835 -14.115 119.165 ;
        RECT -14.445 117.475 -14.115 117.805 ;
        RECT -14.445 116.115 -14.115 116.445 ;
        RECT -14.445 114.755 -14.115 115.085 ;
        RECT -14.445 113.395 -14.115 113.725 ;
        RECT -14.445 112.035 -14.115 112.365 ;
        RECT -14.445 110.675 -14.115 111.005 ;
        RECT -14.445 109.315 -14.115 109.645 ;
        RECT -14.445 107.955 -14.115 108.285 ;
        RECT -14.445 106.595 -14.115 106.925 ;
        RECT -14.445 105.235 -14.115 105.565 ;
        RECT -14.445 103.875 -14.115 104.205 ;
        RECT -14.445 102.515 -14.115 102.845 ;
        RECT -14.445 101.155 -14.115 101.485 ;
        RECT -14.445 99.795 -14.115 100.125 ;
        RECT -14.445 98.435 -14.115 98.765 ;
        RECT -14.445 97.075 -14.115 97.405 ;
        RECT -14.445 95.715 -14.115 96.045 ;
        RECT -14.445 94.355 -14.115 94.685 ;
        RECT -14.445 92.995 -14.115 93.325 ;
        RECT -14.445 91.635 -14.115 91.965 ;
        RECT -14.445 90.275 -14.115 90.605 ;
        RECT -14.445 88.915 -14.115 89.245 ;
        RECT -14.445 87.555 -14.115 87.885 ;
        RECT -14.445 86.195 -14.115 86.525 ;
        RECT -14.445 84.835 -14.115 85.165 ;
        RECT -14.445 83.475 -14.115 83.805 ;
        RECT -14.445 82.115 -14.115 82.445 ;
        RECT -14.445 80.755 -14.115 81.085 ;
        RECT -14.445 79.395 -14.115 79.725 ;
        RECT -14.445 78.035 -14.115 78.365 ;
        RECT -14.445 76.675 -14.115 77.005 ;
        RECT -14.445 75.315 -14.115 75.645 ;
        RECT -14.445 73.955 -14.115 74.285 ;
        RECT -14.445 72.595 -14.115 72.925 ;
        RECT -14.445 71.235 -14.115 71.565 ;
        RECT -14.445 69.875 -14.115 70.205 ;
        RECT -14.445 68.515 -14.115 68.845 ;
        RECT -14.445 67.155 -14.115 67.485 ;
        RECT -14.445 65.795 -14.115 66.125 ;
        RECT -14.445 64.435 -14.115 64.765 ;
        RECT -14.445 63.075 -14.115 63.405 ;
        RECT -14.445 61.715 -14.115 62.045 ;
        RECT -14.445 60.355 -14.115 60.685 ;
        RECT -14.445 58.995 -14.115 59.325 ;
        RECT -14.445 57.635 -14.115 57.965 ;
        RECT -14.445 56.275 -14.115 56.605 ;
        RECT -14.445 54.915 -14.115 55.245 ;
        RECT -14.445 53.555 -14.115 53.885 ;
        RECT -14.445 52.195 -14.115 52.525 ;
        RECT -14.445 50.835 -14.115 51.165 ;
        RECT -14.445 49.475 -14.115 49.805 ;
        RECT -14.445 48.115 -14.115 48.445 ;
        RECT -14.445 46.755 -14.115 47.085 ;
        RECT -14.445 45.395 -14.115 45.725 ;
        RECT -14.445 44.035 -14.115 44.365 ;
        RECT -14.445 42.675 -14.115 43.005 ;
        RECT -14.445 41.315 -14.115 41.645 ;
        RECT -14.445 39.955 -14.115 40.285 ;
        RECT -14.445 38.595 -14.115 38.925 ;
        RECT -14.445 37.235 -14.115 37.565 ;
        RECT -14.445 35.875 -14.115 36.205 ;
        RECT -14.445 34.515 -14.115 34.845 ;
        RECT -14.445 33.155 -14.115 33.485 ;
        RECT -14.445 31.795 -14.115 32.125 ;
        RECT -14.445 30.435 -14.115 30.765 ;
        RECT -14.445 29.075 -14.115 29.405 ;
        RECT -14.445 27.715 -14.115 28.045 ;
        RECT -14.445 26.355 -14.115 26.685 ;
        RECT -14.445 24.995 -14.115 25.325 ;
        RECT -14.445 23.635 -14.115 23.965 ;
        RECT -14.445 22.275 -14.115 22.605 ;
        RECT -14.445 20.915 -14.115 21.245 ;
        RECT -14.445 19.555 -14.115 19.885 ;
        RECT -14.445 18.195 -14.115 18.525 ;
        RECT -14.445 16.835 -14.115 17.165 ;
        RECT -14.445 15.475 -14.115 15.805 ;
        RECT -14.445 14.115 -14.115 14.445 ;
        RECT -14.445 12.755 -14.115 13.085 ;
        RECT -14.445 11.395 -14.115 11.725 ;
        RECT -14.445 10.035 -14.115 10.365 ;
        RECT -14.445 8.675 -14.115 9.005 ;
        RECT -14.445 7.315 -14.115 7.645 ;
        RECT -14.445 5.955 -14.115 6.285 ;
        RECT -14.445 4.595 -14.115 4.925 ;
        RECT -14.445 3.235 -14.115 3.565 ;
        RECT -14.445 1.875 -14.115 2.205 ;
        RECT -14.445 0.515 -14.115 0.845 ;
        RECT -14.445 -2.205 -14.115 -1.875 ;
        RECT -14.445 -3.565 -14.115 -3.235 ;
        RECT -14.445 -4.925 -14.115 -4.595 ;
        RECT -14.445 -7.645 -14.115 -7.315 ;
        RECT -14.445 -10.365 -14.115 -10.035 ;
        RECT -14.445 -11.725 -14.115 -11.395 ;
        RECT -14.445 -13.7 -14.115 -13.37 ;
        RECT -14.445 -14.445 -14.115 -14.115 ;
        RECT -14.445 -15.805 -14.115 -15.475 ;
        RECT -14.445 -18.79 -14.115 -18.46 ;
        RECT -14.445 -19.885 -14.115 -19.555 ;
        RECT -14.445 -23.965 -14.115 -23.635 ;
        RECT -14.445 -25.325 -14.115 -24.995 ;
        RECT -14.445 -26.685 -14.115 -26.355 ;
        RECT -14.445 -29.405 -14.115 -29.075 ;
        RECT -14.445 -32.125 -14.115 -31.795 ;
        RECT -14.445 -33.485 -14.115 -33.155 ;
        RECT -14.445 -34.88 -14.115 -34.55 ;
        RECT -14.445 -36.205 -14.115 -35.875 ;
        RECT -14.445 -38.925 -14.115 -38.595 ;
        RECT -14.445 -39.97 -14.115 -39.64 ;
        RECT -14.445 -47.085 -14.115 -46.755 ;
        RECT -14.445 -48.445 -14.115 -48.115 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.965 244.04 -23.635 245.17 ;
        RECT -23.965 242.595 -23.635 242.925 ;
        RECT -23.965 241.235 -23.635 241.565 ;
        RECT -23.965 239.875 -23.635 240.205 ;
        RECT -23.965 238.515 -23.635 238.845 ;
        RECT -23.965 237.155 -23.635 237.485 ;
        RECT -23.965 235.795 -23.635 236.125 ;
        RECT -23.965 234.435 -23.635 234.765 ;
        RECT -23.965 233.075 -23.635 233.405 ;
        RECT -23.965 231.715 -23.635 232.045 ;
        RECT -23.965 230.355 -23.635 230.685 ;
        RECT -23.965 228.995 -23.635 229.325 ;
        RECT -23.965 227.635 -23.635 227.965 ;
        RECT -23.965 226.275 -23.635 226.605 ;
        RECT -23.965 224.915 -23.635 225.245 ;
        RECT -23.965 223.555 -23.635 223.885 ;
        RECT -23.965 222.195 -23.635 222.525 ;
        RECT -23.965 220.835 -23.635 221.165 ;
        RECT -23.965 219.475 -23.635 219.805 ;
        RECT -23.965 218.115 -23.635 218.445 ;
        RECT -23.965 216.755 -23.635 217.085 ;
        RECT -23.965 215.395 -23.635 215.725 ;
        RECT -23.965 214.035 -23.635 214.365 ;
        RECT -23.965 212.675 -23.635 213.005 ;
        RECT -23.965 211.315 -23.635 211.645 ;
        RECT -23.965 209.955 -23.635 210.285 ;
        RECT -23.965 208.595 -23.635 208.925 ;
        RECT -23.965 207.235 -23.635 207.565 ;
        RECT -23.965 205.875 -23.635 206.205 ;
        RECT -23.965 204.515 -23.635 204.845 ;
        RECT -23.965 203.155 -23.635 203.485 ;
        RECT -23.965 201.795 -23.635 202.125 ;
        RECT -23.965 200.435 -23.635 200.765 ;
        RECT -23.965 199.075 -23.635 199.405 ;
        RECT -23.965 197.715 -23.635 198.045 ;
        RECT -23.965 196.355 -23.635 196.685 ;
        RECT -23.965 194.995 -23.635 195.325 ;
        RECT -23.965 193.635 -23.635 193.965 ;
        RECT -23.965 192.275 -23.635 192.605 ;
        RECT -23.965 190.915 -23.635 191.245 ;
        RECT -23.965 189.555 -23.635 189.885 ;
        RECT -23.965 188.195 -23.635 188.525 ;
        RECT -23.965 186.835 -23.635 187.165 ;
        RECT -23.965 185.475 -23.635 185.805 ;
        RECT -23.965 184.115 -23.635 184.445 ;
        RECT -23.965 182.755 -23.635 183.085 ;
        RECT -23.965 181.395 -23.635 181.725 ;
        RECT -23.965 180.035 -23.635 180.365 ;
        RECT -23.965 178.675 -23.635 179.005 ;
        RECT -23.965 177.315 -23.635 177.645 ;
        RECT -23.965 175.955 -23.635 176.285 ;
        RECT -23.965 174.595 -23.635 174.925 ;
        RECT -23.965 173.235 -23.635 173.565 ;
        RECT -23.965 171.875 -23.635 172.205 ;
        RECT -23.965 170.515 -23.635 170.845 ;
        RECT -23.965 169.155 -23.635 169.485 ;
        RECT -23.965 167.795 -23.635 168.125 ;
        RECT -23.965 166.435 -23.635 166.765 ;
        RECT -23.965 165.075 -23.635 165.405 ;
        RECT -23.965 163.715 -23.635 164.045 ;
        RECT -23.965 162.355 -23.635 162.685 ;
        RECT -23.965 160.995 -23.635 161.325 ;
        RECT -23.965 159.635 -23.635 159.965 ;
        RECT -23.965 158.275 -23.635 158.605 ;
        RECT -23.965 156.915 -23.635 157.245 ;
        RECT -23.965 155.555 -23.635 155.885 ;
        RECT -23.965 154.195 -23.635 154.525 ;
        RECT -23.965 152.835 -23.635 153.165 ;
        RECT -23.965 151.475 -23.635 151.805 ;
        RECT -23.965 150.115 -23.635 150.445 ;
        RECT -23.965 148.755 -23.635 149.085 ;
        RECT -23.965 147.395 -23.635 147.725 ;
        RECT -23.965 146.035 -23.635 146.365 ;
        RECT -23.965 144.675 -23.635 145.005 ;
        RECT -23.965 143.315 -23.635 143.645 ;
        RECT -23.965 141.955 -23.635 142.285 ;
        RECT -23.965 140.595 -23.635 140.925 ;
        RECT -23.965 139.235 -23.635 139.565 ;
        RECT -23.965 137.875 -23.635 138.205 ;
        RECT -23.965 136.515 -23.635 136.845 ;
        RECT -23.965 135.155 -23.635 135.485 ;
        RECT -23.965 133.795 -23.635 134.125 ;
        RECT -23.965 132.435 -23.635 132.765 ;
        RECT -23.965 131.075 -23.635 131.405 ;
        RECT -23.965 129.715 -23.635 130.045 ;
        RECT -23.965 128.355 -23.635 128.685 ;
        RECT -23.965 126.995 -23.635 127.325 ;
        RECT -23.965 125.635 -23.635 125.965 ;
        RECT -23.965 124.275 -23.635 124.605 ;
        RECT -23.965 122.915 -23.635 123.245 ;
        RECT -23.965 121.555 -23.635 121.885 ;
        RECT -23.965 120.195 -23.635 120.525 ;
        RECT -23.965 118.835 -23.635 119.165 ;
        RECT -23.965 117.475 -23.635 117.805 ;
        RECT -23.965 116.115 -23.635 116.445 ;
        RECT -23.965 114.755 -23.635 115.085 ;
        RECT -23.965 113.395 -23.635 113.725 ;
        RECT -23.965 112.035 -23.635 112.365 ;
        RECT -23.965 110.675 -23.635 111.005 ;
        RECT -23.965 109.315 -23.635 109.645 ;
        RECT -23.965 107.955 -23.635 108.285 ;
        RECT -23.965 106.595 -23.635 106.925 ;
        RECT -23.965 105.235 -23.635 105.565 ;
        RECT -23.965 103.875 -23.635 104.205 ;
        RECT -23.965 102.515 -23.635 102.845 ;
        RECT -23.965 101.155 -23.635 101.485 ;
        RECT -23.965 99.795 -23.635 100.125 ;
        RECT -23.965 98.435 -23.635 98.765 ;
        RECT -23.965 97.075 -23.635 97.405 ;
        RECT -23.965 95.715 -23.635 96.045 ;
        RECT -23.965 94.355 -23.635 94.685 ;
        RECT -23.965 92.995 -23.635 93.325 ;
        RECT -23.965 91.635 -23.635 91.965 ;
        RECT -23.965 90.275 -23.635 90.605 ;
        RECT -23.965 88.915 -23.635 89.245 ;
        RECT -23.965 87.555 -23.635 87.885 ;
        RECT -23.965 86.195 -23.635 86.525 ;
        RECT -23.965 84.835 -23.635 85.165 ;
        RECT -23.965 83.475 -23.635 83.805 ;
        RECT -23.965 82.115 -23.635 82.445 ;
        RECT -23.965 80.755 -23.635 81.085 ;
        RECT -23.965 79.395 -23.635 79.725 ;
        RECT -23.965 78.035 -23.635 78.365 ;
        RECT -23.965 76.675 -23.635 77.005 ;
        RECT -23.965 75.315 -23.635 75.645 ;
        RECT -23.965 73.955 -23.635 74.285 ;
        RECT -23.965 72.595 -23.635 72.925 ;
        RECT -23.965 71.235 -23.635 71.565 ;
        RECT -23.965 69.875 -23.635 70.205 ;
        RECT -23.965 68.515 -23.635 68.845 ;
        RECT -23.965 67.155 -23.635 67.485 ;
        RECT -23.965 65.795 -23.635 66.125 ;
        RECT -23.965 64.435 -23.635 64.765 ;
        RECT -23.965 63.075 -23.635 63.405 ;
        RECT -23.965 61.715 -23.635 62.045 ;
        RECT -23.965 60.355 -23.635 60.685 ;
        RECT -23.965 58.995 -23.635 59.325 ;
        RECT -23.965 57.635 -23.635 57.965 ;
        RECT -23.965 56.275 -23.635 56.605 ;
        RECT -23.965 54.915 -23.635 55.245 ;
        RECT -23.965 53.555 -23.635 53.885 ;
        RECT -23.965 52.195 -23.635 52.525 ;
        RECT -23.965 50.835 -23.635 51.165 ;
        RECT -23.965 49.475 -23.635 49.805 ;
        RECT -23.965 48.115 -23.635 48.445 ;
        RECT -23.965 46.755 -23.635 47.085 ;
        RECT -23.965 45.395 -23.635 45.725 ;
        RECT -23.965 44.035 -23.635 44.365 ;
        RECT -23.965 42.675 -23.635 43.005 ;
        RECT -23.965 41.315 -23.635 41.645 ;
        RECT -23.965 39.955 -23.635 40.285 ;
        RECT -23.965 38.595 -23.635 38.925 ;
        RECT -23.965 37.235 -23.635 37.565 ;
        RECT -23.965 35.875 -23.635 36.205 ;
        RECT -23.965 34.515 -23.635 34.845 ;
        RECT -23.965 33.155 -23.635 33.485 ;
        RECT -23.965 31.795 -23.635 32.125 ;
        RECT -23.965 30.435 -23.635 30.765 ;
        RECT -23.965 29.075 -23.635 29.405 ;
        RECT -23.965 27.715 -23.635 28.045 ;
        RECT -23.965 26.355 -23.635 26.685 ;
        RECT -23.965 24.995 -23.635 25.325 ;
        RECT -23.965 23.635 -23.635 23.965 ;
        RECT -23.965 22.275 -23.635 22.605 ;
        RECT -23.965 20.915 -23.635 21.245 ;
        RECT -23.965 19.555 -23.635 19.885 ;
        RECT -23.965 18.195 -23.635 18.525 ;
        RECT -23.965 16.835 -23.635 17.165 ;
        RECT -23.965 15.475 -23.635 15.805 ;
        RECT -23.965 14.115 -23.635 14.445 ;
        RECT -23.965 12.755 -23.635 13.085 ;
        RECT -23.965 11.395 -23.635 11.725 ;
        RECT -23.965 10.035 -23.635 10.365 ;
        RECT -23.965 8.675 -23.635 9.005 ;
        RECT -23.965 7.315 -23.635 7.645 ;
        RECT -23.965 5.955 -23.635 6.285 ;
        RECT -23.965 4.595 -23.635 4.925 ;
        RECT -23.965 3.235 -23.635 3.565 ;
        RECT -23.965 1.875 -23.635 2.205 ;
        RECT -23.965 0.515 -23.635 0.845 ;
        RECT -23.965 -2.205 -23.635 -1.875 ;
        RECT -23.965 -7.645 -23.635 -7.315 ;
        RECT -23.965 -10.365 -23.635 -10.035 ;
        RECT -23.965 -11.725 -23.635 -11.395 ;
        RECT -23.965 -13.7 -23.635 -13.37 ;
        RECT -23.965 -14.445 -23.635 -14.115 ;
        RECT -23.965 -15.805 -23.635 -15.475 ;
        RECT -23.965 -18.79 -23.635 -18.46 ;
        RECT -23.965 -19.885 -23.635 -19.555 ;
        RECT -23.965 -23.965 -23.635 -23.635 ;
        RECT -23.965 -29.405 -23.635 -29.075 ;
        RECT -23.965 -32.125 -23.635 -31.795 ;
        RECT -23.965 -33.485 -23.635 -33.155 ;
        RECT -23.965 -34.88 -23.635 -34.55 ;
        RECT -23.965 -36.205 -23.635 -35.875 ;
        RECT -23.965 -38.925 -23.635 -38.595 ;
        RECT -23.965 -39.97 -23.635 -39.64 ;
        RECT -23.965 -47.085 -23.635 -46.755 ;
        RECT -23.965 -48.445 -23.635 -48.115 ;
        RECT -23.965 -49.805 -23.635 -49.475 ;
        RECT -23.965 -51.165 -23.635 -50.835 ;
        RECT -23.965 -52.525 -23.635 -52.195 ;
        RECT -23.965 -53.885 -23.635 -53.555 ;
        RECT -23.965 -55.245 -23.635 -54.915 ;
        RECT -23.965 -56.605 -23.635 -56.275 ;
        RECT -23.965 -57.965 -23.635 -57.635 ;
        RECT -23.965 -59.325 -23.635 -58.995 ;
        RECT -23.965 -60.685 -23.635 -60.355 ;
        RECT -23.965 -62.045 -23.635 -61.715 ;
        RECT -23.965 -63.405 -23.635 -63.075 ;
        RECT -23.965 -64.765 -23.635 -64.435 ;
        RECT -23.965 -66.125 -23.635 -65.795 ;
        RECT -23.965 -68.845 -23.635 -68.515 ;
        RECT -23.965 -71.565 -23.635 -71.235 ;
        RECT -23.965 -72.925 -23.635 -72.595 ;
        RECT -23.965 -74.285 -23.635 -73.955 ;
        RECT -23.965 -75.645 -23.635 -75.315 ;
        RECT -23.965 -77.005 -23.635 -76.675 ;
        RECT -23.965 -78.365 -23.635 -78.035 ;
        RECT -23.965 -80.31 -23.635 -79.98 ;
        RECT -23.965 -81.085 -23.635 -80.755 ;
        RECT -23.965 -82.445 -23.635 -82.115 ;
        RECT -23.965 -83.805 -23.635 -83.475 ;
        RECT -23.965 -85.165 -23.635 -84.835 ;
        RECT -23.965 -86.525 -23.635 -86.195 ;
        RECT -23.965 -87.885 -23.635 -87.555 ;
        RECT -23.965 -90.605 -23.635 -90.275 ;
        RECT -23.965 -91.965 -23.635 -91.635 ;
        RECT -23.965 -93.325 -23.635 -92.995 ;
        RECT -23.965 -94.685 -23.635 -94.355 ;
        RECT -23.965 -96.045 -23.635 -95.715 ;
        RECT -23.965 -97.405 -23.635 -97.075 ;
        RECT -23.965 -98.85 -23.635 -98.52 ;
        RECT -23.965 -100.125 -23.635 -99.795 ;
        RECT -23.965 -101.485 -23.635 -101.155 ;
        RECT -23.965 -102.845 -23.635 -102.515 ;
        RECT -23.965 -105.565 -23.635 -105.235 ;
        RECT -23.965 -106.925 -23.635 -106.595 ;
        RECT -23.965 -108.285 -23.635 -107.955 ;
        RECT -23.965 -109.645 -23.635 -109.315 ;
        RECT -23.965 -111.005 -23.635 -110.675 ;
        RECT -23.965 -112.365 -23.635 -112.035 ;
        RECT -23.965 -113.725 -23.635 -113.395 ;
        RECT -23.965 -116.445 -23.635 -116.115 ;
        RECT -23.965 -117.805 -23.635 -117.475 ;
        RECT -23.965 -119.165 -23.635 -118.835 ;
        RECT -23.965 -120.525 -23.635 -120.195 ;
        RECT -23.965 -121.885 -23.635 -121.555 ;
        RECT -23.965 -124.49 -23.635 -124.16 ;
        RECT -23.965 -128.685 -23.635 -128.355 ;
        RECT -23.965 -130.045 -23.635 -129.715 ;
        RECT -23.965 -131.405 -23.635 -131.075 ;
        RECT -23.965 -132.765 -23.635 -132.435 ;
        RECT -23.965 -136.845 -23.635 -136.515 ;
        RECT -23.965 -138.205 -23.635 -137.875 ;
        RECT -23.965 -139.565 -23.635 -139.235 ;
        RECT -23.965 -140.925 -23.635 -140.595 ;
        RECT -23.965 -142.285 -23.635 -141.955 ;
        RECT -23.965 -143.03 -23.635 -142.7 ;
        RECT -23.965 -145.005 -23.635 -144.675 ;
        RECT -23.965 -146.365 -23.635 -146.035 ;
        RECT -23.965 -147.725 -23.635 -147.395 ;
        RECT -23.965 -153.165 -23.635 -152.835 ;
        RECT -23.965 -154.525 -23.635 -154.195 ;
        RECT -23.965 -155.885 -23.635 -155.555 ;
        RECT -23.965 -157.245 -23.635 -156.915 ;
        RECT -23.965 -162.685 -23.635 -162.355 ;
        RECT -23.965 -164.045 -23.635 -163.715 ;
        RECT -23.965 -165.405 -23.635 -165.075 ;
        RECT -23.965 -166.765 -23.635 -166.435 ;
        RECT -23.965 -168.125 -23.635 -167.795 ;
        RECT -23.965 -169.485 -23.635 -169.155 ;
        RECT -23.965 -170.845 -23.635 -170.515 ;
        RECT -23.965 -172.205 -23.635 -171.875 ;
        RECT -23.965 -174.925 -23.635 -174.595 ;
        RECT -23.965 -176.285 -23.635 -175.955 ;
        RECT -23.965 -177.645 -23.635 -177.315 ;
        RECT -23.965 -179.005 -23.635 -178.675 ;
        RECT -23.965 -180.365 -23.635 -180.035 ;
        RECT -23.965 -181.725 -23.635 -181.395 ;
        RECT -23.965 -183.085 -23.635 -182.755 ;
        RECT -23.965 -192.605 -23.635 -192.275 ;
        RECT -23.965 -193.965 -23.635 -193.635 ;
        RECT -23.965 -195.325 -23.635 -194.995 ;
        RECT -23.965 -198.045 -23.635 -197.715 ;
        RECT -23.965 -199.405 -23.635 -199.075 ;
        RECT -23.965 -200.765 -23.635 -200.435 ;
        RECT -23.965 -204.845 -23.635 -204.515 ;
        RECT -23.965 -206.205 -23.635 -205.875 ;
        RECT -23.965 -208.925 -23.635 -208.595 ;
        RECT -23.965 -210.285 -23.635 -209.955 ;
        RECT -23.965 -215.725 -23.635 -215.395 ;
        RECT -23.965 -217.085 -23.635 -216.755 ;
        RECT -23.965 -218.445 -23.635 -218.115 ;
        RECT -23.965 -219.805 -23.635 -219.475 ;
        RECT -23.965 -221.165 -23.635 -220.835 ;
        RECT -23.965 -222.525 -23.635 -222.195 ;
        RECT -23.965 -223.885 -23.635 -223.555 ;
        RECT -23.965 -225.245 -23.635 -224.915 ;
        RECT -23.965 -232.045 -23.635 -231.715 ;
        RECT -23.965 -233.225 -23.635 -232.895 ;
        RECT -23.965 -234.765 -23.635 -234.435 ;
        RECT -23.965 -236.125 -23.635 -235.795 ;
        RECT -23.965 -237.485 -23.635 -237.155 ;
        RECT -23.965 -238.845 -23.635 -238.515 ;
        RECT -23.965 -241.09 -23.635 -239.96 ;
        RECT -23.96 -241.205 -23.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.605 244.04 -22.275 245.17 ;
        RECT -22.605 242.595 -22.275 242.925 ;
        RECT -22.605 241.235 -22.275 241.565 ;
        RECT -22.605 239.875 -22.275 240.205 ;
        RECT -22.605 238.515 -22.275 238.845 ;
        RECT -22.605 237.155 -22.275 237.485 ;
        RECT -22.605 235.795 -22.275 236.125 ;
        RECT -22.605 234.435 -22.275 234.765 ;
        RECT -22.605 233.075 -22.275 233.405 ;
        RECT -22.605 231.715 -22.275 232.045 ;
        RECT -22.605 230.355 -22.275 230.685 ;
        RECT -22.605 228.995 -22.275 229.325 ;
        RECT -22.605 227.635 -22.275 227.965 ;
        RECT -22.605 226.275 -22.275 226.605 ;
        RECT -22.605 224.915 -22.275 225.245 ;
        RECT -22.605 223.555 -22.275 223.885 ;
        RECT -22.605 222.195 -22.275 222.525 ;
        RECT -22.605 220.835 -22.275 221.165 ;
        RECT -22.605 219.475 -22.275 219.805 ;
        RECT -22.605 218.115 -22.275 218.445 ;
        RECT -22.605 216.755 -22.275 217.085 ;
        RECT -22.605 215.395 -22.275 215.725 ;
        RECT -22.605 214.035 -22.275 214.365 ;
        RECT -22.605 212.675 -22.275 213.005 ;
        RECT -22.605 211.315 -22.275 211.645 ;
        RECT -22.605 209.955 -22.275 210.285 ;
        RECT -22.605 208.595 -22.275 208.925 ;
        RECT -22.605 207.235 -22.275 207.565 ;
        RECT -22.605 205.875 -22.275 206.205 ;
        RECT -22.605 204.515 -22.275 204.845 ;
        RECT -22.605 203.155 -22.275 203.485 ;
        RECT -22.605 201.795 -22.275 202.125 ;
        RECT -22.605 200.435 -22.275 200.765 ;
        RECT -22.605 199.075 -22.275 199.405 ;
        RECT -22.605 197.715 -22.275 198.045 ;
        RECT -22.605 196.355 -22.275 196.685 ;
        RECT -22.605 194.995 -22.275 195.325 ;
        RECT -22.605 193.635 -22.275 193.965 ;
        RECT -22.605 192.275 -22.275 192.605 ;
        RECT -22.605 190.915 -22.275 191.245 ;
        RECT -22.605 189.555 -22.275 189.885 ;
        RECT -22.605 188.195 -22.275 188.525 ;
        RECT -22.605 186.835 -22.275 187.165 ;
        RECT -22.605 185.475 -22.275 185.805 ;
        RECT -22.605 184.115 -22.275 184.445 ;
        RECT -22.605 182.755 -22.275 183.085 ;
        RECT -22.605 181.395 -22.275 181.725 ;
        RECT -22.605 180.035 -22.275 180.365 ;
        RECT -22.605 178.675 -22.275 179.005 ;
        RECT -22.605 177.315 -22.275 177.645 ;
        RECT -22.605 175.955 -22.275 176.285 ;
        RECT -22.605 174.595 -22.275 174.925 ;
        RECT -22.605 173.235 -22.275 173.565 ;
        RECT -22.605 171.875 -22.275 172.205 ;
        RECT -22.605 170.515 -22.275 170.845 ;
        RECT -22.605 169.155 -22.275 169.485 ;
        RECT -22.605 167.795 -22.275 168.125 ;
        RECT -22.605 166.435 -22.275 166.765 ;
        RECT -22.605 165.075 -22.275 165.405 ;
        RECT -22.605 163.715 -22.275 164.045 ;
        RECT -22.605 162.355 -22.275 162.685 ;
        RECT -22.605 160.995 -22.275 161.325 ;
        RECT -22.605 159.635 -22.275 159.965 ;
        RECT -22.605 158.275 -22.275 158.605 ;
        RECT -22.605 156.915 -22.275 157.245 ;
        RECT -22.605 155.555 -22.275 155.885 ;
        RECT -22.605 154.195 -22.275 154.525 ;
        RECT -22.605 152.835 -22.275 153.165 ;
        RECT -22.605 151.475 -22.275 151.805 ;
        RECT -22.605 150.115 -22.275 150.445 ;
        RECT -22.605 148.755 -22.275 149.085 ;
        RECT -22.605 147.395 -22.275 147.725 ;
        RECT -22.605 146.035 -22.275 146.365 ;
        RECT -22.605 144.675 -22.275 145.005 ;
        RECT -22.605 143.315 -22.275 143.645 ;
        RECT -22.605 141.955 -22.275 142.285 ;
        RECT -22.605 140.595 -22.275 140.925 ;
        RECT -22.605 139.235 -22.275 139.565 ;
        RECT -22.605 137.875 -22.275 138.205 ;
        RECT -22.605 136.515 -22.275 136.845 ;
        RECT -22.605 135.155 -22.275 135.485 ;
        RECT -22.605 133.795 -22.275 134.125 ;
        RECT -22.605 132.435 -22.275 132.765 ;
        RECT -22.605 131.075 -22.275 131.405 ;
        RECT -22.605 129.715 -22.275 130.045 ;
        RECT -22.605 128.355 -22.275 128.685 ;
        RECT -22.605 126.995 -22.275 127.325 ;
        RECT -22.605 125.635 -22.275 125.965 ;
        RECT -22.605 124.275 -22.275 124.605 ;
        RECT -22.605 122.915 -22.275 123.245 ;
        RECT -22.605 121.555 -22.275 121.885 ;
        RECT -22.605 120.195 -22.275 120.525 ;
        RECT -22.605 118.835 -22.275 119.165 ;
        RECT -22.605 117.475 -22.275 117.805 ;
        RECT -22.605 116.115 -22.275 116.445 ;
        RECT -22.605 114.755 -22.275 115.085 ;
        RECT -22.605 113.395 -22.275 113.725 ;
        RECT -22.605 112.035 -22.275 112.365 ;
        RECT -22.605 110.675 -22.275 111.005 ;
        RECT -22.605 109.315 -22.275 109.645 ;
        RECT -22.605 107.955 -22.275 108.285 ;
        RECT -22.605 106.595 -22.275 106.925 ;
        RECT -22.605 105.235 -22.275 105.565 ;
        RECT -22.605 103.875 -22.275 104.205 ;
        RECT -22.605 102.515 -22.275 102.845 ;
        RECT -22.605 101.155 -22.275 101.485 ;
        RECT -22.605 99.795 -22.275 100.125 ;
        RECT -22.605 98.435 -22.275 98.765 ;
        RECT -22.605 97.075 -22.275 97.405 ;
        RECT -22.605 95.715 -22.275 96.045 ;
        RECT -22.605 94.355 -22.275 94.685 ;
        RECT -22.605 92.995 -22.275 93.325 ;
        RECT -22.605 91.635 -22.275 91.965 ;
        RECT -22.605 90.275 -22.275 90.605 ;
        RECT -22.605 88.915 -22.275 89.245 ;
        RECT -22.605 87.555 -22.275 87.885 ;
        RECT -22.605 86.195 -22.275 86.525 ;
        RECT -22.605 84.835 -22.275 85.165 ;
        RECT -22.605 83.475 -22.275 83.805 ;
        RECT -22.605 82.115 -22.275 82.445 ;
        RECT -22.605 80.755 -22.275 81.085 ;
        RECT -22.605 79.395 -22.275 79.725 ;
        RECT -22.605 78.035 -22.275 78.365 ;
        RECT -22.605 76.675 -22.275 77.005 ;
        RECT -22.605 75.315 -22.275 75.645 ;
        RECT -22.605 73.955 -22.275 74.285 ;
        RECT -22.605 72.595 -22.275 72.925 ;
        RECT -22.605 71.235 -22.275 71.565 ;
        RECT -22.605 69.875 -22.275 70.205 ;
        RECT -22.605 68.515 -22.275 68.845 ;
        RECT -22.605 67.155 -22.275 67.485 ;
        RECT -22.605 65.795 -22.275 66.125 ;
        RECT -22.605 64.435 -22.275 64.765 ;
        RECT -22.605 63.075 -22.275 63.405 ;
        RECT -22.605 61.715 -22.275 62.045 ;
        RECT -22.605 60.355 -22.275 60.685 ;
        RECT -22.605 58.995 -22.275 59.325 ;
        RECT -22.605 57.635 -22.275 57.965 ;
        RECT -22.605 56.275 -22.275 56.605 ;
        RECT -22.605 54.915 -22.275 55.245 ;
        RECT -22.605 53.555 -22.275 53.885 ;
        RECT -22.605 52.195 -22.275 52.525 ;
        RECT -22.605 50.835 -22.275 51.165 ;
        RECT -22.605 49.475 -22.275 49.805 ;
        RECT -22.605 48.115 -22.275 48.445 ;
        RECT -22.605 46.755 -22.275 47.085 ;
        RECT -22.605 45.395 -22.275 45.725 ;
        RECT -22.605 44.035 -22.275 44.365 ;
        RECT -22.605 42.675 -22.275 43.005 ;
        RECT -22.605 41.315 -22.275 41.645 ;
        RECT -22.605 39.955 -22.275 40.285 ;
        RECT -22.605 38.595 -22.275 38.925 ;
        RECT -22.605 37.235 -22.275 37.565 ;
        RECT -22.605 35.875 -22.275 36.205 ;
        RECT -22.605 34.515 -22.275 34.845 ;
        RECT -22.605 33.155 -22.275 33.485 ;
        RECT -22.605 31.795 -22.275 32.125 ;
        RECT -22.605 30.435 -22.275 30.765 ;
        RECT -22.605 29.075 -22.275 29.405 ;
        RECT -22.605 27.715 -22.275 28.045 ;
        RECT -22.605 26.355 -22.275 26.685 ;
        RECT -22.605 24.995 -22.275 25.325 ;
        RECT -22.605 23.635 -22.275 23.965 ;
        RECT -22.605 22.275 -22.275 22.605 ;
        RECT -22.605 20.915 -22.275 21.245 ;
        RECT -22.605 19.555 -22.275 19.885 ;
        RECT -22.605 18.195 -22.275 18.525 ;
        RECT -22.605 16.835 -22.275 17.165 ;
        RECT -22.605 15.475 -22.275 15.805 ;
        RECT -22.605 14.115 -22.275 14.445 ;
        RECT -22.605 12.755 -22.275 13.085 ;
        RECT -22.605 11.395 -22.275 11.725 ;
        RECT -22.605 10.035 -22.275 10.365 ;
        RECT -22.605 8.675 -22.275 9.005 ;
        RECT -22.605 7.315 -22.275 7.645 ;
        RECT -22.605 5.955 -22.275 6.285 ;
        RECT -22.605 4.595 -22.275 4.925 ;
        RECT -22.605 3.235 -22.275 3.565 ;
        RECT -22.605 1.875 -22.275 2.205 ;
        RECT -22.605 0.515 -22.275 0.845 ;
        RECT -22.605 -2.205 -22.275 -1.875 ;
        RECT -22.605 -3.565 -22.275 -3.235 ;
        RECT -22.605 -7.645 -22.275 -7.315 ;
        RECT -22.605 -10.365 -22.275 -10.035 ;
        RECT -22.605 -11.725 -22.275 -11.395 ;
        RECT -22.605 -13.7 -22.275 -13.37 ;
        RECT -22.605 -14.445 -22.275 -14.115 ;
        RECT -22.605 -15.805 -22.275 -15.475 ;
        RECT -22.605 -18.79 -22.275 -18.46 ;
        RECT -22.605 -19.885 -22.275 -19.555 ;
        RECT -22.605 -23.965 -22.275 -23.635 ;
        RECT -22.605 -25.325 -22.275 -24.995 ;
        RECT -22.605 -29.405 -22.275 -29.075 ;
        RECT -22.605 -32.125 -22.275 -31.795 ;
        RECT -22.605 -33.485 -22.275 -33.155 ;
        RECT -22.605 -34.88 -22.275 -34.55 ;
        RECT -22.605 -36.205 -22.275 -35.875 ;
        RECT -22.605 -38.925 -22.275 -38.595 ;
        RECT -22.605 -39.97 -22.275 -39.64 ;
        RECT -22.605 -47.085 -22.275 -46.755 ;
        RECT -22.605 -48.445 -22.275 -48.115 ;
        RECT -22.605 -49.805 -22.275 -49.475 ;
        RECT -22.605 -51.165 -22.275 -50.835 ;
        RECT -22.605 -52.525 -22.275 -52.195 ;
        RECT -22.605 -53.885 -22.275 -53.555 ;
        RECT -22.605 -55.245 -22.275 -54.915 ;
        RECT -22.605 -56.605 -22.275 -56.275 ;
        RECT -22.605 -57.965 -22.275 -57.635 ;
        RECT -22.605 -59.325 -22.275 -58.995 ;
        RECT -22.605 -60.685 -22.275 -60.355 ;
        RECT -22.605 -62.045 -22.275 -61.715 ;
        RECT -22.605 -63.405 -22.275 -63.075 ;
        RECT -22.605 -64.765 -22.275 -64.435 ;
        RECT -22.605 -68.845 -22.275 -68.515 ;
        RECT -22.605 -71.565 -22.275 -71.235 ;
        RECT -22.605 -72.925 -22.275 -72.595 ;
        RECT -22.605 -74.285 -22.275 -73.955 ;
        RECT -22.605 -75.645 -22.275 -75.315 ;
        RECT -22.605 -77.005 -22.275 -76.675 ;
        RECT -22.605 -78.365 -22.275 -78.035 ;
        RECT -22.605 -80.31 -22.275 -79.98 ;
        RECT -22.605 -81.085 -22.275 -80.755 ;
        RECT -22.605 -82.445 -22.275 -82.115 ;
        RECT -22.605 -83.805 -22.275 -83.475 ;
        RECT -22.605 -85.165 -22.275 -84.835 ;
        RECT -22.605 -86.525 -22.275 -86.195 ;
        RECT -22.605 -87.885 -22.275 -87.555 ;
        RECT -22.605 -90.605 -22.275 -90.275 ;
        RECT -22.605 -91.965 -22.275 -91.635 ;
        RECT -22.605 -93.325 -22.275 -92.995 ;
        RECT -22.605 -94.685 -22.275 -94.355 ;
        RECT -22.605 -96.045 -22.275 -95.715 ;
        RECT -22.605 -97.405 -22.275 -97.075 ;
        RECT -22.605 -98.85 -22.275 -98.52 ;
        RECT -22.605 -100.125 -22.275 -99.795 ;
        RECT -22.605 -101.485 -22.275 -101.155 ;
        RECT -22.605 -102.845 -22.275 -102.515 ;
        RECT -22.605 -105.565 -22.275 -105.235 ;
        RECT -22.605 -106.925 -22.275 -106.595 ;
        RECT -22.605 -108.285 -22.275 -107.955 ;
        RECT -22.605 -109.645 -22.275 -109.315 ;
        RECT -22.605 -111.005 -22.275 -110.675 ;
        RECT -22.605 -112.365 -22.275 -112.035 ;
        RECT -22.605 -113.725 -22.275 -113.395 ;
        RECT -22.605 -116.445 -22.275 -116.115 ;
        RECT -22.605 -117.805 -22.275 -117.475 ;
        RECT -22.605 -119.165 -22.275 -118.835 ;
        RECT -22.605 -120.525 -22.275 -120.195 ;
        RECT -22.605 -121.885 -22.275 -121.555 ;
        RECT -22.605 -124.49 -22.275 -124.16 ;
        RECT -22.605 -128.685 -22.275 -128.355 ;
        RECT -22.605 -130.045 -22.275 -129.715 ;
        RECT -22.605 -131.405 -22.275 -131.075 ;
        RECT -22.605 -132.765 -22.275 -132.435 ;
        RECT -22.605 -136.845 -22.275 -136.515 ;
        RECT -22.605 -138.205 -22.275 -137.875 ;
        RECT -22.605 -139.565 -22.275 -139.235 ;
        RECT -22.605 -140.925 -22.275 -140.595 ;
        RECT -22.605 -142.285 -22.275 -141.955 ;
        RECT -22.605 -143.03 -22.275 -142.7 ;
        RECT -22.605 -145.005 -22.275 -144.675 ;
        RECT -22.605 -146.365 -22.275 -146.035 ;
        RECT -22.605 -147.725 -22.275 -147.395 ;
        RECT -22.605 -153.165 -22.275 -152.835 ;
        RECT -22.605 -154.525 -22.275 -154.195 ;
        RECT -22.605 -155.885 -22.275 -155.555 ;
        RECT -22.605 -157.245 -22.275 -156.915 ;
        RECT -22.605 -162.685 -22.275 -162.355 ;
        RECT -22.605 -164.045 -22.275 -163.715 ;
        RECT -22.605 -165.405 -22.275 -165.075 ;
        RECT -22.605 -166.765 -22.275 -166.435 ;
        RECT -22.605 -168.125 -22.275 -167.795 ;
        RECT -22.605 -169.485 -22.275 -169.155 ;
        RECT -22.605 -170.845 -22.275 -170.515 ;
        RECT -22.605 -172.205 -22.275 -171.875 ;
        RECT -22.605 -174.925 -22.275 -174.595 ;
        RECT -22.605 -176.285 -22.275 -175.955 ;
        RECT -22.605 -177.645 -22.275 -177.315 ;
        RECT -22.605 -179.005 -22.275 -178.675 ;
        RECT -22.605 -180.365 -22.275 -180.035 ;
        RECT -22.605 -181.725 -22.275 -181.395 ;
        RECT -22.605 -183.085 -22.275 -182.755 ;
        RECT -22.605 -192.605 -22.275 -192.275 ;
        RECT -22.605 -193.965 -22.275 -193.635 ;
        RECT -22.605 -195.325 -22.275 -194.995 ;
        RECT -22.605 -198.045 -22.275 -197.715 ;
        RECT -22.605 -199.405 -22.275 -199.075 ;
        RECT -22.605 -200.765 -22.275 -200.435 ;
        RECT -22.605 -203.485 -22.275 -203.155 ;
        RECT -22.605 -204.845 -22.275 -204.515 ;
        RECT -22.605 -206.205 -22.275 -205.875 ;
        RECT -22.605 -208.925 -22.275 -208.595 ;
        RECT -22.605 -210.285 -22.275 -209.955 ;
        RECT -22.605 -214.365 -22.275 -214.035 ;
        RECT -22.605 -215.725 -22.275 -215.395 ;
        RECT -22.605 -217.085 -22.275 -216.755 ;
        RECT -22.605 -218.445 -22.275 -218.115 ;
        RECT -22.605 -219.805 -22.275 -219.475 ;
        RECT -22.605 -221.165 -22.275 -220.835 ;
        RECT -22.605 -222.525 -22.275 -222.195 ;
        RECT -22.605 -223.885 -22.275 -223.555 ;
        RECT -22.605 -225.245 -22.275 -224.915 ;
        RECT -22.605 -232.045 -22.275 -231.715 ;
        RECT -22.605 -234.765 -22.275 -234.435 ;
        RECT -22.605 -236.125 -22.275 -235.795 ;
        RECT -22.605 -237.485 -22.275 -237.155 ;
        RECT -22.605 -238.845 -22.275 -238.515 ;
        RECT -22.605 -241.09 -22.275 -239.96 ;
        RECT -22.6 -241.205 -22.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 244.04 -20.915 245.17 ;
        RECT -21.245 242.595 -20.915 242.925 ;
        RECT -21.245 241.235 -20.915 241.565 ;
        RECT -21.245 239.875 -20.915 240.205 ;
        RECT -21.245 238.515 -20.915 238.845 ;
        RECT -21.245 237.155 -20.915 237.485 ;
        RECT -21.245 235.795 -20.915 236.125 ;
        RECT -21.245 234.435 -20.915 234.765 ;
        RECT -21.245 233.075 -20.915 233.405 ;
        RECT -21.245 231.715 -20.915 232.045 ;
        RECT -21.245 230.355 -20.915 230.685 ;
        RECT -21.245 228.995 -20.915 229.325 ;
        RECT -21.245 227.635 -20.915 227.965 ;
        RECT -21.245 226.275 -20.915 226.605 ;
        RECT -21.245 224.915 -20.915 225.245 ;
        RECT -21.245 223.555 -20.915 223.885 ;
        RECT -21.245 222.195 -20.915 222.525 ;
        RECT -21.245 220.835 -20.915 221.165 ;
        RECT -21.245 219.475 -20.915 219.805 ;
        RECT -21.245 218.115 -20.915 218.445 ;
        RECT -21.245 216.755 -20.915 217.085 ;
        RECT -21.245 215.395 -20.915 215.725 ;
        RECT -21.245 214.035 -20.915 214.365 ;
        RECT -21.245 212.675 -20.915 213.005 ;
        RECT -21.245 211.315 -20.915 211.645 ;
        RECT -21.245 209.955 -20.915 210.285 ;
        RECT -21.245 208.595 -20.915 208.925 ;
        RECT -21.245 207.235 -20.915 207.565 ;
        RECT -21.245 205.875 -20.915 206.205 ;
        RECT -21.245 204.515 -20.915 204.845 ;
        RECT -21.245 203.155 -20.915 203.485 ;
        RECT -21.245 201.795 -20.915 202.125 ;
        RECT -21.245 200.435 -20.915 200.765 ;
        RECT -21.245 199.075 -20.915 199.405 ;
        RECT -21.245 197.715 -20.915 198.045 ;
        RECT -21.245 196.355 -20.915 196.685 ;
        RECT -21.245 194.995 -20.915 195.325 ;
        RECT -21.245 193.635 -20.915 193.965 ;
        RECT -21.245 192.275 -20.915 192.605 ;
        RECT -21.245 190.915 -20.915 191.245 ;
        RECT -21.245 189.555 -20.915 189.885 ;
        RECT -21.245 188.195 -20.915 188.525 ;
        RECT -21.245 186.835 -20.915 187.165 ;
        RECT -21.245 185.475 -20.915 185.805 ;
        RECT -21.245 184.115 -20.915 184.445 ;
        RECT -21.245 182.755 -20.915 183.085 ;
        RECT -21.245 181.395 -20.915 181.725 ;
        RECT -21.245 180.035 -20.915 180.365 ;
        RECT -21.245 178.675 -20.915 179.005 ;
        RECT -21.245 177.315 -20.915 177.645 ;
        RECT -21.245 175.955 -20.915 176.285 ;
        RECT -21.245 174.595 -20.915 174.925 ;
        RECT -21.245 173.235 -20.915 173.565 ;
        RECT -21.245 171.875 -20.915 172.205 ;
        RECT -21.245 170.515 -20.915 170.845 ;
        RECT -21.245 169.155 -20.915 169.485 ;
        RECT -21.245 167.795 -20.915 168.125 ;
        RECT -21.245 166.435 -20.915 166.765 ;
        RECT -21.245 165.075 -20.915 165.405 ;
        RECT -21.245 163.715 -20.915 164.045 ;
        RECT -21.245 162.355 -20.915 162.685 ;
        RECT -21.245 160.995 -20.915 161.325 ;
        RECT -21.245 159.635 -20.915 159.965 ;
        RECT -21.245 158.275 -20.915 158.605 ;
        RECT -21.245 156.915 -20.915 157.245 ;
        RECT -21.245 155.555 -20.915 155.885 ;
        RECT -21.245 154.195 -20.915 154.525 ;
        RECT -21.245 152.835 -20.915 153.165 ;
        RECT -21.245 151.475 -20.915 151.805 ;
        RECT -21.245 150.115 -20.915 150.445 ;
        RECT -21.245 148.755 -20.915 149.085 ;
        RECT -21.245 147.395 -20.915 147.725 ;
        RECT -21.245 146.035 -20.915 146.365 ;
        RECT -21.245 144.675 -20.915 145.005 ;
        RECT -21.245 143.315 -20.915 143.645 ;
        RECT -21.245 141.955 -20.915 142.285 ;
        RECT -21.245 140.595 -20.915 140.925 ;
        RECT -21.245 139.235 -20.915 139.565 ;
        RECT -21.245 137.875 -20.915 138.205 ;
        RECT -21.245 136.515 -20.915 136.845 ;
        RECT -21.245 135.155 -20.915 135.485 ;
        RECT -21.245 133.795 -20.915 134.125 ;
        RECT -21.245 132.435 -20.915 132.765 ;
        RECT -21.245 131.075 -20.915 131.405 ;
        RECT -21.245 129.715 -20.915 130.045 ;
        RECT -21.245 128.355 -20.915 128.685 ;
        RECT -21.245 126.995 -20.915 127.325 ;
        RECT -21.245 125.635 -20.915 125.965 ;
        RECT -21.245 124.275 -20.915 124.605 ;
        RECT -21.245 122.915 -20.915 123.245 ;
        RECT -21.245 121.555 -20.915 121.885 ;
        RECT -21.245 120.195 -20.915 120.525 ;
        RECT -21.245 118.835 -20.915 119.165 ;
        RECT -21.245 117.475 -20.915 117.805 ;
        RECT -21.245 116.115 -20.915 116.445 ;
        RECT -21.245 114.755 -20.915 115.085 ;
        RECT -21.245 113.395 -20.915 113.725 ;
        RECT -21.245 112.035 -20.915 112.365 ;
        RECT -21.245 110.675 -20.915 111.005 ;
        RECT -21.245 109.315 -20.915 109.645 ;
        RECT -21.245 107.955 -20.915 108.285 ;
        RECT -21.245 106.595 -20.915 106.925 ;
        RECT -21.245 105.235 -20.915 105.565 ;
        RECT -21.245 103.875 -20.915 104.205 ;
        RECT -21.245 102.515 -20.915 102.845 ;
        RECT -21.245 101.155 -20.915 101.485 ;
        RECT -21.245 99.795 -20.915 100.125 ;
        RECT -21.245 98.435 -20.915 98.765 ;
        RECT -21.245 97.075 -20.915 97.405 ;
        RECT -21.245 95.715 -20.915 96.045 ;
        RECT -21.245 94.355 -20.915 94.685 ;
        RECT -21.245 92.995 -20.915 93.325 ;
        RECT -21.245 91.635 -20.915 91.965 ;
        RECT -21.245 90.275 -20.915 90.605 ;
        RECT -21.245 88.915 -20.915 89.245 ;
        RECT -21.245 87.555 -20.915 87.885 ;
        RECT -21.245 86.195 -20.915 86.525 ;
        RECT -21.245 84.835 -20.915 85.165 ;
        RECT -21.245 83.475 -20.915 83.805 ;
        RECT -21.245 82.115 -20.915 82.445 ;
        RECT -21.245 80.755 -20.915 81.085 ;
        RECT -21.245 79.395 -20.915 79.725 ;
        RECT -21.245 78.035 -20.915 78.365 ;
        RECT -21.245 76.675 -20.915 77.005 ;
        RECT -21.245 75.315 -20.915 75.645 ;
        RECT -21.245 73.955 -20.915 74.285 ;
        RECT -21.245 72.595 -20.915 72.925 ;
        RECT -21.245 71.235 -20.915 71.565 ;
        RECT -21.245 69.875 -20.915 70.205 ;
        RECT -21.245 68.515 -20.915 68.845 ;
        RECT -21.245 67.155 -20.915 67.485 ;
        RECT -21.245 65.795 -20.915 66.125 ;
        RECT -21.245 64.435 -20.915 64.765 ;
        RECT -21.245 63.075 -20.915 63.405 ;
        RECT -21.245 61.715 -20.915 62.045 ;
        RECT -21.245 60.355 -20.915 60.685 ;
        RECT -21.245 58.995 -20.915 59.325 ;
        RECT -21.245 57.635 -20.915 57.965 ;
        RECT -21.245 56.275 -20.915 56.605 ;
        RECT -21.245 54.915 -20.915 55.245 ;
        RECT -21.245 53.555 -20.915 53.885 ;
        RECT -21.245 52.195 -20.915 52.525 ;
        RECT -21.245 50.835 -20.915 51.165 ;
        RECT -21.245 49.475 -20.915 49.805 ;
        RECT -21.245 48.115 -20.915 48.445 ;
        RECT -21.245 46.755 -20.915 47.085 ;
        RECT -21.245 45.395 -20.915 45.725 ;
        RECT -21.245 44.035 -20.915 44.365 ;
        RECT -21.245 42.675 -20.915 43.005 ;
        RECT -21.245 41.315 -20.915 41.645 ;
        RECT -21.245 39.955 -20.915 40.285 ;
        RECT -21.245 38.595 -20.915 38.925 ;
        RECT -21.245 37.235 -20.915 37.565 ;
        RECT -21.245 35.875 -20.915 36.205 ;
        RECT -21.245 34.515 -20.915 34.845 ;
        RECT -21.245 33.155 -20.915 33.485 ;
        RECT -21.245 31.795 -20.915 32.125 ;
        RECT -21.245 30.435 -20.915 30.765 ;
        RECT -21.245 29.075 -20.915 29.405 ;
        RECT -21.245 27.715 -20.915 28.045 ;
        RECT -21.245 26.355 -20.915 26.685 ;
        RECT -21.245 24.995 -20.915 25.325 ;
        RECT -21.245 23.635 -20.915 23.965 ;
        RECT -21.245 22.275 -20.915 22.605 ;
        RECT -21.245 20.915 -20.915 21.245 ;
        RECT -21.245 19.555 -20.915 19.885 ;
        RECT -21.245 18.195 -20.915 18.525 ;
        RECT -21.245 16.835 -20.915 17.165 ;
        RECT -21.245 15.475 -20.915 15.805 ;
        RECT -21.245 14.115 -20.915 14.445 ;
        RECT -21.245 12.755 -20.915 13.085 ;
        RECT -21.245 11.395 -20.915 11.725 ;
        RECT -21.245 10.035 -20.915 10.365 ;
        RECT -21.245 8.675 -20.915 9.005 ;
        RECT -21.245 7.315 -20.915 7.645 ;
        RECT -21.245 5.955 -20.915 6.285 ;
        RECT -21.245 4.595 -20.915 4.925 ;
        RECT -21.245 3.235 -20.915 3.565 ;
        RECT -21.245 1.875 -20.915 2.205 ;
        RECT -21.245 0.515 -20.915 0.845 ;
        RECT -21.245 -2.205 -20.915 -1.875 ;
        RECT -21.245 -3.565 -20.915 -3.235 ;
        RECT -21.245 -7.645 -20.915 -7.315 ;
        RECT -21.245 -10.365 -20.915 -10.035 ;
        RECT -21.245 -11.725 -20.915 -11.395 ;
        RECT -21.245 -13.7 -20.915 -13.37 ;
        RECT -21.245 -14.445 -20.915 -14.115 ;
        RECT -21.245 -15.805 -20.915 -15.475 ;
        RECT -21.245 -18.79 -20.915 -18.46 ;
        RECT -21.245 -19.885 -20.915 -19.555 ;
        RECT -21.24 -21.92 -20.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -128.685 -20.915 -128.355 ;
        RECT -21.245 -130.045 -20.915 -129.715 ;
        RECT -21.245 -131.405 -20.915 -131.075 ;
        RECT -21.245 -132.765 -20.915 -132.435 ;
        RECT -21.245 -138.205 -20.915 -137.875 ;
        RECT -21.245 -139.565 -20.915 -139.235 ;
        RECT -21.245 -140.925 -20.915 -140.595 ;
        RECT -21.245 -142.285 -20.915 -141.955 ;
        RECT -21.245 -143.03 -20.915 -142.7 ;
        RECT -21.245 -145.005 -20.915 -144.675 ;
        RECT -21.245 -146.365 -20.915 -146.035 ;
        RECT -21.245 -147.725 -20.915 -147.395 ;
        RECT -21.24 -149.76 -20.92 -125.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -232.045 -20.915 -231.715 ;
        RECT -21.245 -233.225 -20.915 -232.895 ;
        RECT -21.245 -234.765 -20.915 -234.435 ;
        RECT -21.245 -236.125 -20.915 -235.795 ;
        RECT -21.245 -237.485 -20.915 -237.155 ;
        RECT -21.245 -238.845 -20.915 -238.515 ;
        RECT -21.245 -241.09 -20.915 -239.96 ;
        RECT -21.24 -241.205 -20.92 -225.6 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 170.515 -19.555 170.845 ;
        RECT -19.885 169.155 -19.555 169.485 ;
        RECT -19.885 167.795 -19.555 168.125 ;
        RECT -19.885 166.435 -19.555 166.765 ;
        RECT -19.885 165.075 -19.555 165.405 ;
        RECT -19.885 163.715 -19.555 164.045 ;
        RECT -19.885 162.355 -19.555 162.685 ;
        RECT -19.885 160.995 -19.555 161.325 ;
        RECT -19.885 159.635 -19.555 159.965 ;
        RECT -19.885 158.275 -19.555 158.605 ;
        RECT -19.885 156.915 -19.555 157.245 ;
        RECT -19.885 155.555 -19.555 155.885 ;
        RECT -19.885 154.195 -19.555 154.525 ;
        RECT -19.885 152.835 -19.555 153.165 ;
        RECT -19.885 151.475 -19.555 151.805 ;
        RECT -19.885 150.115 -19.555 150.445 ;
        RECT -19.885 148.755 -19.555 149.085 ;
        RECT -19.885 147.395 -19.555 147.725 ;
        RECT -19.885 146.035 -19.555 146.365 ;
        RECT -19.885 144.675 -19.555 145.005 ;
        RECT -19.885 143.315 -19.555 143.645 ;
        RECT -19.885 141.955 -19.555 142.285 ;
        RECT -19.885 140.595 -19.555 140.925 ;
        RECT -19.885 139.235 -19.555 139.565 ;
        RECT -19.885 137.875 -19.555 138.205 ;
        RECT -19.885 136.515 -19.555 136.845 ;
        RECT -19.885 135.155 -19.555 135.485 ;
        RECT -19.885 133.795 -19.555 134.125 ;
        RECT -19.885 132.435 -19.555 132.765 ;
        RECT -19.885 131.075 -19.555 131.405 ;
        RECT -19.885 129.715 -19.555 130.045 ;
        RECT -19.885 128.355 -19.555 128.685 ;
        RECT -19.885 126.995 -19.555 127.325 ;
        RECT -19.885 125.635 -19.555 125.965 ;
        RECT -19.885 124.275 -19.555 124.605 ;
        RECT -19.885 122.915 -19.555 123.245 ;
        RECT -19.885 121.555 -19.555 121.885 ;
        RECT -19.885 120.195 -19.555 120.525 ;
        RECT -19.885 118.835 -19.555 119.165 ;
        RECT -19.885 117.475 -19.555 117.805 ;
        RECT -19.885 116.115 -19.555 116.445 ;
        RECT -19.885 114.755 -19.555 115.085 ;
        RECT -19.885 113.395 -19.555 113.725 ;
        RECT -19.885 112.035 -19.555 112.365 ;
        RECT -19.885 110.675 -19.555 111.005 ;
        RECT -19.885 109.315 -19.555 109.645 ;
        RECT -19.885 107.955 -19.555 108.285 ;
        RECT -19.885 106.595 -19.555 106.925 ;
        RECT -19.885 105.235 -19.555 105.565 ;
        RECT -19.885 103.875 -19.555 104.205 ;
        RECT -19.885 102.515 -19.555 102.845 ;
        RECT -19.885 101.155 -19.555 101.485 ;
        RECT -19.885 99.795 -19.555 100.125 ;
        RECT -19.885 98.435 -19.555 98.765 ;
        RECT -19.885 97.075 -19.555 97.405 ;
        RECT -19.885 95.715 -19.555 96.045 ;
        RECT -19.885 94.355 -19.555 94.685 ;
        RECT -19.885 92.995 -19.555 93.325 ;
        RECT -19.885 91.635 -19.555 91.965 ;
        RECT -19.885 90.275 -19.555 90.605 ;
        RECT -19.885 88.915 -19.555 89.245 ;
        RECT -19.885 87.555 -19.555 87.885 ;
        RECT -19.885 86.195 -19.555 86.525 ;
        RECT -19.885 84.835 -19.555 85.165 ;
        RECT -19.885 83.475 -19.555 83.805 ;
        RECT -19.885 82.115 -19.555 82.445 ;
        RECT -19.885 80.755 -19.555 81.085 ;
        RECT -19.885 79.395 -19.555 79.725 ;
        RECT -19.885 78.035 -19.555 78.365 ;
        RECT -19.885 76.675 -19.555 77.005 ;
        RECT -19.885 75.315 -19.555 75.645 ;
        RECT -19.885 73.955 -19.555 74.285 ;
        RECT -19.885 72.595 -19.555 72.925 ;
        RECT -19.885 71.235 -19.555 71.565 ;
        RECT -19.885 69.875 -19.555 70.205 ;
        RECT -19.885 68.515 -19.555 68.845 ;
        RECT -19.885 67.155 -19.555 67.485 ;
        RECT -19.885 65.795 -19.555 66.125 ;
        RECT -19.885 64.435 -19.555 64.765 ;
        RECT -19.885 63.075 -19.555 63.405 ;
        RECT -19.885 61.715 -19.555 62.045 ;
        RECT -19.885 60.355 -19.555 60.685 ;
        RECT -19.885 58.995 -19.555 59.325 ;
        RECT -19.885 57.635 -19.555 57.965 ;
        RECT -19.885 56.275 -19.555 56.605 ;
        RECT -19.885 54.915 -19.555 55.245 ;
        RECT -19.885 53.555 -19.555 53.885 ;
        RECT -19.885 52.195 -19.555 52.525 ;
        RECT -19.885 50.835 -19.555 51.165 ;
        RECT -19.885 49.475 -19.555 49.805 ;
        RECT -19.885 48.115 -19.555 48.445 ;
        RECT -19.885 46.755 -19.555 47.085 ;
        RECT -19.885 45.395 -19.555 45.725 ;
        RECT -19.885 44.035 -19.555 44.365 ;
        RECT -19.885 42.675 -19.555 43.005 ;
        RECT -19.885 41.315 -19.555 41.645 ;
        RECT -19.885 39.955 -19.555 40.285 ;
        RECT -19.885 38.595 -19.555 38.925 ;
        RECT -19.885 37.235 -19.555 37.565 ;
        RECT -19.885 35.875 -19.555 36.205 ;
        RECT -19.885 34.515 -19.555 34.845 ;
        RECT -19.885 33.155 -19.555 33.485 ;
        RECT -19.885 31.795 -19.555 32.125 ;
        RECT -19.885 30.435 -19.555 30.765 ;
        RECT -19.885 29.075 -19.555 29.405 ;
        RECT -19.885 27.715 -19.555 28.045 ;
        RECT -19.885 26.355 -19.555 26.685 ;
        RECT -19.885 24.995 -19.555 25.325 ;
        RECT -19.885 23.635 -19.555 23.965 ;
        RECT -19.885 22.275 -19.555 22.605 ;
        RECT -19.885 20.915 -19.555 21.245 ;
        RECT -19.885 19.555 -19.555 19.885 ;
        RECT -19.885 18.195 -19.555 18.525 ;
        RECT -19.885 16.835 -19.555 17.165 ;
        RECT -19.885 15.475 -19.555 15.805 ;
        RECT -19.885 14.115 -19.555 14.445 ;
        RECT -19.885 12.755 -19.555 13.085 ;
        RECT -19.885 11.395 -19.555 11.725 ;
        RECT -19.885 10.035 -19.555 10.365 ;
        RECT -19.885 8.675 -19.555 9.005 ;
        RECT -19.885 7.315 -19.555 7.645 ;
        RECT -19.885 5.955 -19.555 6.285 ;
        RECT -19.885 4.595 -19.555 4.925 ;
        RECT -19.885 3.235 -19.555 3.565 ;
        RECT -19.885 1.875 -19.555 2.205 ;
        RECT -19.885 0.515 -19.555 0.845 ;
        RECT -19.885 -2.205 -19.555 -1.875 ;
        RECT -19.885 -3.565 -19.555 -3.235 ;
        RECT -19.885 -7.645 -19.555 -7.315 ;
        RECT -19.885 -10.365 -19.555 -10.035 ;
        RECT -19.885 -11.725 -19.555 -11.395 ;
        RECT -19.885 -13.7 -19.555 -13.37 ;
        RECT -19.885 -14.445 -19.555 -14.115 ;
        RECT -19.885 -15.805 -19.555 -15.475 ;
        RECT -19.885 -18.79 -19.555 -18.46 ;
        RECT -19.885 -19.885 -19.555 -19.555 ;
        RECT -19.88 -20.56 -19.56 245.285 ;
        RECT -19.885 244.04 -19.555 245.17 ;
        RECT -19.885 242.595 -19.555 242.925 ;
        RECT -19.885 241.235 -19.555 241.565 ;
        RECT -19.885 239.875 -19.555 240.205 ;
        RECT -19.885 238.515 -19.555 238.845 ;
        RECT -19.885 237.155 -19.555 237.485 ;
        RECT -19.885 235.795 -19.555 236.125 ;
        RECT -19.885 234.435 -19.555 234.765 ;
        RECT -19.885 233.075 -19.555 233.405 ;
        RECT -19.885 231.715 -19.555 232.045 ;
        RECT -19.885 230.355 -19.555 230.685 ;
        RECT -19.885 228.995 -19.555 229.325 ;
        RECT -19.885 227.635 -19.555 227.965 ;
        RECT -19.885 226.275 -19.555 226.605 ;
        RECT -19.885 224.915 -19.555 225.245 ;
        RECT -19.885 223.555 -19.555 223.885 ;
        RECT -19.885 222.195 -19.555 222.525 ;
        RECT -19.885 220.835 -19.555 221.165 ;
        RECT -19.885 219.475 -19.555 219.805 ;
        RECT -19.885 218.115 -19.555 218.445 ;
        RECT -19.885 216.755 -19.555 217.085 ;
        RECT -19.885 215.395 -19.555 215.725 ;
        RECT -19.885 214.035 -19.555 214.365 ;
        RECT -19.885 212.675 -19.555 213.005 ;
        RECT -19.885 211.315 -19.555 211.645 ;
        RECT -19.885 209.955 -19.555 210.285 ;
        RECT -19.885 208.595 -19.555 208.925 ;
        RECT -19.885 207.235 -19.555 207.565 ;
        RECT -19.885 205.875 -19.555 206.205 ;
        RECT -19.885 204.515 -19.555 204.845 ;
        RECT -19.885 203.155 -19.555 203.485 ;
        RECT -19.885 201.795 -19.555 202.125 ;
        RECT -19.885 200.435 -19.555 200.765 ;
        RECT -19.885 199.075 -19.555 199.405 ;
        RECT -19.885 197.715 -19.555 198.045 ;
        RECT -19.885 196.355 -19.555 196.685 ;
        RECT -19.885 194.995 -19.555 195.325 ;
        RECT -19.885 193.635 -19.555 193.965 ;
        RECT -19.885 192.275 -19.555 192.605 ;
        RECT -19.885 190.915 -19.555 191.245 ;
        RECT -19.885 189.555 -19.555 189.885 ;
        RECT -19.885 188.195 -19.555 188.525 ;
        RECT -19.885 186.835 -19.555 187.165 ;
        RECT -19.885 185.475 -19.555 185.805 ;
        RECT -19.885 184.115 -19.555 184.445 ;
        RECT -19.885 182.755 -19.555 183.085 ;
        RECT -19.885 181.395 -19.555 181.725 ;
        RECT -19.885 180.035 -19.555 180.365 ;
        RECT -19.885 178.675 -19.555 179.005 ;
        RECT -19.885 177.315 -19.555 177.645 ;
        RECT -19.885 175.955 -19.555 176.285 ;
        RECT -19.885 174.595 -19.555 174.925 ;
        RECT -19.885 173.235 -19.555 173.565 ;
        RECT -19.885 171.875 -19.555 172.205 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -124.49 -29.075 -124.16 ;
        RECT -29.405 -128.685 -29.075 -128.355 ;
        RECT -29.405 -130.045 -29.075 -129.715 ;
        RECT -29.405 -131.405 -29.075 -131.075 ;
        RECT -29.405 -132.765 -29.075 -132.435 ;
        RECT -29.405 -135.485 -29.075 -135.155 ;
        RECT -29.405 -136.845 -29.075 -136.515 ;
        RECT -29.405 -138.205 -29.075 -137.875 ;
        RECT -29.405 -139.565 -29.075 -139.235 ;
        RECT -29.405 -140.925 -29.075 -140.595 ;
        RECT -29.405 -142.285 -29.075 -141.955 ;
        RECT -29.405 -143.03 -29.075 -142.7 ;
        RECT -29.405 -145.005 -29.075 -144.675 ;
        RECT -29.405 -146.365 -29.075 -146.035 ;
        RECT -29.405 -147.725 -29.075 -147.395 ;
        RECT -29.405 -153.165 -29.075 -152.835 ;
        RECT -29.405 -154.525 -29.075 -154.195 ;
        RECT -29.405 -155.885 -29.075 -155.555 ;
        RECT -29.405 -157.245 -29.075 -156.915 ;
        RECT -29.405 -162.685 -29.075 -162.355 ;
        RECT -29.405 -164.045 -29.075 -163.715 ;
        RECT -29.405 -165.405 -29.075 -165.075 ;
        RECT -29.405 -166.765 -29.075 -166.435 ;
        RECT -29.405 -168.125 -29.075 -167.795 ;
        RECT -29.405 -169.485 -29.075 -169.155 ;
        RECT -29.405 -170.845 -29.075 -170.515 ;
        RECT -29.405 -172.205 -29.075 -171.875 ;
        RECT -29.405 -173.565 -29.075 -173.235 ;
        RECT -29.405 -174.925 -29.075 -174.595 ;
        RECT -29.405 -176.285 -29.075 -175.955 ;
        RECT -29.405 -177.645 -29.075 -177.315 ;
        RECT -29.405 -179.005 -29.075 -178.675 ;
        RECT -29.405 -180.365 -29.075 -180.035 ;
        RECT -29.405 -181.725 -29.075 -181.395 ;
        RECT -29.405 -183.085 -29.075 -182.755 ;
        RECT -29.405 -184.445 -29.075 -184.115 ;
        RECT -29.405 -185.805 -29.075 -185.475 ;
        RECT -29.405 -187.165 -29.075 -186.835 ;
        RECT -29.405 -191.245 -29.075 -190.915 ;
        RECT -29.405 -192.605 -29.075 -192.275 ;
        RECT -29.405 -193.965 -29.075 -193.635 ;
        RECT -29.405 -195.325 -29.075 -194.995 ;
        RECT -29.405 -198.045 -29.075 -197.715 ;
        RECT -29.405 -199.405 -29.075 -199.075 ;
        RECT -29.405 -200.765 -29.075 -200.435 ;
        RECT -29.405 -202.125 -29.075 -201.795 ;
        RECT -29.405 -203.485 -29.075 -203.155 ;
        RECT -29.405 -204.845 -29.075 -204.515 ;
        RECT -29.405 -206.205 -29.075 -205.875 ;
        RECT -29.405 -208.925 -29.075 -208.595 ;
        RECT -29.405 -210.285 -29.075 -209.955 ;
        RECT -29.405 -215.725 -29.075 -215.395 ;
        RECT -29.405 -217.085 -29.075 -216.755 ;
        RECT -29.405 -218.445 -29.075 -218.115 ;
        RECT -29.405 -219.805 -29.075 -219.475 ;
        RECT -29.405 -221.165 -29.075 -220.835 ;
        RECT -29.405 -222.525 -29.075 -222.195 ;
        RECT -29.405 -223.885 -29.075 -223.555 ;
        RECT -29.405 -225.245 -29.075 -224.915 ;
        RECT -29.4 -227.96 -29.08 -122.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -232.045 -29.075 -231.715 ;
        RECT -29.405 -233.225 -29.075 -232.895 ;
        RECT -29.405 -234.765 -29.075 -234.435 ;
        RECT -29.405 -236.125 -29.075 -235.795 ;
        RECT -29.405 -237.485 -29.075 -237.155 ;
        RECT -29.405 -238.845 -29.075 -238.515 ;
        RECT -29.405 -241.09 -29.075 -239.96 ;
        RECT -29.4 -241.205 -29.08 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.045 244.04 -27.715 245.17 ;
        RECT -28.045 242.595 -27.715 242.925 ;
        RECT -28.045 241.235 -27.715 241.565 ;
        RECT -28.045 239.875 -27.715 240.205 ;
        RECT -28.045 238.515 -27.715 238.845 ;
        RECT -28.045 237.155 -27.715 237.485 ;
        RECT -28.045 235.795 -27.715 236.125 ;
        RECT -28.045 234.435 -27.715 234.765 ;
        RECT -28.045 233.075 -27.715 233.405 ;
        RECT -28.045 231.715 -27.715 232.045 ;
        RECT -28.045 230.355 -27.715 230.685 ;
        RECT -28.045 228.995 -27.715 229.325 ;
        RECT -28.045 227.635 -27.715 227.965 ;
        RECT -28.045 226.275 -27.715 226.605 ;
        RECT -28.045 224.915 -27.715 225.245 ;
        RECT -28.045 223.555 -27.715 223.885 ;
        RECT -28.045 222.195 -27.715 222.525 ;
        RECT -28.045 220.835 -27.715 221.165 ;
        RECT -28.045 219.475 -27.715 219.805 ;
        RECT -28.045 218.115 -27.715 218.445 ;
        RECT -28.045 216.755 -27.715 217.085 ;
        RECT -28.045 215.395 -27.715 215.725 ;
        RECT -28.045 214.035 -27.715 214.365 ;
        RECT -28.045 212.675 -27.715 213.005 ;
        RECT -28.045 211.315 -27.715 211.645 ;
        RECT -28.045 209.955 -27.715 210.285 ;
        RECT -28.045 208.595 -27.715 208.925 ;
        RECT -28.045 207.235 -27.715 207.565 ;
        RECT -28.045 205.875 -27.715 206.205 ;
        RECT -28.045 204.515 -27.715 204.845 ;
        RECT -28.045 203.155 -27.715 203.485 ;
        RECT -28.045 201.795 -27.715 202.125 ;
        RECT -28.045 200.435 -27.715 200.765 ;
        RECT -28.045 199.075 -27.715 199.405 ;
        RECT -28.045 197.715 -27.715 198.045 ;
        RECT -28.045 196.355 -27.715 196.685 ;
        RECT -28.045 194.995 -27.715 195.325 ;
        RECT -28.045 193.635 -27.715 193.965 ;
        RECT -28.045 192.275 -27.715 192.605 ;
        RECT -28.045 190.915 -27.715 191.245 ;
        RECT -28.045 189.555 -27.715 189.885 ;
        RECT -28.045 188.195 -27.715 188.525 ;
        RECT -28.045 186.835 -27.715 187.165 ;
        RECT -28.045 185.475 -27.715 185.805 ;
        RECT -28.045 184.115 -27.715 184.445 ;
        RECT -28.045 182.755 -27.715 183.085 ;
        RECT -28.045 181.395 -27.715 181.725 ;
        RECT -28.045 180.035 -27.715 180.365 ;
        RECT -28.045 178.675 -27.715 179.005 ;
        RECT -28.045 177.315 -27.715 177.645 ;
        RECT -28.045 175.955 -27.715 176.285 ;
        RECT -28.045 174.595 -27.715 174.925 ;
        RECT -28.045 173.235 -27.715 173.565 ;
        RECT -28.045 171.875 -27.715 172.205 ;
        RECT -28.045 170.515 -27.715 170.845 ;
        RECT -28.045 169.155 -27.715 169.485 ;
        RECT -28.045 167.795 -27.715 168.125 ;
        RECT -28.045 166.435 -27.715 166.765 ;
        RECT -28.045 165.075 -27.715 165.405 ;
        RECT -28.045 163.715 -27.715 164.045 ;
        RECT -28.045 162.355 -27.715 162.685 ;
        RECT -28.045 160.995 -27.715 161.325 ;
        RECT -28.045 159.635 -27.715 159.965 ;
        RECT -28.045 158.275 -27.715 158.605 ;
        RECT -28.045 156.915 -27.715 157.245 ;
        RECT -28.045 155.555 -27.715 155.885 ;
        RECT -28.045 154.195 -27.715 154.525 ;
        RECT -28.045 152.835 -27.715 153.165 ;
        RECT -28.045 151.475 -27.715 151.805 ;
        RECT -28.045 150.115 -27.715 150.445 ;
        RECT -28.045 148.755 -27.715 149.085 ;
        RECT -28.045 147.395 -27.715 147.725 ;
        RECT -28.045 146.035 -27.715 146.365 ;
        RECT -28.045 144.675 -27.715 145.005 ;
        RECT -28.045 143.315 -27.715 143.645 ;
        RECT -28.045 141.955 -27.715 142.285 ;
        RECT -28.045 140.595 -27.715 140.925 ;
        RECT -28.045 139.235 -27.715 139.565 ;
        RECT -28.045 137.875 -27.715 138.205 ;
        RECT -28.045 136.515 -27.715 136.845 ;
        RECT -28.045 135.155 -27.715 135.485 ;
        RECT -28.045 133.795 -27.715 134.125 ;
        RECT -28.045 132.435 -27.715 132.765 ;
        RECT -28.045 131.075 -27.715 131.405 ;
        RECT -28.045 129.715 -27.715 130.045 ;
        RECT -28.045 128.355 -27.715 128.685 ;
        RECT -28.045 126.995 -27.715 127.325 ;
        RECT -28.045 125.635 -27.715 125.965 ;
        RECT -28.045 124.275 -27.715 124.605 ;
        RECT -28.045 122.915 -27.715 123.245 ;
        RECT -28.045 121.555 -27.715 121.885 ;
        RECT -28.045 120.195 -27.715 120.525 ;
        RECT -28.045 118.835 -27.715 119.165 ;
        RECT -28.045 117.475 -27.715 117.805 ;
        RECT -28.045 116.115 -27.715 116.445 ;
        RECT -28.045 114.755 -27.715 115.085 ;
        RECT -28.045 113.395 -27.715 113.725 ;
        RECT -28.045 112.035 -27.715 112.365 ;
        RECT -28.045 110.675 -27.715 111.005 ;
        RECT -28.045 109.315 -27.715 109.645 ;
        RECT -28.045 107.955 -27.715 108.285 ;
        RECT -28.045 106.595 -27.715 106.925 ;
        RECT -28.045 105.235 -27.715 105.565 ;
        RECT -28.045 103.875 -27.715 104.205 ;
        RECT -28.045 102.515 -27.715 102.845 ;
        RECT -28.045 101.155 -27.715 101.485 ;
        RECT -28.045 99.795 -27.715 100.125 ;
        RECT -28.045 98.435 -27.715 98.765 ;
        RECT -28.045 97.075 -27.715 97.405 ;
        RECT -28.045 95.715 -27.715 96.045 ;
        RECT -28.045 94.355 -27.715 94.685 ;
        RECT -28.045 92.995 -27.715 93.325 ;
        RECT -28.045 91.635 -27.715 91.965 ;
        RECT -28.045 90.275 -27.715 90.605 ;
        RECT -28.045 88.915 -27.715 89.245 ;
        RECT -28.045 87.555 -27.715 87.885 ;
        RECT -28.045 86.195 -27.715 86.525 ;
        RECT -28.045 84.835 -27.715 85.165 ;
        RECT -28.045 83.475 -27.715 83.805 ;
        RECT -28.045 82.115 -27.715 82.445 ;
        RECT -28.045 80.755 -27.715 81.085 ;
        RECT -28.045 79.395 -27.715 79.725 ;
        RECT -28.045 78.035 -27.715 78.365 ;
        RECT -28.045 76.675 -27.715 77.005 ;
        RECT -28.045 75.315 -27.715 75.645 ;
        RECT -28.045 73.955 -27.715 74.285 ;
        RECT -28.045 72.595 -27.715 72.925 ;
        RECT -28.045 71.235 -27.715 71.565 ;
        RECT -28.045 69.875 -27.715 70.205 ;
        RECT -28.045 68.515 -27.715 68.845 ;
        RECT -28.045 67.155 -27.715 67.485 ;
        RECT -28.045 65.795 -27.715 66.125 ;
        RECT -28.045 64.435 -27.715 64.765 ;
        RECT -28.045 63.075 -27.715 63.405 ;
        RECT -28.045 61.715 -27.715 62.045 ;
        RECT -28.045 60.355 -27.715 60.685 ;
        RECT -28.045 58.995 -27.715 59.325 ;
        RECT -28.045 57.635 -27.715 57.965 ;
        RECT -28.045 56.275 -27.715 56.605 ;
        RECT -28.045 54.915 -27.715 55.245 ;
        RECT -28.045 53.555 -27.715 53.885 ;
        RECT -28.045 52.195 -27.715 52.525 ;
        RECT -28.045 50.835 -27.715 51.165 ;
        RECT -28.045 49.475 -27.715 49.805 ;
        RECT -28.045 48.115 -27.715 48.445 ;
        RECT -28.045 46.755 -27.715 47.085 ;
        RECT -28.045 45.395 -27.715 45.725 ;
        RECT -28.045 44.035 -27.715 44.365 ;
        RECT -28.045 42.675 -27.715 43.005 ;
        RECT -28.045 41.315 -27.715 41.645 ;
        RECT -28.045 39.955 -27.715 40.285 ;
        RECT -28.045 38.595 -27.715 38.925 ;
        RECT -28.045 37.235 -27.715 37.565 ;
        RECT -28.045 35.875 -27.715 36.205 ;
        RECT -28.045 34.515 -27.715 34.845 ;
        RECT -28.045 33.155 -27.715 33.485 ;
        RECT -28.045 31.795 -27.715 32.125 ;
        RECT -28.045 30.435 -27.715 30.765 ;
        RECT -28.045 29.075 -27.715 29.405 ;
        RECT -28.045 27.715 -27.715 28.045 ;
        RECT -28.045 26.355 -27.715 26.685 ;
        RECT -28.045 24.995 -27.715 25.325 ;
        RECT -28.045 23.635 -27.715 23.965 ;
        RECT -28.045 22.275 -27.715 22.605 ;
        RECT -28.045 20.915 -27.715 21.245 ;
        RECT -28.045 19.555 -27.715 19.885 ;
        RECT -28.045 18.195 -27.715 18.525 ;
        RECT -28.045 16.835 -27.715 17.165 ;
        RECT -28.045 15.475 -27.715 15.805 ;
        RECT -28.045 14.115 -27.715 14.445 ;
        RECT -28.045 12.755 -27.715 13.085 ;
        RECT -28.045 11.395 -27.715 11.725 ;
        RECT -28.045 10.035 -27.715 10.365 ;
        RECT -28.045 8.675 -27.715 9.005 ;
        RECT -28.045 7.315 -27.715 7.645 ;
        RECT -28.045 5.955 -27.715 6.285 ;
        RECT -28.045 4.595 -27.715 4.925 ;
        RECT -28.045 3.235 -27.715 3.565 ;
        RECT -28.045 1.875 -27.715 2.205 ;
        RECT -28.045 0.515 -27.715 0.845 ;
        RECT -28.045 -7.645 -27.715 -7.315 ;
        RECT -28.045 -10.365 -27.715 -10.035 ;
        RECT -28.045 -11.725 -27.715 -11.395 ;
        RECT -28.045 -13.7 -27.715 -13.37 ;
        RECT -28.045 -14.445 -27.715 -14.115 ;
        RECT -28.045 -15.805 -27.715 -15.475 ;
        RECT -28.045 -18.79 -27.715 -18.46 ;
        RECT -28.045 -19.885 -27.715 -19.555 ;
        RECT -28.045 -29.405 -27.715 -29.075 ;
        RECT -28.045 -32.125 -27.715 -31.795 ;
        RECT -28.045 -33.485 -27.715 -33.155 ;
        RECT -28.045 -34.88 -27.715 -34.55 ;
        RECT -28.045 -36.205 -27.715 -35.875 ;
        RECT -28.045 -38.925 -27.715 -38.595 ;
        RECT -28.045 -39.97 -27.715 -39.64 ;
        RECT -28.045 -48.445 -27.715 -48.115 ;
        RECT -28.045 -49.805 -27.715 -49.475 ;
        RECT -28.045 -51.165 -27.715 -50.835 ;
        RECT -28.045 -53.885 -27.715 -53.555 ;
        RECT -28.045 -57.965 -27.715 -57.635 ;
        RECT -28.045 -62.045 -27.715 -61.715 ;
        RECT -28.045 -63.405 -27.715 -63.075 ;
        RECT -28.045 -64.765 -27.715 -64.435 ;
        RECT -28.045 -66.125 -27.715 -65.795 ;
        RECT -28.045 -68.845 -27.715 -68.515 ;
        RECT -28.045 -71.565 -27.715 -71.235 ;
        RECT -28.045 -72.925 -27.715 -72.595 ;
        RECT -28.045 -74.285 -27.715 -73.955 ;
        RECT -28.045 -75.645 -27.715 -75.315 ;
        RECT -28.045 -77.005 -27.715 -76.675 ;
        RECT -28.045 -78.365 -27.715 -78.035 ;
        RECT -28.045 -80.31 -27.715 -79.98 ;
        RECT -28.045 -81.085 -27.715 -80.755 ;
        RECT -28.045 -82.445 -27.715 -82.115 ;
        RECT -28.045 -83.805 -27.715 -83.475 ;
        RECT -28.045 -85.165 -27.715 -84.835 ;
        RECT -28.045 -86.525 -27.715 -86.195 ;
        RECT -28.045 -87.885 -27.715 -87.555 ;
        RECT -28.045 -90.605 -27.715 -90.275 ;
        RECT -28.045 -91.965 -27.715 -91.635 ;
        RECT -28.045 -93.325 -27.715 -92.995 ;
        RECT -28.045 -94.685 -27.715 -94.355 ;
        RECT -28.045 -96.045 -27.715 -95.715 ;
        RECT -28.045 -97.405 -27.715 -97.075 ;
        RECT -28.045 -98.85 -27.715 -98.52 ;
        RECT -28.045 -100.125 -27.715 -99.795 ;
        RECT -28.045 -101.485 -27.715 -101.155 ;
        RECT -28.045 -102.845 -27.715 -102.515 ;
        RECT -28.045 -105.565 -27.715 -105.235 ;
        RECT -28.045 -106.925 -27.715 -106.595 ;
        RECT -28.045 -108.285 -27.715 -107.955 ;
        RECT -28.045 -109.645 -27.715 -109.315 ;
        RECT -28.045 -111.005 -27.715 -110.675 ;
        RECT -28.045 -112.365 -27.715 -112.035 ;
        RECT -28.045 -113.725 -27.715 -113.395 ;
        RECT -28.045 -116.445 -27.715 -116.115 ;
        RECT -28.045 -117.805 -27.715 -117.475 ;
        RECT -28.045 -119.165 -27.715 -118.835 ;
        RECT -28.045 -120.525 -27.715 -120.195 ;
        RECT -28.045 -121.885 -27.715 -121.555 ;
        RECT -28.045 -124.49 -27.715 -124.16 ;
        RECT -28.045 -128.685 -27.715 -128.355 ;
        RECT -28.045 -130.045 -27.715 -129.715 ;
        RECT -28.045 -131.405 -27.715 -131.075 ;
        RECT -28.045 -132.765 -27.715 -132.435 ;
        RECT -28.045 -135.485 -27.715 -135.155 ;
        RECT -28.045 -136.845 -27.715 -136.515 ;
        RECT -28.045 -138.205 -27.715 -137.875 ;
        RECT -28.045 -139.565 -27.715 -139.235 ;
        RECT -28.045 -140.925 -27.715 -140.595 ;
        RECT -28.045 -142.285 -27.715 -141.955 ;
        RECT -28.045 -143.03 -27.715 -142.7 ;
        RECT -28.045 -145.005 -27.715 -144.675 ;
        RECT -28.045 -146.365 -27.715 -146.035 ;
        RECT -28.045 -147.725 -27.715 -147.395 ;
        RECT -28.045 -153.165 -27.715 -152.835 ;
        RECT -28.045 -154.525 -27.715 -154.195 ;
        RECT -28.045 -155.885 -27.715 -155.555 ;
        RECT -28.045 -157.245 -27.715 -156.915 ;
        RECT -28.045 -162.685 -27.715 -162.355 ;
        RECT -28.045 -164.045 -27.715 -163.715 ;
        RECT -28.045 -165.405 -27.715 -165.075 ;
        RECT -28.045 -166.765 -27.715 -166.435 ;
        RECT -28.045 -168.125 -27.715 -167.795 ;
        RECT -28.045 -169.485 -27.715 -169.155 ;
        RECT -28.045 -170.845 -27.715 -170.515 ;
        RECT -28.045 -172.205 -27.715 -171.875 ;
        RECT -28.045 -173.565 -27.715 -173.235 ;
        RECT -28.045 -174.925 -27.715 -174.595 ;
        RECT -28.045 -176.285 -27.715 -175.955 ;
        RECT -28.045 -177.645 -27.715 -177.315 ;
        RECT -28.045 -179.005 -27.715 -178.675 ;
        RECT -28.045 -180.365 -27.715 -180.035 ;
        RECT -28.045 -181.725 -27.715 -181.395 ;
        RECT -28.045 -183.085 -27.715 -182.755 ;
        RECT -28.045 -184.445 -27.715 -184.115 ;
        RECT -28.045 -185.805 -27.715 -185.475 ;
        RECT -28.045 -187.165 -27.715 -186.835 ;
        RECT -28.045 -191.245 -27.715 -190.915 ;
        RECT -28.045 -192.605 -27.715 -192.275 ;
        RECT -28.045 -193.965 -27.715 -193.635 ;
        RECT -28.045 -195.325 -27.715 -194.995 ;
        RECT -28.045 -198.045 -27.715 -197.715 ;
        RECT -28.045 -199.405 -27.715 -199.075 ;
        RECT -28.045 -200.765 -27.715 -200.435 ;
        RECT -28.045 -202.125 -27.715 -201.795 ;
        RECT -28.045 -203.485 -27.715 -203.155 ;
        RECT -28.045 -204.845 -27.715 -204.515 ;
        RECT -28.045 -206.205 -27.715 -205.875 ;
        RECT -28.045 -208.925 -27.715 -208.595 ;
        RECT -28.045 -210.285 -27.715 -209.955 ;
        RECT -28.045 -215.725 -27.715 -215.395 ;
        RECT -28.045 -217.085 -27.715 -216.755 ;
        RECT -28.045 -218.445 -27.715 -218.115 ;
        RECT -28.045 -219.805 -27.715 -219.475 ;
        RECT -28.045 -221.165 -27.715 -220.835 ;
        RECT -28.045 -222.525 -27.715 -222.195 ;
        RECT -28.045 -223.885 -27.715 -223.555 ;
        RECT -28.045 -225.245 -27.715 -224.915 ;
        RECT -28.04 -229.32 -27.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 244.04 -26.355 245.17 ;
        RECT -26.685 242.595 -26.355 242.925 ;
        RECT -26.685 241.235 -26.355 241.565 ;
        RECT -26.685 239.875 -26.355 240.205 ;
        RECT -26.685 238.515 -26.355 238.845 ;
        RECT -26.685 237.155 -26.355 237.485 ;
        RECT -26.685 235.795 -26.355 236.125 ;
        RECT -26.685 234.435 -26.355 234.765 ;
        RECT -26.685 233.075 -26.355 233.405 ;
        RECT -26.685 231.715 -26.355 232.045 ;
        RECT -26.685 230.355 -26.355 230.685 ;
        RECT -26.685 228.995 -26.355 229.325 ;
        RECT -26.685 227.635 -26.355 227.965 ;
        RECT -26.685 226.275 -26.355 226.605 ;
        RECT -26.685 224.915 -26.355 225.245 ;
        RECT -26.685 223.555 -26.355 223.885 ;
        RECT -26.685 222.195 -26.355 222.525 ;
        RECT -26.685 220.835 -26.355 221.165 ;
        RECT -26.685 219.475 -26.355 219.805 ;
        RECT -26.685 218.115 -26.355 218.445 ;
        RECT -26.685 216.755 -26.355 217.085 ;
        RECT -26.685 215.395 -26.355 215.725 ;
        RECT -26.685 214.035 -26.355 214.365 ;
        RECT -26.685 212.675 -26.355 213.005 ;
        RECT -26.685 211.315 -26.355 211.645 ;
        RECT -26.685 209.955 -26.355 210.285 ;
        RECT -26.685 208.595 -26.355 208.925 ;
        RECT -26.685 207.235 -26.355 207.565 ;
        RECT -26.685 205.875 -26.355 206.205 ;
        RECT -26.685 204.515 -26.355 204.845 ;
        RECT -26.685 203.155 -26.355 203.485 ;
        RECT -26.685 201.795 -26.355 202.125 ;
        RECT -26.685 200.435 -26.355 200.765 ;
        RECT -26.685 199.075 -26.355 199.405 ;
        RECT -26.685 197.715 -26.355 198.045 ;
        RECT -26.685 196.355 -26.355 196.685 ;
        RECT -26.685 194.995 -26.355 195.325 ;
        RECT -26.685 193.635 -26.355 193.965 ;
        RECT -26.685 192.275 -26.355 192.605 ;
        RECT -26.685 190.915 -26.355 191.245 ;
        RECT -26.685 189.555 -26.355 189.885 ;
        RECT -26.685 188.195 -26.355 188.525 ;
        RECT -26.685 186.835 -26.355 187.165 ;
        RECT -26.685 185.475 -26.355 185.805 ;
        RECT -26.685 184.115 -26.355 184.445 ;
        RECT -26.685 182.755 -26.355 183.085 ;
        RECT -26.685 181.395 -26.355 181.725 ;
        RECT -26.685 180.035 -26.355 180.365 ;
        RECT -26.685 178.675 -26.355 179.005 ;
        RECT -26.685 177.315 -26.355 177.645 ;
        RECT -26.685 175.955 -26.355 176.285 ;
        RECT -26.685 174.595 -26.355 174.925 ;
        RECT -26.685 173.235 -26.355 173.565 ;
        RECT -26.685 171.875 -26.355 172.205 ;
        RECT -26.685 170.515 -26.355 170.845 ;
        RECT -26.685 169.155 -26.355 169.485 ;
        RECT -26.685 167.795 -26.355 168.125 ;
        RECT -26.685 166.435 -26.355 166.765 ;
        RECT -26.685 165.075 -26.355 165.405 ;
        RECT -26.685 163.715 -26.355 164.045 ;
        RECT -26.685 162.355 -26.355 162.685 ;
        RECT -26.685 160.995 -26.355 161.325 ;
        RECT -26.685 159.635 -26.355 159.965 ;
        RECT -26.685 158.275 -26.355 158.605 ;
        RECT -26.685 156.915 -26.355 157.245 ;
        RECT -26.685 155.555 -26.355 155.885 ;
        RECT -26.685 154.195 -26.355 154.525 ;
        RECT -26.685 152.835 -26.355 153.165 ;
        RECT -26.685 151.475 -26.355 151.805 ;
        RECT -26.685 150.115 -26.355 150.445 ;
        RECT -26.685 148.755 -26.355 149.085 ;
        RECT -26.685 147.395 -26.355 147.725 ;
        RECT -26.685 146.035 -26.355 146.365 ;
        RECT -26.685 144.675 -26.355 145.005 ;
        RECT -26.685 143.315 -26.355 143.645 ;
        RECT -26.685 141.955 -26.355 142.285 ;
        RECT -26.685 140.595 -26.355 140.925 ;
        RECT -26.685 139.235 -26.355 139.565 ;
        RECT -26.685 137.875 -26.355 138.205 ;
        RECT -26.685 136.515 -26.355 136.845 ;
        RECT -26.685 135.155 -26.355 135.485 ;
        RECT -26.685 133.795 -26.355 134.125 ;
        RECT -26.685 132.435 -26.355 132.765 ;
        RECT -26.685 131.075 -26.355 131.405 ;
        RECT -26.685 129.715 -26.355 130.045 ;
        RECT -26.685 128.355 -26.355 128.685 ;
        RECT -26.685 126.995 -26.355 127.325 ;
        RECT -26.685 125.635 -26.355 125.965 ;
        RECT -26.685 124.275 -26.355 124.605 ;
        RECT -26.685 122.915 -26.355 123.245 ;
        RECT -26.685 121.555 -26.355 121.885 ;
        RECT -26.685 120.195 -26.355 120.525 ;
        RECT -26.685 118.835 -26.355 119.165 ;
        RECT -26.685 117.475 -26.355 117.805 ;
        RECT -26.685 116.115 -26.355 116.445 ;
        RECT -26.685 114.755 -26.355 115.085 ;
        RECT -26.685 113.395 -26.355 113.725 ;
        RECT -26.685 112.035 -26.355 112.365 ;
        RECT -26.685 110.675 -26.355 111.005 ;
        RECT -26.685 109.315 -26.355 109.645 ;
        RECT -26.685 107.955 -26.355 108.285 ;
        RECT -26.685 106.595 -26.355 106.925 ;
        RECT -26.685 105.235 -26.355 105.565 ;
        RECT -26.685 103.875 -26.355 104.205 ;
        RECT -26.685 102.515 -26.355 102.845 ;
        RECT -26.685 101.155 -26.355 101.485 ;
        RECT -26.685 99.795 -26.355 100.125 ;
        RECT -26.685 98.435 -26.355 98.765 ;
        RECT -26.685 97.075 -26.355 97.405 ;
        RECT -26.685 95.715 -26.355 96.045 ;
        RECT -26.685 94.355 -26.355 94.685 ;
        RECT -26.685 92.995 -26.355 93.325 ;
        RECT -26.685 91.635 -26.355 91.965 ;
        RECT -26.685 90.275 -26.355 90.605 ;
        RECT -26.685 88.915 -26.355 89.245 ;
        RECT -26.685 87.555 -26.355 87.885 ;
        RECT -26.685 86.195 -26.355 86.525 ;
        RECT -26.685 84.835 -26.355 85.165 ;
        RECT -26.685 83.475 -26.355 83.805 ;
        RECT -26.685 82.115 -26.355 82.445 ;
        RECT -26.685 80.755 -26.355 81.085 ;
        RECT -26.685 79.395 -26.355 79.725 ;
        RECT -26.685 78.035 -26.355 78.365 ;
        RECT -26.685 76.675 -26.355 77.005 ;
        RECT -26.685 75.315 -26.355 75.645 ;
        RECT -26.685 73.955 -26.355 74.285 ;
        RECT -26.685 72.595 -26.355 72.925 ;
        RECT -26.685 71.235 -26.355 71.565 ;
        RECT -26.685 69.875 -26.355 70.205 ;
        RECT -26.685 68.515 -26.355 68.845 ;
        RECT -26.685 67.155 -26.355 67.485 ;
        RECT -26.685 65.795 -26.355 66.125 ;
        RECT -26.685 64.435 -26.355 64.765 ;
        RECT -26.685 63.075 -26.355 63.405 ;
        RECT -26.685 61.715 -26.355 62.045 ;
        RECT -26.685 60.355 -26.355 60.685 ;
        RECT -26.685 58.995 -26.355 59.325 ;
        RECT -26.685 57.635 -26.355 57.965 ;
        RECT -26.685 56.275 -26.355 56.605 ;
        RECT -26.685 54.915 -26.355 55.245 ;
        RECT -26.685 53.555 -26.355 53.885 ;
        RECT -26.685 52.195 -26.355 52.525 ;
        RECT -26.685 50.835 -26.355 51.165 ;
        RECT -26.685 49.475 -26.355 49.805 ;
        RECT -26.685 48.115 -26.355 48.445 ;
        RECT -26.685 46.755 -26.355 47.085 ;
        RECT -26.685 45.395 -26.355 45.725 ;
        RECT -26.685 44.035 -26.355 44.365 ;
        RECT -26.685 42.675 -26.355 43.005 ;
        RECT -26.685 41.315 -26.355 41.645 ;
        RECT -26.685 39.955 -26.355 40.285 ;
        RECT -26.685 38.595 -26.355 38.925 ;
        RECT -26.685 37.235 -26.355 37.565 ;
        RECT -26.685 35.875 -26.355 36.205 ;
        RECT -26.685 34.515 -26.355 34.845 ;
        RECT -26.685 33.155 -26.355 33.485 ;
        RECT -26.685 31.795 -26.355 32.125 ;
        RECT -26.685 30.435 -26.355 30.765 ;
        RECT -26.685 29.075 -26.355 29.405 ;
        RECT -26.685 27.715 -26.355 28.045 ;
        RECT -26.685 26.355 -26.355 26.685 ;
        RECT -26.685 24.995 -26.355 25.325 ;
        RECT -26.685 23.635 -26.355 23.965 ;
        RECT -26.685 22.275 -26.355 22.605 ;
        RECT -26.685 20.915 -26.355 21.245 ;
        RECT -26.685 19.555 -26.355 19.885 ;
        RECT -26.685 18.195 -26.355 18.525 ;
        RECT -26.685 16.835 -26.355 17.165 ;
        RECT -26.685 15.475 -26.355 15.805 ;
        RECT -26.685 14.115 -26.355 14.445 ;
        RECT -26.685 12.755 -26.355 13.085 ;
        RECT -26.685 11.395 -26.355 11.725 ;
        RECT -26.685 10.035 -26.355 10.365 ;
        RECT -26.685 8.675 -26.355 9.005 ;
        RECT -26.685 7.315 -26.355 7.645 ;
        RECT -26.685 5.955 -26.355 6.285 ;
        RECT -26.685 4.595 -26.355 4.925 ;
        RECT -26.685 3.235 -26.355 3.565 ;
        RECT -26.685 1.875 -26.355 2.205 ;
        RECT -26.685 0.515 -26.355 0.845 ;
        RECT -26.685 -2.205 -26.355 -1.875 ;
        RECT -26.685 -7.645 -26.355 -7.315 ;
        RECT -26.685 -10.365 -26.355 -10.035 ;
        RECT -26.685 -11.725 -26.355 -11.395 ;
        RECT -26.685 -13.7 -26.355 -13.37 ;
        RECT -26.685 -14.445 -26.355 -14.115 ;
        RECT -26.685 -15.805 -26.355 -15.475 ;
        RECT -26.685 -18.79 -26.355 -18.46 ;
        RECT -26.685 -19.885 -26.355 -19.555 ;
        RECT -26.685 -23.965 -26.355 -23.635 ;
        RECT -26.685 -29.405 -26.355 -29.075 ;
        RECT -26.685 -32.125 -26.355 -31.795 ;
        RECT -26.685 -33.485 -26.355 -33.155 ;
        RECT -26.685 -34.88 -26.355 -34.55 ;
        RECT -26.685 -36.205 -26.355 -35.875 ;
        RECT -26.685 -38.925 -26.355 -38.595 ;
        RECT -26.685 -39.97 -26.355 -39.64 ;
        RECT -26.685 -48.445 -26.355 -48.115 ;
        RECT -26.685 -49.805 -26.355 -49.475 ;
        RECT -26.685 -51.165 -26.355 -50.835 ;
        RECT -26.685 -53.885 -26.355 -53.555 ;
        RECT -26.685 -57.965 -26.355 -57.635 ;
        RECT -26.685 -62.045 -26.355 -61.715 ;
        RECT -26.685 -63.405 -26.355 -63.075 ;
        RECT -26.685 -64.765 -26.355 -64.435 ;
        RECT -26.685 -66.125 -26.355 -65.795 ;
        RECT -26.685 -68.845 -26.355 -68.515 ;
        RECT -26.685 -71.565 -26.355 -71.235 ;
        RECT -26.685 -72.925 -26.355 -72.595 ;
        RECT -26.685 -74.285 -26.355 -73.955 ;
        RECT -26.685 -75.645 -26.355 -75.315 ;
        RECT -26.685 -77.005 -26.355 -76.675 ;
        RECT -26.685 -78.365 -26.355 -78.035 ;
        RECT -26.685 -80.31 -26.355 -79.98 ;
        RECT -26.685 -81.085 -26.355 -80.755 ;
        RECT -26.685 -82.445 -26.355 -82.115 ;
        RECT -26.685 -83.805 -26.355 -83.475 ;
        RECT -26.685 -85.165 -26.355 -84.835 ;
        RECT -26.685 -86.525 -26.355 -86.195 ;
        RECT -26.685 -87.885 -26.355 -87.555 ;
        RECT -26.685 -90.605 -26.355 -90.275 ;
        RECT -26.685 -91.965 -26.355 -91.635 ;
        RECT -26.685 -93.325 -26.355 -92.995 ;
        RECT -26.685 -94.685 -26.355 -94.355 ;
        RECT -26.685 -96.045 -26.355 -95.715 ;
        RECT -26.685 -97.405 -26.355 -97.075 ;
        RECT -26.685 -98.85 -26.355 -98.52 ;
        RECT -26.685 -100.125 -26.355 -99.795 ;
        RECT -26.685 -101.485 -26.355 -101.155 ;
        RECT -26.685 -102.845 -26.355 -102.515 ;
        RECT -26.685 -105.565 -26.355 -105.235 ;
        RECT -26.685 -106.925 -26.355 -106.595 ;
        RECT -26.685 -108.285 -26.355 -107.955 ;
        RECT -26.685 -109.645 -26.355 -109.315 ;
        RECT -26.685 -111.005 -26.355 -110.675 ;
        RECT -26.685 -112.365 -26.355 -112.035 ;
        RECT -26.685 -113.725 -26.355 -113.395 ;
        RECT -26.685 -116.445 -26.355 -116.115 ;
        RECT -26.685 -117.805 -26.355 -117.475 ;
        RECT -26.685 -119.165 -26.355 -118.835 ;
        RECT -26.685 -120.525 -26.355 -120.195 ;
        RECT -26.685 -121.885 -26.355 -121.555 ;
        RECT -26.685 -124.49 -26.355 -124.16 ;
        RECT -26.685 -128.685 -26.355 -128.355 ;
        RECT -26.685 -130.045 -26.355 -129.715 ;
        RECT -26.685 -131.405 -26.355 -131.075 ;
        RECT -26.685 -132.765 -26.355 -132.435 ;
        RECT -26.685 -136.845 -26.355 -136.515 ;
        RECT -26.685 -138.205 -26.355 -137.875 ;
        RECT -26.685 -139.565 -26.355 -139.235 ;
        RECT -26.685 -140.925 -26.355 -140.595 ;
        RECT -26.685 -142.285 -26.355 -141.955 ;
        RECT -26.685 -143.03 -26.355 -142.7 ;
        RECT -26.685 -145.005 -26.355 -144.675 ;
        RECT -26.685 -146.365 -26.355 -146.035 ;
        RECT -26.685 -147.725 -26.355 -147.395 ;
        RECT -26.685 -153.165 -26.355 -152.835 ;
        RECT -26.685 -154.525 -26.355 -154.195 ;
        RECT -26.685 -155.885 -26.355 -155.555 ;
        RECT -26.685 -157.245 -26.355 -156.915 ;
        RECT -26.685 -162.685 -26.355 -162.355 ;
        RECT -26.685 -164.045 -26.355 -163.715 ;
        RECT -26.685 -165.405 -26.355 -165.075 ;
        RECT -26.685 -166.765 -26.355 -166.435 ;
        RECT -26.685 -168.125 -26.355 -167.795 ;
        RECT -26.685 -169.485 -26.355 -169.155 ;
        RECT -26.685 -170.845 -26.355 -170.515 ;
        RECT -26.685 -172.205 -26.355 -171.875 ;
        RECT -26.685 -173.565 -26.355 -173.235 ;
        RECT -26.685 -174.925 -26.355 -174.595 ;
        RECT -26.685 -176.285 -26.355 -175.955 ;
        RECT -26.685 -177.645 -26.355 -177.315 ;
        RECT -26.685 -179.005 -26.355 -178.675 ;
        RECT -26.685 -180.365 -26.355 -180.035 ;
        RECT -26.685 -181.725 -26.355 -181.395 ;
        RECT -26.685 -183.085 -26.355 -182.755 ;
        RECT -26.685 -185.805 -26.355 -185.475 ;
        RECT -26.685 -187.165 -26.355 -186.835 ;
        RECT -26.685 -192.605 -26.355 -192.275 ;
        RECT -26.685 -193.965 -26.355 -193.635 ;
        RECT -26.685 -195.325 -26.355 -194.995 ;
        RECT -26.685 -198.045 -26.355 -197.715 ;
        RECT -26.685 -199.405 -26.355 -199.075 ;
        RECT -26.685 -200.765 -26.355 -200.435 ;
        RECT -26.685 -202.125 -26.355 -201.795 ;
        RECT -26.685 -204.845 -26.355 -204.515 ;
        RECT -26.685 -206.205 -26.355 -205.875 ;
        RECT -26.685 -208.925 -26.355 -208.595 ;
        RECT -26.685 -210.285 -26.355 -209.955 ;
        RECT -26.685 -215.725 -26.355 -215.395 ;
        RECT -26.685 -217.085 -26.355 -216.755 ;
        RECT -26.685 -218.445 -26.355 -218.115 ;
        RECT -26.685 -219.805 -26.355 -219.475 ;
        RECT -26.685 -221.165 -26.355 -220.835 ;
        RECT -26.685 -222.525 -26.355 -222.195 ;
        RECT -26.685 -223.885 -26.355 -223.555 ;
        RECT -26.685 -225.245 -26.355 -224.915 ;
        RECT -26.685 -230.685 -26.355 -230.355 ;
        RECT -26.685 -232.045 -26.355 -231.715 ;
        RECT -26.685 -233.225 -26.355 -232.895 ;
        RECT -26.685 -234.765 -26.355 -234.435 ;
        RECT -26.685 -236.125 -26.355 -235.795 ;
        RECT -26.685 -237.485 -26.355 -237.155 ;
        RECT -26.685 -238.845 -26.355 -238.515 ;
        RECT -26.685 -241.09 -26.355 -239.96 ;
        RECT -26.68 -241.205 -26.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.325 196.355 -24.995 196.685 ;
        RECT -25.325 194.995 -24.995 195.325 ;
        RECT -25.325 193.635 -24.995 193.965 ;
        RECT -25.325 192.275 -24.995 192.605 ;
        RECT -25.325 190.915 -24.995 191.245 ;
        RECT -25.325 189.555 -24.995 189.885 ;
        RECT -25.325 188.195 -24.995 188.525 ;
        RECT -25.325 186.835 -24.995 187.165 ;
        RECT -25.325 185.475 -24.995 185.805 ;
        RECT -25.325 184.115 -24.995 184.445 ;
        RECT -25.325 182.755 -24.995 183.085 ;
        RECT -25.325 181.395 -24.995 181.725 ;
        RECT -25.325 180.035 -24.995 180.365 ;
        RECT -25.325 178.675 -24.995 179.005 ;
        RECT -25.325 177.315 -24.995 177.645 ;
        RECT -25.325 175.955 -24.995 176.285 ;
        RECT -25.325 174.595 -24.995 174.925 ;
        RECT -25.325 173.235 -24.995 173.565 ;
        RECT -25.325 171.875 -24.995 172.205 ;
        RECT -25.325 170.515 -24.995 170.845 ;
        RECT -25.325 169.155 -24.995 169.485 ;
        RECT -25.325 167.795 -24.995 168.125 ;
        RECT -25.325 166.435 -24.995 166.765 ;
        RECT -25.325 165.075 -24.995 165.405 ;
        RECT -25.325 163.715 -24.995 164.045 ;
        RECT -25.325 162.355 -24.995 162.685 ;
        RECT -25.325 160.995 -24.995 161.325 ;
        RECT -25.325 159.635 -24.995 159.965 ;
        RECT -25.325 158.275 -24.995 158.605 ;
        RECT -25.325 156.915 -24.995 157.245 ;
        RECT -25.325 155.555 -24.995 155.885 ;
        RECT -25.325 154.195 -24.995 154.525 ;
        RECT -25.325 152.835 -24.995 153.165 ;
        RECT -25.325 151.475 -24.995 151.805 ;
        RECT -25.325 150.115 -24.995 150.445 ;
        RECT -25.325 148.755 -24.995 149.085 ;
        RECT -25.325 147.395 -24.995 147.725 ;
        RECT -25.325 146.035 -24.995 146.365 ;
        RECT -25.325 144.675 -24.995 145.005 ;
        RECT -25.325 143.315 -24.995 143.645 ;
        RECT -25.325 141.955 -24.995 142.285 ;
        RECT -25.325 140.595 -24.995 140.925 ;
        RECT -25.325 139.235 -24.995 139.565 ;
        RECT -25.325 137.875 -24.995 138.205 ;
        RECT -25.325 136.515 -24.995 136.845 ;
        RECT -25.325 135.155 -24.995 135.485 ;
        RECT -25.325 133.795 -24.995 134.125 ;
        RECT -25.325 132.435 -24.995 132.765 ;
        RECT -25.325 131.075 -24.995 131.405 ;
        RECT -25.325 129.715 -24.995 130.045 ;
        RECT -25.325 128.355 -24.995 128.685 ;
        RECT -25.325 126.995 -24.995 127.325 ;
        RECT -25.325 125.635 -24.995 125.965 ;
        RECT -25.325 124.275 -24.995 124.605 ;
        RECT -25.325 122.915 -24.995 123.245 ;
        RECT -25.325 121.555 -24.995 121.885 ;
        RECT -25.325 120.195 -24.995 120.525 ;
        RECT -25.325 118.835 -24.995 119.165 ;
        RECT -25.325 117.475 -24.995 117.805 ;
        RECT -25.325 116.115 -24.995 116.445 ;
        RECT -25.325 114.755 -24.995 115.085 ;
        RECT -25.325 113.395 -24.995 113.725 ;
        RECT -25.325 112.035 -24.995 112.365 ;
        RECT -25.325 110.675 -24.995 111.005 ;
        RECT -25.325 109.315 -24.995 109.645 ;
        RECT -25.325 107.955 -24.995 108.285 ;
        RECT -25.325 106.595 -24.995 106.925 ;
        RECT -25.325 105.235 -24.995 105.565 ;
        RECT -25.325 103.875 -24.995 104.205 ;
        RECT -25.325 102.515 -24.995 102.845 ;
        RECT -25.325 101.155 -24.995 101.485 ;
        RECT -25.325 99.795 -24.995 100.125 ;
        RECT -25.325 98.435 -24.995 98.765 ;
        RECT -25.325 97.075 -24.995 97.405 ;
        RECT -25.325 95.715 -24.995 96.045 ;
        RECT -25.325 94.355 -24.995 94.685 ;
        RECT -25.325 92.995 -24.995 93.325 ;
        RECT -25.325 91.635 -24.995 91.965 ;
        RECT -25.325 90.275 -24.995 90.605 ;
        RECT -25.325 88.915 -24.995 89.245 ;
        RECT -25.325 87.555 -24.995 87.885 ;
        RECT -25.325 86.195 -24.995 86.525 ;
        RECT -25.325 84.835 -24.995 85.165 ;
        RECT -25.325 83.475 -24.995 83.805 ;
        RECT -25.325 82.115 -24.995 82.445 ;
        RECT -25.325 80.755 -24.995 81.085 ;
        RECT -25.325 79.395 -24.995 79.725 ;
        RECT -25.325 78.035 -24.995 78.365 ;
        RECT -25.325 76.675 -24.995 77.005 ;
        RECT -25.325 75.315 -24.995 75.645 ;
        RECT -25.325 73.955 -24.995 74.285 ;
        RECT -25.325 72.595 -24.995 72.925 ;
        RECT -25.325 71.235 -24.995 71.565 ;
        RECT -25.325 69.875 -24.995 70.205 ;
        RECT -25.325 68.515 -24.995 68.845 ;
        RECT -25.325 67.155 -24.995 67.485 ;
        RECT -25.325 65.795 -24.995 66.125 ;
        RECT -25.325 64.435 -24.995 64.765 ;
        RECT -25.325 63.075 -24.995 63.405 ;
        RECT -25.325 61.715 -24.995 62.045 ;
        RECT -25.325 60.355 -24.995 60.685 ;
        RECT -25.325 58.995 -24.995 59.325 ;
        RECT -25.325 57.635 -24.995 57.965 ;
        RECT -25.325 56.275 -24.995 56.605 ;
        RECT -25.325 54.915 -24.995 55.245 ;
        RECT -25.325 53.555 -24.995 53.885 ;
        RECT -25.325 52.195 -24.995 52.525 ;
        RECT -25.325 50.835 -24.995 51.165 ;
        RECT -25.325 49.475 -24.995 49.805 ;
        RECT -25.325 48.115 -24.995 48.445 ;
        RECT -25.325 46.755 -24.995 47.085 ;
        RECT -25.325 45.395 -24.995 45.725 ;
        RECT -25.325 44.035 -24.995 44.365 ;
        RECT -25.325 42.675 -24.995 43.005 ;
        RECT -25.325 41.315 -24.995 41.645 ;
        RECT -25.325 39.955 -24.995 40.285 ;
        RECT -25.325 38.595 -24.995 38.925 ;
        RECT -25.325 37.235 -24.995 37.565 ;
        RECT -25.325 35.875 -24.995 36.205 ;
        RECT -25.325 34.515 -24.995 34.845 ;
        RECT -25.325 33.155 -24.995 33.485 ;
        RECT -25.325 31.795 -24.995 32.125 ;
        RECT -25.325 30.435 -24.995 30.765 ;
        RECT -25.325 29.075 -24.995 29.405 ;
        RECT -25.325 27.715 -24.995 28.045 ;
        RECT -25.325 26.355 -24.995 26.685 ;
        RECT -25.325 24.995 -24.995 25.325 ;
        RECT -25.325 23.635 -24.995 23.965 ;
        RECT -25.325 22.275 -24.995 22.605 ;
        RECT -25.325 20.915 -24.995 21.245 ;
        RECT -25.325 19.555 -24.995 19.885 ;
        RECT -25.325 18.195 -24.995 18.525 ;
        RECT -25.325 16.835 -24.995 17.165 ;
        RECT -25.325 15.475 -24.995 15.805 ;
        RECT -25.325 14.115 -24.995 14.445 ;
        RECT -25.325 12.755 -24.995 13.085 ;
        RECT -25.325 11.395 -24.995 11.725 ;
        RECT -25.325 10.035 -24.995 10.365 ;
        RECT -25.325 8.675 -24.995 9.005 ;
        RECT -25.325 7.315 -24.995 7.645 ;
        RECT -25.325 5.955 -24.995 6.285 ;
        RECT -25.325 4.595 -24.995 4.925 ;
        RECT -25.325 3.235 -24.995 3.565 ;
        RECT -25.325 1.875 -24.995 2.205 ;
        RECT -25.325 0.515 -24.995 0.845 ;
        RECT -25.325 -2.205 -24.995 -1.875 ;
        RECT -25.325 -7.645 -24.995 -7.315 ;
        RECT -25.325 -10.365 -24.995 -10.035 ;
        RECT -25.325 -11.725 -24.995 -11.395 ;
        RECT -25.325 -13.7 -24.995 -13.37 ;
        RECT -25.325 -14.445 -24.995 -14.115 ;
        RECT -25.325 -15.805 -24.995 -15.475 ;
        RECT -25.325 -18.79 -24.995 -18.46 ;
        RECT -25.325 -19.885 -24.995 -19.555 ;
        RECT -25.325 -23.965 -24.995 -23.635 ;
        RECT -25.325 -29.405 -24.995 -29.075 ;
        RECT -25.325 -32.125 -24.995 -31.795 ;
        RECT -25.325 -33.485 -24.995 -33.155 ;
        RECT -25.325 -34.88 -24.995 -34.55 ;
        RECT -25.325 -36.205 -24.995 -35.875 ;
        RECT -25.325 -38.925 -24.995 -38.595 ;
        RECT -25.325 -39.97 -24.995 -39.64 ;
        RECT -25.325 -48.445 -24.995 -48.115 ;
        RECT -25.325 -49.805 -24.995 -49.475 ;
        RECT -25.325 -51.165 -24.995 -50.835 ;
        RECT -25.325 -53.885 -24.995 -53.555 ;
        RECT -25.325 -57.965 -24.995 -57.635 ;
        RECT -25.325 -62.045 -24.995 -61.715 ;
        RECT -25.325 -63.405 -24.995 -63.075 ;
        RECT -25.325 -64.765 -24.995 -64.435 ;
        RECT -25.325 -66.125 -24.995 -65.795 ;
        RECT -25.325 -68.845 -24.995 -68.515 ;
        RECT -25.325 -71.565 -24.995 -71.235 ;
        RECT -25.325 -72.925 -24.995 -72.595 ;
        RECT -25.325 -74.285 -24.995 -73.955 ;
        RECT -25.325 -75.645 -24.995 -75.315 ;
        RECT -25.325 -77.005 -24.995 -76.675 ;
        RECT -25.325 -78.365 -24.995 -78.035 ;
        RECT -25.325 -80.31 -24.995 -79.98 ;
        RECT -25.325 -81.085 -24.995 -80.755 ;
        RECT -25.325 -82.445 -24.995 -82.115 ;
        RECT -25.325 -83.805 -24.995 -83.475 ;
        RECT -25.325 -85.165 -24.995 -84.835 ;
        RECT -25.325 -86.525 -24.995 -86.195 ;
        RECT -25.325 -87.885 -24.995 -87.555 ;
        RECT -25.325 -90.605 -24.995 -90.275 ;
        RECT -25.325 -91.965 -24.995 -91.635 ;
        RECT -25.325 -93.325 -24.995 -92.995 ;
        RECT -25.325 -94.685 -24.995 -94.355 ;
        RECT -25.325 -96.045 -24.995 -95.715 ;
        RECT -25.325 -97.405 -24.995 -97.075 ;
        RECT -25.325 -98.85 -24.995 -98.52 ;
        RECT -25.325 -100.125 -24.995 -99.795 ;
        RECT -25.325 -101.485 -24.995 -101.155 ;
        RECT -25.325 -102.845 -24.995 -102.515 ;
        RECT -25.325 -105.565 -24.995 -105.235 ;
        RECT -25.325 -106.925 -24.995 -106.595 ;
        RECT -25.325 -108.285 -24.995 -107.955 ;
        RECT -25.325 -109.645 -24.995 -109.315 ;
        RECT -25.325 -111.005 -24.995 -110.675 ;
        RECT -25.325 -112.365 -24.995 -112.035 ;
        RECT -25.325 -113.725 -24.995 -113.395 ;
        RECT -25.325 -116.445 -24.995 -116.115 ;
        RECT -25.325 -117.805 -24.995 -117.475 ;
        RECT -25.325 -119.165 -24.995 -118.835 ;
        RECT -25.325 -120.525 -24.995 -120.195 ;
        RECT -25.325 -121.885 -24.995 -121.555 ;
        RECT -25.325 -124.49 -24.995 -124.16 ;
        RECT -25.325 -128.685 -24.995 -128.355 ;
        RECT -25.325 -130.045 -24.995 -129.715 ;
        RECT -25.325 -131.405 -24.995 -131.075 ;
        RECT -25.325 -132.765 -24.995 -132.435 ;
        RECT -25.325 -136.845 -24.995 -136.515 ;
        RECT -25.325 -138.205 -24.995 -137.875 ;
        RECT -25.325 -139.565 -24.995 -139.235 ;
        RECT -25.325 -140.925 -24.995 -140.595 ;
        RECT -25.325 -142.285 -24.995 -141.955 ;
        RECT -25.325 -143.03 -24.995 -142.7 ;
        RECT -25.325 -145.005 -24.995 -144.675 ;
        RECT -25.325 -146.365 -24.995 -146.035 ;
        RECT -25.325 -147.725 -24.995 -147.395 ;
        RECT -25.325 -153.165 -24.995 -152.835 ;
        RECT -25.325 -154.525 -24.995 -154.195 ;
        RECT -25.325 -155.885 -24.995 -155.555 ;
        RECT -25.325 -157.245 -24.995 -156.915 ;
        RECT -25.325 -162.685 -24.995 -162.355 ;
        RECT -25.325 -164.045 -24.995 -163.715 ;
        RECT -25.325 -165.405 -24.995 -165.075 ;
        RECT -25.325 -166.765 -24.995 -166.435 ;
        RECT -25.325 -168.125 -24.995 -167.795 ;
        RECT -25.325 -169.485 -24.995 -169.155 ;
        RECT -25.325 -170.845 -24.995 -170.515 ;
        RECT -25.325 -172.205 -24.995 -171.875 ;
        RECT -25.325 -173.565 -24.995 -173.235 ;
        RECT -25.325 -174.925 -24.995 -174.595 ;
        RECT -25.325 -176.285 -24.995 -175.955 ;
        RECT -25.325 -177.645 -24.995 -177.315 ;
        RECT -25.325 -179.005 -24.995 -178.675 ;
        RECT -25.325 -180.365 -24.995 -180.035 ;
        RECT -25.325 -181.725 -24.995 -181.395 ;
        RECT -25.325 -183.085 -24.995 -182.755 ;
        RECT -25.325 -185.805 -24.995 -185.475 ;
        RECT -25.325 -187.165 -24.995 -186.835 ;
        RECT -25.325 -192.605 -24.995 -192.275 ;
        RECT -25.325 -193.965 -24.995 -193.635 ;
        RECT -25.325 -195.325 -24.995 -194.995 ;
        RECT -25.325 -198.045 -24.995 -197.715 ;
        RECT -25.325 -199.405 -24.995 -199.075 ;
        RECT -25.325 -200.765 -24.995 -200.435 ;
        RECT -25.325 -202.125 -24.995 -201.795 ;
        RECT -25.325 -204.845 -24.995 -204.515 ;
        RECT -25.325 -206.205 -24.995 -205.875 ;
        RECT -25.325 -208.925 -24.995 -208.595 ;
        RECT -25.325 -210.285 -24.995 -209.955 ;
        RECT -25.325 -215.725 -24.995 -215.395 ;
        RECT -25.325 -217.085 -24.995 -216.755 ;
        RECT -25.325 -218.445 -24.995 -218.115 ;
        RECT -25.325 -219.805 -24.995 -219.475 ;
        RECT -25.325 -221.165 -24.995 -220.835 ;
        RECT -25.325 -222.525 -24.995 -222.195 ;
        RECT -25.325 -223.885 -24.995 -223.555 ;
        RECT -25.325 -225.245 -24.995 -224.915 ;
        RECT -25.325 -230.685 -24.995 -230.355 ;
        RECT -25.325 -232.045 -24.995 -231.715 ;
        RECT -25.325 -233.225 -24.995 -232.895 ;
        RECT -25.325 -234.765 -24.995 -234.435 ;
        RECT -25.325 -236.125 -24.995 -235.795 ;
        RECT -25.325 -237.485 -24.995 -237.155 ;
        RECT -25.325 -238.845 -24.995 -238.515 ;
        RECT -25.325 -241.09 -24.995 -239.96 ;
        RECT -25.32 -241.205 -25 245.285 ;
        RECT -25.325 244.04 -24.995 245.17 ;
        RECT -25.325 242.595 -24.995 242.925 ;
        RECT -25.325 241.235 -24.995 241.565 ;
        RECT -25.325 239.875 -24.995 240.205 ;
        RECT -25.325 238.515 -24.995 238.845 ;
        RECT -25.325 237.155 -24.995 237.485 ;
        RECT -25.325 235.795 -24.995 236.125 ;
        RECT -25.325 234.435 -24.995 234.765 ;
        RECT -25.325 233.075 -24.995 233.405 ;
        RECT -25.325 231.715 -24.995 232.045 ;
        RECT -25.325 230.355 -24.995 230.685 ;
        RECT -25.325 228.995 -24.995 229.325 ;
        RECT -25.325 227.635 -24.995 227.965 ;
        RECT -25.325 226.275 -24.995 226.605 ;
        RECT -25.325 224.915 -24.995 225.245 ;
        RECT -25.325 223.555 -24.995 223.885 ;
        RECT -25.325 222.195 -24.995 222.525 ;
        RECT -25.325 220.835 -24.995 221.165 ;
        RECT -25.325 219.475 -24.995 219.805 ;
        RECT -25.325 218.115 -24.995 218.445 ;
        RECT -25.325 216.755 -24.995 217.085 ;
        RECT -25.325 215.395 -24.995 215.725 ;
        RECT -25.325 214.035 -24.995 214.365 ;
        RECT -25.325 212.675 -24.995 213.005 ;
        RECT -25.325 211.315 -24.995 211.645 ;
        RECT -25.325 209.955 -24.995 210.285 ;
        RECT -25.325 208.595 -24.995 208.925 ;
        RECT -25.325 207.235 -24.995 207.565 ;
        RECT -25.325 205.875 -24.995 206.205 ;
        RECT -25.325 204.515 -24.995 204.845 ;
        RECT -25.325 203.155 -24.995 203.485 ;
        RECT -25.325 201.795 -24.995 202.125 ;
        RECT -25.325 200.435 -24.995 200.765 ;
        RECT -25.325 199.075 -24.995 199.405 ;
        RECT -25.325 197.715 -24.995 198.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.125 244.04 -31.795 245.17 ;
        RECT -32.125 242.595 -31.795 242.925 ;
        RECT -32.125 241.235 -31.795 241.565 ;
        RECT -32.125 239.875 -31.795 240.205 ;
        RECT -32.125 238.515 -31.795 238.845 ;
        RECT -32.125 237.155 -31.795 237.485 ;
        RECT -32.125 235.795 -31.795 236.125 ;
        RECT -32.125 234.435 -31.795 234.765 ;
        RECT -32.125 233.075 -31.795 233.405 ;
        RECT -32.125 231.715 -31.795 232.045 ;
        RECT -32.125 230.355 -31.795 230.685 ;
        RECT -32.125 228.995 -31.795 229.325 ;
        RECT -32.125 227.635 -31.795 227.965 ;
        RECT -32.125 226.275 -31.795 226.605 ;
        RECT -32.125 224.915 -31.795 225.245 ;
        RECT -32.125 223.555 -31.795 223.885 ;
        RECT -32.125 222.195 -31.795 222.525 ;
        RECT -32.125 220.835 -31.795 221.165 ;
        RECT -32.125 219.475 -31.795 219.805 ;
        RECT -32.125 218.115 -31.795 218.445 ;
        RECT -32.125 216.755 -31.795 217.085 ;
        RECT -32.125 215.395 -31.795 215.725 ;
        RECT -32.125 214.035 -31.795 214.365 ;
        RECT -32.125 212.675 -31.795 213.005 ;
        RECT -32.125 211.315 -31.795 211.645 ;
        RECT -32.125 209.955 -31.795 210.285 ;
        RECT -32.125 208.595 -31.795 208.925 ;
        RECT -32.125 207.235 -31.795 207.565 ;
        RECT -32.125 205.875 -31.795 206.205 ;
        RECT -32.125 204.515 -31.795 204.845 ;
        RECT -32.125 203.155 -31.795 203.485 ;
        RECT -32.125 201.795 -31.795 202.125 ;
        RECT -32.125 200.435 -31.795 200.765 ;
        RECT -32.125 199.075 -31.795 199.405 ;
        RECT -32.125 197.715 -31.795 198.045 ;
        RECT -32.125 196.355 -31.795 196.685 ;
        RECT -32.125 194.995 -31.795 195.325 ;
        RECT -32.125 193.635 -31.795 193.965 ;
        RECT -32.125 192.275 -31.795 192.605 ;
        RECT -32.125 190.915 -31.795 191.245 ;
        RECT -32.125 189.555 -31.795 189.885 ;
        RECT -32.125 188.195 -31.795 188.525 ;
        RECT -32.125 186.835 -31.795 187.165 ;
        RECT -32.125 185.475 -31.795 185.805 ;
        RECT -32.125 184.115 -31.795 184.445 ;
        RECT -32.125 182.755 -31.795 183.085 ;
        RECT -32.125 181.395 -31.795 181.725 ;
        RECT -32.125 180.035 -31.795 180.365 ;
        RECT -32.125 178.675 -31.795 179.005 ;
        RECT -32.125 177.315 -31.795 177.645 ;
        RECT -32.125 175.955 -31.795 176.285 ;
        RECT -32.125 174.595 -31.795 174.925 ;
        RECT -32.125 173.235 -31.795 173.565 ;
        RECT -32.125 171.875 -31.795 172.205 ;
        RECT -32.125 170.515 -31.795 170.845 ;
        RECT -32.125 169.155 -31.795 169.485 ;
        RECT -32.125 167.795 -31.795 168.125 ;
        RECT -32.125 166.435 -31.795 166.765 ;
        RECT -32.125 165.075 -31.795 165.405 ;
        RECT -32.125 163.715 -31.795 164.045 ;
        RECT -32.125 162.355 -31.795 162.685 ;
        RECT -32.125 160.995 -31.795 161.325 ;
        RECT -32.125 159.635 -31.795 159.965 ;
        RECT -32.125 158.275 -31.795 158.605 ;
        RECT -32.125 156.915 -31.795 157.245 ;
        RECT -32.125 155.555 -31.795 155.885 ;
        RECT -32.125 154.195 -31.795 154.525 ;
        RECT -32.125 152.835 -31.795 153.165 ;
        RECT -32.125 151.475 -31.795 151.805 ;
        RECT -32.125 150.115 -31.795 150.445 ;
        RECT -32.125 148.755 -31.795 149.085 ;
        RECT -32.125 147.395 -31.795 147.725 ;
        RECT -32.125 146.035 -31.795 146.365 ;
        RECT -32.125 144.675 -31.795 145.005 ;
        RECT -32.125 143.315 -31.795 143.645 ;
        RECT -32.125 141.955 -31.795 142.285 ;
        RECT -32.125 140.595 -31.795 140.925 ;
        RECT -32.125 139.235 -31.795 139.565 ;
        RECT -32.125 137.875 -31.795 138.205 ;
        RECT -32.125 136.515 -31.795 136.845 ;
        RECT -32.125 135.155 -31.795 135.485 ;
        RECT -32.125 133.795 -31.795 134.125 ;
        RECT -32.125 132.435 -31.795 132.765 ;
        RECT -32.125 131.075 -31.795 131.405 ;
        RECT -32.125 129.715 -31.795 130.045 ;
        RECT -32.125 128.355 -31.795 128.685 ;
        RECT -32.125 126.995 -31.795 127.325 ;
        RECT -32.125 125.635 -31.795 125.965 ;
        RECT -32.125 124.275 -31.795 124.605 ;
        RECT -32.125 122.915 -31.795 123.245 ;
        RECT -32.125 121.555 -31.795 121.885 ;
        RECT -32.125 120.195 -31.795 120.525 ;
        RECT -32.125 118.835 -31.795 119.165 ;
        RECT -32.125 117.475 -31.795 117.805 ;
        RECT -32.125 116.115 -31.795 116.445 ;
        RECT -32.125 114.755 -31.795 115.085 ;
        RECT -32.125 113.395 -31.795 113.725 ;
        RECT -32.125 112.035 -31.795 112.365 ;
        RECT -32.125 110.675 -31.795 111.005 ;
        RECT -32.125 109.315 -31.795 109.645 ;
        RECT -32.125 107.955 -31.795 108.285 ;
        RECT -32.125 106.595 -31.795 106.925 ;
        RECT -32.125 105.235 -31.795 105.565 ;
        RECT -32.125 103.875 -31.795 104.205 ;
        RECT -32.125 102.515 -31.795 102.845 ;
        RECT -32.125 101.155 -31.795 101.485 ;
        RECT -32.125 99.795 -31.795 100.125 ;
        RECT -32.125 98.435 -31.795 98.765 ;
        RECT -32.125 97.075 -31.795 97.405 ;
        RECT -32.125 95.715 -31.795 96.045 ;
        RECT -32.125 94.355 -31.795 94.685 ;
        RECT -32.125 92.995 -31.795 93.325 ;
        RECT -32.125 91.635 -31.795 91.965 ;
        RECT -32.125 90.275 -31.795 90.605 ;
        RECT -32.125 88.915 -31.795 89.245 ;
        RECT -32.125 87.555 -31.795 87.885 ;
        RECT -32.125 86.195 -31.795 86.525 ;
        RECT -32.125 84.835 -31.795 85.165 ;
        RECT -32.125 83.475 -31.795 83.805 ;
        RECT -32.125 82.115 -31.795 82.445 ;
        RECT -32.125 80.755 -31.795 81.085 ;
        RECT -32.125 79.395 -31.795 79.725 ;
        RECT -32.125 78.035 -31.795 78.365 ;
        RECT -32.125 76.675 -31.795 77.005 ;
        RECT -32.125 75.315 -31.795 75.645 ;
        RECT -32.125 73.955 -31.795 74.285 ;
        RECT -32.125 72.595 -31.795 72.925 ;
        RECT -32.125 71.235 -31.795 71.565 ;
        RECT -32.125 69.875 -31.795 70.205 ;
        RECT -32.125 68.515 -31.795 68.845 ;
        RECT -32.125 67.155 -31.795 67.485 ;
        RECT -32.125 65.795 -31.795 66.125 ;
        RECT -32.125 64.435 -31.795 64.765 ;
        RECT -32.125 63.075 -31.795 63.405 ;
        RECT -32.125 61.715 -31.795 62.045 ;
        RECT -32.125 60.355 -31.795 60.685 ;
        RECT -32.125 58.995 -31.795 59.325 ;
        RECT -32.125 57.635 -31.795 57.965 ;
        RECT -32.125 56.275 -31.795 56.605 ;
        RECT -32.125 54.915 -31.795 55.245 ;
        RECT -32.125 53.555 -31.795 53.885 ;
        RECT -32.125 52.195 -31.795 52.525 ;
        RECT -32.125 50.835 -31.795 51.165 ;
        RECT -32.125 49.475 -31.795 49.805 ;
        RECT -32.125 48.115 -31.795 48.445 ;
        RECT -32.125 46.755 -31.795 47.085 ;
        RECT -32.125 45.395 -31.795 45.725 ;
        RECT -32.125 44.035 -31.795 44.365 ;
        RECT -32.125 42.675 -31.795 43.005 ;
        RECT -32.125 41.315 -31.795 41.645 ;
        RECT -32.125 39.955 -31.795 40.285 ;
        RECT -32.125 38.595 -31.795 38.925 ;
        RECT -32.125 37.235 -31.795 37.565 ;
        RECT -32.125 35.875 -31.795 36.205 ;
        RECT -32.125 34.515 -31.795 34.845 ;
        RECT -32.125 33.155 -31.795 33.485 ;
        RECT -32.125 31.795 -31.795 32.125 ;
        RECT -32.125 30.435 -31.795 30.765 ;
        RECT -32.125 29.075 -31.795 29.405 ;
        RECT -32.125 27.715 -31.795 28.045 ;
        RECT -32.125 26.355 -31.795 26.685 ;
        RECT -32.125 24.995 -31.795 25.325 ;
        RECT -32.125 23.635 -31.795 23.965 ;
        RECT -32.125 22.275 -31.795 22.605 ;
        RECT -32.125 20.915 -31.795 21.245 ;
        RECT -32.125 19.555 -31.795 19.885 ;
        RECT -32.125 18.195 -31.795 18.525 ;
        RECT -32.125 16.835 -31.795 17.165 ;
        RECT -32.125 15.475 -31.795 15.805 ;
        RECT -32.125 14.115 -31.795 14.445 ;
        RECT -32.125 12.755 -31.795 13.085 ;
        RECT -32.125 11.395 -31.795 11.725 ;
        RECT -32.125 10.035 -31.795 10.365 ;
        RECT -32.125 8.675 -31.795 9.005 ;
        RECT -32.125 7.315 -31.795 7.645 ;
        RECT -32.125 5.955 -31.795 6.285 ;
        RECT -32.125 4.595 -31.795 4.925 ;
        RECT -32.125 3.235 -31.795 3.565 ;
        RECT -32.125 1.875 -31.795 2.205 ;
        RECT -32.125 0.515 -31.795 0.845 ;
        RECT -32.125 -7.645 -31.795 -7.315 ;
        RECT -32.125 -9.005 -31.795 -8.675 ;
        RECT -32.125 -10.365 -31.795 -10.035 ;
        RECT -32.125 -11.725 -31.795 -11.395 ;
        RECT -32.125 -13.085 -31.795 -12.755 ;
        RECT -32.125 -14.445 -31.795 -14.115 ;
        RECT -32.125 -15.805 -31.795 -15.475 ;
        RECT -32.125 -17.165 -31.795 -16.835 ;
        RECT -32.125 -18.525 -31.795 -18.195 ;
        RECT -32.125 -19.885 -31.795 -19.555 ;
        RECT -32.125 -21.245 -31.795 -20.915 ;
        RECT -32.125 -22.605 -31.795 -22.275 ;
        RECT -32.125 -29.405 -31.795 -29.075 ;
        RECT -32.125 -32.125 -31.795 -31.795 ;
        RECT -32.125 -33.485 -31.795 -33.155 ;
        RECT -32.125 -34.88 -31.795 -34.55 ;
        RECT -32.125 -36.205 -31.795 -35.875 ;
        RECT -32.125 -38.925 -31.795 -38.595 ;
        RECT -32.125 -39.97 -31.795 -39.64 ;
        RECT -32.125 -48.445 -31.795 -48.115 ;
        RECT -32.125 -49.805 -31.795 -49.475 ;
        RECT -32.125 -51.165 -31.795 -50.835 ;
        RECT -32.125 -53.885 -31.795 -53.555 ;
        RECT -32.125 -57.965 -31.795 -57.635 ;
        RECT -32.125 -62.045 -31.795 -61.715 ;
        RECT -32.125 -63.405 -31.795 -63.075 ;
        RECT -32.125 -64.765 -31.795 -64.435 ;
        RECT -32.125 -66.125 -31.795 -65.795 ;
        RECT -32.125 -67.485 -31.795 -67.155 ;
        RECT -32.125 -68.845 -31.795 -68.515 ;
        RECT -32.125 -70.205 -31.795 -69.875 ;
        RECT -32.125 -71.565 -31.795 -71.235 ;
        RECT -32.125 -72.925 -31.795 -72.595 ;
        RECT -32.125 -74.285 -31.795 -73.955 ;
        RECT -32.125 -75.645 -31.795 -75.315 ;
        RECT -32.125 -77.005 -31.795 -76.675 ;
        RECT -32.125 -78.365 -31.795 -78.035 ;
        RECT -32.125 -79.725 -31.795 -79.395 ;
        RECT -32.125 -81.085 -31.795 -80.755 ;
        RECT -32.125 -82.445 -31.795 -82.115 ;
        RECT -32.125 -83.805 -31.795 -83.475 ;
        RECT -32.125 -85.165 -31.795 -84.835 ;
        RECT -32.125 -86.525 -31.795 -86.195 ;
        RECT -32.125 -87.885 -31.795 -87.555 ;
        RECT -32.125 -89.245 -31.795 -88.915 ;
        RECT -32.125 -90.605 -31.795 -90.275 ;
        RECT -32.125 -91.965 -31.795 -91.635 ;
        RECT -32.125 -93.325 -31.795 -92.995 ;
        RECT -32.125 -94.685 -31.795 -94.355 ;
        RECT -32.125 -96.045 -31.795 -95.715 ;
        RECT -32.125 -97.405 -31.795 -97.075 ;
        RECT -32.125 -98.765 -31.795 -98.435 ;
        RECT -32.125 -100.125 -31.795 -99.795 ;
        RECT -32.125 -101.485 -31.795 -101.155 ;
        RECT -32.125 -102.845 -31.795 -102.515 ;
        RECT -32.125 -104.205 -31.795 -103.875 ;
        RECT -32.125 -105.565 -31.795 -105.235 ;
        RECT -32.125 -106.925 -31.795 -106.595 ;
        RECT -32.125 -108.285 -31.795 -107.955 ;
        RECT -32.125 -109.645 -31.795 -109.315 ;
        RECT -32.125 -111.005 -31.795 -110.675 ;
        RECT -32.125 -112.365 -31.795 -112.035 ;
        RECT -32.125 -113.725 -31.795 -113.395 ;
        RECT -32.125 -115.085 -31.795 -114.755 ;
        RECT -32.125 -116.445 -31.795 -116.115 ;
        RECT -32.125 -117.805 -31.795 -117.475 ;
        RECT -32.125 -119.165 -31.795 -118.835 ;
        RECT -32.125 -124.605 -31.795 -124.275 ;
        RECT -32.125 -128.685 -31.795 -128.355 ;
        RECT -32.125 -130.045 -31.795 -129.715 ;
        RECT -32.125 -131.405 -31.795 -131.075 ;
        RECT -32.125 -132.765 -31.795 -132.435 ;
        RECT -32.125 -134.125 -31.795 -133.795 ;
        RECT -32.125 -135.485 -31.795 -135.155 ;
        RECT -32.125 -136.845 -31.795 -136.515 ;
        RECT -32.125 -138.205 -31.795 -137.875 ;
        RECT -32.125 -139.565 -31.795 -139.235 ;
        RECT -32.125 -140.925 -31.795 -140.595 ;
        RECT -32.125 -142.285 -31.795 -141.955 ;
        RECT -32.125 -143.645 -31.795 -143.315 ;
        RECT -32.125 -145.005 -31.795 -144.675 ;
        RECT -32.125 -146.365 -31.795 -146.035 ;
        RECT -32.125 -147.725 -31.795 -147.395 ;
        RECT -32.125 -149.085 -31.795 -148.755 ;
        RECT -32.125 -150.445 -31.795 -150.115 ;
        RECT -32.125 -151.805 -31.795 -151.475 ;
        RECT -32.125 -153.165 -31.795 -152.835 ;
        RECT -32.125 -154.525 -31.795 -154.195 ;
        RECT -32.125 -155.885 -31.795 -155.555 ;
        RECT -32.125 -157.245 -31.795 -156.915 ;
        RECT -32.125 -159.965 -31.795 -159.635 ;
        RECT -32.125 -162.685 -31.795 -162.355 ;
        RECT -32.125 -164.045 -31.795 -163.715 ;
        RECT -32.125 -165.405 -31.795 -165.075 ;
        RECT -32.125 -166.765 -31.795 -166.435 ;
        RECT -32.125 -168.125 -31.795 -167.795 ;
        RECT -32.125 -169.485 -31.795 -169.155 ;
        RECT -32.125 -170.845 -31.795 -170.515 ;
        RECT -32.125 -172.205 -31.795 -171.875 ;
        RECT -32.125 -173.565 -31.795 -173.235 ;
        RECT -32.125 -174.925 -31.795 -174.595 ;
        RECT -32.125 -176.285 -31.795 -175.955 ;
        RECT -32.125 -177.645 -31.795 -177.315 ;
        RECT -32.125 -179.005 -31.795 -178.675 ;
        RECT -32.125 -180.365 -31.795 -180.035 ;
        RECT -32.125 -181.725 -31.795 -181.395 ;
        RECT -32.125 -183.085 -31.795 -182.755 ;
        RECT -32.125 -184.445 -31.795 -184.115 ;
        RECT -32.125 -185.805 -31.795 -185.475 ;
        RECT -32.125 -187.165 -31.795 -186.835 ;
        RECT -32.125 -191.245 -31.795 -190.915 ;
        RECT -32.125 -192.605 -31.795 -192.275 ;
        RECT -32.125 -193.965 -31.795 -193.635 ;
        RECT -32.125 -195.325 -31.795 -194.995 ;
        RECT -32.125 -196.685 -31.795 -196.355 ;
        RECT -32.125 -198.045 -31.795 -197.715 ;
        RECT -32.125 -199.405 -31.795 -199.075 ;
        RECT -32.125 -200.765 -31.795 -200.435 ;
        RECT -32.125 -202.125 -31.795 -201.795 ;
        RECT -32.125 -203.485 -31.795 -203.155 ;
        RECT -32.125 -204.845 -31.795 -204.515 ;
        RECT -32.125 -206.205 -31.795 -205.875 ;
        RECT -32.125 -208.925 -31.795 -208.595 ;
        RECT -32.125 -210.285 -31.795 -209.955 ;
        RECT -32.125 -214.365 -31.795 -214.035 ;
        RECT -32.125 -215.725 -31.795 -215.395 ;
        RECT -32.125 -217.085 -31.795 -216.755 ;
        RECT -32.125 -218.445 -31.795 -218.115 ;
        RECT -32.125 -219.805 -31.795 -219.475 ;
        RECT -32.125 -221.165 -31.795 -220.835 ;
        RECT -32.125 -222.525 -31.795 -222.195 ;
        RECT -32.125 -223.885 -31.795 -223.555 ;
        RECT -32.125 -225.245 -31.795 -224.915 ;
        RECT -32.125 -227.965 -31.795 -227.635 ;
        RECT -32.125 -230.685 -31.795 -230.355 ;
        RECT -32.125 -232.045 -31.795 -231.715 ;
        RECT -32.125 -233.225 -31.795 -232.895 ;
        RECT -32.125 -234.765 -31.795 -234.435 ;
        RECT -32.125 -236.125 -31.795 -235.795 ;
        RECT -32.125 -237.485 -31.795 -237.155 ;
        RECT -32.125 -238.845 -31.795 -238.515 ;
        RECT -32.125 -241.09 -31.795 -239.96 ;
        RECT -32.12 -241.205 -31.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 244.04 -30.435 245.17 ;
        RECT -30.765 242.595 -30.435 242.925 ;
        RECT -30.765 241.235 -30.435 241.565 ;
        RECT -30.765 239.875 -30.435 240.205 ;
        RECT -30.765 238.515 -30.435 238.845 ;
        RECT -30.765 237.155 -30.435 237.485 ;
        RECT -30.765 235.795 -30.435 236.125 ;
        RECT -30.765 234.435 -30.435 234.765 ;
        RECT -30.765 233.075 -30.435 233.405 ;
        RECT -30.765 231.715 -30.435 232.045 ;
        RECT -30.765 230.355 -30.435 230.685 ;
        RECT -30.765 228.995 -30.435 229.325 ;
        RECT -30.765 227.635 -30.435 227.965 ;
        RECT -30.765 226.275 -30.435 226.605 ;
        RECT -30.765 224.915 -30.435 225.245 ;
        RECT -30.765 223.555 -30.435 223.885 ;
        RECT -30.765 222.195 -30.435 222.525 ;
        RECT -30.765 220.835 -30.435 221.165 ;
        RECT -30.765 219.475 -30.435 219.805 ;
        RECT -30.765 218.115 -30.435 218.445 ;
        RECT -30.765 216.755 -30.435 217.085 ;
        RECT -30.765 215.395 -30.435 215.725 ;
        RECT -30.765 214.035 -30.435 214.365 ;
        RECT -30.765 212.675 -30.435 213.005 ;
        RECT -30.765 211.315 -30.435 211.645 ;
        RECT -30.765 209.955 -30.435 210.285 ;
        RECT -30.765 208.595 -30.435 208.925 ;
        RECT -30.765 207.235 -30.435 207.565 ;
        RECT -30.765 205.875 -30.435 206.205 ;
        RECT -30.765 204.515 -30.435 204.845 ;
        RECT -30.765 203.155 -30.435 203.485 ;
        RECT -30.765 201.795 -30.435 202.125 ;
        RECT -30.765 200.435 -30.435 200.765 ;
        RECT -30.765 199.075 -30.435 199.405 ;
        RECT -30.765 197.715 -30.435 198.045 ;
        RECT -30.765 196.355 -30.435 196.685 ;
        RECT -30.765 194.995 -30.435 195.325 ;
        RECT -30.765 193.635 -30.435 193.965 ;
        RECT -30.765 192.275 -30.435 192.605 ;
        RECT -30.765 190.915 -30.435 191.245 ;
        RECT -30.765 189.555 -30.435 189.885 ;
        RECT -30.765 188.195 -30.435 188.525 ;
        RECT -30.765 186.835 -30.435 187.165 ;
        RECT -30.765 185.475 -30.435 185.805 ;
        RECT -30.765 184.115 -30.435 184.445 ;
        RECT -30.765 182.755 -30.435 183.085 ;
        RECT -30.765 181.395 -30.435 181.725 ;
        RECT -30.765 180.035 -30.435 180.365 ;
        RECT -30.765 178.675 -30.435 179.005 ;
        RECT -30.765 177.315 -30.435 177.645 ;
        RECT -30.765 175.955 -30.435 176.285 ;
        RECT -30.765 174.595 -30.435 174.925 ;
        RECT -30.765 173.235 -30.435 173.565 ;
        RECT -30.765 171.875 -30.435 172.205 ;
        RECT -30.765 170.515 -30.435 170.845 ;
        RECT -30.765 169.155 -30.435 169.485 ;
        RECT -30.765 167.795 -30.435 168.125 ;
        RECT -30.765 166.435 -30.435 166.765 ;
        RECT -30.765 165.075 -30.435 165.405 ;
        RECT -30.765 163.715 -30.435 164.045 ;
        RECT -30.765 162.355 -30.435 162.685 ;
        RECT -30.765 160.995 -30.435 161.325 ;
        RECT -30.765 159.635 -30.435 159.965 ;
        RECT -30.765 158.275 -30.435 158.605 ;
        RECT -30.765 156.915 -30.435 157.245 ;
        RECT -30.765 155.555 -30.435 155.885 ;
        RECT -30.765 154.195 -30.435 154.525 ;
        RECT -30.765 152.835 -30.435 153.165 ;
        RECT -30.765 151.475 -30.435 151.805 ;
        RECT -30.765 150.115 -30.435 150.445 ;
        RECT -30.765 148.755 -30.435 149.085 ;
        RECT -30.765 147.395 -30.435 147.725 ;
        RECT -30.765 146.035 -30.435 146.365 ;
        RECT -30.765 144.675 -30.435 145.005 ;
        RECT -30.765 143.315 -30.435 143.645 ;
        RECT -30.765 141.955 -30.435 142.285 ;
        RECT -30.765 140.595 -30.435 140.925 ;
        RECT -30.765 139.235 -30.435 139.565 ;
        RECT -30.765 137.875 -30.435 138.205 ;
        RECT -30.765 136.515 -30.435 136.845 ;
        RECT -30.765 135.155 -30.435 135.485 ;
        RECT -30.765 133.795 -30.435 134.125 ;
        RECT -30.765 132.435 -30.435 132.765 ;
        RECT -30.765 131.075 -30.435 131.405 ;
        RECT -30.765 129.715 -30.435 130.045 ;
        RECT -30.765 128.355 -30.435 128.685 ;
        RECT -30.765 126.995 -30.435 127.325 ;
        RECT -30.765 125.635 -30.435 125.965 ;
        RECT -30.765 124.275 -30.435 124.605 ;
        RECT -30.765 122.915 -30.435 123.245 ;
        RECT -30.765 121.555 -30.435 121.885 ;
        RECT -30.765 120.195 -30.435 120.525 ;
        RECT -30.765 118.835 -30.435 119.165 ;
        RECT -30.765 117.475 -30.435 117.805 ;
        RECT -30.765 116.115 -30.435 116.445 ;
        RECT -30.765 114.755 -30.435 115.085 ;
        RECT -30.765 113.395 -30.435 113.725 ;
        RECT -30.765 112.035 -30.435 112.365 ;
        RECT -30.765 110.675 -30.435 111.005 ;
        RECT -30.765 109.315 -30.435 109.645 ;
        RECT -30.765 107.955 -30.435 108.285 ;
        RECT -30.765 106.595 -30.435 106.925 ;
        RECT -30.765 105.235 -30.435 105.565 ;
        RECT -30.765 103.875 -30.435 104.205 ;
        RECT -30.765 102.515 -30.435 102.845 ;
        RECT -30.765 101.155 -30.435 101.485 ;
        RECT -30.765 99.795 -30.435 100.125 ;
        RECT -30.765 98.435 -30.435 98.765 ;
        RECT -30.765 97.075 -30.435 97.405 ;
        RECT -30.765 95.715 -30.435 96.045 ;
        RECT -30.765 94.355 -30.435 94.685 ;
        RECT -30.765 92.995 -30.435 93.325 ;
        RECT -30.765 91.635 -30.435 91.965 ;
        RECT -30.765 90.275 -30.435 90.605 ;
        RECT -30.765 88.915 -30.435 89.245 ;
        RECT -30.765 87.555 -30.435 87.885 ;
        RECT -30.765 86.195 -30.435 86.525 ;
        RECT -30.765 84.835 -30.435 85.165 ;
        RECT -30.765 83.475 -30.435 83.805 ;
        RECT -30.765 82.115 -30.435 82.445 ;
        RECT -30.765 80.755 -30.435 81.085 ;
        RECT -30.765 79.395 -30.435 79.725 ;
        RECT -30.765 78.035 -30.435 78.365 ;
        RECT -30.765 76.675 -30.435 77.005 ;
        RECT -30.765 75.315 -30.435 75.645 ;
        RECT -30.765 73.955 -30.435 74.285 ;
        RECT -30.765 72.595 -30.435 72.925 ;
        RECT -30.765 71.235 -30.435 71.565 ;
        RECT -30.765 69.875 -30.435 70.205 ;
        RECT -30.765 68.515 -30.435 68.845 ;
        RECT -30.765 67.155 -30.435 67.485 ;
        RECT -30.765 65.795 -30.435 66.125 ;
        RECT -30.765 64.435 -30.435 64.765 ;
        RECT -30.765 63.075 -30.435 63.405 ;
        RECT -30.765 61.715 -30.435 62.045 ;
        RECT -30.765 60.355 -30.435 60.685 ;
        RECT -30.765 58.995 -30.435 59.325 ;
        RECT -30.765 57.635 -30.435 57.965 ;
        RECT -30.765 56.275 -30.435 56.605 ;
        RECT -30.765 54.915 -30.435 55.245 ;
        RECT -30.765 53.555 -30.435 53.885 ;
        RECT -30.765 52.195 -30.435 52.525 ;
        RECT -30.765 50.835 -30.435 51.165 ;
        RECT -30.765 49.475 -30.435 49.805 ;
        RECT -30.765 48.115 -30.435 48.445 ;
        RECT -30.765 46.755 -30.435 47.085 ;
        RECT -30.765 45.395 -30.435 45.725 ;
        RECT -30.765 44.035 -30.435 44.365 ;
        RECT -30.765 42.675 -30.435 43.005 ;
        RECT -30.765 41.315 -30.435 41.645 ;
        RECT -30.765 39.955 -30.435 40.285 ;
        RECT -30.765 38.595 -30.435 38.925 ;
        RECT -30.765 37.235 -30.435 37.565 ;
        RECT -30.765 35.875 -30.435 36.205 ;
        RECT -30.765 34.515 -30.435 34.845 ;
        RECT -30.765 33.155 -30.435 33.485 ;
        RECT -30.765 31.795 -30.435 32.125 ;
        RECT -30.765 30.435 -30.435 30.765 ;
        RECT -30.765 29.075 -30.435 29.405 ;
        RECT -30.765 27.715 -30.435 28.045 ;
        RECT -30.765 26.355 -30.435 26.685 ;
        RECT -30.765 24.995 -30.435 25.325 ;
        RECT -30.765 23.635 -30.435 23.965 ;
        RECT -30.765 22.275 -30.435 22.605 ;
        RECT -30.765 20.915 -30.435 21.245 ;
        RECT -30.765 19.555 -30.435 19.885 ;
        RECT -30.765 18.195 -30.435 18.525 ;
        RECT -30.765 16.835 -30.435 17.165 ;
        RECT -30.765 15.475 -30.435 15.805 ;
        RECT -30.765 14.115 -30.435 14.445 ;
        RECT -30.765 12.755 -30.435 13.085 ;
        RECT -30.765 11.395 -30.435 11.725 ;
        RECT -30.765 10.035 -30.435 10.365 ;
        RECT -30.765 8.675 -30.435 9.005 ;
        RECT -30.765 7.315 -30.435 7.645 ;
        RECT -30.765 5.955 -30.435 6.285 ;
        RECT -30.765 4.595 -30.435 4.925 ;
        RECT -30.765 3.235 -30.435 3.565 ;
        RECT -30.765 1.875 -30.435 2.205 ;
        RECT -30.765 0.515 -30.435 0.845 ;
        RECT -30.765 -7.645 -30.435 -7.315 ;
        RECT -30.765 -10.365 -30.435 -10.035 ;
        RECT -30.765 -11.725 -30.435 -11.395 ;
        RECT -30.765 -14.445 -30.435 -14.115 ;
        RECT -30.765 -15.805 -30.435 -15.475 ;
        RECT -30.765 -19.885 -30.435 -19.555 ;
        RECT -30.765 -29.405 -30.435 -29.075 ;
        RECT -30.765 -32.125 -30.435 -31.795 ;
        RECT -30.765 -33.485 -30.435 -33.155 ;
        RECT -30.765 -34.88 -30.435 -34.55 ;
        RECT -30.765 -36.205 -30.435 -35.875 ;
        RECT -30.765 -38.925 -30.435 -38.595 ;
        RECT -30.765 -39.97 -30.435 -39.64 ;
        RECT -30.765 -48.445 -30.435 -48.115 ;
        RECT -30.765 -49.805 -30.435 -49.475 ;
        RECT -30.765 -51.165 -30.435 -50.835 ;
        RECT -30.765 -53.885 -30.435 -53.555 ;
        RECT -30.765 -57.965 -30.435 -57.635 ;
        RECT -30.76 -59.32 -30.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 -128.685 -30.435 -128.355 ;
        RECT -30.765 -130.045 -30.435 -129.715 ;
        RECT -30.765 -131.405 -30.435 -131.075 ;
        RECT -30.765 -132.765 -30.435 -132.435 ;
        RECT -30.765 -135.485 -30.435 -135.155 ;
        RECT -30.765 -136.845 -30.435 -136.515 ;
        RECT -30.765 -138.205 -30.435 -137.875 ;
        RECT -30.765 -139.565 -30.435 -139.235 ;
        RECT -30.765 -140.925 -30.435 -140.595 ;
        RECT -30.765 -142.285 -30.435 -141.955 ;
        RECT -30.765 -145.005 -30.435 -144.675 ;
        RECT -30.765 -146.365 -30.435 -146.035 ;
        RECT -30.765 -147.725 -30.435 -147.395 ;
        RECT -30.765 -153.165 -30.435 -152.835 ;
        RECT -30.765 -154.525 -30.435 -154.195 ;
        RECT -30.765 -155.885 -30.435 -155.555 ;
        RECT -30.765 -157.245 -30.435 -156.915 ;
        RECT -30.765 -162.685 -30.435 -162.355 ;
        RECT -30.765 -164.045 -30.435 -163.715 ;
        RECT -30.765 -165.405 -30.435 -165.075 ;
        RECT -30.765 -166.765 -30.435 -166.435 ;
        RECT -30.765 -168.125 -30.435 -167.795 ;
        RECT -30.765 -169.485 -30.435 -169.155 ;
        RECT -30.765 -170.845 -30.435 -170.515 ;
        RECT -30.765 -172.205 -30.435 -171.875 ;
        RECT -30.765 -173.565 -30.435 -173.235 ;
        RECT -30.765 -174.925 -30.435 -174.595 ;
        RECT -30.765 -176.285 -30.435 -175.955 ;
        RECT -30.765 -177.645 -30.435 -177.315 ;
        RECT -30.765 -179.005 -30.435 -178.675 ;
        RECT -30.765 -180.365 -30.435 -180.035 ;
        RECT -30.765 -181.725 -30.435 -181.395 ;
        RECT -30.765 -183.085 -30.435 -182.755 ;
        RECT -30.765 -184.445 -30.435 -184.115 ;
        RECT -30.765 -185.805 -30.435 -185.475 ;
        RECT -30.765 -187.165 -30.435 -186.835 ;
        RECT -30.765 -191.245 -30.435 -190.915 ;
        RECT -30.765 -192.605 -30.435 -192.275 ;
        RECT -30.765 -193.965 -30.435 -193.635 ;
        RECT -30.765 -195.325 -30.435 -194.995 ;
        RECT -30.765 -196.685 -30.435 -196.355 ;
        RECT -30.765 -198.045 -30.435 -197.715 ;
        RECT -30.765 -199.405 -30.435 -199.075 ;
        RECT -30.765 -200.765 -30.435 -200.435 ;
        RECT -30.765 -202.125 -30.435 -201.795 ;
        RECT -30.765 -203.485 -30.435 -203.155 ;
        RECT -30.765 -204.845 -30.435 -204.515 ;
        RECT -30.765 -206.205 -30.435 -205.875 ;
        RECT -30.765 -208.925 -30.435 -208.595 ;
        RECT -30.765 -210.285 -30.435 -209.955 ;
        RECT -30.765 -214.365 -30.435 -214.035 ;
        RECT -30.765 -215.725 -30.435 -215.395 ;
        RECT -30.765 -217.085 -30.435 -216.755 ;
        RECT -30.765 -218.445 -30.435 -218.115 ;
        RECT -30.765 -219.805 -30.435 -219.475 ;
        RECT -30.765 -221.165 -30.435 -220.835 ;
        RECT -30.765 -222.525 -30.435 -222.195 ;
        RECT -30.765 -223.885 -30.435 -223.555 ;
        RECT -30.765 -225.245 -30.435 -224.915 ;
        RECT -30.765 -227.965 -30.435 -227.635 ;
        RECT -30.765 -230.685 -30.435 -230.355 ;
        RECT -30.765 -232.045 -30.435 -231.715 ;
        RECT -30.765 -233.225 -30.435 -232.895 ;
        RECT -30.765 -234.765 -30.435 -234.435 ;
        RECT -30.765 -236.125 -30.435 -235.795 ;
        RECT -30.765 -237.485 -30.435 -237.155 ;
        RECT -30.765 -238.845 -30.435 -238.515 ;
        RECT -30.765 -241.09 -30.435 -239.96 ;
        RECT -30.76 -241.205 -30.44 -120.88 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 169.155 -29.075 169.485 ;
        RECT -29.405 167.795 -29.075 168.125 ;
        RECT -29.405 166.435 -29.075 166.765 ;
        RECT -29.405 165.075 -29.075 165.405 ;
        RECT -29.405 163.715 -29.075 164.045 ;
        RECT -29.405 162.355 -29.075 162.685 ;
        RECT -29.405 160.995 -29.075 161.325 ;
        RECT -29.405 159.635 -29.075 159.965 ;
        RECT -29.405 158.275 -29.075 158.605 ;
        RECT -29.405 156.915 -29.075 157.245 ;
        RECT -29.405 155.555 -29.075 155.885 ;
        RECT -29.405 154.195 -29.075 154.525 ;
        RECT -29.405 152.835 -29.075 153.165 ;
        RECT -29.405 151.475 -29.075 151.805 ;
        RECT -29.405 150.115 -29.075 150.445 ;
        RECT -29.405 148.755 -29.075 149.085 ;
        RECT -29.405 147.395 -29.075 147.725 ;
        RECT -29.405 146.035 -29.075 146.365 ;
        RECT -29.405 144.675 -29.075 145.005 ;
        RECT -29.405 143.315 -29.075 143.645 ;
        RECT -29.405 141.955 -29.075 142.285 ;
        RECT -29.405 140.595 -29.075 140.925 ;
        RECT -29.405 139.235 -29.075 139.565 ;
        RECT -29.405 137.875 -29.075 138.205 ;
        RECT -29.405 136.515 -29.075 136.845 ;
        RECT -29.405 135.155 -29.075 135.485 ;
        RECT -29.405 133.795 -29.075 134.125 ;
        RECT -29.405 132.435 -29.075 132.765 ;
        RECT -29.405 131.075 -29.075 131.405 ;
        RECT -29.405 129.715 -29.075 130.045 ;
        RECT -29.405 128.355 -29.075 128.685 ;
        RECT -29.405 126.995 -29.075 127.325 ;
        RECT -29.405 125.635 -29.075 125.965 ;
        RECT -29.405 124.275 -29.075 124.605 ;
        RECT -29.405 122.915 -29.075 123.245 ;
        RECT -29.405 121.555 -29.075 121.885 ;
        RECT -29.405 120.195 -29.075 120.525 ;
        RECT -29.405 118.835 -29.075 119.165 ;
        RECT -29.405 117.475 -29.075 117.805 ;
        RECT -29.405 116.115 -29.075 116.445 ;
        RECT -29.405 114.755 -29.075 115.085 ;
        RECT -29.405 113.395 -29.075 113.725 ;
        RECT -29.405 112.035 -29.075 112.365 ;
        RECT -29.405 110.675 -29.075 111.005 ;
        RECT -29.405 109.315 -29.075 109.645 ;
        RECT -29.405 107.955 -29.075 108.285 ;
        RECT -29.405 106.595 -29.075 106.925 ;
        RECT -29.405 105.235 -29.075 105.565 ;
        RECT -29.405 103.875 -29.075 104.205 ;
        RECT -29.405 102.515 -29.075 102.845 ;
        RECT -29.405 101.155 -29.075 101.485 ;
        RECT -29.405 99.795 -29.075 100.125 ;
        RECT -29.405 98.435 -29.075 98.765 ;
        RECT -29.405 97.075 -29.075 97.405 ;
        RECT -29.405 95.715 -29.075 96.045 ;
        RECT -29.405 94.355 -29.075 94.685 ;
        RECT -29.405 92.995 -29.075 93.325 ;
        RECT -29.405 91.635 -29.075 91.965 ;
        RECT -29.405 90.275 -29.075 90.605 ;
        RECT -29.405 88.915 -29.075 89.245 ;
        RECT -29.405 87.555 -29.075 87.885 ;
        RECT -29.405 86.195 -29.075 86.525 ;
        RECT -29.405 84.835 -29.075 85.165 ;
        RECT -29.405 83.475 -29.075 83.805 ;
        RECT -29.405 82.115 -29.075 82.445 ;
        RECT -29.405 80.755 -29.075 81.085 ;
        RECT -29.405 79.395 -29.075 79.725 ;
        RECT -29.405 78.035 -29.075 78.365 ;
        RECT -29.405 76.675 -29.075 77.005 ;
        RECT -29.405 75.315 -29.075 75.645 ;
        RECT -29.405 73.955 -29.075 74.285 ;
        RECT -29.405 72.595 -29.075 72.925 ;
        RECT -29.405 71.235 -29.075 71.565 ;
        RECT -29.405 69.875 -29.075 70.205 ;
        RECT -29.405 68.515 -29.075 68.845 ;
        RECT -29.405 67.155 -29.075 67.485 ;
        RECT -29.405 65.795 -29.075 66.125 ;
        RECT -29.405 64.435 -29.075 64.765 ;
        RECT -29.405 63.075 -29.075 63.405 ;
        RECT -29.405 61.715 -29.075 62.045 ;
        RECT -29.405 60.355 -29.075 60.685 ;
        RECT -29.405 58.995 -29.075 59.325 ;
        RECT -29.405 57.635 -29.075 57.965 ;
        RECT -29.405 56.275 -29.075 56.605 ;
        RECT -29.405 54.915 -29.075 55.245 ;
        RECT -29.405 53.555 -29.075 53.885 ;
        RECT -29.405 52.195 -29.075 52.525 ;
        RECT -29.405 50.835 -29.075 51.165 ;
        RECT -29.405 49.475 -29.075 49.805 ;
        RECT -29.405 48.115 -29.075 48.445 ;
        RECT -29.405 46.755 -29.075 47.085 ;
        RECT -29.405 45.395 -29.075 45.725 ;
        RECT -29.405 44.035 -29.075 44.365 ;
        RECT -29.405 42.675 -29.075 43.005 ;
        RECT -29.405 41.315 -29.075 41.645 ;
        RECT -29.405 39.955 -29.075 40.285 ;
        RECT -29.405 38.595 -29.075 38.925 ;
        RECT -29.405 37.235 -29.075 37.565 ;
        RECT -29.405 35.875 -29.075 36.205 ;
        RECT -29.405 34.515 -29.075 34.845 ;
        RECT -29.405 33.155 -29.075 33.485 ;
        RECT -29.405 31.795 -29.075 32.125 ;
        RECT -29.405 30.435 -29.075 30.765 ;
        RECT -29.405 29.075 -29.075 29.405 ;
        RECT -29.405 27.715 -29.075 28.045 ;
        RECT -29.405 26.355 -29.075 26.685 ;
        RECT -29.405 24.995 -29.075 25.325 ;
        RECT -29.405 23.635 -29.075 23.965 ;
        RECT -29.405 22.275 -29.075 22.605 ;
        RECT -29.405 20.915 -29.075 21.245 ;
        RECT -29.405 19.555 -29.075 19.885 ;
        RECT -29.405 18.195 -29.075 18.525 ;
        RECT -29.405 16.835 -29.075 17.165 ;
        RECT -29.405 15.475 -29.075 15.805 ;
        RECT -29.405 14.115 -29.075 14.445 ;
        RECT -29.405 12.755 -29.075 13.085 ;
        RECT -29.405 11.395 -29.075 11.725 ;
        RECT -29.405 10.035 -29.075 10.365 ;
        RECT -29.405 8.675 -29.075 9.005 ;
        RECT -29.405 7.315 -29.075 7.645 ;
        RECT -29.405 5.955 -29.075 6.285 ;
        RECT -29.405 4.595 -29.075 4.925 ;
        RECT -29.405 3.235 -29.075 3.565 ;
        RECT -29.405 1.875 -29.075 2.205 ;
        RECT -29.405 0.515 -29.075 0.845 ;
        RECT -29.405 -7.645 -29.075 -7.315 ;
        RECT -29.405 -10.365 -29.075 -10.035 ;
        RECT -29.405 -11.725 -29.075 -11.395 ;
        RECT -29.405 -13.7 -29.075 -13.37 ;
        RECT -29.405 -14.445 -29.075 -14.115 ;
        RECT -29.405 -15.805 -29.075 -15.475 ;
        RECT -29.405 -18.79 -29.075 -18.46 ;
        RECT -29.405 -19.885 -29.075 -19.555 ;
        RECT -29.405 -29.405 -29.075 -29.075 ;
        RECT -29.405 -32.125 -29.075 -31.795 ;
        RECT -29.405 -33.485 -29.075 -33.155 ;
        RECT -29.405 -34.88 -29.075 -34.55 ;
        RECT -29.405 -36.205 -29.075 -35.875 ;
        RECT -29.405 -38.925 -29.075 -38.595 ;
        RECT -29.405 -39.97 -29.075 -39.64 ;
        RECT -29.405 -48.445 -29.075 -48.115 ;
        RECT -29.405 -49.805 -29.075 -49.475 ;
        RECT -29.405 -51.165 -29.075 -50.835 ;
        RECT -29.405 -53.885 -29.075 -53.555 ;
        RECT -29.405 -57.965 -29.075 -57.635 ;
        RECT -29.4 -58.64 -29.08 245.285 ;
        RECT -29.405 244.04 -29.075 245.17 ;
        RECT -29.405 242.595 -29.075 242.925 ;
        RECT -29.405 241.235 -29.075 241.565 ;
        RECT -29.405 239.875 -29.075 240.205 ;
        RECT -29.405 238.515 -29.075 238.845 ;
        RECT -29.405 237.155 -29.075 237.485 ;
        RECT -29.405 235.795 -29.075 236.125 ;
        RECT -29.405 234.435 -29.075 234.765 ;
        RECT -29.405 233.075 -29.075 233.405 ;
        RECT -29.405 231.715 -29.075 232.045 ;
        RECT -29.405 230.355 -29.075 230.685 ;
        RECT -29.405 228.995 -29.075 229.325 ;
        RECT -29.405 227.635 -29.075 227.965 ;
        RECT -29.405 226.275 -29.075 226.605 ;
        RECT -29.405 224.915 -29.075 225.245 ;
        RECT -29.405 223.555 -29.075 223.885 ;
        RECT -29.405 222.195 -29.075 222.525 ;
        RECT -29.405 220.835 -29.075 221.165 ;
        RECT -29.405 219.475 -29.075 219.805 ;
        RECT -29.405 218.115 -29.075 218.445 ;
        RECT -29.405 216.755 -29.075 217.085 ;
        RECT -29.405 215.395 -29.075 215.725 ;
        RECT -29.405 214.035 -29.075 214.365 ;
        RECT -29.405 212.675 -29.075 213.005 ;
        RECT -29.405 211.315 -29.075 211.645 ;
        RECT -29.405 209.955 -29.075 210.285 ;
        RECT -29.405 208.595 -29.075 208.925 ;
        RECT -29.405 207.235 -29.075 207.565 ;
        RECT -29.405 205.875 -29.075 206.205 ;
        RECT -29.405 204.515 -29.075 204.845 ;
        RECT -29.405 203.155 -29.075 203.485 ;
        RECT -29.405 201.795 -29.075 202.125 ;
        RECT -29.405 200.435 -29.075 200.765 ;
        RECT -29.405 199.075 -29.075 199.405 ;
        RECT -29.405 197.715 -29.075 198.045 ;
        RECT -29.405 196.355 -29.075 196.685 ;
        RECT -29.405 194.995 -29.075 195.325 ;
        RECT -29.405 193.635 -29.075 193.965 ;
        RECT -29.405 192.275 -29.075 192.605 ;
        RECT -29.405 190.915 -29.075 191.245 ;
        RECT -29.405 189.555 -29.075 189.885 ;
        RECT -29.405 188.195 -29.075 188.525 ;
        RECT -29.405 186.835 -29.075 187.165 ;
        RECT -29.405 185.475 -29.075 185.805 ;
        RECT -29.405 184.115 -29.075 184.445 ;
        RECT -29.405 182.755 -29.075 183.085 ;
        RECT -29.405 181.395 -29.075 181.725 ;
        RECT -29.405 180.035 -29.075 180.365 ;
        RECT -29.405 178.675 -29.075 179.005 ;
        RECT -29.405 177.315 -29.075 177.645 ;
        RECT -29.405 175.955 -29.075 176.285 ;
        RECT -29.405 174.595 -29.075 174.925 ;
        RECT -29.405 173.235 -29.075 173.565 ;
        RECT -29.405 171.875 -29.075 172.205 ;
        RECT -29.405 170.515 -29.075 170.845 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.205 244.04 -35.875 245.17 ;
        RECT -36.205 242.595 -35.875 242.925 ;
        RECT -36.205 241.235 -35.875 241.565 ;
        RECT -36.205 239.875 -35.875 240.205 ;
        RECT -36.205 238.515 -35.875 238.845 ;
        RECT -36.205 237.155 -35.875 237.485 ;
        RECT -36.205 235.795 -35.875 236.125 ;
        RECT -36.205 234.435 -35.875 234.765 ;
        RECT -36.205 233.075 -35.875 233.405 ;
        RECT -36.205 231.715 -35.875 232.045 ;
        RECT -36.205 230.355 -35.875 230.685 ;
        RECT -36.205 228.995 -35.875 229.325 ;
        RECT -36.205 227.635 -35.875 227.965 ;
        RECT -36.205 226.275 -35.875 226.605 ;
        RECT -36.205 224.915 -35.875 225.245 ;
        RECT -36.205 223.555 -35.875 223.885 ;
        RECT -36.205 222.195 -35.875 222.525 ;
        RECT -36.205 220.835 -35.875 221.165 ;
        RECT -36.205 219.475 -35.875 219.805 ;
        RECT -36.205 218.115 -35.875 218.445 ;
        RECT -36.205 216.755 -35.875 217.085 ;
        RECT -36.205 215.395 -35.875 215.725 ;
        RECT -36.205 214.035 -35.875 214.365 ;
        RECT -36.205 212.675 -35.875 213.005 ;
        RECT -36.205 211.315 -35.875 211.645 ;
        RECT -36.205 209.955 -35.875 210.285 ;
        RECT -36.205 208.595 -35.875 208.925 ;
        RECT -36.205 207.235 -35.875 207.565 ;
        RECT -36.205 205.875 -35.875 206.205 ;
        RECT -36.205 204.515 -35.875 204.845 ;
        RECT -36.205 203.155 -35.875 203.485 ;
        RECT -36.205 201.795 -35.875 202.125 ;
        RECT -36.205 200.435 -35.875 200.765 ;
        RECT -36.205 199.075 -35.875 199.405 ;
        RECT -36.205 197.715 -35.875 198.045 ;
        RECT -36.205 196.355 -35.875 196.685 ;
        RECT -36.205 194.995 -35.875 195.325 ;
        RECT -36.205 193.635 -35.875 193.965 ;
        RECT -36.205 192.275 -35.875 192.605 ;
        RECT -36.205 190.915 -35.875 191.245 ;
        RECT -36.205 189.555 -35.875 189.885 ;
        RECT -36.205 188.195 -35.875 188.525 ;
        RECT -36.205 186.835 -35.875 187.165 ;
        RECT -36.205 185.475 -35.875 185.805 ;
        RECT -36.205 184.115 -35.875 184.445 ;
        RECT -36.205 182.755 -35.875 183.085 ;
        RECT -36.205 181.395 -35.875 181.725 ;
        RECT -36.205 180.035 -35.875 180.365 ;
        RECT -36.205 178.675 -35.875 179.005 ;
        RECT -36.205 177.315 -35.875 177.645 ;
        RECT -36.205 175.955 -35.875 176.285 ;
        RECT -36.205 174.595 -35.875 174.925 ;
        RECT -36.205 173.235 -35.875 173.565 ;
        RECT -36.205 171.875 -35.875 172.205 ;
        RECT -36.205 170.515 -35.875 170.845 ;
        RECT -36.205 169.155 -35.875 169.485 ;
        RECT -36.205 167.795 -35.875 168.125 ;
        RECT -36.205 166.435 -35.875 166.765 ;
        RECT -36.205 165.075 -35.875 165.405 ;
        RECT -36.205 163.715 -35.875 164.045 ;
        RECT -36.205 162.355 -35.875 162.685 ;
        RECT -36.205 160.995 -35.875 161.325 ;
        RECT -36.205 159.635 -35.875 159.965 ;
        RECT -36.205 158.275 -35.875 158.605 ;
        RECT -36.205 156.915 -35.875 157.245 ;
        RECT -36.205 155.555 -35.875 155.885 ;
        RECT -36.205 154.195 -35.875 154.525 ;
        RECT -36.205 152.835 -35.875 153.165 ;
        RECT -36.205 151.475 -35.875 151.805 ;
        RECT -36.205 150.115 -35.875 150.445 ;
        RECT -36.205 148.755 -35.875 149.085 ;
        RECT -36.205 147.395 -35.875 147.725 ;
        RECT -36.205 146.035 -35.875 146.365 ;
        RECT -36.205 144.675 -35.875 145.005 ;
        RECT -36.205 143.315 -35.875 143.645 ;
        RECT -36.205 141.955 -35.875 142.285 ;
        RECT -36.205 140.595 -35.875 140.925 ;
        RECT -36.205 139.235 -35.875 139.565 ;
        RECT -36.205 137.875 -35.875 138.205 ;
        RECT -36.205 136.515 -35.875 136.845 ;
        RECT -36.205 135.155 -35.875 135.485 ;
        RECT -36.205 133.795 -35.875 134.125 ;
        RECT -36.205 132.435 -35.875 132.765 ;
        RECT -36.205 131.075 -35.875 131.405 ;
        RECT -36.205 129.715 -35.875 130.045 ;
        RECT -36.205 128.355 -35.875 128.685 ;
        RECT -36.205 126.995 -35.875 127.325 ;
        RECT -36.205 125.635 -35.875 125.965 ;
        RECT -36.205 124.275 -35.875 124.605 ;
        RECT -36.205 122.915 -35.875 123.245 ;
        RECT -36.205 121.555 -35.875 121.885 ;
        RECT -36.205 120.195 -35.875 120.525 ;
        RECT -36.205 118.835 -35.875 119.165 ;
        RECT -36.205 117.475 -35.875 117.805 ;
        RECT -36.205 116.115 -35.875 116.445 ;
        RECT -36.205 114.755 -35.875 115.085 ;
        RECT -36.205 113.395 -35.875 113.725 ;
        RECT -36.205 112.035 -35.875 112.365 ;
        RECT -36.205 110.675 -35.875 111.005 ;
        RECT -36.205 109.315 -35.875 109.645 ;
        RECT -36.205 107.955 -35.875 108.285 ;
        RECT -36.205 106.595 -35.875 106.925 ;
        RECT -36.205 105.235 -35.875 105.565 ;
        RECT -36.205 103.875 -35.875 104.205 ;
        RECT -36.205 102.515 -35.875 102.845 ;
        RECT -36.205 101.155 -35.875 101.485 ;
        RECT -36.205 99.795 -35.875 100.125 ;
        RECT -36.205 98.435 -35.875 98.765 ;
        RECT -36.205 97.075 -35.875 97.405 ;
        RECT -36.205 95.715 -35.875 96.045 ;
        RECT -36.205 94.355 -35.875 94.685 ;
        RECT -36.205 92.995 -35.875 93.325 ;
        RECT -36.205 91.635 -35.875 91.965 ;
        RECT -36.205 90.275 -35.875 90.605 ;
        RECT -36.205 88.915 -35.875 89.245 ;
        RECT -36.205 87.555 -35.875 87.885 ;
        RECT -36.205 86.195 -35.875 86.525 ;
        RECT -36.205 84.835 -35.875 85.165 ;
        RECT -36.205 83.475 -35.875 83.805 ;
        RECT -36.205 82.115 -35.875 82.445 ;
        RECT -36.205 80.755 -35.875 81.085 ;
        RECT -36.205 79.395 -35.875 79.725 ;
        RECT -36.205 78.035 -35.875 78.365 ;
        RECT -36.205 76.675 -35.875 77.005 ;
        RECT -36.205 75.315 -35.875 75.645 ;
        RECT -36.205 73.955 -35.875 74.285 ;
        RECT -36.205 72.595 -35.875 72.925 ;
        RECT -36.205 71.235 -35.875 71.565 ;
        RECT -36.205 69.875 -35.875 70.205 ;
        RECT -36.205 68.515 -35.875 68.845 ;
        RECT -36.205 67.155 -35.875 67.485 ;
        RECT -36.205 65.795 -35.875 66.125 ;
        RECT -36.205 64.435 -35.875 64.765 ;
        RECT -36.205 63.075 -35.875 63.405 ;
        RECT -36.205 61.715 -35.875 62.045 ;
        RECT -36.205 60.355 -35.875 60.685 ;
        RECT -36.205 58.995 -35.875 59.325 ;
        RECT -36.205 57.635 -35.875 57.965 ;
        RECT -36.205 56.275 -35.875 56.605 ;
        RECT -36.205 54.915 -35.875 55.245 ;
        RECT -36.205 53.555 -35.875 53.885 ;
        RECT -36.205 52.195 -35.875 52.525 ;
        RECT -36.205 50.835 -35.875 51.165 ;
        RECT -36.205 49.475 -35.875 49.805 ;
        RECT -36.205 48.115 -35.875 48.445 ;
        RECT -36.205 46.755 -35.875 47.085 ;
        RECT -36.205 45.395 -35.875 45.725 ;
        RECT -36.205 44.035 -35.875 44.365 ;
        RECT -36.205 42.675 -35.875 43.005 ;
        RECT -36.205 41.315 -35.875 41.645 ;
        RECT -36.205 39.955 -35.875 40.285 ;
        RECT -36.205 38.595 -35.875 38.925 ;
        RECT -36.205 37.235 -35.875 37.565 ;
        RECT -36.205 35.875 -35.875 36.205 ;
        RECT -36.205 34.515 -35.875 34.845 ;
        RECT -36.205 33.155 -35.875 33.485 ;
        RECT -36.205 31.795 -35.875 32.125 ;
        RECT -36.205 30.435 -35.875 30.765 ;
        RECT -36.205 29.075 -35.875 29.405 ;
        RECT -36.205 27.715 -35.875 28.045 ;
        RECT -36.205 26.355 -35.875 26.685 ;
        RECT -36.205 24.995 -35.875 25.325 ;
        RECT -36.205 23.635 -35.875 23.965 ;
        RECT -36.205 22.275 -35.875 22.605 ;
        RECT -36.205 20.915 -35.875 21.245 ;
        RECT -36.205 19.555 -35.875 19.885 ;
        RECT -36.205 18.195 -35.875 18.525 ;
        RECT -36.205 16.835 -35.875 17.165 ;
        RECT -36.205 15.475 -35.875 15.805 ;
        RECT -36.205 14.115 -35.875 14.445 ;
        RECT -36.205 12.755 -35.875 13.085 ;
        RECT -36.205 11.395 -35.875 11.725 ;
        RECT -36.205 10.035 -35.875 10.365 ;
        RECT -36.205 8.675 -35.875 9.005 ;
        RECT -36.205 7.315 -35.875 7.645 ;
        RECT -36.205 5.955 -35.875 6.285 ;
        RECT -36.205 4.595 -35.875 4.925 ;
        RECT -36.205 3.235 -35.875 3.565 ;
        RECT -36.205 1.875 -35.875 2.205 ;
        RECT -36.205 0.515 -35.875 0.845 ;
        RECT -36.205 -2.205 -35.875 -1.875 ;
        RECT -36.205 -3.565 -35.875 -3.235 ;
        RECT -36.205 -4.925 -35.875 -4.595 ;
        RECT -36.205 -7.645 -35.875 -7.315 ;
        RECT -36.205 -9.005 -35.875 -8.675 ;
        RECT -36.205 -10.365 -35.875 -10.035 ;
        RECT -36.205 -11.725 -35.875 -11.395 ;
        RECT -36.205 -13.085 -35.875 -12.755 ;
        RECT -36.205 -14.445 -35.875 -14.115 ;
        RECT -36.205 -15.805 -35.875 -15.475 ;
        RECT -36.205 -17.165 -35.875 -16.835 ;
        RECT -36.205 -18.525 -35.875 -18.195 ;
        RECT -36.205 -19.885 -35.875 -19.555 ;
        RECT -36.205 -21.245 -35.875 -20.915 ;
        RECT -36.205 -22.605 -35.875 -22.275 ;
        RECT -36.205 -29.405 -35.875 -29.075 ;
        RECT -36.205 -32.125 -35.875 -31.795 ;
        RECT -36.205 -33.485 -35.875 -33.155 ;
        RECT -36.205 -34.88 -35.875 -34.55 ;
        RECT -36.205 -36.205 -35.875 -35.875 ;
        RECT -36.205 -38.925 -35.875 -38.595 ;
        RECT -36.205 -39.97 -35.875 -39.64 ;
        RECT -36.205 -47.085 -35.875 -46.755 ;
        RECT -36.205 -48.445 -35.875 -48.115 ;
        RECT -36.205 -49.805 -35.875 -49.475 ;
        RECT -36.205 -51.165 -35.875 -50.835 ;
        RECT -36.205 -52.525 -35.875 -52.195 ;
        RECT -36.205 -53.885 -35.875 -53.555 ;
        RECT -36.205 -55.245 -35.875 -54.915 ;
        RECT -36.205 -56.605 -35.875 -56.275 ;
        RECT -36.205 -57.965 -35.875 -57.635 ;
        RECT -36.205 -59.325 -35.875 -58.995 ;
        RECT -36.205 -60.685 -35.875 -60.355 ;
        RECT -36.205 -62.045 -35.875 -61.715 ;
        RECT -36.205 -63.405 -35.875 -63.075 ;
        RECT -36.205 -64.765 -35.875 -64.435 ;
        RECT -36.205 -66.125 -35.875 -65.795 ;
        RECT -36.205 -67.485 -35.875 -67.155 ;
        RECT -36.205 -68.845 -35.875 -68.515 ;
        RECT -36.205 -70.205 -35.875 -69.875 ;
        RECT -36.205 -71.565 -35.875 -71.235 ;
        RECT -36.205 -72.925 -35.875 -72.595 ;
        RECT -36.205 -74.285 -35.875 -73.955 ;
        RECT -36.205 -75.645 -35.875 -75.315 ;
        RECT -36.205 -77.005 -35.875 -76.675 ;
        RECT -36.205 -78.365 -35.875 -78.035 ;
        RECT -36.205 -79.725 -35.875 -79.395 ;
        RECT -36.205 -81.085 -35.875 -80.755 ;
        RECT -36.205 -82.445 -35.875 -82.115 ;
        RECT -36.205 -83.805 -35.875 -83.475 ;
        RECT -36.205 -85.165 -35.875 -84.835 ;
        RECT -36.205 -86.525 -35.875 -86.195 ;
        RECT -36.205 -87.885 -35.875 -87.555 ;
        RECT -36.205 -89.245 -35.875 -88.915 ;
        RECT -36.205 -90.605 -35.875 -90.275 ;
        RECT -36.205 -91.965 -35.875 -91.635 ;
        RECT -36.205 -93.325 -35.875 -92.995 ;
        RECT -36.205 -94.685 -35.875 -94.355 ;
        RECT -36.205 -96.045 -35.875 -95.715 ;
        RECT -36.205 -97.405 -35.875 -97.075 ;
        RECT -36.205 -98.765 -35.875 -98.435 ;
        RECT -36.205 -100.125 -35.875 -99.795 ;
        RECT -36.205 -101.485 -35.875 -101.155 ;
        RECT -36.205 -102.845 -35.875 -102.515 ;
        RECT -36.205 -104.205 -35.875 -103.875 ;
        RECT -36.205 -105.565 -35.875 -105.235 ;
        RECT -36.205 -106.925 -35.875 -106.595 ;
        RECT -36.205 -108.285 -35.875 -107.955 ;
        RECT -36.205 -109.645 -35.875 -109.315 ;
        RECT -36.205 -111.005 -35.875 -110.675 ;
        RECT -36.205 -112.365 -35.875 -112.035 ;
        RECT -36.205 -113.725 -35.875 -113.395 ;
        RECT -36.205 -115.085 -35.875 -114.755 ;
        RECT -36.205 -116.445 -35.875 -116.115 ;
        RECT -36.205 -117.805 -35.875 -117.475 ;
        RECT -36.205 -119.165 -35.875 -118.835 ;
        RECT -36.205 -124.605 -35.875 -124.275 ;
        RECT -36.205 -128.685 -35.875 -128.355 ;
        RECT -36.205 -130.045 -35.875 -129.715 ;
        RECT -36.205 -132.765 -35.875 -132.435 ;
        RECT -36.205 -134.125 -35.875 -133.795 ;
        RECT -36.205 -135.485 -35.875 -135.155 ;
        RECT -36.205 -136.845 -35.875 -136.515 ;
        RECT -36.205 -138.205 -35.875 -137.875 ;
        RECT -36.205 -140.925 -35.875 -140.595 ;
        RECT -36.205 -142.285 -35.875 -141.955 ;
        RECT -36.205 -145.005 -35.875 -144.675 ;
        RECT -36.205 -146.365 -35.875 -146.035 ;
        RECT -36.205 -149.085 -35.875 -148.755 ;
        RECT -36.205 -150.445 -35.875 -150.115 ;
        RECT -36.205 -153.165 -35.875 -152.835 ;
        RECT -36.205 -154.525 -35.875 -154.195 ;
        RECT -36.205 -155.885 -35.875 -155.555 ;
        RECT -36.205 -157.245 -35.875 -156.915 ;
        RECT -36.205 -159.965 -35.875 -159.635 ;
        RECT -36.205 -162.685 -35.875 -162.355 ;
        RECT -36.205 -164.045 -35.875 -163.715 ;
        RECT -36.205 -165.405 -35.875 -165.075 ;
        RECT -36.205 -166.765 -35.875 -166.435 ;
        RECT -36.205 -168.125 -35.875 -167.795 ;
        RECT -36.205 -169.485 -35.875 -169.155 ;
        RECT -36.205 -170.845 -35.875 -170.515 ;
        RECT -36.205 -172.205 -35.875 -171.875 ;
        RECT -36.205 -173.565 -35.875 -173.235 ;
        RECT -36.205 -174.925 -35.875 -174.595 ;
        RECT -36.205 -176.285 -35.875 -175.955 ;
        RECT -36.205 -177.645 -35.875 -177.315 ;
        RECT -36.205 -179.005 -35.875 -178.675 ;
        RECT -36.205 -180.365 -35.875 -180.035 ;
        RECT -36.205 -181.725 -35.875 -181.395 ;
        RECT -36.205 -183.085 -35.875 -182.755 ;
        RECT -36.205 -184.445 -35.875 -184.115 ;
        RECT -36.205 -185.805 -35.875 -185.475 ;
        RECT -36.205 -187.165 -35.875 -186.835 ;
        RECT -36.205 -188.525 -35.875 -188.195 ;
        RECT -36.205 -189.885 -35.875 -189.555 ;
        RECT -36.205 -191.245 -35.875 -190.915 ;
        RECT -36.205 -192.605 -35.875 -192.275 ;
        RECT -36.205 -193.965 -35.875 -193.635 ;
        RECT -36.205 -195.325 -35.875 -194.995 ;
        RECT -36.205 -196.685 -35.875 -196.355 ;
        RECT -36.205 -198.045 -35.875 -197.715 ;
        RECT -36.205 -199.405 -35.875 -199.075 ;
        RECT -36.205 -200.765 -35.875 -200.435 ;
        RECT -36.205 -202.125 -35.875 -201.795 ;
        RECT -36.205 -203.485 -35.875 -203.155 ;
        RECT -36.205 -204.845 -35.875 -204.515 ;
        RECT -36.205 -206.205 -35.875 -205.875 ;
        RECT -36.205 -207.565 -35.875 -207.235 ;
        RECT -36.205 -208.925 -35.875 -208.595 ;
        RECT -36.205 -210.285 -35.875 -209.955 ;
        RECT -36.205 -211.645 -35.875 -211.315 ;
        RECT -36.205 -213.005 -35.875 -212.675 ;
        RECT -36.205 -214.365 -35.875 -214.035 ;
        RECT -36.205 -215.725 -35.875 -215.395 ;
        RECT -36.205 -217.085 -35.875 -216.755 ;
        RECT -36.205 -218.445 -35.875 -218.115 ;
        RECT -36.205 -219.805 -35.875 -219.475 ;
        RECT -36.205 -221.165 -35.875 -220.835 ;
        RECT -36.205 -222.525 -35.875 -222.195 ;
        RECT -36.205 -223.885 -35.875 -223.555 ;
        RECT -36.205 -225.245 -35.875 -224.915 ;
        RECT -36.205 -227.965 -35.875 -227.635 ;
        RECT -36.205 -232.045 -35.875 -231.715 ;
        RECT -36.205 -233.225 -35.875 -232.895 ;
        RECT -36.205 -234.765 -35.875 -234.435 ;
        RECT -36.205 -236.125 -35.875 -235.795 ;
        RECT -36.205 -237.485 -35.875 -237.155 ;
        RECT -36.205 -238.845 -35.875 -238.515 ;
        RECT -36.205 -241.09 -35.875 -239.96 ;
        RECT -36.2 -241.205 -35.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 244.04 -34.515 245.17 ;
        RECT -34.845 242.595 -34.515 242.925 ;
        RECT -34.845 241.235 -34.515 241.565 ;
        RECT -34.845 239.875 -34.515 240.205 ;
        RECT -34.845 238.515 -34.515 238.845 ;
        RECT -34.845 237.155 -34.515 237.485 ;
        RECT -34.845 235.795 -34.515 236.125 ;
        RECT -34.845 234.435 -34.515 234.765 ;
        RECT -34.845 233.075 -34.515 233.405 ;
        RECT -34.845 231.715 -34.515 232.045 ;
        RECT -34.845 230.355 -34.515 230.685 ;
        RECT -34.845 228.995 -34.515 229.325 ;
        RECT -34.845 227.635 -34.515 227.965 ;
        RECT -34.845 226.275 -34.515 226.605 ;
        RECT -34.845 224.915 -34.515 225.245 ;
        RECT -34.845 223.555 -34.515 223.885 ;
        RECT -34.845 222.195 -34.515 222.525 ;
        RECT -34.845 220.835 -34.515 221.165 ;
        RECT -34.845 219.475 -34.515 219.805 ;
        RECT -34.845 218.115 -34.515 218.445 ;
        RECT -34.845 216.755 -34.515 217.085 ;
        RECT -34.845 215.395 -34.515 215.725 ;
        RECT -34.845 214.035 -34.515 214.365 ;
        RECT -34.845 212.675 -34.515 213.005 ;
        RECT -34.845 211.315 -34.515 211.645 ;
        RECT -34.845 209.955 -34.515 210.285 ;
        RECT -34.845 208.595 -34.515 208.925 ;
        RECT -34.845 207.235 -34.515 207.565 ;
        RECT -34.845 205.875 -34.515 206.205 ;
        RECT -34.845 204.515 -34.515 204.845 ;
        RECT -34.845 203.155 -34.515 203.485 ;
        RECT -34.845 201.795 -34.515 202.125 ;
        RECT -34.845 200.435 -34.515 200.765 ;
        RECT -34.845 199.075 -34.515 199.405 ;
        RECT -34.845 197.715 -34.515 198.045 ;
        RECT -34.845 196.355 -34.515 196.685 ;
        RECT -34.845 194.995 -34.515 195.325 ;
        RECT -34.845 193.635 -34.515 193.965 ;
        RECT -34.845 192.275 -34.515 192.605 ;
        RECT -34.845 190.915 -34.515 191.245 ;
        RECT -34.845 189.555 -34.515 189.885 ;
        RECT -34.845 188.195 -34.515 188.525 ;
        RECT -34.845 186.835 -34.515 187.165 ;
        RECT -34.845 185.475 -34.515 185.805 ;
        RECT -34.845 184.115 -34.515 184.445 ;
        RECT -34.845 182.755 -34.515 183.085 ;
        RECT -34.845 181.395 -34.515 181.725 ;
        RECT -34.845 180.035 -34.515 180.365 ;
        RECT -34.845 178.675 -34.515 179.005 ;
        RECT -34.845 177.315 -34.515 177.645 ;
        RECT -34.845 175.955 -34.515 176.285 ;
        RECT -34.845 174.595 -34.515 174.925 ;
        RECT -34.845 173.235 -34.515 173.565 ;
        RECT -34.845 171.875 -34.515 172.205 ;
        RECT -34.845 170.515 -34.515 170.845 ;
        RECT -34.845 169.155 -34.515 169.485 ;
        RECT -34.845 167.795 -34.515 168.125 ;
        RECT -34.845 166.435 -34.515 166.765 ;
        RECT -34.845 165.075 -34.515 165.405 ;
        RECT -34.845 163.715 -34.515 164.045 ;
        RECT -34.845 162.355 -34.515 162.685 ;
        RECT -34.845 160.995 -34.515 161.325 ;
        RECT -34.845 159.635 -34.515 159.965 ;
        RECT -34.845 158.275 -34.515 158.605 ;
        RECT -34.845 156.915 -34.515 157.245 ;
        RECT -34.845 155.555 -34.515 155.885 ;
        RECT -34.845 154.195 -34.515 154.525 ;
        RECT -34.845 152.835 -34.515 153.165 ;
        RECT -34.845 151.475 -34.515 151.805 ;
        RECT -34.845 150.115 -34.515 150.445 ;
        RECT -34.845 148.755 -34.515 149.085 ;
        RECT -34.845 147.395 -34.515 147.725 ;
        RECT -34.845 146.035 -34.515 146.365 ;
        RECT -34.845 144.675 -34.515 145.005 ;
        RECT -34.845 143.315 -34.515 143.645 ;
        RECT -34.845 141.955 -34.515 142.285 ;
        RECT -34.845 140.595 -34.515 140.925 ;
        RECT -34.845 139.235 -34.515 139.565 ;
        RECT -34.845 137.875 -34.515 138.205 ;
        RECT -34.845 136.515 -34.515 136.845 ;
        RECT -34.845 135.155 -34.515 135.485 ;
        RECT -34.845 133.795 -34.515 134.125 ;
        RECT -34.845 132.435 -34.515 132.765 ;
        RECT -34.845 131.075 -34.515 131.405 ;
        RECT -34.845 129.715 -34.515 130.045 ;
        RECT -34.845 128.355 -34.515 128.685 ;
        RECT -34.845 126.995 -34.515 127.325 ;
        RECT -34.845 125.635 -34.515 125.965 ;
        RECT -34.845 124.275 -34.515 124.605 ;
        RECT -34.845 122.915 -34.515 123.245 ;
        RECT -34.845 121.555 -34.515 121.885 ;
        RECT -34.845 120.195 -34.515 120.525 ;
        RECT -34.845 118.835 -34.515 119.165 ;
        RECT -34.845 117.475 -34.515 117.805 ;
        RECT -34.845 116.115 -34.515 116.445 ;
        RECT -34.845 114.755 -34.515 115.085 ;
        RECT -34.845 113.395 -34.515 113.725 ;
        RECT -34.845 112.035 -34.515 112.365 ;
        RECT -34.845 110.675 -34.515 111.005 ;
        RECT -34.845 109.315 -34.515 109.645 ;
        RECT -34.845 107.955 -34.515 108.285 ;
        RECT -34.845 106.595 -34.515 106.925 ;
        RECT -34.845 105.235 -34.515 105.565 ;
        RECT -34.845 103.875 -34.515 104.205 ;
        RECT -34.845 102.515 -34.515 102.845 ;
        RECT -34.845 101.155 -34.515 101.485 ;
        RECT -34.845 99.795 -34.515 100.125 ;
        RECT -34.845 98.435 -34.515 98.765 ;
        RECT -34.845 97.075 -34.515 97.405 ;
        RECT -34.845 95.715 -34.515 96.045 ;
        RECT -34.845 94.355 -34.515 94.685 ;
        RECT -34.845 92.995 -34.515 93.325 ;
        RECT -34.845 91.635 -34.515 91.965 ;
        RECT -34.845 90.275 -34.515 90.605 ;
        RECT -34.845 88.915 -34.515 89.245 ;
        RECT -34.845 87.555 -34.515 87.885 ;
        RECT -34.845 86.195 -34.515 86.525 ;
        RECT -34.845 84.835 -34.515 85.165 ;
        RECT -34.845 83.475 -34.515 83.805 ;
        RECT -34.845 82.115 -34.515 82.445 ;
        RECT -34.845 80.755 -34.515 81.085 ;
        RECT -34.845 79.395 -34.515 79.725 ;
        RECT -34.845 78.035 -34.515 78.365 ;
        RECT -34.845 76.675 -34.515 77.005 ;
        RECT -34.845 75.315 -34.515 75.645 ;
        RECT -34.845 73.955 -34.515 74.285 ;
        RECT -34.845 72.595 -34.515 72.925 ;
        RECT -34.845 71.235 -34.515 71.565 ;
        RECT -34.845 69.875 -34.515 70.205 ;
        RECT -34.845 68.515 -34.515 68.845 ;
        RECT -34.845 67.155 -34.515 67.485 ;
        RECT -34.845 65.795 -34.515 66.125 ;
        RECT -34.845 64.435 -34.515 64.765 ;
        RECT -34.845 63.075 -34.515 63.405 ;
        RECT -34.845 61.715 -34.515 62.045 ;
        RECT -34.845 60.355 -34.515 60.685 ;
        RECT -34.845 58.995 -34.515 59.325 ;
        RECT -34.845 57.635 -34.515 57.965 ;
        RECT -34.845 56.275 -34.515 56.605 ;
        RECT -34.845 54.915 -34.515 55.245 ;
        RECT -34.845 53.555 -34.515 53.885 ;
        RECT -34.845 52.195 -34.515 52.525 ;
        RECT -34.845 50.835 -34.515 51.165 ;
        RECT -34.845 49.475 -34.515 49.805 ;
        RECT -34.845 48.115 -34.515 48.445 ;
        RECT -34.845 46.755 -34.515 47.085 ;
        RECT -34.845 45.395 -34.515 45.725 ;
        RECT -34.845 44.035 -34.515 44.365 ;
        RECT -34.845 42.675 -34.515 43.005 ;
        RECT -34.845 41.315 -34.515 41.645 ;
        RECT -34.845 39.955 -34.515 40.285 ;
        RECT -34.845 38.595 -34.515 38.925 ;
        RECT -34.845 37.235 -34.515 37.565 ;
        RECT -34.845 35.875 -34.515 36.205 ;
        RECT -34.845 34.515 -34.515 34.845 ;
        RECT -34.845 33.155 -34.515 33.485 ;
        RECT -34.845 31.795 -34.515 32.125 ;
        RECT -34.845 30.435 -34.515 30.765 ;
        RECT -34.845 29.075 -34.515 29.405 ;
        RECT -34.845 27.715 -34.515 28.045 ;
        RECT -34.845 26.355 -34.515 26.685 ;
        RECT -34.845 24.995 -34.515 25.325 ;
        RECT -34.845 23.635 -34.515 23.965 ;
        RECT -34.845 22.275 -34.515 22.605 ;
        RECT -34.845 20.915 -34.515 21.245 ;
        RECT -34.845 19.555 -34.515 19.885 ;
        RECT -34.845 18.195 -34.515 18.525 ;
        RECT -34.845 16.835 -34.515 17.165 ;
        RECT -34.845 15.475 -34.515 15.805 ;
        RECT -34.845 14.115 -34.515 14.445 ;
        RECT -34.845 12.755 -34.515 13.085 ;
        RECT -34.845 11.395 -34.515 11.725 ;
        RECT -34.845 10.035 -34.515 10.365 ;
        RECT -34.845 8.675 -34.515 9.005 ;
        RECT -34.845 7.315 -34.515 7.645 ;
        RECT -34.845 5.955 -34.515 6.285 ;
        RECT -34.845 4.595 -34.515 4.925 ;
        RECT -34.845 3.235 -34.515 3.565 ;
        RECT -34.845 1.875 -34.515 2.205 ;
        RECT -34.845 0.515 -34.515 0.845 ;
        RECT -34.845 -2.205 -34.515 -1.875 ;
        RECT -34.845 -3.565 -34.515 -3.235 ;
        RECT -34.845 -7.645 -34.515 -7.315 ;
        RECT -34.845 -9.005 -34.515 -8.675 ;
        RECT -34.845 -10.365 -34.515 -10.035 ;
        RECT -34.845 -11.725 -34.515 -11.395 ;
        RECT -34.845 -13.085 -34.515 -12.755 ;
        RECT -34.845 -14.445 -34.515 -14.115 ;
        RECT -34.845 -15.805 -34.515 -15.475 ;
        RECT -34.845 -17.165 -34.515 -16.835 ;
        RECT -34.845 -18.525 -34.515 -18.195 ;
        RECT -34.845 -19.885 -34.515 -19.555 ;
        RECT -34.845 -21.245 -34.515 -20.915 ;
        RECT -34.845 -22.605 -34.515 -22.275 ;
        RECT -34.845 -29.405 -34.515 -29.075 ;
        RECT -34.845 -32.125 -34.515 -31.795 ;
        RECT -34.845 -33.485 -34.515 -33.155 ;
        RECT -34.845 -34.88 -34.515 -34.55 ;
        RECT -34.845 -36.205 -34.515 -35.875 ;
        RECT -34.845 -38.925 -34.515 -38.595 ;
        RECT -34.845 -39.97 -34.515 -39.64 ;
        RECT -34.845 -48.445 -34.515 -48.115 ;
        RECT -34.845 -49.805 -34.515 -49.475 ;
        RECT -34.845 -51.165 -34.515 -50.835 ;
        RECT -34.845 -53.885 -34.515 -53.555 ;
        RECT -34.845 -57.965 -34.515 -57.635 ;
        RECT -34.845 -62.045 -34.515 -61.715 ;
        RECT -34.845 -63.405 -34.515 -63.075 ;
        RECT -34.845 -64.765 -34.515 -64.435 ;
        RECT -34.845 -66.125 -34.515 -65.795 ;
        RECT -34.845 -67.485 -34.515 -67.155 ;
        RECT -34.845 -68.845 -34.515 -68.515 ;
        RECT -34.845 -70.205 -34.515 -69.875 ;
        RECT -34.845 -71.565 -34.515 -71.235 ;
        RECT -34.845 -72.925 -34.515 -72.595 ;
        RECT -34.845 -74.285 -34.515 -73.955 ;
        RECT -34.845 -75.645 -34.515 -75.315 ;
        RECT -34.845 -77.005 -34.515 -76.675 ;
        RECT -34.845 -78.365 -34.515 -78.035 ;
        RECT -34.845 -79.725 -34.515 -79.395 ;
        RECT -34.845 -81.085 -34.515 -80.755 ;
        RECT -34.845 -82.445 -34.515 -82.115 ;
        RECT -34.845 -83.805 -34.515 -83.475 ;
        RECT -34.845 -85.165 -34.515 -84.835 ;
        RECT -34.845 -86.525 -34.515 -86.195 ;
        RECT -34.845 -87.885 -34.515 -87.555 ;
        RECT -34.845 -89.245 -34.515 -88.915 ;
        RECT -34.845 -90.605 -34.515 -90.275 ;
        RECT -34.845 -91.965 -34.515 -91.635 ;
        RECT -34.845 -93.325 -34.515 -92.995 ;
        RECT -34.845 -94.685 -34.515 -94.355 ;
        RECT -34.845 -96.045 -34.515 -95.715 ;
        RECT -34.845 -97.405 -34.515 -97.075 ;
        RECT -34.845 -98.765 -34.515 -98.435 ;
        RECT -34.845 -100.125 -34.515 -99.795 ;
        RECT -34.845 -101.485 -34.515 -101.155 ;
        RECT -34.845 -102.845 -34.515 -102.515 ;
        RECT -34.845 -104.205 -34.515 -103.875 ;
        RECT -34.845 -105.565 -34.515 -105.235 ;
        RECT -34.845 -106.925 -34.515 -106.595 ;
        RECT -34.845 -108.285 -34.515 -107.955 ;
        RECT -34.845 -109.645 -34.515 -109.315 ;
        RECT -34.845 -111.005 -34.515 -110.675 ;
        RECT -34.845 -112.365 -34.515 -112.035 ;
        RECT -34.845 -113.725 -34.515 -113.395 ;
        RECT -34.845 -115.085 -34.515 -114.755 ;
        RECT -34.845 -116.445 -34.515 -116.115 ;
        RECT -34.845 -117.805 -34.515 -117.475 ;
        RECT -34.845 -119.165 -34.515 -118.835 ;
        RECT -34.845 -124.605 -34.515 -124.275 ;
        RECT -34.845 -128.685 -34.515 -128.355 ;
        RECT -34.845 -130.045 -34.515 -129.715 ;
        RECT -34.845 -131.405 -34.515 -131.075 ;
        RECT -34.845 -132.765 -34.515 -132.435 ;
        RECT -34.845 -134.125 -34.515 -133.795 ;
        RECT -34.845 -135.485 -34.515 -135.155 ;
        RECT -34.845 -136.845 -34.515 -136.515 ;
        RECT -34.845 -138.205 -34.515 -137.875 ;
        RECT -34.845 -139.565 -34.515 -139.235 ;
        RECT -34.845 -140.925 -34.515 -140.595 ;
        RECT -34.845 -142.285 -34.515 -141.955 ;
        RECT -34.845 -143.645 -34.515 -143.315 ;
        RECT -34.845 -145.005 -34.515 -144.675 ;
        RECT -34.845 -146.365 -34.515 -146.035 ;
        RECT -34.845 -147.725 -34.515 -147.395 ;
        RECT -34.845 -149.085 -34.515 -148.755 ;
        RECT -34.845 -150.445 -34.515 -150.115 ;
        RECT -34.845 -151.805 -34.515 -151.475 ;
        RECT -34.845 -153.165 -34.515 -152.835 ;
        RECT -34.845 -154.525 -34.515 -154.195 ;
        RECT -34.845 -155.885 -34.515 -155.555 ;
        RECT -34.845 -157.245 -34.515 -156.915 ;
        RECT -34.845 -159.965 -34.515 -159.635 ;
        RECT -34.845 -162.685 -34.515 -162.355 ;
        RECT -34.845 -164.045 -34.515 -163.715 ;
        RECT -34.845 -165.405 -34.515 -165.075 ;
        RECT -34.845 -166.765 -34.515 -166.435 ;
        RECT -34.845 -168.125 -34.515 -167.795 ;
        RECT -34.845 -169.485 -34.515 -169.155 ;
        RECT -34.845 -170.845 -34.515 -170.515 ;
        RECT -34.845 -172.205 -34.515 -171.875 ;
        RECT -34.845 -173.565 -34.515 -173.235 ;
        RECT -34.845 -174.925 -34.515 -174.595 ;
        RECT -34.845 -176.285 -34.515 -175.955 ;
        RECT -34.845 -177.645 -34.515 -177.315 ;
        RECT -34.845 -179.005 -34.515 -178.675 ;
        RECT -34.845 -180.365 -34.515 -180.035 ;
        RECT -34.845 -181.725 -34.515 -181.395 ;
        RECT -34.845 -183.085 -34.515 -182.755 ;
        RECT -34.845 -184.445 -34.515 -184.115 ;
        RECT -34.845 -185.805 -34.515 -185.475 ;
        RECT -34.845 -187.165 -34.515 -186.835 ;
        RECT -34.845 -188.525 -34.515 -188.195 ;
        RECT -34.845 -189.885 -34.515 -189.555 ;
        RECT -34.845 -191.245 -34.515 -190.915 ;
        RECT -34.845 -192.605 -34.515 -192.275 ;
        RECT -34.845 -193.965 -34.515 -193.635 ;
        RECT -34.845 -195.325 -34.515 -194.995 ;
        RECT -34.845 -196.685 -34.515 -196.355 ;
        RECT -34.845 -198.045 -34.515 -197.715 ;
        RECT -34.845 -199.405 -34.515 -199.075 ;
        RECT -34.845 -200.765 -34.515 -200.435 ;
        RECT -34.845 -202.125 -34.515 -201.795 ;
        RECT -34.845 -203.485 -34.515 -203.155 ;
        RECT -34.845 -204.845 -34.515 -204.515 ;
        RECT -34.845 -206.205 -34.515 -205.875 ;
        RECT -34.845 -208.925 -34.515 -208.595 ;
        RECT -34.845 -210.285 -34.515 -209.955 ;
        RECT -34.845 -211.645 -34.515 -211.315 ;
        RECT -34.845 -213.005 -34.515 -212.675 ;
        RECT -34.845 -215.725 -34.515 -215.395 ;
        RECT -34.845 -217.085 -34.515 -216.755 ;
        RECT -34.845 -218.445 -34.515 -218.115 ;
        RECT -34.845 -219.805 -34.515 -219.475 ;
        RECT -34.845 -221.165 -34.515 -220.835 ;
        RECT -34.845 -222.525 -34.515 -222.195 ;
        RECT -34.845 -223.885 -34.515 -223.555 ;
        RECT -34.845 -225.245 -34.515 -224.915 ;
        RECT -34.845 -227.965 -34.515 -227.635 ;
        RECT -34.845 -232.045 -34.515 -231.715 ;
        RECT -34.845 -233.225 -34.515 -232.895 ;
        RECT -34.845 -234.765 -34.515 -234.435 ;
        RECT -34.845 -236.125 -34.515 -235.795 ;
        RECT -34.845 -237.485 -34.515 -237.155 ;
        RECT -34.845 -238.845 -34.515 -238.515 ;
        RECT -34.845 -241.09 -34.515 -239.96 ;
        RECT -34.84 -241.205 -34.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.485 -147.725 -33.155 -147.395 ;
        RECT -33.485 -149.085 -33.155 -148.755 ;
        RECT -33.485 -150.445 -33.155 -150.115 ;
        RECT -33.485 -151.805 -33.155 -151.475 ;
        RECT -33.485 -153.165 -33.155 -152.835 ;
        RECT -33.485 -154.525 -33.155 -154.195 ;
        RECT -33.485 -155.885 -33.155 -155.555 ;
        RECT -33.485 -157.245 -33.155 -156.915 ;
        RECT -33.485 -159.965 -33.155 -159.635 ;
        RECT -33.485 -162.685 -33.155 -162.355 ;
        RECT -33.485 -164.045 -33.155 -163.715 ;
        RECT -33.485 -165.405 -33.155 -165.075 ;
        RECT -33.485 -166.765 -33.155 -166.435 ;
        RECT -33.485 -168.125 -33.155 -167.795 ;
        RECT -33.485 -169.485 -33.155 -169.155 ;
        RECT -33.485 -170.845 -33.155 -170.515 ;
        RECT -33.485 -172.205 -33.155 -171.875 ;
        RECT -33.485 -173.565 -33.155 -173.235 ;
        RECT -33.485 -174.925 -33.155 -174.595 ;
        RECT -33.485 -176.285 -33.155 -175.955 ;
        RECT -33.485 -177.645 -33.155 -177.315 ;
        RECT -33.485 -179.005 -33.155 -178.675 ;
        RECT -33.485 -180.365 -33.155 -180.035 ;
        RECT -33.485 -181.725 -33.155 -181.395 ;
        RECT -33.485 -183.085 -33.155 -182.755 ;
        RECT -33.485 -184.445 -33.155 -184.115 ;
        RECT -33.485 -185.805 -33.155 -185.475 ;
        RECT -33.485 -187.165 -33.155 -186.835 ;
        RECT -33.485 -188.525 -33.155 -188.195 ;
        RECT -33.485 -191.245 -33.155 -190.915 ;
        RECT -33.485 -192.605 -33.155 -192.275 ;
        RECT -33.485 -193.965 -33.155 -193.635 ;
        RECT -33.485 -195.325 -33.155 -194.995 ;
        RECT -33.485 -196.685 -33.155 -196.355 ;
        RECT -33.485 -198.045 -33.155 -197.715 ;
        RECT -33.485 -199.405 -33.155 -199.075 ;
        RECT -33.485 -200.765 -33.155 -200.435 ;
        RECT -33.485 -202.125 -33.155 -201.795 ;
        RECT -33.485 -203.485 -33.155 -203.155 ;
        RECT -33.485 -204.845 -33.155 -204.515 ;
        RECT -33.485 -206.205 -33.155 -205.875 ;
        RECT -33.485 -208.925 -33.155 -208.595 ;
        RECT -33.485 -210.285 -33.155 -209.955 ;
        RECT -33.485 -213.005 -33.155 -212.675 ;
        RECT -33.485 -215.725 -33.155 -215.395 ;
        RECT -33.485 -217.085 -33.155 -216.755 ;
        RECT -33.485 -218.445 -33.155 -218.115 ;
        RECT -33.485 -219.805 -33.155 -219.475 ;
        RECT -33.485 -221.165 -33.155 -220.835 ;
        RECT -33.485 -222.525 -33.155 -222.195 ;
        RECT -33.485 -223.885 -33.155 -223.555 ;
        RECT -33.485 -225.245 -33.155 -224.915 ;
        RECT -33.485 -227.965 -33.155 -227.635 ;
        RECT -33.485 -232.045 -33.155 -231.715 ;
        RECT -33.485 -233.225 -33.155 -232.895 ;
        RECT -33.485 -234.765 -33.155 -234.435 ;
        RECT -33.485 -236.125 -33.155 -235.795 ;
        RECT -33.485 -237.485 -33.155 -237.155 ;
        RECT -33.485 -238.845 -33.155 -238.515 ;
        RECT -33.485 -241.09 -33.155 -239.96 ;
        RECT -33.48 -241.205 -33.16 245.285 ;
        RECT -33.485 244.04 -33.155 245.17 ;
        RECT -33.485 242.595 -33.155 242.925 ;
        RECT -33.485 241.235 -33.155 241.565 ;
        RECT -33.485 239.875 -33.155 240.205 ;
        RECT -33.485 238.515 -33.155 238.845 ;
        RECT -33.485 237.155 -33.155 237.485 ;
        RECT -33.485 235.795 -33.155 236.125 ;
        RECT -33.485 234.435 -33.155 234.765 ;
        RECT -33.485 233.075 -33.155 233.405 ;
        RECT -33.485 231.715 -33.155 232.045 ;
        RECT -33.485 230.355 -33.155 230.685 ;
        RECT -33.485 228.995 -33.155 229.325 ;
        RECT -33.485 227.635 -33.155 227.965 ;
        RECT -33.485 226.275 -33.155 226.605 ;
        RECT -33.485 224.915 -33.155 225.245 ;
        RECT -33.485 223.555 -33.155 223.885 ;
        RECT -33.485 222.195 -33.155 222.525 ;
        RECT -33.485 220.835 -33.155 221.165 ;
        RECT -33.485 219.475 -33.155 219.805 ;
        RECT -33.485 218.115 -33.155 218.445 ;
        RECT -33.485 216.755 -33.155 217.085 ;
        RECT -33.485 215.395 -33.155 215.725 ;
        RECT -33.485 214.035 -33.155 214.365 ;
        RECT -33.485 212.675 -33.155 213.005 ;
        RECT -33.485 211.315 -33.155 211.645 ;
        RECT -33.485 209.955 -33.155 210.285 ;
        RECT -33.485 208.595 -33.155 208.925 ;
        RECT -33.485 207.235 -33.155 207.565 ;
        RECT -33.485 205.875 -33.155 206.205 ;
        RECT -33.485 204.515 -33.155 204.845 ;
        RECT -33.485 203.155 -33.155 203.485 ;
        RECT -33.485 201.795 -33.155 202.125 ;
        RECT -33.485 200.435 -33.155 200.765 ;
        RECT -33.485 199.075 -33.155 199.405 ;
        RECT -33.485 197.715 -33.155 198.045 ;
        RECT -33.485 196.355 -33.155 196.685 ;
        RECT -33.485 194.995 -33.155 195.325 ;
        RECT -33.485 193.635 -33.155 193.965 ;
        RECT -33.485 192.275 -33.155 192.605 ;
        RECT -33.485 190.915 -33.155 191.245 ;
        RECT -33.485 189.555 -33.155 189.885 ;
        RECT -33.485 188.195 -33.155 188.525 ;
        RECT -33.485 186.835 -33.155 187.165 ;
        RECT -33.485 185.475 -33.155 185.805 ;
        RECT -33.485 184.115 -33.155 184.445 ;
        RECT -33.485 182.755 -33.155 183.085 ;
        RECT -33.485 181.395 -33.155 181.725 ;
        RECT -33.485 180.035 -33.155 180.365 ;
        RECT -33.485 178.675 -33.155 179.005 ;
        RECT -33.485 177.315 -33.155 177.645 ;
        RECT -33.485 175.955 -33.155 176.285 ;
        RECT -33.485 174.595 -33.155 174.925 ;
        RECT -33.485 173.235 -33.155 173.565 ;
        RECT -33.485 171.875 -33.155 172.205 ;
        RECT -33.485 170.515 -33.155 170.845 ;
        RECT -33.485 169.155 -33.155 169.485 ;
        RECT -33.485 167.795 -33.155 168.125 ;
        RECT -33.485 166.435 -33.155 166.765 ;
        RECT -33.485 165.075 -33.155 165.405 ;
        RECT -33.485 163.715 -33.155 164.045 ;
        RECT -33.485 162.355 -33.155 162.685 ;
        RECT -33.485 160.995 -33.155 161.325 ;
        RECT -33.485 159.635 -33.155 159.965 ;
        RECT -33.485 158.275 -33.155 158.605 ;
        RECT -33.485 156.915 -33.155 157.245 ;
        RECT -33.485 155.555 -33.155 155.885 ;
        RECT -33.485 154.195 -33.155 154.525 ;
        RECT -33.485 152.835 -33.155 153.165 ;
        RECT -33.485 151.475 -33.155 151.805 ;
        RECT -33.485 150.115 -33.155 150.445 ;
        RECT -33.485 148.755 -33.155 149.085 ;
        RECT -33.485 147.395 -33.155 147.725 ;
        RECT -33.485 146.035 -33.155 146.365 ;
        RECT -33.485 144.675 -33.155 145.005 ;
        RECT -33.485 143.315 -33.155 143.645 ;
        RECT -33.485 141.955 -33.155 142.285 ;
        RECT -33.485 140.595 -33.155 140.925 ;
        RECT -33.485 139.235 -33.155 139.565 ;
        RECT -33.485 137.875 -33.155 138.205 ;
        RECT -33.485 136.515 -33.155 136.845 ;
        RECT -33.485 135.155 -33.155 135.485 ;
        RECT -33.485 133.795 -33.155 134.125 ;
        RECT -33.485 132.435 -33.155 132.765 ;
        RECT -33.485 131.075 -33.155 131.405 ;
        RECT -33.485 129.715 -33.155 130.045 ;
        RECT -33.485 128.355 -33.155 128.685 ;
        RECT -33.485 126.995 -33.155 127.325 ;
        RECT -33.485 125.635 -33.155 125.965 ;
        RECT -33.485 124.275 -33.155 124.605 ;
        RECT -33.485 122.915 -33.155 123.245 ;
        RECT -33.485 121.555 -33.155 121.885 ;
        RECT -33.485 120.195 -33.155 120.525 ;
        RECT -33.485 118.835 -33.155 119.165 ;
        RECT -33.485 117.475 -33.155 117.805 ;
        RECT -33.485 116.115 -33.155 116.445 ;
        RECT -33.485 114.755 -33.155 115.085 ;
        RECT -33.485 113.395 -33.155 113.725 ;
        RECT -33.485 112.035 -33.155 112.365 ;
        RECT -33.485 110.675 -33.155 111.005 ;
        RECT -33.485 109.315 -33.155 109.645 ;
        RECT -33.485 107.955 -33.155 108.285 ;
        RECT -33.485 106.595 -33.155 106.925 ;
        RECT -33.485 105.235 -33.155 105.565 ;
        RECT -33.485 103.875 -33.155 104.205 ;
        RECT -33.485 102.515 -33.155 102.845 ;
        RECT -33.485 101.155 -33.155 101.485 ;
        RECT -33.485 99.795 -33.155 100.125 ;
        RECT -33.485 98.435 -33.155 98.765 ;
        RECT -33.485 97.075 -33.155 97.405 ;
        RECT -33.485 95.715 -33.155 96.045 ;
        RECT -33.485 94.355 -33.155 94.685 ;
        RECT -33.485 92.995 -33.155 93.325 ;
        RECT -33.485 91.635 -33.155 91.965 ;
        RECT -33.485 90.275 -33.155 90.605 ;
        RECT -33.485 88.915 -33.155 89.245 ;
        RECT -33.485 87.555 -33.155 87.885 ;
        RECT -33.485 86.195 -33.155 86.525 ;
        RECT -33.485 84.835 -33.155 85.165 ;
        RECT -33.485 83.475 -33.155 83.805 ;
        RECT -33.485 82.115 -33.155 82.445 ;
        RECT -33.485 80.755 -33.155 81.085 ;
        RECT -33.485 79.395 -33.155 79.725 ;
        RECT -33.485 78.035 -33.155 78.365 ;
        RECT -33.485 76.675 -33.155 77.005 ;
        RECT -33.485 75.315 -33.155 75.645 ;
        RECT -33.485 73.955 -33.155 74.285 ;
        RECT -33.485 72.595 -33.155 72.925 ;
        RECT -33.485 71.235 -33.155 71.565 ;
        RECT -33.485 69.875 -33.155 70.205 ;
        RECT -33.485 68.515 -33.155 68.845 ;
        RECT -33.485 67.155 -33.155 67.485 ;
        RECT -33.485 65.795 -33.155 66.125 ;
        RECT -33.485 64.435 -33.155 64.765 ;
        RECT -33.485 63.075 -33.155 63.405 ;
        RECT -33.485 61.715 -33.155 62.045 ;
        RECT -33.485 60.355 -33.155 60.685 ;
        RECT -33.485 58.995 -33.155 59.325 ;
        RECT -33.485 57.635 -33.155 57.965 ;
        RECT -33.485 56.275 -33.155 56.605 ;
        RECT -33.485 54.915 -33.155 55.245 ;
        RECT -33.485 53.555 -33.155 53.885 ;
        RECT -33.485 52.195 -33.155 52.525 ;
        RECT -33.485 50.835 -33.155 51.165 ;
        RECT -33.485 49.475 -33.155 49.805 ;
        RECT -33.485 48.115 -33.155 48.445 ;
        RECT -33.485 46.755 -33.155 47.085 ;
        RECT -33.485 45.395 -33.155 45.725 ;
        RECT -33.485 44.035 -33.155 44.365 ;
        RECT -33.485 42.675 -33.155 43.005 ;
        RECT -33.485 41.315 -33.155 41.645 ;
        RECT -33.485 39.955 -33.155 40.285 ;
        RECT -33.485 38.595 -33.155 38.925 ;
        RECT -33.485 37.235 -33.155 37.565 ;
        RECT -33.485 35.875 -33.155 36.205 ;
        RECT -33.485 34.515 -33.155 34.845 ;
        RECT -33.485 33.155 -33.155 33.485 ;
        RECT -33.485 31.795 -33.155 32.125 ;
        RECT -33.485 30.435 -33.155 30.765 ;
        RECT -33.485 29.075 -33.155 29.405 ;
        RECT -33.485 27.715 -33.155 28.045 ;
        RECT -33.485 26.355 -33.155 26.685 ;
        RECT -33.485 24.995 -33.155 25.325 ;
        RECT -33.485 23.635 -33.155 23.965 ;
        RECT -33.485 22.275 -33.155 22.605 ;
        RECT -33.485 20.915 -33.155 21.245 ;
        RECT -33.485 19.555 -33.155 19.885 ;
        RECT -33.485 18.195 -33.155 18.525 ;
        RECT -33.485 16.835 -33.155 17.165 ;
        RECT -33.485 15.475 -33.155 15.805 ;
        RECT -33.485 14.115 -33.155 14.445 ;
        RECT -33.485 12.755 -33.155 13.085 ;
        RECT -33.485 11.395 -33.155 11.725 ;
        RECT -33.485 10.035 -33.155 10.365 ;
        RECT -33.485 8.675 -33.155 9.005 ;
        RECT -33.485 7.315 -33.155 7.645 ;
        RECT -33.485 5.955 -33.155 6.285 ;
        RECT -33.485 4.595 -33.155 4.925 ;
        RECT -33.485 3.235 -33.155 3.565 ;
        RECT -33.485 1.875 -33.155 2.205 ;
        RECT -33.485 0.515 -33.155 0.845 ;
        RECT -33.485 -2.205 -33.155 -1.875 ;
        RECT -33.485 -7.645 -33.155 -7.315 ;
        RECT -33.485 -9.005 -33.155 -8.675 ;
        RECT -33.485 -10.365 -33.155 -10.035 ;
        RECT -33.485 -11.725 -33.155 -11.395 ;
        RECT -33.485 -13.085 -33.155 -12.755 ;
        RECT -33.485 -14.445 -33.155 -14.115 ;
        RECT -33.485 -15.805 -33.155 -15.475 ;
        RECT -33.485 -17.165 -33.155 -16.835 ;
        RECT -33.485 -18.525 -33.155 -18.195 ;
        RECT -33.485 -19.885 -33.155 -19.555 ;
        RECT -33.485 -21.245 -33.155 -20.915 ;
        RECT -33.485 -22.605 -33.155 -22.275 ;
        RECT -33.485 -29.405 -33.155 -29.075 ;
        RECT -33.485 -32.125 -33.155 -31.795 ;
        RECT -33.485 -33.485 -33.155 -33.155 ;
        RECT -33.485 -34.88 -33.155 -34.55 ;
        RECT -33.485 -36.205 -33.155 -35.875 ;
        RECT -33.485 -38.925 -33.155 -38.595 ;
        RECT -33.485 -39.97 -33.155 -39.64 ;
        RECT -33.485 -48.445 -33.155 -48.115 ;
        RECT -33.485 -49.805 -33.155 -49.475 ;
        RECT -33.485 -51.165 -33.155 -50.835 ;
        RECT -33.485 -53.885 -33.155 -53.555 ;
        RECT -33.485 -57.965 -33.155 -57.635 ;
        RECT -33.485 -62.045 -33.155 -61.715 ;
        RECT -33.485 -63.405 -33.155 -63.075 ;
        RECT -33.485 -64.765 -33.155 -64.435 ;
        RECT -33.485 -66.125 -33.155 -65.795 ;
        RECT -33.485 -67.485 -33.155 -67.155 ;
        RECT -33.485 -68.845 -33.155 -68.515 ;
        RECT -33.485 -70.205 -33.155 -69.875 ;
        RECT -33.485 -71.565 -33.155 -71.235 ;
        RECT -33.485 -72.925 -33.155 -72.595 ;
        RECT -33.485 -74.285 -33.155 -73.955 ;
        RECT -33.485 -75.645 -33.155 -75.315 ;
        RECT -33.485 -77.005 -33.155 -76.675 ;
        RECT -33.485 -78.365 -33.155 -78.035 ;
        RECT -33.485 -79.725 -33.155 -79.395 ;
        RECT -33.485 -81.085 -33.155 -80.755 ;
        RECT -33.485 -82.445 -33.155 -82.115 ;
        RECT -33.485 -83.805 -33.155 -83.475 ;
        RECT -33.485 -85.165 -33.155 -84.835 ;
        RECT -33.485 -86.525 -33.155 -86.195 ;
        RECT -33.485 -87.885 -33.155 -87.555 ;
        RECT -33.485 -89.245 -33.155 -88.915 ;
        RECT -33.485 -90.605 -33.155 -90.275 ;
        RECT -33.485 -91.965 -33.155 -91.635 ;
        RECT -33.485 -93.325 -33.155 -92.995 ;
        RECT -33.485 -94.685 -33.155 -94.355 ;
        RECT -33.485 -96.045 -33.155 -95.715 ;
        RECT -33.485 -97.405 -33.155 -97.075 ;
        RECT -33.485 -98.765 -33.155 -98.435 ;
        RECT -33.485 -100.125 -33.155 -99.795 ;
        RECT -33.485 -101.485 -33.155 -101.155 ;
        RECT -33.485 -102.845 -33.155 -102.515 ;
        RECT -33.485 -104.205 -33.155 -103.875 ;
        RECT -33.485 -105.565 -33.155 -105.235 ;
        RECT -33.485 -106.925 -33.155 -106.595 ;
        RECT -33.485 -108.285 -33.155 -107.955 ;
        RECT -33.485 -109.645 -33.155 -109.315 ;
        RECT -33.485 -111.005 -33.155 -110.675 ;
        RECT -33.485 -112.365 -33.155 -112.035 ;
        RECT -33.485 -113.725 -33.155 -113.395 ;
        RECT -33.485 -115.085 -33.155 -114.755 ;
        RECT -33.485 -116.445 -33.155 -116.115 ;
        RECT -33.485 -117.805 -33.155 -117.475 ;
        RECT -33.485 -119.165 -33.155 -118.835 ;
        RECT -33.485 -124.605 -33.155 -124.275 ;
        RECT -33.485 -128.685 -33.155 -128.355 ;
        RECT -33.485 -130.045 -33.155 -129.715 ;
        RECT -33.485 -131.405 -33.155 -131.075 ;
        RECT -33.485 -132.765 -33.155 -132.435 ;
        RECT -33.485 -134.125 -33.155 -133.795 ;
        RECT -33.485 -135.485 -33.155 -135.155 ;
        RECT -33.485 -136.845 -33.155 -136.515 ;
        RECT -33.485 -138.205 -33.155 -137.875 ;
        RECT -33.485 -139.565 -33.155 -139.235 ;
        RECT -33.485 -140.925 -33.155 -140.595 ;
        RECT -33.485 -142.285 -33.155 -141.955 ;
        RECT -33.485 -143.645 -33.155 -143.315 ;
        RECT -33.485 -145.005 -33.155 -144.675 ;
        RECT -33.485 -146.365 -33.155 -146.035 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 -128.685 -42.675 -128.355 ;
        RECT -43.005 -130.045 -42.675 -129.715 ;
        RECT -43.005 -132.765 -42.675 -132.435 ;
        RECT -43.005 -134.125 -42.675 -133.795 ;
        RECT -43.005 -135.485 -42.675 -135.155 ;
        RECT -43.005 -136.845 -42.675 -136.515 ;
        RECT -43.005 -138.205 -42.675 -137.875 ;
        RECT -43.005 -139.39 -42.675 -139.06 ;
        RECT -43.005 -140.925 -42.675 -140.595 ;
        RECT -43.005 -142.285 -42.675 -141.955 ;
        RECT -43.005 -145.005 -42.675 -144.675 ;
        RECT -43.005 -146.365 -42.675 -146.035 ;
        RECT -43.005 -148.03 -42.675 -147.7 ;
        RECT -43.005 -149.085 -42.675 -148.755 ;
        RECT -43.005 -150.445 -42.675 -150.115 ;
        RECT -43.005 -153.165 -42.675 -152.835 ;
        RECT -43.005 -154.525 -42.675 -154.195 ;
        RECT -43.005 -155.885 -42.675 -155.555 ;
        RECT -43.005 -157.245 -42.675 -156.915 ;
        RECT -43.005 -159.965 -42.675 -159.635 ;
        RECT -43.005 -162.685 -42.675 -162.355 ;
        RECT -43.005 -164.045 -42.675 -163.715 ;
        RECT -43.005 -165.405 -42.675 -165.075 ;
        RECT -43.005 -166.765 -42.675 -166.435 ;
        RECT -43.005 -168.125 -42.675 -167.795 ;
        RECT -43.005 -169.485 -42.675 -169.155 ;
        RECT -43.005 -170.845 -42.675 -170.515 ;
        RECT -43.005 -172.205 -42.675 -171.875 ;
        RECT -43.005 -173.565 -42.675 -173.235 ;
        RECT -43.005 -174.925 -42.675 -174.595 ;
        RECT -43.005 -176.285 -42.675 -175.955 ;
        RECT -43.005 -177.645 -42.675 -177.315 ;
        RECT -43.005 -179.005 -42.675 -178.675 ;
        RECT -43.005 -180.365 -42.675 -180.035 ;
        RECT -43.005 -181.725 -42.675 -181.395 ;
        RECT -43.005 -183.085 -42.675 -182.755 ;
        RECT -43.005 -184.445 -42.675 -184.115 ;
        RECT -43.005 -185.805 -42.675 -185.475 ;
        RECT -43.005 -187.165 -42.675 -186.835 ;
        RECT -43.005 -188.525 -42.675 -188.195 ;
        RECT -43.005 -189.885 -42.675 -189.555 ;
        RECT -43.005 -191.245 -42.675 -190.915 ;
        RECT -43.005 -192.605 -42.675 -192.275 ;
        RECT -43.005 -193.965 -42.675 -193.635 ;
        RECT -43.005 -195.325 -42.675 -194.995 ;
        RECT -43.005 -196.685 -42.675 -196.355 ;
        RECT -43.005 -198.045 -42.675 -197.715 ;
        RECT -43.005 -199.405 -42.675 -199.075 ;
        RECT -43.005 -200.765 -42.675 -200.435 ;
        RECT -43.005 -202.125 -42.675 -201.795 ;
        RECT -43.005 -203.485 -42.675 -203.155 ;
        RECT -43.005 -204.845 -42.675 -204.515 ;
        RECT -43.005 -206.205 -42.675 -205.875 ;
        RECT -43.005 -207.565 -42.675 -207.235 ;
        RECT -43.005 -208.925 -42.675 -208.595 ;
        RECT -43.005 -210.285 -42.675 -209.955 ;
        RECT -43.005 -211.645 -42.675 -211.315 ;
        RECT -43.005 -213.005 -42.675 -212.675 ;
        RECT -43.005 -214.365 -42.675 -214.035 ;
        RECT -43.005 -215.725 -42.675 -215.395 ;
        RECT -43.005 -217.085 -42.675 -216.755 ;
        RECT -43.005 -218.445 -42.675 -218.115 ;
        RECT -43.005 -219.805 -42.675 -219.475 ;
        RECT -43.005 -221.165 -42.675 -220.835 ;
        RECT -43.005 -222.525 -42.675 -222.195 ;
        RECT -43.005 -223.885 -42.675 -223.555 ;
        RECT -43.005 -225.245 -42.675 -224.915 ;
        RECT -43.005 -227.965 -42.675 -227.635 ;
        RECT -43.005 -230.685 -42.675 -230.355 ;
        RECT -43.005 -232.045 -42.675 -231.715 ;
        RECT -43.005 -233.225 -42.675 -232.895 ;
        RECT -43.005 -234.765 -42.675 -234.435 ;
        RECT -43.005 -236.125 -42.675 -235.795 ;
        RECT -43.005 -237.485 -42.675 -237.155 ;
        RECT -43.005 -238.845 -42.675 -238.515 ;
        RECT -43.005 -241.09 -42.675 -239.96 ;
        RECT -43 -241.205 -42.68 -124.96 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 244.04 -41.315 245.17 ;
        RECT -41.645 242.595 -41.315 242.925 ;
        RECT -41.645 241.235 -41.315 241.565 ;
        RECT -41.645 239.875 -41.315 240.205 ;
        RECT -41.645 238.515 -41.315 238.845 ;
        RECT -41.645 237.155 -41.315 237.485 ;
        RECT -41.645 235.795 -41.315 236.125 ;
        RECT -41.645 234.435 -41.315 234.765 ;
        RECT -41.645 233.075 -41.315 233.405 ;
        RECT -41.645 231.715 -41.315 232.045 ;
        RECT -41.645 230.355 -41.315 230.685 ;
        RECT -41.645 228.995 -41.315 229.325 ;
        RECT -41.645 227.635 -41.315 227.965 ;
        RECT -41.645 226.275 -41.315 226.605 ;
        RECT -41.645 224.915 -41.315 225.245 ;
        RECT -41.645 223.555 -41.315 223.885 ;
        RECT -41.645 222.195 -41.315 222.525 ;
        RECT -41.645 220.835 -41.315 221.165 ;
        RECT -41.645 219.475 -41.315 219.805 ;
        RECT -41.645 218.115 -41.315 218.445 ;
        RECT -41.645 216.755 -41.315 217.085 ;
        RECT -41.645 215.395 -41.315 215.725 ;
        RECT -41.645 214.035 -41.315 214.365 ;
        RECT -41.645 212.675 -41.315 213.005 ;
        RECT -41.645 211.315 -41.315 211.645 ;
        RECT -41.645 209.955 -41.315 210.285 ;
        RECT -41.645 208.595 -41.315 208.925 ;
        RECT -41.645 207.235 -41.315 207.565 ;
        RECT -41.645 205.875 -41.315 206.205 ;
        RECT -41.645 204.515 -41.315 204.845 ;
        RECT -41.645 203.155 -41.315 203.485 ;
        RECT -41.645 201.795 -41.315 202.125 ;
        RECT -41.645 200.435 -41.315 200.765 ;
        RECT -41.645 199.075 -41.315 199.405 ;
        RECT -41.645 197.715 -41.315 198.045 ;
        RECT -41.645 196.355 -41.315 196.685 ;
        RECT -41.645 194.995 -41.315 195.325 ;
        RECT -41.645 193.635 -41.315 193.965 ;
        RECT -41.645 192.275 -41.315 192.605 ;
        RECT -41.645 190.915 -41.315 191.245 ;
        RECT -41.645 189.555 -41.315 189.885 ;
        RECT -41.645 188.195 -41.315 188.525 ;
        RECT -41.645 186.835 -41.315 187.165 ;
        RECT -41.645 185.475 -41.315 185.805 ;
        RECT -41.645 184.115 -41.315 184.445 ;
        RECT -41.645 182.755 -41.315 183.085 ;
        RECT -41.645 181.395 -41.315 181.725 ;
        RECT -41.645 180.035 -41.315 180.365 ;
        RECT -41.645 178.675 -41.315 179.005 ;
        RECT -41.645 177.315 -41.315 177.645 ;
        RECT -41.645 175.955 -41.315 176.285 ;
        RECT -41.645 174.595 -41.315 174.925 ;
        RECT -41.645 173.235 -41.315 173.565 ;
        RECT -41.645 171.875 -41.315 172.205 ;
        RECT -41.645 170.515 -41.315 170.845 ;
        RECT -41.645 169.155 -41.315 169.485 ;
        RECT -41.645 167.795 -41.315 168.125 ;
        RECT -41.645 166.435 -41.315 166.765 ;
        RECT -41.645 165.075 -41.315 165.405 ;
        RECT -41.645 163.715 -41.315 164.045 ;
        RECT -41.645 162.355 -41.315 162.685 ;
        RECT -41.645 160.995 -41.315 161.325 ;
        RECT -41.645 159.635 -41.315 159.965 ;
        RECT -41.645 158.275 -41.315 158.605 ;
        RECT -41.645 156.915 -41.315 157.245 ;
        RECT -41.645 155.555 -41.315 155.885 ;
        RECT -41.645 154.195 -41.315 154.525 ;
        RECT -41.645 152.835 -41.315 153.165 ;
        RECT -41.645 151.475 -41.315 151.805 ;
        RECT -41.645 150.115 -41.315 150.445 ;
        RECT -41.645 148.755 -41.315 149.085 ;
        RECT -41.645 147.395 -41.315 147.725 ;
        RECT -41.645 146.035 -41.315 146.365 ;
        RECT -41.645 144.675 -41.315 145.005 ;
        RECT -41.645 143.315 -41.315 143.645 ;
        RECT -41.645 141.955 -41.315 142.285 ;
        RECT -41.645 140.595 -41.315 140.925 ;
        RECT -41.645 139.235 -41.315 139.565 ;
        RECT -41.645 137.875 -41.315 138.205 ;
        RECT -41.645 136.515 -41.315 136.845 ;
        RECT -41.645 135.155 -41.315 135.485 ;
        RECT -41.645 133.795 -41.315 134.125 ;
        RECT -41.645 132.435 -41.315 132.765 ;
        RECT -41.645 131.075 -41.315 131.405 ;
        RECT -41.645 129.715 -41.315 130.045 ;
        RECT -41.645 128.355 -41.315 128.685 ;
        RECT -41.645 126.995 -41.315 127.325 ;
        RECT -41.645 125.635 -41.315 125.965 ;
        RECT -41.645 124.275 -41.315 124.605 ;
        RECT -41.645 122.915 -41.315 123.245 ;
        RECT -41.645 121.555 -41.315 121.885 ;
        RECT -41.645 120.195 -41.315 120.525 ;
        RECT -41.645 118.835 -41.315 119.165 ;
        RECT -41.645 117.475 -41.315 117.805 ;
        RECT -41.645 116.115 -41.315 116.445 ;
        RECT -41.645 114.755 -41.315 115.085 ;
        RECT -41.645 113.395 -41.315 113.725 ;
        RECT -41.645 112.035 -41.315 112.365 ;
        RECT -41.645 110.675 -41.315 111.005 ;
        RECT -41.645 109.315 -41.315 109.645 ;
        RECT -41.645 107.955 -41.315 108.285 ;
        RECT -41.645 106.595 -41.315 106.925 ;
        RECT -41.645 105.235 -41.315 105.565 ;
        RECT -41.645 103.875 -41.315 104.205 ;
        RECT -41.645 102.515 -41.315 102.845 ;
        RECT -41.645 101.155 -41.315 101.485 ;
        RECT -41.645 99.795 -41.315 100.125 ;
        RECT -41.645 98.435 -41.315 98.765 ;
        RECT -41.645 97.075 -41.315 97.405 ;
        RECT -41.645 95.715 -41.315 96.045 ;
        RECT -41.645 94.355 -41.315 94.685 ;
        RECT -41.645 92.995 -41.315 93.325 ;
        RECT -41.645 91.635 -41.315 91.965 ;
        RECT -41.645 90.275 -41.315 90.605 ;
        RECT -41.645 88.915 -41.315 89.245 ;
        RECT -41.645 87.555 -41.315 87.885 ;
        RECT -41.645 86.195 -41.315 86.525 ;
        RECT -41.645 84.835 -41.315 85.165 ;
        RECT -41.645 83.475 -41.315 83.805 ;
        RECT -41.645 82.115 -41.315 82.445 ;
        RECT -41.645 80.755 -41.315 81.085 ;
        RECT -41.645 79.395 -41.315 79.725 ;
        RECT -41.645 78.035 -41.315 78.365 ;
        RECT -41.645 76.675 -41.315 77.005 ;
        RECT -41.645 75.315 -41.315 75.645 ;
        RECT -41.645 73.955 -41.315 74.285 ;
        RECT -41.645 72.595 -41.315 72.925 ;
        RECT -41.645 71.235 -41.315 71.565 ;
        RECT -41.645 69.875 -41.315 70.205 ;
        RECT -41.645 68.515 -41.315 68.845 ;
        RECT -41.645 67.155 -41.315 67.485 ;
        RECT -41.645 65.795 -41.315 66.125 ;
        RECT -41.645 64.435 -41.315 64.765 ;
        RECT -41.645 63.075 -41.315 63.405 ;
        RECT -41.645 61.715 -41.315 62.045 ;
        RECT -41.645 60.355 -41.315 60.685 ;
        RECT -41.645 58.995 -41.315 59.325 ;
        RECT -41.645 57.635 -41.315 57.965 ;
        RECT -41.645 56.275 -41.315 56.605 ;
        RECT -41.645 54.915 -41.315 55.245 ;
        RECT -41.645 53.555 -41.315 53.885 ;
        RECT -41.645 52.195 -41.315 52.525 ;
        RECT -41.645 50.835 -41.315 51.165 ;
        RECT -41.645 49.475 -41.315 49.805 ;
        RECT -41.645 48.115 -41.315 48.445 ;
        RECT -41.645 46.755 -41.315 47.085 ;
        RECT -41.645 45.395 -41.315 45.725 ;
        RECT -41.645 44.035 -41.315 44.365 ;
        RECT -41.645 42.675 -41.315 43.005 ;
        RECT -41.645 41.315 -41.315 41.645 ;
        RECT -41.645 39.955 -41.315 40.285 ;
        RECT -41.645 38.595 -41.315 38.925 ;
        RECT -41.645 37.235 -41.315 37.565 ;
        RECT -41.645 35.875 -41.315 36.205 ;
        RECT -41.645 34.515 -41.315 34.845 ;
        RECT -41.645 33.155 -41.315 33.485 ;
        RECT -41.645 31.795 -41.315 32.125 ;
        RECT -41.645 30.435 -41.315 30.765 ;
        RECT -41.645 29.075 -41.315 29.405 ;
        RECT -41.645 27.715 -41.315 28.045 ;
        RECT -41.645 26.355 -41.315 26.685 ;
        RECT -41.645 24.995 -41.315 25.325 ;
        RECT -41.645 23.635 -41.315 23.965 ;
        RECT -41.645 22.275 -41.315 22.605 ;
        RECT -41.645 20.915 -41.315 21.245 ;
        RECT -41.645 19.555 -41.315 19.885 ;
        RECT -41.645 18.195 -41.315 18.525 ;
        RECT -41.645 16.835 -41.315 17.165 ;
        RECT -41.645 15.475 -41.315 15.805 ;
        RECT -41.645 14.115 -41.315 14.445 ;
        RECT -41.645 12.755 -41.315 13.085 ;
        RECT -41.645 11.395 -41.315 11.725 ;
        RECT -41.645 10.035 -41.315 10.365 ;
        RECT -41.645 8.675 -41.315 9.005 ;
        RECT -41.645 7.315 -41.315 7.645 ;
        RECT -41.645 5.955 -41.315 6.285 ;
        RECT -41.645 4.595 -41.315 4.925 ;
        RECT -41.645 3.235 -41.315 3.565 ;
        RECT -41.645 1.875 -41.315 2.205 ;
        RECT -41.645 0.515 -41.315 0.845 ;
        RECT -41.645 -0.845 -41.315 -0.515 ;
        RECT -41.645 -6.285 -41.315 -5.955 ;
        RECT -41.645 -7.645 -41.315 -7.315 ;
        RECT -41.645 -9.005 -41.315 -8.675 ;
        RECT -41.645 -10.365 -41.315 -10.035 ;
        RECT -41.645 -11.725 -41.315 -11.395 ;
        RECT -41.645 -13.085 -41.315 -12.755 ;
        RECT -41.645 -14.445 -41.315 -14.115 ;
        RECT -41.645 -15.805 -41.315 -15.475 ;
        RECT -41.645 -17.165 -41.315 -16.835 ;
        RECT -41.645 -18.525 -41.315 -18.195 ;
        RECT -41.645 -19.885 -41.315 -19.555 ;
        RECT -41.645 -21.245 -41.315 -20.915 ;
        RECT -41.645 -22.605 -41.315 -22.275 ;
        RECT -41.645 -29.405 -41.315 -29.075 ;
        RECT -41.645 -32.125 -41.315 -31.795 ;
        RECT -41.645 -33.485 -41.315 -33.155 ;
        RECT -41.645 -34.88 -41.315 -34.55 ;
        RECT -41.645 -36.205 -41.315 -35.875 ;
        RECT -41.645 -38.925 -41.315 -38.595 ;
        RECT -41.645 -39.97 -41.315 -39.64 ;
        RECT -41.645 -48.445 -41.315 -48.115 ;
        RECT -41.645 -49.805 -41.315 -49.475 ;
        RECT -41.645 -51.165 -41.315 -50.835 ;
        RECT -41.645 -53.885 -41.315 -53.555 ;
        RECT -41.645 -57.965 -41.315 -57.635 ;
        RECT -41.645 -62.045 -41.315 -61.715 ;
        RECT -41.645 -63.405 -41.315 -63.075 ;
        RECT -41.645 -64.765 -41.315 -64.435 ;
        RECT -41.645 -66.125 -41.315 -65.795 ;
        RECT -41.645 -67.485 -41.315 -67.155 ;
        RECT -41.645 -68.845 -41.315 -68.515 ;
        RECT -41.645 -70.205 -41.315 -69.875 ;
        RECT -41.645 -71.565 -41.315 -71.235 ;
        RECT -41.645 -72.925 -41.315 -72.595 ;
        RECT -41.645 -74.285 -41.315 -73.955 ;
        RECT -41.645 -75.645 -41.315 -75.315 ;
        RECT -41.645 -77.005 -41.315 -76.675 ;
        RECT -41.645 -78.365 -41.315 -78.035 ;
        RECT -41.645 -79.725 -41.315 -79.395 ;
        RECT -41.645 -81.085 -41.315 -80.755 ;
        RECT -41.645 -82.445 -41.315 -82.115 ;
        RECT -41.645 -83.805 -41.315 -83.475 ;
        RECT -41.645 -85.165 -41.315 -84.835 ;
        RECT -41.645 -86.525 -41.315 -86.195 ;
        RECT -41.645 -87.885 -41.315 -87.555 ;
        RECT -41.645 -89.245 -41.315 -88.915 ;
        RECT -41.645 -90.605 -41.315 -90.275 ;
        RECT -41.645 -91.965 -41.315 -91.635 ;
        RECT -41.645 -93.325 -41.315 -92.995 ;
        RECT -41.645 -94.685 -41.315 -94.355 ;
        RECT -41.645 -96.045 -41.315 -95.715 ;
        RECT -41.645 -97.405 -41.315 -97.075 ;
        RECT -41.645 -98.765 -41.315 -98.435 ;
        RECT -41.645 -100.125 -41.315 -99.795 ;
        RECT -41.645 -101.485 -41.315 -101.155 ;
        RECT -41.645 -102.845 -41.315 -102.515 ;
        RECT -41.645 -104.205 -41.315 -103.875 ;
        RECT -41.645 -105.565 -41.315 -105.235 ;
        RECT -41.645 -106.925 -41.315 -106.595 ;
        RECT -41.645 -108.285 -41.315 -107.955 ;
        RECT -41.645 -109.645 -41.315 -109.315 ;
        RECT -41.645 -111.005 -41.315 -110.675 ;
        RECT -41.645 -112.365 -41.315 -112.035 ;
        RECT -41.645 -113.725 -41.315 -113.395 ;
        RECT -41.645 -115.085 -41.315 -114.755 ;
        RECT -41.645 -116.445 -41.315 -116.115 ;
        RECT -41.645 -117.805 -41.315 -117.475 ;
        RECT -41.645 -119.165 -41.315 -118.835 ;
        RECT -41.645 -120.525 -41.315 -120.195 ;
        RECT -41.645 -124.605 -41.315 -124.275 ;
        RECT -41.645 -128.685 -41.315 -128.355 ;
        RECT -41.645 -130.045 -41.315 -129.715 ;
        RECT -41.645 -132.765 -41.315 -132.435 ;
        RECT -41.645 -134.125 -41.315 -133.795 ;
        RECT -41.645 -135.485 -41.315 -135.155 ;
        RECT -41.645 -136.845 -41.315 -136.515 ;
        RECT -41.645 -138.205 -41.315 -137.875 ;
        RECT -41.645 -139.39 -41.315 -139.06 ;
        RECT -41.645 -140.925 -41.315 -140.595 ;
        RECT -41.645 -142.285 -41.315 -141.955 ;
        RECT -41.645 -145.005 -41.315 -144.675 ;
        RECT -41.645 -146.365 -41.315 -146.035 ;
        RECT -41.645 -148.03 -41.315 -147.7 ;
        RECT -41.645 -149.085 -41.315 -148.755 ;
        RECT -41.645 -150.445 -41.315 -150.115 ;
        RECT -41.64 -151.8 -41.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 -232.045 -41.315 -231.715 ;
        RECT -41.645 -234.765 -41.315 -234.435 ;
        RECT -41.645 -236.125 -41.315 -235.795 ;
        RECT -41.645 -237.485 -41.315 -237.155 ;
        RECT -41.645 -238.845 -41.315 -238.515 ;
        RECT -41.645 -241.09 -41.315 -239.96 ;
        RECT -41.64 -241.205 -41.32 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.285 244.04 -39.955 245.17 ;
        RECT -40.285 242.595 -39.955 242.925 ;
        RECT -40.285 241.235 -39.955 241.565 ;
        RECT -40.285 239.875 -39.955 240.205 ;
        RECT -40.285 238.515 -39.955 238.845 ;
        RECT -40.285 237.155 -39.955 237.485 ;
        RECT -40.285 235.795 -39.955 236.125 ;
        RECT -40.285 234.435 -39.955 234.765 ;
        RECT -40.285 233.075 -39.955 233.405 ;
        RECT -40.285 231.715 -39.955 232.045 ;
        RECT -40.285 230.355 -39.955 230.685 ;
        RECT -40.285 228.995 -39.955 229.325 ;
        RECT -40.285 227.635 -39.955 227.965 ;
        RECT -40.285 226.275 -39.955 226.605 ;
        RECT -40.285 224.915 -39.955 225.245 ;
        RECT -40.285 223.555 -39.955 223.885 ;
        RECT -40.285 222.195 -39.955 222.525 ;
        RECT -40.285 220.835 -39.955 221.165 ;
        RECT -40.285 219.475 -39.955 219.805 ;
        RECT -40.285 218.115 -39.955 218.445 ;
        RECT -40.285 216.755 -39.955 217.085 ;
        RECT -40.285 215.395 -39.955 215.725 ;
        RECT -40.285 214.035 -39.955 214.365 ;
        RECT -40.285 212.675 -39.955 213.005 ;
        RECT -40.285 211.315 -39.955 211.645 ;
        RECT -40.285 209.955 -39.955 210.285 ;
        RECT -40.285 208.595 -39.955 208.925 ;
        RECT -40.285 207.235 -39.955 207.565 ;
        RECT -40.285 205.875 -39.955 206.205 ;
        RECT -40.285 204.515 -39.955 204.845 ;
        RECT -40.285 203.155 -39.955 203.485 ;
        RECT -40.285 201.795 -39.955 202.125 ;
        RECT -40.285 200.435 -39.955 200.765 ;
        RECT -40.285 199.075 -39.955 199.405 ;
        RECT -40.285 197.715 -39.955 198.045 ;
        RECT -40.285 196.355 -39.955 196.685 ;
        RECT -40.285 194.995 -39.955 195.325 ;
        RECT -40.285 193.635 -39.955 193.965 ;
        RECT -40.285 192.275 -39.955 192.605 ;
        RECT -40.285 190.915 -39.955 191.245 ;
        RECT -40.285 189.555 -39.955 189.885 ;
        RECT -40.285 188.195 -39.955 188.525 ;
        RECT -40.285 186.835 -39.955 187.165 ;
        RECT -40.285 185.475 -39.955 185.805 ;
        RECT -40.285 184.115 -39.955 184.445 ;
        RECT -40.285 182.755 -39.955 183.085 ;
        RECT -40.285 181.395 -39.955 181.725 ;
        RECT -40.285 180.035 -39.955 180.365 ;
        RECT -40.285 178.675 -39.955 179.005 ;
        RECT -40.285 177.315 -39.955 177.645 ;
        RECT -40.285 175.955 -39.955 176.285 ;
        RECT -40.285 174.595 -39.955 174.925 ;
        RECT -40.285 173.235 -39.955 173.565 ;
        RECT -40.285 171.875 -39.955 172.205 ;
        RECT -40.285 170.515 -39.955 170.845 ;
        RECT -40.285 169.155 -39.955 169.485 ;
        RECT -40.285 167.795 -39.955 168.125 ;
        RECT -40.285 166.435 -39.955 166.765 ;
        RECT -40.285 165.075 -39.955 165.405 ;
        RECT -40.285 163.715 -39.955 164.045 ;
        RECT -40.285 162.355 -39.955 162.685 ;
        RECT -40.285 160.995 -39.955 161.325 ;
        RECT -40.285 159.635 -39.955 159.965 ;
        RECT -40.285 158.275 -39.955 158.605 ;
        RECT -40.285 156.915 -39.955 157.245 ;
        RECT -40.285 155.555 -39.955 155.885 ;
        RECT -40.285 154.195 -39.955 154.525 ;
        RECT -40.285 152.835 -39.955 153.165 ;
        RECT -40.285 151.475 -39.955 151.805 ;
        RECT -40.285 150.115 -39.955 150.445 ;
        RECT -40.285 148.755 -39.955 149.085 ;
        RECT -40.285 147.395 -39.955 147.725 ;
        RECT -40.285 146.035 -39.955 146.365 ;
        RECT -40.285 144.675 -39.955 145.005 ;
        RECT -40.285 143.315 -39.955 143.645 ;
        RECT -40.285 141.955 -39.955 142.285 ;
        RECT -40.285 140.595 -39.955 140.925 ;
        RECT -40.285 139.235 -39.955 139.565 ;
        RECT -40.285 137.875 -39.955 138.205 ;
        RECT -40.285 136.515 -39.955 136.845 ;
        RECT -40.285 135.155 -39.955 135.485 ;
        RECT -40.285 133.795 -39.955 134.125 ;
        RECT -40.285 132.435 -39.955 132.765 ;
        RECT -40.285 131.075 -39.955 131.405 ;
        RECT -40.285 129.715 -39.955 130.045 ;
        RECT -40.285 128.355 -39.955 128.685 ;
        RECT -40.285 126.995 -39.955 127.325 ;
        RECT -40.285 125.635 -39.955 125.965 ;
        RECT -40.285 124.275 -39.955 124.605 ;
        RECT -40.285 122.915 -39.955 123.245 ;
        RECT -40.285 121.555 -39.955 121.885 ;
        RECT -40.285 120.195 -39.955 120.525 ;
        RECT -40.285 118.835 -39.955 119.165 ;
        RECT -40.285 117.475 -39.955 117.805 ;
        RECT -40.285 116.115 -39.955 116.445 ;
        RECT -40.285 114.755 -39.955 115.085 ;
        RECT -40.285 113.395 -39.955 113.725 ;
        RECT -40.285 112.035 -39.955 112.365 ;
        RECT -40.285 110.675 -39.955 111.005 ;
        RECT -40.285 109.315 -39.955 109.645 ;
        RECT -40.285 107.955 -39.955 108.285 ;
        RECT -40.285 106.595 -39.955 106.925 ;
        RECT -40.285 105.235 -39.955 105.565 ;
        RECT -40.285 103.875 -39.955 104.205 ;
        RECT -40.285 102.515 -39.955 102.845 ;
        RECT -40.285 101.155 -39.955 101.485 ;
        RECT -40.285 99.795 -39.955 100.125 ;
        RECT -40.285 98.435 -39.955 98.765 ;
        RECT -40.285 97.075 -39.955 97.405 ;
        RECT -40.285 95.715 -39.955 96.045 ;
        RECT -40.285 94.355 -39.955 94.685 ;
        RECT -40.285 92.995 -39.955 93.325 ;
        RECT -40.285 91.635 -39.955 91.965 ;
        RECT -40.285 90.275 -39.955 90.605 ;
        RECT -40.285 88.915 -39.955 89.245 ;
        RECT -40.285 87.555 -39.955 87.885 ;
        RECT -40.285 86.195 -39.955 86.525 ;
        RECT -40.285 84.835 -39.955 85.165 ;
        RECT -40.285 83.475 -39.955 83.805 ;
        RECT -40.285 82.115 -39.955 82.445 ;
        RECT -40.285 80.755 -39.955 81.085 ;
        RECT -40.285 79.395 -39.955 79.725 ;
        RECT -40.285 78.035 -39.955 78.365 ;
        RECT -40.285 76.675 -39.955 77.005 ;
        RECT -40.285 75.315 -39.955 75.645 ;
        RECT -40.285 73.955 -39.955 74.285 ;
        RECT -40.285 72.595 -39.955 72.925 ;
        RECT -40.285 71.235 -39.955 71.565 ;
        RECT -40.285 69.875 -39.955 70.205 ;
        RECT -40.285 68.515 -39.955 68.845 ;
        RECT -40.285 67.155 -39.955 67.485 ;
        RECT -40.285 65.795 -39.955 66.125 ;
        RECT -40.285 64.435 -39.955 64.765 ;
        RECT -40.285 63.075 -39.955 63.405 ;
        RECT -40.285 61.715 -39.955 62.045 ;
        RECT -40.285 60.355 -39.955 60.685 ;
        RECT -40.285 58.995 -39.955 59.325 ;
        RECT -40.285 57.635 -39.955 57.965 ;
        RECT -40.285 56.275 -39.955 56.605 ;
        RECT -40.285 54.915 -39.955 55.245 ;
        RECT -40.285 53.555 -39.955 53.885 ;
        RECT -40.285 52.195 -39.955 52.525 ;
        RECT -40.285 50.835 -39.955 51.165 ;
        RECT -40.285 49.475 -39.955 49.805 ;
        RECT -40.285 48.115 -39.955 48.445 ;
        RECT -40.285 46.755 -39.955 47.085 ;
        RECT -40.285 45.395 -39.955 45.725 ;
        RECT -40.285 44.035 -39.955 44.365 ;
        RECT -40.285 42.675 -39.955 43.005 ;
        RECT -40.285 41.315 -39.955 41.645 ;
        RECT -40.285 39.955 -39.955 40.285 ;
        RECT -40.285 38.595 -39.955 38.925 ;
        RECT -40.285 37.235 -39.955 37.565 ;
        RECT -40.285 35.875 -39.955 36.205 ;
        RECT -40.285 34.515 -39.955 34.845 ;
        RECT -40.285 33.155 -39.955 33.485 ;
        RECT -40.285 31.795 -39.955 32.125 ;
        RECT -40.285 30.435 -39.955 30.765 ;
        RECT -40.285 29.075 -39.955 29.405 ;
        RECT -40.285 27.715 -39.955 28.045 ;
        RECT -40.285 26.355 -39.955 26.685 ;
        RECT -40.285 24.995 -39.955 25.325 ;
        RECT -40.285 23.635 -39.955 23.965 ;
        RECT -40.285 22.275 -39.955 22.605 ;
        RECT -40.285 20.915 -39.955 21.245 ;
        RECT -40.285 19.555 -39.955 19.885 ;
        RECT -40.285 18.195 -39.955 18.525 ;
        RECT -40.285 16.835 -39.955 17.165 ;
        RECT -40.285 15.475 -39.955 15.805 ;
        RECT -40.285 14.115 -39.955 14.445 ;
        RECT -40.285 12.755 -39.955 13.085 ;
        RECT -40.285 11.395 -39.955 11.725 ;
        RECT -40.285 10.035 -39.955 10.365 ;
        RECT -40.285 8.675 -39.955 9.005 ;
        RECT -40.285 7.315 -39.955 7.645 ;
        RECT -40.285 5.955 -39.955 6.285 ;
        RECT -40.285 4.595 -39.955 4.925 ;
        RECT -40.285 3.235 -39.955 3.565 ;
        RECT -40.285 1.875 -39.955 2.205 ;
        RECT -40.285 0.515 -39.955 0.845 ;
        RECT -40.285 -0.845 -39.955 -0.515 ;
        RECT -40.285 -7.645 -39.955 -7.315 ;
        RECT -40.285 -9.005 -39.955 -8.675 ;
        RECT -40.285 -10.365 -39.955 -10.035 ;
        RECT -40.285 -11.725 -39.955 -11.395 ;
        RECT -40.285 -13.085 -39.955 -12.755 ;
        RECT -40.285 -14.445 -39.955 -14.115 ;
        RECT -40.285 -15.805 -39.955 -15.475 ;
        RECT -40.285 -17.165 -39.955 -16.835 ;
        RECT -40.285 -18.525 -39.955 -18.195 ;
        RECT -40.285 -19.885 -39.955 -19.555 ;
        RECT -40.285 -21.245 -39.955 -20.915 ;
        RECT -40.285 -22.605 -39.955 -22.275 ;
        RECT -40.285 -29.405 -39.955 -29.075 ;
        RECT -40.285 -32.125 -39.955 -31.795 ;
        RECT -40.285 -33.485 -39.955 -33.155 ;
        RECT -40.285 -34.88 -39.955 -34.55 ;
        RECT -40.285 -36.205 -39.955 -35.875 ;
        RECT -40.285 -38.925 -39.955 -38.595 ;
        RECT -40.285 -39.97 -39.955 -39.64 ;
        RECT -40.285 -48.445 -39.955 -48.115 ;
        RECT -40.285 -49.805 -39.955 -49.475 ;
        RECT -40.285 -51.165 -39.955 -50.835 ;
        RECT -40.285 -53.885 -39.955 -53.555 ;
        RECT -40.285 -57.965 -39.955 -57.635 ;
        RECT -40.285 -62.045 -39.955 -61.715 ;
        RECT -40.285 -63.405 -39.955 -63.075 ;
        RECT -40.285 -64.765 -39.955 -64.435 ;
        RECT -40.285 -66.125 -39.955 -65.795 ;
        RECT -40.285 -67.485 -39.955 -67.155 ;
        RECT -40.285 -68.845 -39.955 -68.515 ;
        RECT -40.285 -70.205 -39.955 -69.875 ;
        RECT -40.285 -71.565 -39.955 -71.235 ;
        RECT -40.285 -72.925 -39.955 -72.595 ;
        RECT -40.285 -74.285 -39.955 -73.955 ;
        RECT -40.285 -75.645 -39.955 -75.315 ;
        RECT -40.285 -77.005 -39.955 -76.675 ;
        RECT -40.285 -78.365 -39.955 -78.035 ;
        RECT -40.285 -79.725 -39.955 -79.395 ;
        RECT -40.285 -81.085 -39.955 -80.755 ;
        RECT -40.285 -82.445 -39.955 -82.115 ;
        RECT -40.285 -83.805 -39.955 -83.475 ;
        RECT -40.285 -85.165 -39.955 -84.835 ;
        RECT -40.285 -86.525 -39.955 -86.195 ;
        RECT -40.285 -87.885 -39.955 -87.555 ;
        RECT -40.285 -89.245 -39.955 -88.915 ;
        RECT -40.285 -90.605 -39.955 -90.275 ;
        RECT -40.285 -91.965 -39.955 -91.635 ;
        RECT -40.285 -93.325 -39.955 -92.995 ;
        RECT -40.285 -94.685 -39.955 -94.355 ;
        RECT -40.285 -96.045 -39.955 -95.715 ;
        RECT -40.285 -97.405 -39.955 -97.075 ;
        RECT -40.285 -98.765 -39.955 -98.435 ;
        RECT -40.285 -100.125 -39.955 -99.795 ;
        RECT -40.285 -101.485 -39.955 -101.155 ;
        RECT -40.285 -102.845 -39.955 -102.515 ;
        RECT -40.285 -104.205 -39.955 -103.875 ;
        RECT -40.285 -105.565 -39.955 -105.235 ;
        RECT -40.285 -106.925 -39.955 -106.595 ;
        RECT -40.285 -108.285 -39.955 -107.955 ;
        RECT -40.285 -109.645 -39.955 -109.315 ;
        RECT -40.285 -111.005 -39.955 -110.675 ;
        RECT -40.285 -112.365 -39.955 -112.035 ;
        RECT -40.285 -113.725 -39.955 -113.395 ;
        RECT -40.285 -115.085 -39.955 -114.755 ;
        RECT -40.285 -116.445 -39.955 -116.115 ;
        RECT -40.285 -117.805 -39.955 -117.475 ;
        RECT -40.285 -119.165 -39.955 -118.835 ;
        RECT -40.285 -120.525 -39.955 -120.195 ;
        RECT -40.285 -124.605 -39.955 -124.275 ;
        RECT -40.285 -128.685 -39.955 -128.355 ;
        RECT -40.285 -130.045 -39.955 -129.715 ;
        RECT -40.285 -132.765 -39.955 -132.435 ;
        RECT -40.285 -134.125 -39.955 -133.795 ;
        RECT -40.285 -135.485 -39.955 -135.155 ;
        RECT -40.285 -136.845 -39.955 -136.515 ;
        RECT -40.285 -138.205 -39.955 -137.875 ;
        RECT -40.285 -139.39 -39.955 -139.06 ;
        RECT -40.285 -140.925 -39.955 -140.595 ;
        RECT -40.285 -142.285 -39.955 -141.955 ;
        RECT -40.285 -145.005 -39.955 -144.675 ;
        RECT -40.285 -146.365 -39.955 -146.035 ;
        RECT -40.285 -148.03 -39.955 -147.7 ;
        RECT -40.285 -149.085 -39.955 -148.755 ;
        RECT -40.285 -150.445 -39.955 -150.115 ;
        RECT -40.285 -153.165 -39.955 -152.835 ;
        RECT -40.285 -154.525 -39.955 -154.195 ;
        RECT -40.285 -155.885 -39.955 -155.555 ;
        RECT -40.285 -157.245 -39.955 -156.915 ;
        RECT -40.285 -159.965 -39.955 -159.635 ;
        RECT -40.285 -162.685 -39.955 -162.355 ;
        RECT -40.285 -164.045 -39.955 -163.715 ;
        RECT -40.285 -165.405 -39.955 -165.075 ;
        RECT -40.285 -166.765 -39.955 -166.435 ;
        RECT -40.285 -168.125 -39.955 -167.795 ;
        RECT -40.285 -169.485 -39.955 -169.155 ;
        RECT -40.285 -170.845 -39.955 -170.515 ;
        RECT -40.285 -172.205 -39.955 -171.875 ;
        RECT -40.285 -173.565 -39.955 -173.235 ;
        RECT -40.285 -174.925 -39.955 -174.595 ;
        RECT -40.285 -176.285 -39.955 -175.955 ;
        RECT -40.285 -177.645 -39.955 -177.315 ;
        RECT -40.285 -179.005 -39.955 -178.675 ;
        RECT -40.285 -180.365 -39.955 -180.035 ;
        RECT -40.285 -181.725 -39.955 -181.395 ;
        RECT -40.285 -183.085 -39.955 -182.755 ;
        RECT -40.285 -184.445 -39.955 -184.115 ;
        RECT -40.285 -185.805 -39.955 -185.475 ;
        RECT -40.285 -187.165 -39.955 -186.835 ;
        RECT -40.285 -188.525 -39.955 -188.195 ;
        RECT -40.285 -189.885 -39.955 -189.555 ;
        RECT -40.285 -191.245 -39.955 -190.915 ;
        RECT -40.285 -192.605 -39.955 -192.275 ;
        RECT -40.285 -193.965 -39.955 -193.635 ;
        RECT -40.285 -195.325 -39.955 -194.995 ;
        RECT -40.285 -196.685 -39.955 -196.355 ;
        RECT -40.285 -198.045 -39.955 -197.715 ;
        RECT -40.285 -199.405 -39.955 -199.075 ;
        RECT -40.285 -200.765 -39.955 -200.435 ;
        RECT -40.285 -202.125 -39.955 -201.795 ;
        RECT -40.285 -203.485 -39.955 -203.155 ;
        RECT -40.285 -204.845 -39.955 -204.515 ;
        RECT -40.285 -206.205 -39.955 -205.875 ;
        RECT -40.285 -207.565 -39.955 -207.235 ;
        RECT -40.285 -208.925 -39.955 -208.595 ;
        RECT -40.285 -210.285 -39.955 -209.955 ;
        RECT -40.285 -211.645 -39.955 -211.315 ;
        RECT -40.285 -213.005 -39.955 -212.675 ;
        RECT -40.285 -214.365 -39.955 -214.035 ;
        RECT -40.285 -215.725 -39.955 -215.395 ;
        RECT -40.285 -217.085 -39.955 -216.755 ;
        RECT -40.285 -218.445 -39.955 -218.115 ;
        RECT -40.285 -219.805 -39.955 -219.475 ;
        RECT -40.285 -221.165 -39.955 -220.835 ;
        RECT -40.285 -222.525 -39.955 -222.195 ;
        RECT -40.285 -223.885 -39.955 -223.555 ;
        RECT -40.285 -225.245 -39.955 -224.915 ;
        RECT -40.285 -227.965 -39.955 -227.635 ;
        RECT -40.28 -229.32 -39.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 244.04 -38.595 245.17 ;
        RECT -38.925 242.595 -38.595 242.925 ;
        RECT -38.925 241.235 -38.595 241.565 ;
        RECT -38.925 239.875 -38.595 240.205 ;
        RECT -38.925 238.515 -38.595 238.845 ;
        RECT -38.925 237.155 -38.595 237.485 ;
        RECT -38.925 235.795 -38.595 236.125 ;
        RECT -38.925 234.435 -38.595 234.765 ;
        RECT -38.925 233.075 -38.595 233.405 ;
        RECT -38.925 231.715 -38.595 232.045 ;
        RECT -38.925 230.355 -38.595 230.685 ;
        RECT -38.925 228.995 -38.595 229.325 ;
        RECT -38.925 227.635 -38.595 227.965 ;
        RECT -38.925 226.275 -38.595 226.605 ;
        RECT -38.925 224.915 -38.595 225.245 ;
        RECT -38.925 223.555 -38.595 223.885 ;
        RECT -38.925 222.195 -38.595 222.525 ;
        RECT -38.925 220.835 -38.595 221.165 ;
        RECT -38.925 219.475 -38.595 219.805 ;
        RECT -38.925 218.115 -38.595 218.445 ;
        RECT -38.925 216.755 -38.595 217.085 ;
        RECT -38.925 215.395 -38.595 215.725 ;
        RECT -38.925 214.035 -38.595 214.365 ;
        RECT -38.925 212.675 -38.595 213.005 ;
        RECT -38.925 211.315 -38.595 211.645 ;
        RECT -38.925 209.955 -38.595 210.285 ;
        RECT -38.925 208.595 -38.595 208.925 ;
        RECT -38.925 207.235 -38.595 207.565 ;
        RECT -38.925 205.875 -38.595 206.205 ;
        RECT -38.925 204.515 -38.595 204.845 ;
        RECT -38.925 203.155 -38.595 203.485 ;
        RECT -38.925 201.795 -38.595 202.125 ;
        RECT -38.925 200.435 -38.595 200.765 ;
        RECT -38.925 199.075 -38.595 199.405 ;
        RECT -38.925 197.715 -38.595 198.045 ;
        RECT -38.925 196.355 -38.595 196.685 ;
        RECT -38.925 194.995 -38.595 195.325 ;
        RECT -38.925 193.635 -38.595 193.965 ;
        RECT -38.925 192.275 -38.595 192.605 ;
        RECT -38.925 190.915 -38.595 191.245 ;
        RECT -38.925 189.555 -38.595 189.885 ;
        RECT -38.925 188.195 -38.595 188.525 ;
        RECT -38.925 186.835 -38.595 187.165 ;
        RECT -38.925 185.475 -38.595 185.805 ;
        RECT -38.925 184.115 -38.595 184.445 ;
        RECT -38.925 182.755 -38.595 183.085 ;
        RECT -38.925 181.395 -38.595 181.725 ;
        RECT -38.925 180.035 -38.595 180.365 ;
        RECT -38.925 178.675 -38.595 179.005 ;
        RECT -38.925 177.315 -38.595 177.645 ;
        RECT -38.925 175.955 -38.595 176.285 ;
        RECT -38.925 174.595 -38.595 174.925 ;
        RECT -38.925 173.235 -38.595 173.565 ;
        RECT -38.925 171.875 -38.595 172.205 ;
        RECT -38.925 170.515 -38.595 170.845 ;
        RECT -38.925 169.155 -38.595 169.485 ;
        RECT -38.925 167.795 -38.595 168.125 ;
        RECT -38.925 166.435 -38.595 166.765 ;
        RECT -38.925 165.075 -38.595 165.405 ;
        RECT -38.925 163.715 -38.595 164.045 ;
        RECT -38.925 162.355 -38.595 162.685 ;
        RECT -38.925 160.995 -38.595 161.325 ;
        RECT -38.925 159.635 -38.595 159.965 ;
        RECT -38.925 158.275 -38.595 158.605 ;
        RECT -38.925 156.915 -38.595 157.245 ;
        RECT -38.925 155.555 -38.595 155.885 ;
        RECT -38.925 154.195 -38.595 154.525 ;
        RECT -38.925 152.835 -38.595 153.165 ;
        RECT -38.925 151.475 -38.595 151.805 ;
        RECT -38.925 150.115 -38.595 150.445 ;
        RECT -38.925 148.755 -38.595 149.085 ;
        RECT -38.925 147.395 -38.595 147.725 ;
        RECT -38.925 146.035 -38.595 146.365 ;
        RECT -38.925 144.675 -38.595 145.005 ;
        RECT -38.925 143.315 -38.595 143.645 ;
        RECT -38.925 141.955 -38.595 142.285 ;
        RECT -38.925 140.595 -38.595 140.925 ;
        RECT -38.925 139.235 -38.595 139.565 ;
        RECT -38.925 137.875 -38.595 138.205 ;
        RECT -38.925 136.515 -38.595 136.845 ;
        RECT -38.925 135.155 -38.595 135.485 ;
        RECT -38.925 133.795 -38.595 134.125 ;
        RECT -38.925 132.435 -38.595 132.765 ;
        RECT -38.925 131.075 -38.595 131.405 ;
        RECT -38.925 129.715 -38.595 130.045 ;
        RECT -38.925 128.355 -38.595 128.685 ;
        RECT -38.925 126.995 -38.595 127.325 ;
        RECT -38.925 125.635 -38.595 125.965 ;
        RECT -38.925 124.275 -38.595 124.605 ;
        RECT -38.925 122.915 -38.595 123.245 ;
        RECT -38.925 121.555 -38.595 121.885 ;
        RECT -38.925 120.195 -38.595 120.525 ;
        RECT -38.925 118.835 -38.595 119.165 ;
        RECT -38.925 117.475 -38.595 117.805 ;
        RECT -38.925 116.115 -38.595 116.445 ;
        RECT -38.925 114.755 -38.595 115.085 ;
        RECT -38.925 113.395 -38.595 113.725 ;
        RECT -38.925 112.035 -38.595 112.365 ;
        RECT -38.925 110.675 -38.595 111.005 ;
        RECT -38.925 109.315 -38.595 109.645 ;
        RECT -38.925 107.955 -38.595 108.285 ;
        RECT -38.925 106.595 -38.595 106.925 ;
        RECT -38.925 105.235 -38.595 105.565 ;
        RECT -38.925 103.875 -38.595 104.205 ;
        RECT -38.925 102.515 -38.595 102.845 ;
        RECT -38.925 101.155 -38.595 101.485 ;
        RECT -38.925 99.795 -38.595 100.125 ;
        RECT -38.925 98.435 -38.595 98.765 ;
        RECT -38.925 97.075 -38.595 97.405 ;
        RECT -38.925 95.715 -38.595 96.045 ;
        RECT -38.925 94.355 -38.595 94.685 ;
        RECT -38.925 92.995 -38.595 93.325 ;
        RECT -38.925 91.635 -38.595 91.965 ;
        RECT -38.925 90.275 -38.595 90.605 ;
        RECT -38.925 88.915 -38.595 89.245 ;
        RECT -38.925 87.555 -38.595 87.885 ;
        RECT -38.925 86.195 -38.595 86.525 ;
        RECT -38.925 84.835 -38.595 85.165 ;
        RECT -38.925 83.475 -38.595 83.805 ;
        RECT -38.925 82.115 -38.595 82.445 ;
        RECT -38.925 80.755 -38.595 81.085 ;
        RECT -38.925 79.395 -38.595 79.725 ;
        RECT -38.925 78.035 -38.595 78.365 ;
        RECT -38.925 76.675 -38.595 77.005 ;
        RECT -38.925 75.315 -38.595 75.645 ;
        RECT -38.925 73.955 -38.595 74.285 ;
        RECT -38.925 72.595 -38.595 72.925 ;
        RECT -38.925 71.235 -38.595 71.565 ;
        RECT -38.925 69.875 -38.595 70.205 ;
        RECT -38.925 68.515 -38.595 68.845 ;
        RECT -38.925 67.155 -38.595 67.485 ;
        RECT -38.925 65.795 -38.595 66.125 ;
        RECT -38.925 64.435 -38.595 64.765 ;
        RECT -38.925 63.075 -38.595 63.405 ;
        RECT -38.925 61.715 -38.595 62.045 ;
        RECT -38.925 60.355 -38.595 60.685 ;
        RECT -38.925 58.995 -38.595 59.325 ;
        RECT -38.925 57.635 -38.595 57.965 ;
        RECT -38.925 56.275 -38.595 56.605 ;
        RECT -38.925 54.915 -38.595 55.245 ;
        RECT -38.925 53.555 -38.595 53.885 ;
        RECT -38.925 52.195 -38.595 52.525 ;
        RECT -38.925 50.835 -38.595 51.165 ;
        RECT -38.925 49.475 -38.595 49.805 ;
        RECT -38.925 48.115 -38.595 48.445 ;
        RECT -38.925 46.755 -38.595 47.085 ;
        RECT -38.925 45.395 -38.595 45.725 ;
        RECT -38.925 44.035 -38.595 44.365 ;
        RECT -38.925 42.675 -38.595 43.005 ;
        RECT -38.925 41.315 -38.595 41.645 ;
        RECT -38.925 39.955 -38.595 40.285 ;
        RECT -38.925 38.595 -38.595 38.925 ;
        RECT -38.925 37.235 -38.595 37.565 ;
        RECT -38.925 35.875 -38.595 36.205 ;
        RECT -38.925 34.515 -38.595 34.845 ;
        RECT -38.925 33.155 -38.595 33.485 ;
        RECT -38.925 31.795 -38.595 32.125 ;
        RECT -38.925 30.435 -38.595 30.765 ;
        RECT -38.925 29.075 -38.595 29.405 ;
        RECT -38.925 27.715 -38.595 28.045 ;
        RECT -38.925 26.355 -38.595 26.685 ;
        RECT -38.925 24.995 -38.595 25.325 ;
        RECT -38.925 23.635 -38.595 23.965 ;
        RECT -38.925 22.275 -38.595 22.605 ;
        RECT -38.925 20.915 -38.595 21.245 ;
        RECT -38.925 19.555 -38.595 19.885 ;
        RECT -38.925 18.195 -38.595 18.525 ;
        RECT -38.925 16.835 -38.595 17.165 ;
        RECT -38.925 15.475 -38.595 15.805 ;
        RECT -38.925 14.115 -38.595 14.445 ;
        RECT -38.925 12.755 -38.595 13.085 ;
        RECT -38.925 11.395 -38.595 11.725 ;
        RECT -38.925 10.035 -38.595 10.365 ;
        RECT -38.925 8.675 -38.595 9.005 ;
        RECT -38.925 7.315 -38.595 7.645 ;
        RECT -38.925 5.955 -38.595 6.285 ;
        RECT -38.925 4.595 -38.595 4.925 ;
        RECT -38.925 3.235 -38.595 3.565 ;
        RECT -38.925 1.875 -38.595 2.205 ;
        RECT -38.925 0.515 -38.595 0.845 ;
        RECT -38.925 -0.845 -38.595 -0.515 ;
        RECT -38.925 -4.925 -38.595 -4.595 ;
        RECT -38.925 -7.645 -38.595 -7.315 ;
        RECT -38.925 -9.005 -38.595 -8.675 ;
        RECT -38.925 -10.365 -38.595 -10.035 ;
        RECT -38.925 -11.725 -38.595 -11.395 ;
        RECT -38.925 -13.085 -38.595 -12.755 ;
        RECT -38.925 -14.445 -38.595 -14.115 ;
        RECT -38.925 -15.805 -38.595 -15.475 ;
        RECT -38.925 -17.165 -38.595 -16.835 ;
        RECT -38.925 -18.525 -38.595 -18.195 ;
        RECT -38.925 -19.885 -38.595 -19.555 ;
        RECT -38.925 -21.245 -38.595 -20.915 ;
        RECT -38.925 -22.605 -38.595 -22.275 ;
        RECT -38.925 -29.405 -38.595 -29.075 ;
        RECT -38.925 -32.125 -38.595 -31.795 ;
        RECT -38.925 -33.485 -38.595 -33.155 ;
        RECT -38.925 -34.88 -38.595 -34.55 ;
        RECT -38.925 -36.205 -38.595 -35.875 ;
        RECT -38.925 -38.925 -38.595 -38.595 ;
        RECT -38.925 -39.97 -38.595 -39.64 ;
        RECT -38.925 -48.445 -38.595 -48.115 ;
        RECT -38.925 -49.805 -38.595 -49.475 ;
        RECT -38.925 -51.165 -38.595 -50.835 ;
        RECT -38.925 -53.885 -38.595 -53.555 ;
        RECT -38.925 -57.965 -38.595 -57.635 ;
        RECT -38.925 -62.045 -38.595 -61.715 ;
        RECT -38.925 -63.405 -38.595 -63.075 ;
        RECT -38.925 -64.765 -38.595 -64.435 ;
        RECT -38.925 -66.125 -38.595 -65.795 ;
        RECT -38.925 -67.485 -38.595 -67.155 ;
        RECT -38.925 -68.845 -38.595 -68.515 ;
        RECT -38.925 -70.205 -38.595 -69.875 ;
        RECT -38.925 -71.565 -38.595 -71.235 ;
        RECT -38.925 -72.925 -38.595 -72.595 ;
        RECT -38.925 -74.285 -38.595 -73.955 ;
        RECT -38.925 -75.645 -38.595 -75.315 ;
        RECT -38.925 -77.005 -38.595 -76.675 ;
        RECT -38.925 -78.365 -38.595 -78.035 ;
        RECT -38.925 -79.725 -38.595 -79.395 ;
        RECT -38.925 -81.085 -38.595 -80.755 ;
        RECT -38.925 -82.445 -38.595 -82.115 ;
        RECT -38.925 -83.805 -38.595 -83.475 ;
        RECT -38.925 -85.165 -38.595 -84.835 ;
        RECT -38.925 -86.525 -38.595 -86.195 ;
        RECT -38.925 -87.885 -38.595 -87.555 ;
        RECT -38.925 -89.245 -38.595 -88.915 ;
        RECT -38.925 -90.605 -38.595 -90.275 ;
        RECT -38.925 -91.965 -38.595 -91.635 ;
        RECT -38.925 -93.325 -38.595 -92.995 ;
        RECT -38.925 -94.685 -38.595 -94.355 ;
        RECT -38.925 -96.045 -38.595 -95.715 ;
        RECT -38.925 -97.405 -38.595 -97.075 ;
        RECT -38.925 -98.765 -38.595 -98.435 ;
        RECT -38.925 -100.125 -38.595 -99.795 ;
        RECT -38.925 -101.485 -38.595 -101.155 ;
        RECT -38.925 -102.845 -38.595 -102.515 ;
        RECT -38.925 -104.205 -38.595 -103.875 ;
        RECT -38.925 -105.565 -38.595 -105.235 ;
        RECT -38.925 -106.925 -38.595 -106.595 ;
        RECT -38.925 -108.285 -38.595 -107.955 ;
        RECT -38.925 -109.645 -38.595 -109.315 ;
        RECT -38.925 -111.005 -38.595 -110.675 ;
        RECT -38.925 -112.365 -38.595 -112.035 ;
        RECT -38.925 -113.725 -38.595 -113.395 ;
        RECT -38.925 -115.085 -38.595 -114.755 ;
        RECT -38.925 -116.445 -38.595 -116.115 ;
        RECT -38.925 -117.805 -38.595 -117.475 ;
        RECT -38.925 -119.165 -38.595 -118.835 ;
        RECT -38.925 -124.605 -38.595 -124.275 ;
        RECT -38.925 -128.685 -38.595 -128.355 ;
        RECT -38.925 -130.045 -38.595 -129.715 ;
        RECT -38.925 -132.765 -38.595 -132.435 ;
        RECT -38.925 -134.125 -38.595 -133.795 ;
        RECT -38.925 -135.485 -38.595 -135.155 ;
        RECT -38.925 -136.845 -38.595 -136.515 ;
        RECT -38.925 -138.205 -38.595 -137.875 ;
        RECT -38.925 -139.39 -38.595 -139.06 ;
        RECT -38.925 -140.925 -38.595 -140.595 ;
        RECT -38.925 -142.285 -38.595 -141.955 ;
        RECT -38.925 -145.005 -38.595 -144.675 ;
        RECT -38.925 -146.365 -38.595 -146.035 ;
        RECT -38.925 -148.03 -38.595 -147.7 ;
        RECT -38.925 -149.085 -38.595 -148.755 ;
        RECT -38.925 -150.445 -38.595 -150.115 ;
        RECT -38.92 -152.48 -38.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 -232.045 -38.595 -231.715 ;
        RECT -38.925 -233.225 -38.595 -232.895 ;
        RECT -38.925 -234.765 -38.595 -234.435 ;
        RECT -38.925 -236.125 -38.595 -235.795 ;
        RECT -38.925 -237.485 -38.595 -237.155 ;
        RECT -38.925 -238.845 -38.595 -238.515 ;
        RECT -38.925 -241.09 -38.595 -239.96 ;
        RECT -38.92 -241.205 -38.6 -231.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.565 -168.125 -37.235 -167.795 ;
        RECT -37.565 -169.485 -37.235 -169.155 ;
        RECT -37.565 -170.845 -37.235 -170.515 ;
        RECT -37.565 -172.205 -37.235 -171.875 ;
        RECT -37.565 -173.565 -37.235 -173.235 ;
        RECT -37.565 -174.925 -37.235 -174.595 ;
        RECT -37.565 -176.285 -37.235 -175.955 ;
        RECT -37.565 -177.645 -37.235 -177.315 ;
        RECT -37.565 -179.005 -37.235 -178.675 ;
        RECT -37.565 -180.365 -37.235 -180.035 ;
        RECT -37.565 -181.725 -37.235 -181.395 ;
        RECT -37.565 -183.085 -37.235 -182.755 ;
        RECT -37.565 -184.445 -37.235 -184.115 ;
        RECT -37.565 -185.805 -37.235 -185.475 ;
        RECT -37.565 -187.165 -37.235 -186.835 ;
        RECT -37.565 -188.525 -37.235 -188.195 ;
        RECT -37.565 -189.885 -37.235 -189.555 ;
        RECT -37.565 -191.245 -37.235 -190.915 ;
        RECT -37.565 -192.605 -37.235 -192.275 ;
        RECT -37.565 -193.965 -37.235 -193.635 ;
        RECT -37.565 -195.325 -37.235 -194.995 ;
        RECT -37.565 -196.685 -37.235 -196.355 ;
        RECT -37.565 -198.045 -37.235 -197.715 ;
        RECT -37.565 -199.405 -37.235 -199.075 ;
        RECT -37.565 -200.765 -37.235 -200.435 ;
        RECT -37.565 -202.125 -37.235 -201.795 ;
        RECT -37.565 -203.485 -37.235 -203.155 ;
        RECT -37.565 -204.845 -37.235 -204.515 ;
        RECT -37.565 -206.205 -37.235 -205.875 ;
        RECT -37.565 -207.565 -37.235 -207.235 ;
        RECT -37.565 -208.925 -37.235 -208.595 ;
        RECT -37.565 -210.285 -37.235 -209.955 ;
        RECT -37.565 -211.645 -37.235 -211.315 ;
        RECT -37.565 -213.005 -37.235 -212.675 ;
        RECT -37.565 -214.365 -37.235 -214.035 ;
        RECT -37.565 -215.725 -37.235 -215.395 ;
        RECT -37.565 -217.085 -37.235 -216.755 ;
        RECT -37.565 -218.445 -37.235 -218.115 ;
        RECT -37.565 -219.805 -37.235 -219.475 ;
        RECT -37.565 -221.165 -37.235 -220.835 ;
        RECT -37.565 -222.525 -37.235 -222.195 ;
        RECT -37.565 -223.885 -37.235 -223.555 ;
        RECT -37.565 -225.245 -37.235 -224.915 ;
        RECT -37.565 -227.965 -37.235 -227.635 ;
        RECT -37.565 -230.685 -37.235 -230.355 ;
        RECT -37.565 -232.045 -37.235 -231.715 ;
        RECT -37.565 -233.225 -37.235 -232.895 ;
        RECT -37.565 -234.765 -37.235 -234.435 ;
        RECT -37.565 -236.125 -37.235 -235.795 ;
        RECT -37.565 -237.485 -37.235 -237.155 ;
        RECT -37.565 -238.845 -37.235 -238.515 ;
        RECT -37.565 -241.09 -37.235 -239.96 ;
        RECT -37.56 -241.205 -37.24 245.285 ;
        RECT -37.565 244.04 -37.235 245.17 ;
        RECT -37.565 242.595 -37.235 242.925 ;
        RECT -37.565 241.235 -37.235 241.565 ;
        RECT -37.565 239.875 -37.235 240.205 ;
        RECT -37.565 238.515 -37.235 238.845 ;
        RECT -37.565 237.155 -37.235 237.485 ;
        RECT -37.565 235.795 -37.235 236.125 ;
        RECT -37.565 234.435 -37.235 234.765 ;
        RECT -37.565 233.075 -37.235 233.405 ;
        RECT -37.565 231.715 -37.235 232.045 ;
        RECT -37.565 230.355 -37.235 230.685 ;
        RECT -37.565 228.995 -37.235 229.325 ;
        RECT -37.565 227.635 -37.235 227.965 ;
        RECT -37.565 226.275 -37.235 226.605 ;
        RECT -37.565 224.915 -37.235 225.245 ;
        RECT -37.565 223.555 -37.235 223.885 ;
        RECT -37.565 222.195 -37.235 222.525 ;
        RECT -37.565 220.835 -37.235 221.165 ;
        RECT -37.565 219.475 -37.235 219.805 ;
        RECT -37.565 218.115 -37.235 218.445 ;
        RECT -37.565 216.755 -37.235 217.085 ;
        RECT -37.565 215.395 -37.235 215.725 ;
        RECT -37.565 214.035 -37.235 214.365 ;
        RECT -37.565 212.675 -37.235 213.005 ;
        RECT -37.565 211.315 -37.235 211.645 ;
        RECT -37.565 209.955 -37.235 210.285 ;
        RECT -37.565 208.595 -37.235 208.925 ;
        RECT -37.565 207.235 -37.235 207.565 ;
        RECT -37.565 205.875 -37.235 206.205 ;
        RECT -37.565 204.515 -37.235 204.845 ;
        RECT -37.565 203.155 -37.235 203.485 ;
        RECT -37.565 201.795 -37.235 202.125 ;
        RECT -37.565 200.435 -37.235 200.765 ;
        RECT -37.565 199.075 -37.235 199.405 ;
        RECT -37.565 197.715 -37.235 198.045 ;
        RECT -37.565 196.355 -37.235 196.685 ;
        RECT -37.565 194.995 -37.235 195.325 ;
        RECT -37.565 193.635 -37.235 193.965 ;
        RECT -37.565 192.275 -37.235 192.605 ;
        RECT -37.565 190.915 -37.235 191.245 ;
        RECT -37.565 189.555 -37.235 189.885 ;
        RECT -37.565 188.195 -37.235 188.525 ;
        RECT -37.565 186.835 -37.235 187.165 ;
        RECT -37.565 185.475 -37.235 185.805 ;
        RECT -37.565 184.115 -37.235 184.445 ;
        RECT -37.565 182.755 -37.235 183.085 ;
        RECT -37.565 181.395 -37.235 181.725 ;
        RECT -37.565 180.035 -37.235 180.365 ;
        RECT -37.565 178.675 -37.235 179.005 ;
        RECT -37.565 177.315 -37.235 177.645 ;
        RECT -37.565 175.955 -37.235 176.285 ;
        RECT -37.565 174.595 -37.235 174.925 ;
        RECT -37.565 173.235 -37.235 173.565 ;
        RECT -37.565 171.875 -37.235 172.205 ;
        RECT -37.565 170.515 -37.235 170.845 ;
        RECT -37.565 169.155 -37.235 169.485 ;
        RECT -37.565 167.795 -37.235 168.125 ;
        RECT -37.565 166.435 -37.235 166.765 ;
        RECT -37.565 165.075 -37.235 165.405 ;
        RECT -37.565 163.715 -37.235 164.045 ;
        RECT -37.565 162.355 -37.235 162.685 ;
        RECT -37.565 160.995 -37.235 161.325 ;
        RECT -37.565 159.635 -37.235 159.965 ;
        RECT -37.565 158.275 -37.235 158.605 ;
        RECT -37.565 156.915 -37.235 157.245 ;
        RECT -37.565 155.555 -37.235 155.885 ;
        RECT -37.565 154.195 -37.235 154.525 ;
        RECT -37.565 152.835 -37.235 153.165 ;
        RECT -37.565 151.475 -37.235 151.805 ;
        RECT -37.565 150.115 -37.235 150.445 ;
        RECT -37.565 148.755 -37.235 149.085 ;
        RECT -37.565 147.395 -37.235 147.725 ;
        RECT -37.565 146.035 -37.235 146.365 ;
        RECT -37.565 144.675 -37.235 145.005 ;
        RECT -37.565 143.315 -37.235 143.645 ;
        RECT -37.565 141.955 -37.235 142.285 ;
        RECT -37.565 140.595 -37.235 140.925 ;
        RECT -37.565 139.235 -37.235 139.565 ;
        RECT -37.565 137.875 -37.235 138.205 ;
        RECT -37.565 136.515 -37.235 136.845 ;
        RECT -37.565 135.155 -37.235 135.485 ;
        RECT -37.565 133.795 -37.235 134.125 ;
        RECT -37.565 132.435 -37.235 132.765 ;
        RECT -37.565 131.075 -37.235 131.405 ;
        RECT -37.565 129.715 -37.235 130.045 ;
        RECT -37.565 128.355 -37.235 128.685 ;
        RECT -37.565 126.995 -37.235 127.325 ;
        RECT -37.565 125.635 -37.235 125.965 ;
        RECT -37.565 124.275 -37.235 124.605 ;
        RECT -37.565 122.915 -37.235 123.245 ;
        RECT -37.565 121.555 -37.235 121.885 ;
        RECT -37.565 120.195 -37.235 120.525 ;
        RECT -37.565 118.835 -37.235 119.165 ;
        RECT -37.565 117.475 -37.235 117.805 ;
        RECT -37.565 116.115 -37.235 116.445 ;
        RECT -37.565 114.755 -37.235 115.085 ;
        RECT -37.565 113.395 -37.235 113.725 ;
        RECT -37.565 112.035 -37.235 112.365 ;
        RECT -37.565 110.675 -37.235 111.005 ;
        RECT -37.565 109.315 -37.235 109.645 ;
        RECT -37.565 107.955 -37.235 108.285 ;
        RECT -37.565 106.595 -37.235 106.925 ;
        RECT -37.565 105.235 -37.235 105.565 ;
        RECT -37.565 103.875 -37.235 104.205 ;
        RECT -37.565 102.515 -37.235 102.845 ;
        RECT -37.565 101.155 -37.235 101.485 ;
        RECT -37.565 99.795 -37.235 100.125 ;
        RECT -37.565 98.435 -37.235 98.765 ;
        RECT -37.565 97.075 -37.235 97.405 ;
        RECT -37.565 95.715 -37.235 96.045 ;
        RECT -37.565 94.355 -37.235 94.685 ;
        RECT -37.565 92.995 -37.235 93.325 ;
        RECT -37.565 91.635 -37.235 91.965 ;
        RECT -37.565 90.275 -37.235 90.605 ;
        RECT -37.565 88.915 -37.235 89.245 ;
        RECT -37.565 87.555 -37.235 87.885 ;
        RECT -37.565 86.195 -37.235 86.525 ;
        RECT -37.565 84.835 -37.235 85.165 ;
        RECT -37.565 83.475 -37.235 83.805 ;
        RECT -37.565 82.115 -37.235 82.445 ;
        RECT -37.565 80.755 -37.235 81.085 ;
        RECT -37.565 79.395 -37.235 79.725 ;
        RECT -37.565 78.035 -37.235 78.365 ;
        RECT -37.565 76.675 -37.235 77.005 ;
        RECT -37.565 75.315 -37.235 75.645 ;
        RECT -37.565 73.955 -37.235 74.285 ;
        RECT -37.565 72.595 -37.235 72.925 ;
        RECT -37.565 71.235 -37.235 71.565 ;
        RECT -37.565 69.875 -37.235 70.205 ;
        RECT -37.565 68.515 -37.235 68.845 ;
        RECT -37.565 67.155 -37.235 67.485 ;
        RECT -37.565 65.795 -37.235 66.125 ;
        RECT -37.565 64.435 -37.235 64.765 ;
        RECT -37.565 63.075 -37.235 63.405 ;
        RECT -37.565 61.715 -37.235 62.045 ;
        RECT -37.565 60.355 -37.235 60.685 ;
        RECT -37.565 58.995 -37.235 59.325 ;
        RECT -37.565 57.635 -37.235 57.965 ;
        RECT -37.565 56.275 -37.235 56.605 ;
        RECT -37.565 54.915 -37.235 55.245 ;
        RECT -37.565 53.555 -37.235 53.885 ;
        RECT -37.565 52.195 -37.235 52.525 ;
        RECT -37.565 50.835 -37.235 51.165 ;
        RECT -37.565 49.475 -37.235 49.805 ;
        RECT -37.565 48.115 -37.235 48.445 ;
        RECT -37.565 46.755 -37.235 47.085 ;
        RECT -37.565 45.395 -37.235 45.725 ;
        RECT -37.565 44.035 -37.235 44.365 ;
        RECT -37.565 42.675 -37.235 43.005 ;
        RECT -37.565 41.315 -37.235 41.645 ;
        RECT -37.565 39.955 -37.235 40.285 ;
        RECT -37.565 38.595 -37.235 38.925 ;
        RECT -37.565 37.235 -37.235 37.565 ;
        RECT -37.565 35.875 -37.235 36.205 ;
        RECT -37.565 34.515 -37.235 34.845 ;
        RECT -37.565 33.155 -37.235 33.485 ;
        RECT -37.565 31.795 -37.235 32.125 ;
        RECT -37.565 30.435 -37.235 30.765 ;
        RECT -37.565 29.075 -37.235 29.405 ;
        RECT -37.565 27.715 -37.235 28.045 ;
        RECT -37.565 26.355 -37.235 26.685 ;
        RECT -37.565 24.995 -37.235 25.325 ;
        RECT -37.565 23.635 -37.235 23.965 ;
        RECT -37.565 22.275 -37.235 22.605 ;
        RECT -37.565 20.915 -37.235 21.245 ;
        RECT -37.565 19.555 -37.235 19.885 ;
        RECT -37.565 18.195 -37.235 18.525 ;
        RECT -37.565 16.835 -37.235 17.165 ;
        RECT -37.565 15.475 -37.235 15.805 ;
        RECT -37.565 14.115 -37.235 14.445 ;
        RECT -37.565 12.755 -37.235 13.085 ;
        RECT -37.565 11.395 -37.235 11.725 ;
        RECT -37.565 10.035 -37.235 10.365 ;
        RECT -37.565 8.675 -37.235 9.005 ;
        RECT -37.565 7.315 -37.235 7.645 ;
        RECT -37.565 5.955 -37.235 6.285 ;
        RECT -37.565 4.595 -37.235 4.925 ;
        RECT -37.565 3.235 -37.235 3.565 ;
        RECT -37.565 1.875 -37.235 2.205 ;
        RECT -37.565 0.515 -37.235 0.845 ;
        RECT -37.565 -0.845 -37.235 -0.515 ;
        RECT -37.565 -3.565 -37.235 -3.235 ;
        RECT -37.565 -4.925 -37.235 -4.595 ;
        RECT -37.565 -7.645 -37.235 -7.315 ;
        RECT -37.565 -9.005 -37.235 -8.675 ;
        RECT -37.565 -10.365 -37.235 -10.035 ;
        RECT -37.565 -11.725 -37.235 -11.395 ;
        RECT -37.565 -13.085 -37.235 -12.755 ;
        RECT -37.565 -14.445 -37.235 -14.115 ;
        RECT -37.565 -15.805 -37.235 -15.475 ;
        RECT -37.565 -17.165 -37.235 -16.835 ;
        RECT -37.565 -18.525 -37.235 -18.195 ;
        RECT -37.565 -19.885 -37.235 -19.555 ;
        RECT -37.565 -21.245 -37.235 -20.915 ;
        RECT -37.565 -22.605 -37.235 -22.275 ;
        RECT -37.565 -29.405 -37.235 -29.075 ;
        RECT -37.565 -32.125 -37.235 -31.795 ;
        RECT -37.565 -33.485 -37.235 -33.155 ;
        RECT -37.565 -34.88 -37.235 -34.55 ;
        RECT -37.565 -36.205 -37.235 -35.875 ;
        RECT -37.565 -38.925 -37.235 -38.595 ;
        RECT -37.565 -39.97 -37.235 -39.64 ;
        RECT -37.565 -47.085 -37.235 -46.755 ;
        RECT -37.565 -48.445 -37.235 -48.115 ;
        RECT -37.565 -49.805 -37.235 -49.475 ;
        RECT -37.565 -51.165 -37.235 -50.835 ;
        RECT -37.565 -52.525 -37.235 -52.195 ;
        RECT -37.565 -53.885 -37.235 -53.555 ;
        RECT -37.565 -55.245 -37.235 -54.915 ;
        RECT -37.565 -56.605 -37.235 -56.275 ;
        RECT -37.565 -57.965 -37.235 -57.635 ;
        RECT -37.565 -59.325 -37.235 -58.995 ;
        RECT -37.565 -60.685 -37.235 -60.355 ;
        RECT -37.565 -62.045 -37.235 -61.715 ;
        RECT -37.565 -63.405 -37.235 -63.075 ;
        RECT -37.565 -64.765 -37.235 -64.435 ;
        RECT -37.565 -66.125 -37.235 -65.795 ;
        RECT -37.565 -67.485 -37.235 -67.155 ;
        RECT -37.565 -68.845 -37.235 -68.515 ;
        RECT -37.565 -70.205 -37.235 -69.875 ;
        RECT -37.565 -71.565 -37.235 -71.235 ;
        RECT -37.565 -72.925 -37.235 -72.595 ;
        RECT -37.565 -74.285 -37.235 -73.955 ;
        RECT -37.565 -75.645 -37.235 -75.315 ;
        RECT -37.565 -77.005 -37.235 -76.675 ;
        RECT -37.565 -78.365 -37.235 -78.035 ;
        RECT -37.565 -79.725 -37.235 -79.395 ;
        RECT -37.565 -81.085 -37.235 -80.755 ;
        RECT -37.565 -82.445 -37.235 -82.115 ;
        RECT -37.565 -83.805 -37.235 -83.475 ;
        RECT -37.565 -85.165 -37.235 -84.835 ;
        RECT -37.565 -86.525 -37.235 -86.195 ;
        RECT -37.565 -87.885 -37.235 -87.555 ;
        RECT -37.565 -89.245 -37.235 -88.915 ;
        RECT -37.565 -90.605 -37.235 -90.275 ;
        RECT -37.565 -91.965 -37.235 -91.635 ;
        RECT -37.565 -93.325 -37.235 -92.995 ;
        RECT -37.565 -94.685 -37.235 -94.355 ;
        RECT -37.565 -96.045 -37.235 -95.715 ;
        RECT -37.565 -97.405 -37.235 -97.075 ;
        RECT -37.565 -98.765 -37.235 -98.435 ;
        RECT -37.565 -100.125 -37.235 -99.795 ;
        RECT -37.565 -101.485 -37.235 -101.155 ;
        RECT -37.565 -102.845 -37.235 -102.515 ;
        RECT -37.565 -104.205 -37.235 -103.875 ;
        RECT -37.565 -105.565 -37.235 -105.235 ;
        RECT -37.565 -106.925 -37.235 -106.595 ;
        RECT -37.565 -108.285 -37.235 -107.955 ;
        RECT -37.565 -109.645 -37.235 -109.315 ;
        RECT -37.565 -111.005 -37.235 -110.675 ;
        RECT -37.565 -112.365 -37.235 -112.035 ;
        RECT -37.565 -113.725 -37.235 -113.395 ;
        RECT -37.565 -115.085 -37.235 -114.755 ;
        RECT -37.565 -116.445 -37.235 -116.115 ;
        RECT -37.565 -117.805 -37.235 -117.475 ;
        RECT -37.565 -119.165 -37.235 -118.835 ;
        RECT -37.565 -124.605 -37.235 -124.275 ;
        RECT -37.565 -128.685 -37.235 -128.355 ;
        RECT -37.565 -130.045 -37.235 -129.715 ;
        RECT -37.565 -132.765 -37.235 -132.435 ;
        RECT -37.565 -134.125 -37.235 -133.795 ;
        RECT -37.565 -135.485 -37.235 -135.155 ;
        RECT -37.565 -136.845 -37.235 -136.515 ;
        RECT -37.565 -138.205 -37.235 -137.875 ;
        RECT -37.565 -139.39 -37.235 -139.06 ;
        RECT -37.565 -140.925 -37.235 -140.595 ;
        RECT -37.565 -142.285 -37.235 -141.955 ;
        RECT -37.565 -145.005 -37.235 -144.675 ;
        RECT -37.565 -146.365 -37.235 -146.035 ;
        RECT -37.565 -148.03 -37.235 -147.7 ;
        RECT -37.565 -149.085 -37.235 -148.755 ;
        RECT -37.565 -150.445 -37.235 -150.115 ;
        RECT -37.565 -153.165 -37.235 -152.835 ;
        RECT -37.565 -154.525 -37.235 -154.195 ;
        RECT -37.565 -155.885 -37.235 -155.555 ;
        RECT -37.565 -157.245 -37.235 -156.915 ;
        RECT -37.565 -159.965 -37.235 -159.635 ;
        RECT -37.565 -162.685 -37.235 -162.355 ;
        RECT -37.565 -164.045 -37.235 -163.715 ;
        RECT -37.565 -165.405 -37.235 -165.075 ;
        RECT -37.565 -166.765 -37.235 -166.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 -29.405 -46.755 -29.075 ;
        RECT -47.085 -32.125 -46.755 -31.795 ;
        RECT -47.085 -33.485 -46.755 -33.155 ;
        RECT -47.085 -34.88 -46.755 -34.55 ;
        RECT -47.085 -36.205 -46.755 -35.875 ;
        RECT -47.085 -38.925 -46.755 -38.595 ;
        RECT -47.085 -39.97 -46.755 -39.64 ;
        RECT -47.085 -48.445 -46.755 -48.115 ;
        RECT -47.085 -49.805 -46.755 -49.475 ;
        RECT -47.085 -51.165 -46.755 -50.835 ;
        RECT -47.085 -53.885 -46.755 -53.555 ;
        RECT -47.085 -57.965 -46.755 -57.635 ;
        RECT -47.085 -62.045 -46.755 -61.715 ;
        RECT -47.085 -63.405 -46.755 -63.075 ;
        RECT -47.085 -64.765 -46.755 -64.435 ;
        RECT -47.085 -66.125 -46.755 -65.795 ;
        RECT -47.085 -67.485 -46.755 -67.155 ;
        RECT -47.085 -68.845 -46.755 -68.515 ;
        RECT -47.085 -70.205 -46.755 -69.875 ;
        RECT -47.085 -71.565 -46.755 -71.235 ;
        RECT -47.085 -72.925 -46.755 -72.595 ;
        RECT -47.085 -74.285 -46.755 -73.955 ;
        RECT -47.085 -75.645 -46.755 -75.315 ;
        RECT -47.085 -77.005 -46.755 -76.675 ;
        RECT -47.085 -78.365 -46.755 -78.035 ;
        RECT -47.085 -79.725 -46.755 -79.395 ;
        RECT -47.085 -81.085 -46.755 -80.755 ;
        RECT -47.085 -82.445 -46.755 -82.115 ;
        RECT -47.085 -83.805 -46.755 -83.475 ;
        RECT -47.085 -85.165 -46.755 -84.835 ;
        RECT -47.085 -86.525 -46.755 -86.195 ;
        RECT -47.085 -87.885 -46.755 -87.555 ;
        RECT -47.085 -89.245 -46.755 -88.915 ;
        RECT -47.085 -90.605 -46.755 -90.275 ;
        RECT -47.085 -91.965 -46.755 -91.635 ;
        RECT -47.085 -93.325 -46.755 -92.995 ;
        RECT -47.085 -94.685 -46.755 -94.355 ;
        RECT -47.085 -96.045 -46.755 -95.715 ;
        RECT -47.085 -97.405 -46.755 -97.075 ;
        RECT -47.085 -98.765 -46.755 -98.435 ;
        RECT -47.085 -100.125 -46.755 -99.795 ;
        RECT -47.085 -101.485 -46.755 -101.155 ;
        RECT -47.085 -102.845 -46.755 -102.515 ;
        RECT -47.085 -104.205 -46.755 -103.875 ;
        RECT -47.085 -105.565 -46.755 -105.235 ;
        RECT -47.085 -106.925 -46.755 -106.595 ;
        RECT -47.085 -108.285 -46.755 -107.955 ;
        RECT -47.085 -109.645 -46.755 -109.315 ;
        RECT -47.085 -111.005 -46.755 -110.675 ;
        RECT -47.085 -112.365 -46.755 -112.035 ;
        RECT -47.085 -113.725 -46.755 -113.395 ;
        RECT -47.085 -115.085 -46.755 -114.755 ;
        RECT -47.085 -116.445 -46.755 -116.115 ;
        RECT -47.085 -117.805 -46.755 -117.475 ;
        RECT -47.085 -119.165 -46.755 -118.835 ;
        RECT -47.085 -120.525 -46.755 -120.195 ;
        RECT -47.085 -128.685 -46.755 -128.355 ;
        RECT -47.085 -130.045 -46.755 -129.715 ;
        RECT -47.085 -132.765 -46.755 -132.435 ;
        RECT -47.085 -134.125 -46.755 -133.795 ;
        RECT -47.085 -135.485 -46.755 -135.155 ;
        RECT -47.085 -136.845 -46.755 -136.515 ;
        RECT -47.085 -138.205 -46.755 -137.875 ;
        RECT -47.085 -139.39 -46.755 -139.06 ;
        RECT -47.085 -140.925 -46.755 -140.595 ;
        RECT -47.085 -142.285 -46.755 -141.955 ;
        RECT -47.085 -145.005 -46.755 -144.675 ;
        RECT -47.085 -146.365 -46.755 -146.035 ;
        RECT -47.085 -148.03 -46.755 -147.7 ;
        RECT -47.085 -149.085 -46.755 -148.755 ;
        RECT -47.085 -150.445 -46.755 -150.115 ;
        RECT -47.085 -153.165 -46.755 -152.835 ;
        RECT -47.085 -154.525 -46.755 -154.195 ;
        RECT -47.085 -155.885 -46.755 -155.555 ;
        RECT -47.085 -157.245 -46.755 -156.915 ;
        RECT -47.085 -159.965 -46.755 -159.635 ;
        RECT -47.085 -162.685 -46.755 -162.355 ;
        RECT -47.085 -164.045 -46.755 -163.715 ;
        RECT -47.085 -165.405 -46.755 -165.075 ;
        RECT -47.085 -166.765 -46.755 -166.435 ;
        RECT -47.085 -168.125 -46.755 -167.795 ;
        RECT -47.085 -169.485 -46.755 -169.155 ;
        RECT -47.085 -170.845 -46.755 -170.515 ;
        RECT -47.085 -172.205 -46.755 -171.875 ;
        RECT -47.085 -173.565 -46.755 -173.235 ;
        RECT -47.085 -174.925 -46.755 -174.595 ;
        RECT -47.085 -176.285 -46.755 -175.955 ;
        RECT -47.085 -177.645 -46.755 -177.315 ;
        RECT -47.085 -179.005 -46.755 -178.675 ;
        RECT -47.085 -180.365 -46.755 -180.035 ;
        RECT -47.085 -181.725 -46.755 -181.395 ;
        RECT -47.085 -183.085 -46.755 -182.755 ;
        RECT -47.085 -184.445 -46.755 -184.115 ;
        RECT -47.085 -185.805 -46.755 -185.475 ;
        RECT -47.085 -187.165 -46.755 -186.835 ;
        RECT -47.085 -188.525 -46.755 -188.195 ;
        RECT -47.085 -189.885 -46.755 -189.555 ;
        RECT -47.085 -191.245 -46.755 -190.915 ;
        RECT -47.085 -192.605 -46.755 -192.275 ;
        RECT -47.085 -193.965 -46.755 -193.635 ;
        RECT -47.085 -195.325 -46.755 -194.995 ;
        RECT -47.085 -196.685 -46.755 -196.355 ;
        RECT -47.085 -198.045 -46.755 -197.715 ;
        RECT -47.085 -199.405 -46.755 -199.075 ;
        RECT -47.085 -200.765 -46.755 -200.435 ;
        RECT -47.085 -202.125 -46.755 -201.795 ;
        RECT -47.085 -203.485 -46.755 -203.155 ;
        RECT -47.085 -204.845 -46.755 -204.515 ;
        RECT -47.085 -206.205 -46.755 -205.875 ;
        RECT -47.085 -207.565 -46.755 -207.235 ;
        RECT -47.085 -208.925 -46.755 -208.595 ;
        RECT -47.085 -210.285 -46.755 -209.955 ;
        RECT -47.085 -211.645 -46.755 -211.315 ;
        RECT -47.085 -213.005 -46.755 -212.675 ;
        RECT -47.085 -214.365 -46.755 -214.035 ;
        RECT -47.085 -215.725 -46.755 -215.395 ;
        RECT -47.085 -217.085 -46.755 -216.755 ;
        RECT -47.085 -218.445 -46.755 -218.115 ;
        RECT -47.085 -219.805 -46.755 -219.475 ;
        RECT -47.085 -221.165 -46.755 -220.835 ;
        RECT -47.085 -222.525 -46.755 -222.195 ;
        RECT -47.085 -223.885 -46.755 -223.555 ;
        RECT -47.085 -225.245 -46.755 -224.915 ;
        RECT -47.085 -227.965 -46.755 -227.635 ;
        RECT -47.085 -232.045 -46.755 -231.715 ;
        RECT -47.085 -233.225 -46.755 -232.895 ;
        RECT -47.085 -234.765 -46.755 -234.435 ;
        RECT -47.085 -236.125 -46.755 -235.795 ;
        RECT -47.085 -237.485 -46.755 -237.155 ;
        RECT -47.085 -238.845 -46.755 -238.515 ;
        RECT -47.085 -241.09 -46.755 -239.96 ;
        RECT -47.08 -241.205 -46.76 -28.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 244.04 -45.395 245.17 ;
        RECT -45.725 242.595 -45.395 242.925 ;
        RECT -45.725 241.235 -45.395 241.565 ;
        RECT -45.725 239.875 -45.395 240.205 ;
        RECT -45.725 238.515 -45.395 238.845 ;
        RECT -45.725 237.155 -45.395 237.485 ;
        RECT -45.725 235.795 -45.395 236.125 ;
        RECT -45.725 234.435 -45.395 234.765 ;
        RECT -45.725 233.075 -45.395 233.405 ;
        RECT -45.725 231.715 -45.395 232.045 ;
        RECT -45.725 230.355 -45.395 230.685 ;
        RECT -45.725 228.995 -45.395 229.325 ;
        RECT -45.725 227.635 -45.395 227.965 ;
        RECT -45.725 226.275 -45.395 226.605 ;
        RECT -45.725 224.915 -45.395 225.245 ;
        RECT -45.725 223.555 -45.395 223.885 ;
        RECT -45.725 222.195 -45.395 222.525 ;
        RECT -45.725 220.835 -45.395 221.165 ;
        RECT -45.725 219.475 -45.395 219.805 ;
        RECT -45.725 218.115 -45.395 218.445 ;
        RECT -45.725 216.755 -45.395 217.085 ;
        RECT -45.725 215.395 -45.395 215.725 ;
        RECT -45.725 214.035 -45.395 214.365 ;
        RECT -45.725 212.675 -45.395 213.005 ;
        RECT -45.725 211.315 -45.395 211.645 ;
        RECT -45.725 209.955 -45.395 210.285 ;
        RECT -45.725 208.595 -45.395 208.925 ;
        RECT -45.725 207.235 -45.395 207.565 ;
        RECT -45.725 205.875 -45.395 206.205 ;
        RECT -45.725 204.515 -45.395 204.845 ;
        RECT -45.725 203.155 -45.395 203.485 ;
        RECT -45.725 201.795 -45.395 202.125 ;
        RECT -45.725 200.435 -45.395 200.765 ;
        RECT -45.725 199.075 -45.395 199.405 ;
        RECT -45.725 197.715 -45.395 198.045 ;
        RECT -45.725 196.355 -45.395 196.685 ;
        RECT -45.725 194.995 -45.395 195.325 ;
        RECT -45.725 193.635 -45.395 193.965 ;
        RECT -45.725 192.275 -45.395 192.605 ;
        RECT -45.725 190.915 -45.395 191.245 ;
        RECT -45.725 189.555 -45.395 189.885 ;
        RECT -45.725 188.195 -45.395 188.525 ;
        RECT -45.725 186.835 -45.395 187.165 ;
        RECT -45.725 185.475 -45.395 185.805 ;
        RECT -45.725 184.115 -45.395 184.445 ;
        RECT -45.725 182.755 -45.395 183.085 ;
        RECT -45.725 181.395 -45.395 181.725 ;
        RECT -45.725 180.035 -45.395 180.365 ;
        RECT -45.725 178.675 -45.395 179.005 ;
        RECT -45.725 177.315 -45.395 177.645 ;
        RECT -45.725 175.955 -45.395 176.285 ;
        RECT -45.725 174.595 -45.395 174.925 ;
        RECT -45.725 173.235 -45.395 173.565 ;
        RECT -45.725 171.875 -45.395 172.205 ;
        RECT -45.725 170.515 -45.395 170.845 ;
        RECT -45.725 169.155 -45.395 169.485 ;
        RECT -45.725 167.795 -45.395 168.125 ;
        RECT -45.725 166.435 -45.395 166.765 ;
        RECT -45.725 165.075 -45.395 165.405 ;
        RECT -45.725 163.715 -45.395 164.045 ;
        RECT -45.725 162.355 -45.395 162.685 ;
        RECT -45.725 160.995 -45.395 161.325 ;
        RECT -45.725 159.635 -45.395 159.965 ;
        RECT -45.725 158.275 -45.395 158.605 ;
        RECT -45.725 156.915 -45.395 157.245 ;
        RECT -45.725 155.555 -45.395 155.885 ;
        RECT -45.725 154.195 -45.395 154.525 ;
        RECT -45.725 152.835 -45.395 153.165 ;
        RECT -45.725 151.475 -45.395 151.805 ;
        RECT -45.725 150.115 -45.395 150.445 ;
        RECT -45.725 148.755 -45.395 149.085 ;
        RECT -45.725 147.395 -45.395 147.725 ;
        RECT -45.725 146.035 -45.395 146.365 ;
        RECT -45.725 144.675 -45.395 145.005 ;
        RECT -45.725 143.315 -45.395 143.645 ;
        RECT -45.725 141.955 -45.395 142.285 ;
        RECT -45.725 140.595 -45.395 140.925 ;
        RECT -45.725 139.235 -45.395 139.565 ;
        RECT -45.725 137.225 -45.395 137.555 ;
        RECT -45.725 135.175 -45.395 135.505 ;
        RECT -45.725 132.815 -45.395 133.145 ;
        RECT -45.725 131.665 -45.395 131.995 ;
        RECT -45.725 129.655 -45.395 129.985 ;
        RECT -45.725 128.505 -45.395 128.835 ;
        RECT -45.725 126.495 -45.395 126.825 ;
        RECT -45.725 125.345 -45.395 125.675 ;
        RECT -45.725 123.335 -45.395 123.665 ;
        RECT -45.725 122.185 -45.395 122.515 ;
        RECT -45.725 120.175 -45.395 120.505 ;
        RECT -45.725 119.025 -45.395 119.355 ;
        RECT -45.725 117.185 -45.395 117.515 ;
        RECT -45.725 115.865 -45.395 116.195 ;
        RECT -45.725 113.855 -45.395 114.185 ;
        RECT -45.725 112.705 -45.395 113.035 ;
        RECT -45.725 110.695 -45.395 111.025 ;
        RECT -45.725 109.545 -45.395 109.875 ;
        RECT -45.725 107.535 -45.395 107.865 ;
        RECT -45.725 106.385 -45.395 106.715 ;
        RECT -45.725 104.375 -45.395 104.705 ;
        RECT -45.725 103.225 -45.395 103.555 ;
        RECT -45.725 100.865 -45.395 101.195 ;
        RECT -45.725 98.81 -45.395 99.14 ;
        RECT -45.725 97.075 -45.395 97.405 ;
        RECT -45.725 95.715 -45.395 96.045 ;
        RECT -45.725 94.355 -45.395 94.685 ;
        RECT -45.725 92.995 -45.395 93.325 ;
        RECT -45.725 91.635 -45.395 91.965 ;
        RECT -45.725 90.275 -45.395 90.605 ;
        RECT -45.725 88.915 -45.395 89.245 ;
        RECT -45.725 87.555 -45.395 87.885 ;
        RECT -45.725 86.195 -45.395 86.525 ;
        RECT -45.725 84.835 -45.395 85.165 ;
        RECT -45.725 83.475 -45.395 83.805 ;
        RECT -45.725 82.115 -45.395 82.445 ;
        RECT -45.725 80.755 -45.395 81.085 ;
        RECT -45.725 79.395 -45.395 79.725 ;
        RECT -45.725 78.035 -45.395 78.365 ;
        RECT -45.725 76.675 -45.395 77.005 ;
        RECT -45.725 75.315 -45.395 75.645 ;
        RECT -45.725 73.955 -45.395 74.285 ;
        RECT -45.725 72.595 -45.395 72.925 ;
        RECT -45.725 71.235 -45.395 71.565 ;
        RECT -45.725 69.875 -45.395 70.205 ;
        RECT -45.725 68.515 -45.395 68.845 ;
        RECT -45.725 67.155 -45.395 67.485 ;
        RECT -45.725 65.795 -45.395 66.125 ;
        RECT -45.725 64.435 -45.395 64.765 ;
        RECT -45.725 63.075 -45.395 63.405 ;
        RECT -45.725 61.715 -45.395 62.045 ;
        RECT -45.725 60.355 -45.395 60.685 ;
        RECT -45.725 58.995 -45.395 59.325 ;
        RECT -45.725 57.635 -45.395 57.965 ;
        RECT -45.725 56.275 -45.395 56.605 ;
        RECT -45.725 54.915 -45.395 55.245 ;
        RECT -45.725 53.555 -45.395 53.885 ;
        RECT -45.725 52.195 -45.395 52.525 ;
        RECT -45.725 50.835 -45.395 51.165 ;
        RECT -45.725 49.475 -45.395 49.805 ;
        RECT -45.725 48.115 -45.395 48.445 ;
        RECT -45.725 46.755 -45.395 47.085 ;
        RECT -45.725 45.395 -45.395 45.725 ;
        RECT -45.725 44.035 -45.395 44.365 ;
        RECT -45.725 42.675 -45.395 43.005 ;
        RECT -45.725 41.315 -45.395 41.645 ;
        RECT -45.725 39.955 -45.395 40.285 ;
        RECT -45.725 38.595 -45.395 38.925 ;
        RECT -45.725 37.235 -45.395 37.565 ;
        RECT -45.725 35.875 -45.395 36.205 ;
        RECT -45.725 34.515 -45.395 34.845 ;
        RECT -45.725 33.155 -45.395 33.485 ;
        RECT -45.725 31.795 -45.395 32.125 ;
        RECT -45.725 30.435 -45.395 30.765 ;
        RECT -45.725 29.075 -45.395 29.405 ;
        RECT -45.725 27.715 -45.395 28.045 ;
        RECT -45.725 26.355 -45.395 26.685 ;
        RECT -45.725 24.995 -45.395 25.325 ;
        RECT -45.725 23.635 -45.395 23.965 ;
        RECT -45.725 22.275 -45.395 22.605 ;
        RECT -45.725 20.915 -45.395 21.245 ;
        RECT -45.725 19.555 -45.395 19.885 ;
        RECT -45.725 18.195 -45.395 18.525 ;
        RECT -45.725 16.835 -45.395 17.165 ;
        RECT -45.725 15.475 -45.395 15.805 ;
        RECT -45.725 14.115 -45.395 14.445 ;
        RECT -45.725 12.755 -45.395 13.085 ;
        RECT -45.725 11.395 -45.395 11.725 ;
        RECT -45.725 10.035 -45.395 10.365 ;
        RECT -45.725 8.675 -45.395 9.005 ;
        RECT -45.725 7.315 -45.395 7.645 ;
        RECT -45.725 5.955 -45.395 6.285 ;
        RECT -45.725 4.595 -45.395 4.925 ;
        RECT -45.725 3.235 -45.395 3.565 ;
        RECT -45.725 1.875 -45.395 2.205 ;
        RECT -45.725 0.515 -45.395 0.845 ;
        RECT -45.725 -0.845 -45.395 -0.515 ;
        RECT -45.725 -2.205 -45.395 -1.875 ;
        RECT -45.725 -4.925 -45.395 -4.595 ;
        RECT -45.725 -6.285 -45.395 -5.955 ;
        RECT -45.725 -7.645 -45.395 -7.315 ;
        RECT -45.725 -9.005 -45.395 -8.675 ;
        RECT -45.725 -10.365 -45.395 -10.035 ;
        RECT -45.725 -11.725 -45.395 -11.395 ;
        RECT -45.725 -13.085 -45.395 -12.755 ;
        RECT -45.725 -14.445 -45.395 -14.115 ;
        RECT -45.725 -15.805 -45.395 -15.475 ;
        RECT -45.725 -17.165 -45.395 -16.835 ;
        RECT -45.725 -18.525 -45.395 -18.195 ;
        RECT -45.725 -19.885 -45.395 -19.555 ;
        RECT -45.725 -21.245 -45.395 -20.915 ;
        RECT -45.725 -22.605 -45.395 -22.275 ;
        RECT -45.725 -23.965 -45.395 -23.635 ;
        RECT -45.725 -25.325 -45.395 -24.995 ;
        RECT -45.725 -29.405 -45.395 -29.075 ;
        RECT -45.725 -32.125 -45.395 -31.795 ;
        RECT -45.725 -33.485 -45.395 -33.155 ;
        RECT -45.725 -34.88 -45.395 -34.55 ;
        RECT -45.725 -36.205 -45.395 -35.875 ;
        RECT -45.725 -38.925 -45.395 -38.595 ;
        RECT -45.725 -39.97 -45.395 -39.64 ;
        RECT -45.725 -48.445 -45.395 -48.115 ;
        RECT -45.725 -49.805 -45.395 -49.475 ;
        RECT -45.725 -51.165 -45.395 -50.835 ;
        RECT -45.725 -53.885 -45.395 -53.555 ;
        RECT -45.725 -57.965 -45.395 -57.635 ;
        RECT -45.725 -62.045 -45.395 -61.715 ;
        RECT -45.725 -63.405 -45.395 -63.075 ;
        RECT -45.725 -64.765 -45.395 -64.435 ;
        RECT -45.725 -66.125 -45.395 -65.795 ;
        RECT -45.725 -67.485 -45.395 -67.155 ;
        RECT -45.725 -68.845 -45.395 -68.515 ;
        RECT -45.725 -70.205 -45.395 -69.875 ;
        RECT -45.725 -71.565 -45.395 -71.235 ;
        RECT -45.725 -72.925 -45.395 -72.595 ;
        RECT -45.725 -74.285 -45.395 -73.955 ;
        RECT -45.725 -75.645 -45.395 -75.315 ;
        RECT -45.725 -77.005 -45.395 -76.675 ;
        RECT -45.725 -78.365 -45.395 -78.035 ;
        RECT -45.725 -79.725 -45.395 -79.395 ;
        RECT -45.725 -81.085 -45.395 -80.755 ;
        RECT -45.725 -82.445 -45.395 -82.115 ;
        RECT -45.725 -83.805 -45.395 -83.475 ;
        RECT -45.725 -85.165 -45.395 -84.835 ;
        RECT -45.725 -86.525 -45.395 -86.195 ;
        RECT -45.725 -87.885 -45.395 -87.555 ;
        RECT -45.725 -89.245 -45.395 -88.915 ;
        RECT -45.725 -90.605 -45.395 -90.275 ;
        RECT -45.725 -91.965 -45.395 -91.635 ;
        RECT -45.725 -93.325 -45.395 -92.995 ;
        RECT -45.725 -94.685 -45.395 -94.355 ;
        RECT -45.725 -96.045 -45.395 -95.715 ;
        RECT -45.725 -97.405 -45.395 -97.075 ;
        RECT -45.725 -98.765 -45.395 -98.435 ;
        RECT -45.725 -100.125 -45.395 -99.795 ;
        RECT -45.725 -101.485 -45.395 -101.155 ;
        RECT -45.725 -102.845 -45.395 -102.515 ;
        RECT -45.725 -104.205 -45.395 -103.875 ;
        RECT -45.725 -105.565 -45.395 -105.235 ;
        RECT -45.725 -106.925 -45.395 -106.595 ;
        RECT -45.725 -108.285 -45.395 -107.955 ;
        RECT -45.725 -109.645 -45.395 -109.315 ;
        RECT -45.725 -111.005 -45.395 -110.675 ;
        RECT -45.725 -112.365 -45.395 -112.035 ;
        RECT -45.725 -113.725 -45.395 -113.395 ;
        RECT -45.725 -115.085 -45.395 -114.755 ;
        RECT -45.725 -116.445 -45.395 -116.115 ;
        RECT -45.725 -117.805 -45.395 -117.475 ;
        RECT -45.725 -119.165 -45.395 -118.835 ;
        RECT -45.725 -120.525 -45.395 -120.195 ;
        RECT -45.725 -128.685 -45.395 -128.355 ;
        RECT -45.725 -130.045 -45.395 -129.715 ;
        RECT -45.725 -132.765 -45.395 -132.435 ;
        RECT -45.725 -134.125 -45.395 -133.795 ;
        RECT -45.725 -135.485 -45.395 -135.155 ;
        RECT -45.725 -136.845 -45.395 -136.515 ;
        RECT -45.725 -138.205 -45.395 -137.875 ;
        RECT -45.725 -139.39 -45.395 -139.06 ;
        RECT -45.725 -140.925 -45.395 -140.595 ;
        RECT -45.725 -142.285 -45.395 -141.955 ;
        RECT -45.725 -145.005 -45.395 -144.675 ;
        RECT -45.725 -146.365 -45.395 -146.035 ;
        RECT -45.725 -148.03 -45.395 -147.7 ;
        RECT -45.725 -149.085 -45.395 -148.755 ;
        RECT -45.725 -150.445 -45.395 -150.115 ;
        RECT -45.725 -153.165 -45.395 -152.835 ;
        RECT -45.725 -154.525 -45.395 -154.195 ;
        RECT -45.725 -155.885 -45.395 -155.555 ;
        RECT -45.725 -157.245 -45.395 -156.915 ;
        RECT -45.725 -159.965 -45.395 -159.635 ;
        RECT -45.725 -162.685 -45.395 -162.355 ;
        RECT -45.725 -164.045 -45.395 -163.715 ;
        RECT -45.725 -165.405 -45.395 -165.075 ;
        RECT -45.725 -166.765 -45.395 -166.435 ;
        RECT -45.725 -168.125 -45.395 -167.795 ;
        RECT -45.725 -169.485 -45.395 -169.155 ;
        RECT -45.725 -170.845 -45.395 -170.515 ;
        RECT -45.725 -172.205 -45.395 -171.875 ;
        RECT -45.725 -173.565 -45.395 -173.235 ;
        RECT -45.725 -174.925 -45.395 -174.595 ;
        RECT -45.725 -176.285 -45.395 -175.955 ;
        RECT -45.725 -177.645 -45.395 -177.315 ;
        RECT -45.725 -179.005 -45.395 -178.675 ;
        RECT -45.725 -180.365 -45.395 -180.035 ;
        RECT -45.725 -181.725 -45.395 -181.395 ;
        RECT -45.725 -183.085 -45.395 -182.755 ;
        RECT -45.725 -184.445 -45.395 -184.115 ;
        RECT -45.725 -185.805 -45.395 -185.475 ;
        RECT -45.725 -187.165 -45.395 -186.835 ;
        RECT -45.725 -188.525 -45.395 -188.195 ;
        RECT -45.725 -189.885 -45.395 -189.555 ;
        RECT -45.725 -191.245 -45.395 -190.915 ;
        RECT -45.725 -192.605 -45.395 -192.275 ;
        RECT -45.725 -193.965 -45.395 -193.635 ;
        RECT -45.725 -195.325 -45.395 -194.995 ;
        RECT -45.725 -196.685 -45.395 -196.355 ;
        RECT -45.725 -198.045 -45.395 -197.715 ;
        RECT -45.725 -199.405 -45.395 -199.075 ;
        RECT -45.725 -200.765 -45.395 -200.435 ;
        RECT -45.725 -202.125 -45.395 -201.795 ;
        RECT -45.725 -203.485 -45.395 -203.155 ;
        RECT -45.725 -204.845 -45.395 -204.515 ;
        RECT -45.725 -206.205 -45.395 -205.875 ;
        RECT -45.725 -207.565 -45.395 -207.235 ;
        RECT -45.725 -208.925 -45.395 -208.595 ;
        RECT -45.725 -210.285 -45.395 -209.955 ;
        RECT -45.725 -211.645 -45.395 -211.315 ;
        RECT -45.725 -213.005 -45.395 -212.675 ;
        RECT -45.725 -214.365 -45.395 -214.035 ;
        RECT -45.725 -215.725 -45.395 -215.395 ;
        RECT -45.725 -217.085 -45.395 -216.755 ;
        RECT -45.725 -218.445 -45.395 -218.115 ;
        RECT -45.725 -219.805 -45.395 -219.475 ;
        RECT -45.725 -221.165 -45.395 -220.835 ;
        RECT -45.725 -222.525 -45.395 -222.195 ;
        RECT -45.725 -223.885 -45.395 -223.555 ;
        RECT -45.725 -225.245 -45.395 -224.915 ;
        RECT -45.725 -227.965 -45.395 -227.635 ;
        RECT -45.725 -230.685 -45.395 -230.355 ;
        RECT -45.725 -232.045 -45.395 -231.715 ;
        RECT -45.725 -233.225 -45.395 -232.895 ;
        RECT -45.725 -234.765 -45.395 -234.435 ;
        RECT -45.725 -236.125 -45.395 -235.795 ;
        RECT -45.725 -237.485 -45.395 -237.155 ;
        RECT -45.725 -238.845 -45.395 -238.515 ;
        RECT -45.725 -241.09 -45.395 -239.96 ;
        RECT -45.72 -241.205 -45.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 244.04 -44.035 245.17 ;
        RECT -44.365 242.595 -44.035 242.925 ;
        RECT -44.365 241.235 -44.035 241.565 ;
        RECT -44.365 239.875 -44.035 240.205 ;
        RECT -44.365 238.515 -44.035 238.845 ;
        RECT -44.365 237.155 -44.035 237.485 ;
        RECT -44.365 235.795 -44.035 236.125 ;
        RECT -44.365 234.435 -44.035 234.765 ;
        RECT -44.365 233.075 -44.035 233.405 ;
        RECT -44.365 231.715 -44.035 232.045 ;
        RECT -44.365 230.355 -44.035 230.685 ;
        RECT -44.365 228.995 -44.035 229.325 ;
        RECT -44.365 227.635 -44.035 227.965 ;
        RECT -44.365 226.275 -44.035 226.605 ;
        RECT -44.365 224.915 -44.035 225.245 ;
        RECT -44.365 223.555 -44.035 223.885 ;
        RECT -44.365 222.195 -44.035 222.525 ;
        RECT -44.365 220.835 -44.035 221.165 ;
        RECT -44.365 219.475 -44.035 219.805 ;
        RECT -44.365 218.115 -44.035 218.445 ;
        RECT -44.365 216.755 -44.035 217.085 ;
        RECT -44.365 215.395 -44.035 215.725 ;
        RECT -44.365 214.035 -44.035 214.365 ;
        RECT -44.365 212.675 -44.035 213.005 ;
        RECT -44.365 211.315 -44.035 211.645 ;
        RECT -44.365 209.955 -44.035 210.285 ;
        RECT -44.365 208.595 -44.035 208.925 ;
        RECT -44.365 207.235 -44.035 207.565 ;
        RECT -44.365 205.875 -44.035 206.205 ;
        RECT -44.365 204.515 -44.035 204.845 ;
        RECT -44.365 203.155 -44.035 203.485 ;
        RECT -44.365 201.795 -44.035 202.125 ;
        RECT -44.365 200.435 -44.035 200.765 ;
        RECT -44.365 199.075 -44.035 199.405 ;
        RECT -44.365 197.715 -44.035 198.045 ;
        RECT -44.365 196.355 -44.035 196.685 ;
        RECT -44.365 194.995 -44.035 195.325 ;
        RECT -44.365 193.635 -44.035 193.965 ;
        RECT -44.365 192.275 -44.035 192.605 ;
        RECT -44.365 190.915 -44.035 191.245 ;
        RECT -44.365 189.555 -44.035 189.885 ;
        RECT -44.365 188.195 -44.035 188.525 ;
        RECT -44.365 186.835 -44.035 187.165 ;
        RECT -44.365 185.475 -44.035 185.805 ;
        RECT -44.365 184.115 -44.035 184.445 ;
        RECT -44.365 182.755 -44.035 183.085 ;
        RECT -44.365 181.395 -44.035 181.725 ;
        RECT -44.365 180.035 -44.035 180.365 ;
        RECT -44.365 178.675 -44.035 179.005 ;
        RECT -44.365 177.315 -44.035 177.645 ;
        RECT -44.365 175.955 -44.035 176.285 ;
        RECT -44.365 174.595 -44.035 174.925 ;
        RECT -44.365 173.235 -44.035 173.565 ;
        RECT -44.365 171.875 -44.035 172.205 ;
        RECT -44.365 170.515 -44.035 170.845 ;
        RECT -44.365 169.155 -44.035 169.485 ;
        RECT -44.365 167.795 -44.035 168.125 ;
        RECT -44.365 166.435 -44.035 166.765 ;
        RECT -44.365 165.075 -44.035 165.405 ;
        RECT -44.365 163.715 -44.035 164.045 ;
        RECT -44.365 162.355 -44.035 162.685 ;
        RECT -44.365 160.995 -44.035 161.325 ;
        RECT -44.365 159.635 -44.035 159.965 ;
        RECT -44.365 158.275 -44.035 158.605 ;
        RECT -44.365 156.915 -44.035 157.245 ;
        RECT -44.365 155.555 -44.035 155.885 ;
        RECT -44.365 154.195 -44.035 154.525 ;
        RECT -44.365 152.835 -44.035 153.165 ;
        RECT -44.365 151.475 -44.035 151.805 ;
        RECT -44.365 150.115 -44.035 150.445 ;
        RECT -44.365 148.755 -44.035 149.085 ;
        RECT -44.365 147.395 -44.035 147.725 ;
        RECT -44.365 146.035 -44.035 146.365 ;
        RECT -44.365 144.675 -44.035 145.005 ;
        RECT -44.365 143.315 -44.035 143.645 ;
        RECT -44.365 141.955 -44.035 142.285 ;
        RECT -44.365 140.595 -44.035 140.925 ;
        RECT -44.365 139.235 -44.035 139.565 ;
        RECT -44.365 97.075 -44.035 97.405 ;
        RECT -44.365 95.715 -44.035 96.045 ;
        RECT -44.365 94.355 -44.035 94.685 ;
        RECT -44.365 92.995 -44.035 93.325 ;
        RECT -44.365 91.635 -44.035 91.965 ;
        RECT -44.365 90.275 -44.035 90.605 ;
        RECT -44.365 88.915 -44.035 89.245 ;
        RECT -44.365 87.555 -44.035 87.885 ;
        RECT -44.365 86.195 -44.035 86.525 ;
        RECT -44.365 84.835 -44.035 85.165 ;
        RECT -44.365 83.475 -44.035 83.805 ;
        RECT -44.365 82.115 -44.035 82.445 ;
        RECT -44.365 80.755 -44.035 81.085 ;
        RECT -44.365 79.395 -44.035 79.725 ;
        RECT -44.365 78.035 -44.035 78.365 ;
        RECT -44.365 76.675 -44.035 77.005 ;
        RECT -44.365 75.315 -44.035 75.645 ;
        RECT -44.365 73.955 -44.035 74.285 ;
        RECT -44.365 72.595 -44.035 72.925 ;
        RECT -44.365 71.235 -44.035 71.565 ;
        RECT -44.365 69.875 -44.035 70.205 ;
        RECT -44.365 68.515 -44.035 68.845 ;
        RECT -44.365 67.155 -44.035 67.485 ;
        RECT -44.365 65.795 -44.035 66.125 ;
        RECT -44.365 64.435 -44.035 64.765 ;
        RECT -44.365 63.075 -44.035 63.405 ;
        RECT -44.365 61.715 -44.035 62.045 ;
        RECT -44.365 60.355 -44.035 60.685 ;
        RECT -44.365 58.995 -44.035 59.325 ;
        RECT -44.365 57.635 -44.035 57.965 ;
        RECT -44.365 56.275 -44.035 56.605 ;
        RECT -44.365 54.915 -44.035 55.245 ;
        RECT -44.365 53.555 -44.035 53.885 ;
        RECT -44.365 52.195 -44.035 52.525 ;
        RECT -44.365 50.835 -44.035 51.165 ;
        RECT -44.365 49.475 -44.035 49.805 ;
        RECT -44.365 48.115 -44.035 48.445 ;
        RECT -44.365 46.755 -44.035 47.085 ;
        RECT -44.365 45.395 -44.035 45.725 ;
        RECT -44.365 44.035 -44.035 44.365 ;
        RECT -44.365 42.675 -44.035 43.005 ;
        RECT -44.365 41.315 -44.035 41.645 ;
        RECT -44.365 39.955 -44.035 40.285 ;
        RECT -44.365 38.595 -44.035 38.925 ;
        RECT -44.365 37.235 -44.035 37.565 ;
        RECT -44.365 35.875 -44.035 36.205 ;
        RECT -44.365 34.515 -44.035 34.845 ;
        RECT -44.365 33.155 -44.035 33.485 ;
        RECT -44.365 31.795 -44.035 32.125 ;
        RECT -44.365 30.435 -44.035 30.765 ;
        RECT -44.365 29.075 -44.035 29.405 ;
        RECT -44.365 27.715 -44.035 28.045 ;
        RECT -44.365 26.355 -44.035 26.685 ;
        RECT -44.365 24.995 -44.035 25.325 ;
        RECT -44.365 23.635 -44.035 23.965 ;
        RECT -44.365 22.275 -44.035 22.605 ;
        RECT -44.365 20.915 -44.035 21.245 ;
        RECT -44.365 19.555 -44.035 19.885 ;
        RECT -44.365 18.195 -44.035 18.525 ;
        RECT -44.365 16.835 -44.035 17.165 ;
        RECT -44.365 15.475 -44.035 15.805 ;
        RECT -44.365 14.115 -44.035 14.445 ;
        RECT -44.365 12.755 -44.035 13.085 ;
        RECT -44.365 11.395 -44.035 11.725 ;
        RECT -44.365 10.035 -44.035 10.365 ;
        RECT -44.365 8.675 -44.035 9.005 ;
        RECT -44.365 7.315 -44.035 7.645 ;
        RECT -44.365 5.955 -44.035 6.285 ;
        RECT -44.365 4.595 -44.035 4.925 ;
        RECT -44.365 3.235 -44.035 3.565 ;
        RECT -44.365 1.875 -44.035 2.205 ;
        RECT -44.365 0.515 -44.035 0.845 ;
        RECT -44.365 -0.845 -44.035 -0.515 ;
        RECT -44.365 -2.205 -44.035 -1.875 ;
        RECT -44.365 -4.925 -44.035 -4.595 ;
        RECT -44.365 -6.285 -44.035 -5.955 ;
        RECT -44.365 -7.645 -44.035 -7.315 ;
        RECT -44.365 -9.005 -44.035 -8.675 ;
        RECT -44.365 -10.365 -44.035 -10.035 ;
        RECT -44.365 -11.725 -44.035 -11.395 ;
        RECT -44.365 -13.085 -44.035 -12.755 ;
        RECT -44.365 -14.445 -44.035 -14.115 ;
        RECT -44.365 -15.805 -44.035 -15.475 ;
        RECT -44.365 -17.165 -44.035 -16.835 ;
        RECT -44.365 -18.525 -44.035 -18.195 ;
        RECT -44.365 -19.885 -44.035 -19.555 ;
        RECT -44.365 -21.245 -44.035 -20.915 ;
        RECT -44.365 -22.605 -44.035 -22.275 ;
        RECT -44.365 -23.965 -44.035 -23.635 ;
        RECT -44.365 -29.405 -44.035 -29.075 ;
        RECT -44.365 -32.125 -44.035 -31.795 ;
        RECT -44.365 -33.485 -44.035 -33.155 ;
        RECT -44.365 -34.88 -44.035 -34.55 ;
        RECT -44.365 -36.205 -44.035 -35.875 ;
        RECT -44.365 -38.925 -44.035 -38.595 ;
        RECT -44.365 -39.97 -44.035 -39.64 ;
        RECT -44.365 -48.445 -44.035 -48.115 ;
        RECT -44.365 -49.805 -44.035 -49.475 ;
        RECT -44.365 -51.165 -44.035 -50.835 ;
        RECT -44.365 -53.885 -44.035 -53.555 ;
        RECT -44.365 -57.965 -44.035 -57.635 ;
        RECT -44.36 -58.64 -44.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 -128.685 -44.035 -128.355 ;
        RECT -44.365 -130.045 -44.035 -129.715 ;
        RECT -44.365 -132.765 -44.035 -132.435 ;
        RECT -44.365 -134.125 -44.035 -133.795 ;
        RECT -44.365 -135.485 -44.035 -135.155 ;
        RECT -44.365 -136.845 -44.035 -136.515 ;
        RECT -44.365 -138.205 -44.035 -137.875 ;
        RECT -44.365 -139.39 -44.035 -139.06 ;
        RECT -44.365 -140.925 -44.035 -140.595 ;
        RECT -44.365 -142.285 -44.035 -141.955 ;
        RECT -44.365 -145.005 -44.035 -144.675 ;
        RECT -44.365 -146.365 -44.035 -146.035 ;
        RECT -44.365 -148.03 -44.035 -147.7 ;
        RECT -44.365 -149.085 -44.035 -148.755 ;
        RECT -44.365 -150.445 -44.035 -150.115 ;
        RECT -44.365 -153.165 -44.035 -152.835 ;
        RECT -44.365 -154.525 -44.035 -154.195 ;
        RECT -44.365 -155.885 -44.035 -155.555 ;
        RECT -44.365 -157.245 -44.035 -156.915 ;
        RECT -44.365 -159.965 -44.035 -159.635 ;
        RECT -44.365 -162.685 -44.035 -162.355 ;
        RECT -44.365 -164.045 -44.035 -163.715 ;
        RECT -44.365 -165.405 -44.035 -165.075 ;
        RECT -44.365 -166.765 -44.035 -166.435 ;
        RECT -44.365 -168.125 -44.035 -167.795 ;
        RECT -44.365 -169.485 -44.035 -169.155 ;
        RECT -44.365 -170.845 -44.035 -170.515 ;
        RECT -44.365 -172.205 -44.035 -171.875 ;
        RECT -44.365 -173.565 -44.035 -173.235 ;
        RECT -44.365 -174.925 -44.035 -174.595 ;
        RECT -44.365 -176.285 -44.035 -175.955 ;
        RECT -44.365 -177.645 -44.035 -177.315 ;
        RECT -44.365 -179.005 -44.035 -178.675 ;
        RECT -44.365 -180.365 -44.035 -180.035 ;
        RECT -44.365 -181.725 -44.035 -181.395 ;
        RECT -44.365 -183.085 -44.035 -182.755 ;
        RECT -44.365 -184.445 -44.035 -184.115 ;
        RECT -44.365 -185.805 -44.035 -185.475 ;
        RECT -44.365 -187.165 -44.035 -186.835 ;
        RECT -44.365 -188.525 -44.035 -188.195 ;
        RECT -44.365 -189.885 -44.035 -189.555 ;
        RECT -44.365 -191.245 -44.035 -190.915 ;
        RECT -44.365 -192.605 -44.035 -192.275 ;
        RECT -44.365 -193.965 -44.035 -193.635 ;
        RECT -44.365 -195.325 -44.035 -194.995 ;
        RECT -44.365 -196.685 -44.035 -196.355 ;
        RECT -44.365 -198.045 -44.035 -197.715 ;
        RECT -44.365 -199.405 -44.035 -199.075 ;
        RECT -44.365 -200.765 -44.035 -200.435 ;
        RECT -44.365 -202.125 -44.035 -201.795 ;
        RECT -44.365 -203.485 -44.035 -203.155 ;
        RECT -44.365 -204.845 -44.035 -204.515 ;
        RECT -44.365 -206.205 -44.035 -205.875 ;
        RECT -44.365 -207.565 -44.035 -207.235 ;
        RECT -44.365 -208.925 -44.035 -208.595 ;
        RECT -44.365 -210.285 -44.035 -209.955 ;
        RECT -44.365 -211.645 -44.035 -211.315 ;
        RECT -44.365 -213.005 -44.035 -212.675 ;
        RECT -44.365 -214.365 -44.035 -214.035 ;
        RECT -44.365 -215.725 -44.035 -215.395 ;
        RECT -44.365 -217.085 -44.035 -216.755 ;
        RECT -44.365 -218.445 -44.035 -218.115 ;
        RECT -44.365 -219.805 -44.035 -219.475 ;
        RECT -44.365 -221.165 -44.035 -220.835 ;
        RECT -44.365 -222.525 -44.035 -222.195 ;
        RECT -44.365 -223.885 -44.035 -223.555 ;
        RECT -44.365 -225.245 -44.035 -224.915 ;
        RECT -44.365 -227.965 -44.035 -227.635 ;
        RECT -44.365 -230.685 -44.035 -230.355 ;
        RECT -44.365 -232.045 -44.035 -231.715 ;
        RECT -44.365 -233.225 -44.035 -232.895 ;
        RECT -44.365 -234.765 -44.035 -234.435 ;
        RECT -44.365 -236.125 -44.035 -235.795 ;
        RECT -44.365 -237.485 -44.035 -237.155 ;
        RECT -44.365 -238.845 -44.035 -238.515 ;
        RECT -44.365 -241.09 -44.035 -239.96 ;
        RECT -44.36 -241.205 -44.04 -122.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 239.875 -42.675 240.205 ;
        RECT -43.005 238.515 -42.675 238.845 ;
        RECT -43.005 237.155 -42.675 237.485 ;
        RECT -43.005 235.795 -42.675 236.125 ;
        RECT -43.005 234.435 -42.675 234.765 ;
        RECT -43.005 233.075 -42.675 233.405 ;
        RECT -43.005 231.715 -42.675 232.045 ;
        RECT -43.005 230.355 -42.675 230.685 ;
        RECT -43.005 228.995 -42.675 229.325 ;
        RECT -43.005 227.635 -42.675 227.965 ;
        RECT -43.005 226.275 -42.675 226.605 ;
        RECT -43.005 224.915 -42.675 225.245 ;
        RECT -43.005 223.555 -42.675 223.885 ;
        RECT -43.005 222.195 -42.675 222.525 ;
        RECT -43.005 220.835 -42.675 221.165 ;
        RECT -43.005 219.475 -42.675 219.805 ;
        RECT -43.005 218.115 -42.675 218.445 ;
        RECT -43.005 216.755 -42.675 217.085 ;
        RECT -43.005 215.395 -42.675 215.725 ;
        RECT -43.005 214.035 -42.675 214.365 ;
        RECT -43.005 212.675 -42.675 213.005 ;
        RECT -43.005 211.315 -42.675 211.645 ;
        RECT -43.005 209.955 -42.675 210.285 ;
        RECT -43.005 208.595 -42.675 208.925 ;
        RECT -43.005 207.235 -42.675 207.565 ;
        RECT -43.005 205.875 -42.675 206.205 ;
        RECT -43.005 204.515 -42.675 204.845 ;
        RECT -43.005 203.155 -42.675 203.485 ;
        RECT -43.005 201.795 -42.675 202.125 ;
        RECT -43.005 200.435 -42.675 200.765 ;
        RECT -43.005 199.075 -42.675 199.405 ;
        RECT -43.005 197.715 -42.675 198.045 ;
        RECT -43.005 196.355 -42.675 196.685 ;
        RECT -43.005 194.995 -42.675 195.325 ;
        RECT -43.005 193.635 -42.675 193.965 ;
        RECT -43.005 192.275 -42.675 192.605 ;
        RECT -43.005 190.915 -42.675 191.245 ;
        RECT -43.005 189.555 -42.675 189.885 ;
        RECT -43.005 188.195 -42.675 188.525 ;
        RECT -43.005 186.835 -42.675 187.165 ;
        RECT -43.005 185.475 -42.675 185.805 ;
        RECT -43.005 184.115 -42.675 184.445 ;
        RECT -43.005 182.755 -42.675 183.085 ;
        RECT -43.005 181.395 -42.675 181.725 ;
        RECT -43.005 180.035 -42.675 180.365 ;
        RECT -43.005 178.675 -42.675 179.005 ;
        RECT -43.005 177.315 -42.675 177.645 ;
        RECT -43.005 175.955 -42.675 176.285 ;
        RECT -43.005 174.595 -42.675 174.925 ;
        RECT -43.005 173.235 -42.675 173.565 ;
        RECT -43.005 171.875 -42.675 172.205 ;
        RECT -43.005 170.515 -42.675 170.845 ;
        RECT -43.005 169.155 -42.675 169.485 ;
        RECT -43.005 167.795 -42.675 168.125 ;
        RECT -43.005 166.435 -42.675 166.765 ;
        RECT -43.005 165.075 -42.675 165.405 ;
        RECT -43.005 163.715 -42.675 164.045 ;
        RECT -43.005 162.355 -42.675 162.685 ;
        RECT -43.005 160.995 -42.675 161.325 ;
        RECT -43.005 159.635 -42.675 159.965 ;
        RECT -43.005 158.275 -42.675 158.605 ;
        RECT -43.005 156.915 -42.675 157.245 ;
        RECT -43.005 155.555 -42.675 155.885 ;
        RECT -43.005 154.195 -42.675 154.525 ;
        RECT -43.005 152.835 -42.675 153.165 ;
        RECT -43.005 151.475 -42.675 151.805 ;
        RECT -43.005 150.115 -42.675 150.445 ;
        RECT -43.005 148.755 -42.675 149.085 ;
        RECT -43.005 147.395 -42.675 147.725 ;
        RECT -43.005 146.035 -42.675 146.365 ;
        RECT -43.005 144.675 -42.675 145.005 ;
        RECT -43.005 143.315 -42.675 143.645 ;
        RECT -43.005 141.955 -42.675 142.285 ;
        RECT -43.005 140.595 -42.675 140.925 ;
        RECT -43.005 139.235 -42.675 139.565 ;
        RECT -43.005 137.875 -42.675 138.205 ;
        RECT -43.005 136.515 -42.675 136.845 ;
        RECT -43.005 135.155 -42.675 135.485 ;
        RECT -43.005 133.795 -42.675 134.125 ;
        RECT -43.005 132.435 -42.675 132.765 ;
        RECT -43.005 131.075 -42.675 131.405 ;
        RECT -43.005 129.715 -42.675 130.045 ;
        RECT -43.005 128.355 -42.675 128.685 ;
        RECT -43.005 126.995 -42.675 127.325 ;
        RECT -43.005 125.635 -42.675 125.965 ;
        RECT -43.005 124.275 -42.675 124.605 ;
        RECT -43.005 122.915 -42.675 123.245 ;
        RECT -43.005 121.555 -42.675 121.885 ;
        RECT -43.005 120.195 -42.675 120.525 ;
        RECT -43.005 118.835 -42.675 119.165 ;
        RECT -43.005 117.475 -42.675 117.805 ;
        RECT -43.005 116.115 -42.675 116.445 ;
        RECT -43.005 114.755 -42.675 115.085 ;
        RECT -43.005 113.395 -42.675 113.725 ;
        RECT -43.005 112.035 -42.675 112.365 ;
        RECT -43.005 110.675 -42.675 111.005 ;
        RECT -43.005 109.315 -42.675 109.645 ;
        RECT -43.005 107.955 -42.675 108.285 ;
        RECT -43.005 106.595 -42.675 106.925 ;
        RECT -43.005 105.235 -42.675 105.565 ;
        RECT -43.005 103.875 -42.675 104.205 ;
        RECT -43.005 102.515 -42.675 102.845 ;
        RECT -43.005 101.155 -42.675 101.485 ;
        RECT -43.005 99.795 -42.675 100.125 ;
        RECT -43.005 98.435 -42.675 98.765 ;
        RECT -43.005 97.075 -42.675 97.405 ;
        RECT -43.005 95.715 -42.675 96.045 ;
        RECT -43.005 94.355 -42.675 94.685 ;
        RECT -43.005 92.995 -42.675 93.325 ;
        RECT -43.005 91.635 -42.675 91.965 ;
        RECT -43.005 90.275 -42.675 90.605 ;
        RECT -43.005 88.915 -42.675 89.245 ;
        RECT -43.005 87.555 -42.675 87.885 ;
        RECT -43.005 86.195 -42.675 86.525 ;
        RECT -43.005 84.835 -42.675 85.165 ;
        RECT -43.005 83.475 -42.675 83.805 ;
        RECT -43.005 82.115 -42.675 82.445 ;
        RECT -43.005 80.755 -42.675 81.085 ;
        RECT -43.005 79.395 -42.675 79.725 ;
        RECT -43.005 78.035 -42.675 78.365 ;
        RECT -43.005 76.675 -42.675 77.005 ;
        RECT -43.005 75.315 -42.675 75.645 ;
        RECT -43.005 73.955 -42.675 74.285 ;
        RECT -43.005 72.595 -42.675 72.925 ;
        RECT -43.005 71.235 -42.675 71.565 ;
        RECT -43.005 69.875 -42.675 70.205 ;
        RECT -43.005 68.515 -42.675 68.845 ;
        RECT -43.005 67.155 -42.675 67.485 ;
        RECT -43.005 65.795 -42.675 66.125 ;
        RECT -43.005 64.435 -42.675 64.765 ;
        RECT -43.005 63.075 -42.675 63.405 ;
        RECT -43.005 61.715 -42.675 62.045 ;
        RECT -43.005 60.355 -42.675 60.685 ;
        RECT -43.005 58.995 -42.675 59.325 ;
        RECT -43.005 57.635 -42.675 57.965 ;
        RECT -43.005 56.275 -42.675 56.605 ;
        RECT -43.005 54.915 -42.675 55.245 ;
        RECT -43.005 53.555 -42.675 53.885 ;
        RECT -43.005 52.195 -42.675 52.525 ;
        RECT -43.005 50.835 -42.675 51.165 ;
        RECT -43.005 49.475 -42.675 49.805 ;
        RECT -43.005 48.115 -42.675 48.445 ;
        RECT -43.005 46.755 -42.675 47.085 ;
        RECT -43.005 45.395 -42.675 45.725 ;
        RECT -43.005 44.035 -42.675 44.365 ;
        RECT -43.005 42.675 -42.675 43.005 ;
        RECT -43.005 41.315 -42.675 41.645 ;
        RECT -43.005 39.955 -42.675 40.285 ;
        RECT -43.005 38.595 -42.675 38.925 ;
        RECT -43.005 37.235 -42.675 37.565 ;
        RECT -43.005 35.875 -42.675 36.205 ;
        RECT -43.005 34.515 -42.675 34.845 ;
        RECT -43.005 33.155 -42.675 33.485 ;
        RECT -43.005 31.795 -42.675 32.125 ;
        RECT -43.005 30.435 -42.675 30.765 ;
        RECT -43.005 29.075 -42.675 29.405 ;
        RECT -43.005 27.715 -42.675 28.045 ;
        RECT -43.005 26.355 -42.675 26.685 ;
        RECT -43.005 24.995 -42.675 25.325 ;
        RECT -43.005 23.635 -42.675 23.965 ;
        RECT -43.005 22.275 -42.675 22.605 ;
        RECT -43.005 20.915 -42.675 21.245 ;
        RECT -43.005 19.555 -42.675 19.885 ;
        RECT -43.005 18.195 -42.675 18.525 ;
        RECT -43.005 16.835 -42.675 17.165 ;
        RECT -43.005 15.475 -42.675 15.805 ;
        RECT -43.005 14.115 -42.675 14.445 ;
        RECT -43.005 12.755 -42.675 13.085 ;
        RECT -43.005 11.395 -42.675 11.725 ;
        RECT -43.005 10.035 -42.675 10.365 ;
        RECT -43.005 8.675 -42.675 9.005 ;
        RECT -43.005 7.315 -42.675 7.645 ;
        RECT -43.005 5.955 -42.675 6.285 ;
        RECT -43.005 4.595 -42.675 4.925 ;
        RECT -43.005 3.235 -42.675 3.565 ;
        RECT -43.005 1.875 -42.675 2.205 ;
        RECT -43.005 0.515 -42.675 0.845 ;
        RECT -43.005 -0.845 -42.675 -0.515 ;
        RECT -43.005 -2.205 -42.675 -1.875 ;
        RECT -43.005 -4.925 -42.675 -4.595 ;
        RECT -43.005 -6.285 -42.675 -5.955 ;
        RECT -43.005 -7.645 -42.675 -7.315 ;
        RECT -43.005 -9.005 -42.675 -8.675 ;
        RECT -43.005 -10.365 -42.675 -10.035 ;
        RECT -43.005 -11.725 -42.675 -11.395 ;
        RECT -43.005 -13.085 -42.675 -12.755 ;
        RECT -43.005 -14.445 -42.675 -14.115 ;
        RECT -43.005 -15.805 -42.675 -15.475 ;
        RECT -43.005 -17.165 -42.675 -16.835 ;
        RECT -43.005 -18.525 -42.675 -18.195 ;
        RECT -43.005 -19.885 -42.675 -19.555 ;
        RECT -43.005 -21.245 -42.675 -20.915 ;
        RECT -43.005 -22.605 -42.675 -22.275 ;
        RECT -43.005 -29.405 -42.675 -29.075 ;
        RECT -43.005 -32.125 -42.675 -31.795 ;
        RECT -43.005 -33.485 -42.675 -33.155 ;
        RECT -43.005 -34.88 -42.675 -34.55 ;
        RECT -43.005 -36.205 -42.675 -35.875 ;
        RECT -43.005 -38.925 -42.675 -38.595 ;
        RECT -43.005 -39.97 -42.675 -39.64 ;
        RECT -43.005 -48.445 -42.675 -48.115 ;
        RECT -43.005 -49.805 -42.675 -49.475 ;
        RECT -43.005 -51.165 -42.675 -50.835 ;
        RECT -43.005 -53.885 -42.675 -53.555 ;
        RECT -43.005 -57.965 -42.675 -57.635 ;
        RECT -43 -57.965 -42.68 245.285 ;
        RECT -43.005 244.04 -42.675 245.17 ;
        RECT -43.005 242.595 -42.675 242.925 ;
        RECT -43.005 241.235 -42.675 241.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 244.04 -50.835 245.17 ;
        RECT -51.165 242.595 -50.835 242.925 ;
        RECT -51.165 241.235 -50.835 241.565 ;
        RECT -51.165 239.875 -50.835 240.205 ;
        RECT -51.165 238.515 -50.835 238.845 ;
        RECT -51.165 237.155 -50.835 237.485 ;
        RECT -51.165 235.795 -50.835 236.125 ;
        RECT -51.165 234.435 -50.835 234.765 ;
        RECT -51.165 233.075 -50.835 233.405 ;
        RECT -51.165 231.715 -50.835 232.045 ;
        RECT -51.165 230.355 -50.835 230.685 ;
        RECT -51.165 228.995 -50.835 229.325 ;
        RECT -51.165 227.635 -50.835 227.965 ;
        RECT -51.165 226.275 -50.835 226.605 ;
        RECT -51.165 224.915 -50.835 225.245 ;
        RECT -51.165 223.555 -50.835 223.885 ;
        RECT -51.165 222.195 -50.835 222.525 ;
        RECT -51.165 220.835 -50.835 221.165 ;
        RECT -51.165 219.475 -50.835 219.805 ;
        RECT -51.165 218.115 -50.835 218.445 ;
        RECT -51.165 216.755 -50.835 217.085 ;
        RECT -51.165 215.395 -50.835 215.725 ;
        RECT -51.165 214.035 -50.835 214.365 ;
        RECT -51.165 212.675 -50.835 213.005 ;
        RECT -51.165 211.315 -50.835 211.645 ;
        RECT -51.165 209.955 -50.835 210.285 ;
        RECT -51.165 208.595 -50.835 208.925 ;
        RECT -51.165 207.235 -50.835 207.565 ;
        RECT -51.165 205.875 -50.835 206.205 ;
        RECT -51.165 204.515 -50.835 204.845 ;
        RECT -51.165 203.155 -50.835 203.485 ;
        RECT -51.165 201.795 -50.835 202.125 ;
        RECT -51.165 200.435 -50.835 200.765 ;
        RECT -51.165 199.075 -50.835 199.405 ;
        RECT -51.165 197.715 -50.835 198.045 ;
        RECT -51.165 196.355 -50.835 196.685 ;
        RECT -51.165 194.995 -50.835 195.325 ;
        RECT -51.165 193.635 -50.835 193.965 ;
        RECT -51.165 192.275 -50.835 192.605 ;
        RECT -51.165 190.915 -50.835 191.245 ;
        RECT -51.165 189.555 -50.835 189.885 ;
        RECT -51.165 188.195 -50.835 188.525 ;
        RECT -51.165 186.835 -50.835 187.165 ;
        RECT -51.165 185.475 -50.835 185.805 ;
        RECT -51.165 184.115 -50.835 184.445 ;
        RECT -51.165 182.755 -50.835 183.085 ;
        RECT -51.165 181.395 -50.835 181.725 ;
        RECT -51.165 180.035 -50.835 180.365 ;
        RECT -51.165 178.675 -50.835 179.005 ;
        RECT -51.165 177.315 -50.835 177.645 ;
        RECT -51.165 175.955 -50.835 176.285 ;
        RECT -51.165 174.595 -50.835 174.925 ;
        RECT -51.165 173.235 -50.835 173.565 ;
        RECT -51.165 171.875 -50.835 172.205 ;
        RECT -51.165 170.515 -50.835 170.845 ;
        RECT -51.165 169.155 -50.835 169.485 ;
        RECT -51.165 167.795 -50.835 168.125 ;
        RECT -51.165 166.435 -50.835 166.765 ;
        RECT -51.165 165.075 -50.835 165.405 ;
        RECT -51.165 163.715 -50.835 164.045 ;
        RECT -51.165 162.355 -50.835 162.685 ;
        RECT -51.165 160.995 -50.835 161.325 ;
        RECT -51.165 159.635 -50.835 159.965 ;
        RECT -51.165 158.275 -50.835 158.605 ;
        RECT -51.165 156.915 -50.835 157.245 ;
        RECT -51.165 155.555 -50.835 155.885 ;
        RECT -51.165 154.195 -50.835 154.525 ;
        RECT -51.165 152.835 -50.835 153.165 ;
        RECT -51.165 151.475 -50.835 151.805 ;
        RECT -51.165 150.115 -50.835 150.445 ;
        RECT -51.165 148.755 -50.835 149.085 ;
        RECT -51.165 147.395 -50.835 147.725 ;
        RECT -51.165 146.035 -50.835 146.365 ;
        RECT -51.165 144.675 -50.835 145.005 ;
        RECT -51.165 143.315 -50.835 143.645 ;
        RECT -51.165 141.955 -50.835 142.285 ;
        RECT -51.165 140.595 -50.835 140.925 ;
        RECT -51.165 139.235 -50.835 139.565 ;
        RECT -51.16 138.56 -50.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 97.075 -50.835 97.405 ;
        RECT -51.165 95.715 -50.835 96.045 ;
        RECT -51.165 94.355 -50.835 94.685 ;
        RECT -51.165 92.995 -50.835 93.325 ;
        RECT -51.165 88.915 -50.835 89.245 ;
        RECT -51.165 84.835 -50.835 85.165 ;
        RECT -51.165 83.475 -50.835 83.805 ;
        RECT -51.165 82.115 -50.835 82.445 ;
        RECT -51.165 80.755 -50.835 81.085 ;
        RECT -51.165 79.395 -50.835 79.725 ;
        RECT -51.165 78.035 -50.835 78.365 ;
        RECT -51.165 76.675 -50.835 77.005 ;
        RECT -51.165 75.315 -50.835 75.645 ;
        RECT -51.165 73.955 -50.835 74.285 ;
        RECT -51.165 72.595 -50.835 72.925 ;
        RECT -51.165 71.235 -50.835 71.565 ;
        RECT -51.165 69.875 -50.835 70.205 ;
        RECT -51.165 68.515 -50.835 68.845 ;
        RECT -51.165 67.155 -50.835 67.485 ;
        RECT -51.165 65.795 -50.835 66.125 ;
        RECT -51.165 64.435 -50.835 64.765 ;
        RECT -51.165 63.075 -50.835 63.405 ;
        RECT -51.165 61.715 -50.835 62.045 ;
        RECT -51.165 60.355 -50.835 60.685 ;
        RECT -51.165 58.995 -50.835 59.325 ;
        RECT -51.165 57.635 -50.835 57.965 ;
        RECT -51.165 56.275 -50.835 56.605 ;
        RECT -51.165 54.915 -50.835 55.245 ;
        RECT -51.165 53.555 -50.835 53.885 ;
        RECT -51.165 52.195 -50.835 52.525 ;
        RECT -51.165 50.835 -50.835 51.165 ;
        RECT -51.165 49.475 -50.835 49.805 ;
        RECT -51.165 48.115 -50.835 48.445 ;
        RECT -51.165 46.755 -50.835 47.085 ;
        RECT -51.165 45.395 -50.835 45.725 ;
        RECT -51.165 44.035 -50.835 44.365 ;
        RECT -51.165 42.675 -50.835 43.005 ;
        RECT -51.165 41.315 -50.835 41.645 ;
        RECT -51.165 39.955 -50.835 40.285 ;
        RECT -51.165 38.595 -50.835 38.925 ;
        RECT -51.165 37.235 -50.835 37.565 ;
        RECT -51.165 35.875 -50.835 36.205 ;
        RECT -51.165 34.515 -50.835 34.845 ;
        RECT -51.165 33.155 -50.835 33.485 ;
        RECT -51.165 31.795 -50.835 32.125 ;
        RECT -51.165 30.435 -50.835 30.765 ;
        RECT -51.165 29.075 -50.835 29.405 ;
        RECT -51.165 27.715 -50.835 28.045 ;
        RECT -51.165 26.355 -50.835 26.685 ;
        RECT -51.165 24.995 -50.835 25.325 ;
        RECT -51.165 23.635 -50.835 23.965 ;
        RECT -51.165 22.275 -50.835 22.605 ;
        RECT -51.165 20.915 -50.835 21.245 ;
        RECT -51.165 19.555 -50.835 19.885 ;
        RECT -51.165 18.195 -50.835 18.525 ;
        RECT -51.165 16.835 -50.835 17.165 ;
        RECT -51.165 15.475 -50.835 15.805 ;
        RECT -51.165 14.115 -50.835 14.445 ;
        RECT -51.165 12.755 -50.835 13.085 ;
        RECT -51.165 11.395 -50.835 11.725 ;
        RECT -51.165 10.035 -50.835 10.365 ;
        RECT -51.165 8.675 -50.835 9.005 ;
        RECT -51.165 7.315 -50.835 7.645 ;
        RECT -51.165 5.955 -50.835 6.285 ;
        RECT -51.165 4.595 -50.835 4.925 ;
        RECT -51.165 3.235 -50.835 3.565 ;
        RECT -51.165 1.875 -50.835 2.205 ;
        RECT -51.165 0.515 -50.835 0.845 ;
        RECT -51.165 -0.845 -50.835 -0.515 ;
        RECT -51.165 -2.205 -50.835 -1.875 ;
        RECT -51.165 -3.565 -50.835 -3.235 ;
        RECT -51.165 -4.925 -50.835 -4.595 ;
        RECT -51.165 -6.285 -50.835 -5.955 ;
        RECT -51.165 -7.645 -50.835 -7.315 ;
        RECT -51.165 -9.005 -50.835 -8.675 ;
        RECT -51.165 -10.365 -50.835 -10.035 ;
        RECT -51.165 -11.725 -50.835 -11.395 ;
        RECT -51.165 -13.085 -50.835 -12.755 ;
        RECT -51.165 -14.445 -50.835 -14.115 ;
        RECT -51.165 -15.805 -50.835 -15.475 ;
        RECT -51.165 -17.165 -50.835 -16.835 ;
        RECT -51.165 -18.525 -50.835 -18.195 ;
        RECT -51.165 -19.885 -50.835 -19.555 ;
        RECT -51.165 -21.245 -50.835 -20.915 ;
        RECT -51.165 -22.605 -50.835 -22.275 ;
        RECT -51.165 -23.965 -50.835 -23.635 ;
        RECT -51.165 -25.325 -50.835 -24.995 ;
        RECT -51.165 -26.685 -50.835 -26.355 ;
        RECT -51.165 -28.045 -50.835 -27.715 ;
        RECT -51.165 -29.405 -50.835 -29.075 ;
        RECT -51.165 -30.765 -50.835 -30.435 ;
        RECT -51.165 -32.125 -50.835 -31.795 ;
        RECT -51.165 -33.485 -50.835 -33.155 ;
        RECT -51.165 -34.845 -50.835 -34.515 ;
        RECT -51.165 -36.205 -50.835 -35.875 ;
        RECT -51.165 -37.565 -50.835 -37.235 ;
        RECT -51.165 -38.925 -50.835 -38.595 ;
        RECT -51.165 -40.285 -50.835 -39.955 ;
        RECT -51.165 -41.645 -50.835 -41.315 ;
        RECT -51.165 -43.005 -50.835 -42.675 ;
        RECT -51.165 -44.365 -50.835 -44.035 ;
        RECT -51.165 -45.725 -50.835 -45.395 ;
        RECT -51.165 -47.085 -50.835 -46.755 ;
        RECT -51.165 -48.445 -50.835 -48.115 ;
        RECT -51.165 -49.805 -50.835 -49.475 ;
        RECT -51.165 -51.165 -50.835 -50.835 ;
        RECT -51.165 -52.525 -50.835 -52.195 ;
        RECT -51.165 -53.885 -50.835 -53.555 ;
        RECT -51.165 -55.245 -50.835 -54.915 ;
        RECT -51.165 -56.605 -50.835 -56.275 ;
        RECT -51.165 -57.965 -50.835 -57.635 ;
        RECT -51.165 -59.325 -50.835 -58.995 ;
        RECT -51.165 -60.685 -50.835 -60.355 ;
        RECT -51.165 -62.045 -50.835 -61.715 ;
        RECT -51.165 -63.405 -50.835 -63.075 ;
        RECT -51.165 -64.765 -50.835 -64.435 ;
        RECT -51.165 -66.125 -50.835 -65.795 ;
        RECT -51.165 -67.485 -50.835 -67.155 ;
        RECT -51.165 -68.845 -50.835 -68.515 ;
        RECT -51.165 -70.205 -50.835 -69.875 ;
        RECT -51.165 -71.565 -50.835 -71.235 ;
        RECT -51.165 -72.925 -50.835 -72.595 ;
        RECT -51.165 -74.285 -50.835 -73.955 ;
        RECT -51.165 -75.645 -50.835 -75.315 ;
        RECT -51.165 -77.005 -50.835 -76.675 ;
        RECT -51.165 -78.365 -50.835 -78.035 ;
        RECT -51.165 -79.725 -50.835 -79.395 ;
        RECT -51.165 -81.085 -50.835 -80.755 ;
        RECT -51.165 -82.445 -50.835 -82.115 ;
        RECT -51.165 -83.805 -50.835 -83.475 ;
        RECT -51.165 -85.165 -50.835 -84.835 ;
        RECT -51.165 -86.525 -50.835 -86.195 ;
        RECT -51.165 -87.885 -50.835 -87.555 ;
        RECT -51.165 -89.245 -50.835 -88.915 ;
        RECT -51.165 -90.605 -50.835 -90.275 ;
        RECT -51.165 -91.965 -50.835 -91.635 ;
        RECT -51.165 -93.325 -50.835 -92.995 ;
        RECT -51.165 -94.685 -50.835 -94.355 ;
        RECT -51.165 -96.045 -50.835 -95.715 ;
        RECT -51.165 -97.405 -50.835 -97.075 ;
        RECT -51.165 -98.765 -50.835 -98.435 ;
        RECT -51.165 -100.125 -50.835 -99.795 ;
        RECT -51.165 -101.485 -50.835 -101.155 ;
        RECT -51.165 -102.845 -50.835 -102.515 ;
        RECT -51.165 -104.205 -50.835 -103.875 ;
        RECT -51.165 -105.565 -50.835 -105.235 ;
        RECT -51.165 -106.925 -50.835 -106.595 ;
        RECT -51.165 -108.285 -50.835 -107.955 ;
        RECT -51.165 -109.645 -50.835 -109.315 ;
        RECT -51.165 -111.005 -50.835 -110.675 ;
        RECT -51.165 -112.365 -50.835 -112.035 ;
        RECT -51.165 -113.725 -50.835 -113.395 ;
        RECT -51.165 -115.085 -50.835 -114.755 ;
        RECT -51.165 -116.445 -50.835 -116.115 ;
        RECT -51.165 -117.805 -50.835 -117.475 ;
        RECT -51.165 -119.165 -50.835 -118.835 ;
        RECT -51.165 -120.525 -50.835 -120.195 ;
        RECT -51.165 -121.885 -50.835 -121.555 ;
        RECT -51.165 -128.685 -50.835 -128.355 ;
        RECT -51.165 -130.045 -50.835 -129.715 ;
        RECT -51.165 -132.765 -50.835 -132.435 ;
        RECT -51.165 -134.125 -50.835 -133.795 ;
        RECT -51.165 -135.485 -50.835 -135.155 ;
        RECT -51.165 -136.845 -50.835 -136.515 ;
        RECT -51.165 -138.205 -50.835 -137.875 ;
        RECT -51.165 -139.39 -50.835 -139.06 ;
        RECT -51.165 -140.925 -50.835 -140.595 ;
        RECT -51.165 -142.285 -50.835 -141.955 ;
        RECT -51.165 -145.005 -50.835 -144.675 ;
        RECT -51.165 -146.365 -50.835 -146.035 ;
        RECT -51.165 -148.03 -50.835 -147.7 ;
        RECT -51.165 -149.085 -50.835 -148.755 ;
        RECT -51.165 -150.445 -50.835 -150.115 ;
        RECT -51.165 -153.165 -50.835 -152.835 ;
        RECT -51.165 -154.525 -50.835 -154.195 ;
        RECT -51.165 -155.885 -50.835 -155.555 ;
        RECT -51.165 -157.245 -50.835 -156.915 ;
        RECT -51.165 -158.605 -50.835 -158.275 ;
        RECT -51.165 -159.965 -50.835 -159.635 ;
        RECT -51.165 -162.685 -50.835 -162.355 ;
        RECT -51.165 -164.045 -50.835 -163.715 ;
        RECT -51.165 -165.405 -50.835 -165.075 ;
        RECT -51.165 -166.765 -50.835 -166.435 ;
        RECT -51.165 -168.125 -50.835 -167.795 ;
        RECT -51.165 -169.485 -50.835 -169.155 ;
        RECT -51.165 -170.845 -50.835 -170.515 ;
        RECT -51.165 -172.205 -50.835 -171.875 ;
        RECT -51.165 -173.565 -50.835 -173.235 ;
        RECT -51.165 -174.925 -50.835 -174.595 ;
        RECT -51.165 -176.285 -50.835 -175.955 ;
        RECT -51.165 -177.645 -50.835 -177.315 ;
        RECT -51.165 -179.005 -50.835 -178.675 ;
        RECT -51.165 -180.365 -50.835 -180.035 ;
        RECT -51.165 -181.725 -50.835 -181.395 ;
        RECT -51.165 -183.085 -50.835 -182.755 ;
        RECT -51.165 -184.445 -50.835 -184.115 ;
        RECT -51.165 -185.805 -50.835 -185.475 ;
        RECT -51.165 -187.165 -50.835 -186.835 ;
        RECT -51.165 -188.525 -50.835 -188.195 ;
        RECT -51.165 -189.885 -50.835 -189.555 ;
        RECT -51.165 -191.245 -50.835 -190.915 ;
        RECT -51.165 -192.605 -50.835 -192.275 ;
        RECT -51.165 -193.965 -50.835 -193.635 ;
        RECT -51.165 -195.325 -50.835 -194.995 ;
        RECT -51.165 -196.685 -50.835 -196.355 ;
        RECT -51.165 -198.045 -50.835 -197.715 ;
        RECT -51.165 -199.405 -50.835 -199.075 ;
        RECT -51.165 -200.765 -50.835 -200.435 ;
        RECT -51.165 -202.125 -50.835 -201.795 ;
        RECT -51.165 -203.485 -50.835 -203.155 ;
        RECT -51.165 -204.845 -50.835 -204.515 ;
        RECT -51.165 -206.205 -50.835 -205.875 ;
        RECT -51.165 -207.565 -50.835 -207.235 ;
        RECT -51.165 -208.925 -50.835 -208.595 ;
        RECT -51.165 -210.285 -50.835 -209.955 ;
        RECT -51.165 -211.645 -50.835 -211.315 ;
        RECT -51.165 -213.005 -50.835 -212.675 ;
        RECT -51.165 -214.365 -50.835 -214.035 ;
        RECT -51.165 -215.725 -50.835 -215.395 ;
        RECT -51.165 -217.085 -50.835 -216.755 ;
        RECT -51.165 -218.445 -50.835 -218.115 ;
        RECT -51.165 -219.805 -50.835 -219.475 ;
        RECT -51.165 -221.165 -50.835 -220.835 ;
        RECT -51.165 -222.525 -50.835 -222.195 ;
        RECT -51.165 -223.885 -50.835 -223.555 ;
        RECT -51.165 -225.245 -50.835 -224.915 ;
        RECT -51.165 -227.965 -50.835 -227.635 ;
        RECT -51.165 -230.685 -50.835 -230.355 ;
        RECT -51.165 -232.045 -50.835 -231.715 ;
        RECT -51.165 -233.225 -50.835 -232.895 ;
        RECT -51.165 -234.765 -50.835 -234.435 ;
        RECT -51.165 -236.125 -50.835 -235.795 ;
        RECT -51.165 -237.485 -50.835 -237.155 ;
        RECT -51.165 -238.845 -50.835 -238.515 ;
        RECT -51.165 -241.09 -50.835 -239.96 ;
        RECT -51.16 -241.205 -50.84 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 244.04 -49.475 245.17 ;
        RECT -49.805 242.595 -49.475 242.925 ;
        RECT -49.805 241.235 -49.475 241.565 ;
        RECT -49.805 239.875 -49.475 240.205 ;
        RECT -49.805 238.515 -49.475 238.845 ;
        RECT -49.805 237.155 -49.475 237.485 ;
        RECT -49.805 235.795 -49.475 236.125 ;
        RECT -49.805 234.435 -49.475 234.765 ;
        RECT -49.805 233.075 -49.475 233.405 ;
        RECT -49.805 231.715 -49.475 232.045 ;
        RECT -49.805 230.355 -49.475 230.685 ;
        RECT -49.805 228.995 -49.475 229.325 ;
        RECT -49.805 227.635 -49.475 227.965 ;
        RECT -49.805 226.275 -49.475 226.605 ;
        RECT -49.805 224.915 -49.475 225.245 ;
        RECT -49.805 223.555 -49.475 223.885 ;
        RECT -49.805 222.195 -49.475 222.525 ;
        RECT -49.805 220.835 -49.475 221.165 ;
        RECT -49.805 219.475 -49.475 219.805 ;
        RECT -49.805 218.115 -49.475 218.445 ;
        RECT -49.805 216.755 -49.475 217.085 ;
        RECT -49.805 215.395 -49.475 215.725 ;
        RECT -49.805 214.035 -49.475 214.365 ;
        RECT -49.805 212.675 -49.475 213.005 ;
        RECT -49.805 211.315 -49.475 211.645 ;
        RECT -49.805 209.955 -49.475 210.285 ;
        RECT -49.805 208.595 -49.475 208.925 ;
        RECT -49.805 207.235 -49.475 207.565 ;
        RECT -49.805 205.875 -49.475 206.205 ;
        RECT -49.805 204.515 -49.475 204.845 ;
        RECT -49.805 203.155 -49.475 203.485 ;
        RECT -49.805 201.795 -49.475 202.125 ;
        RECT -49.805 200.435 -49.475 200.765 ;
        RECT -49.805 199.075 -49.475 199.405 ;
        RECT -49.805 197.715 -49.475 198.045 ;
        RECT -49.805 196.355 -49.475 196.685 ;
        RECT -49.805 194.995 -49.475 195.325 ;
        RECT -49.805 193.635 -49.475 193.965 ;
        RECT -49.805 192.275 -49.475 192.605 ;
        RECT -49.805 190.915 -49.475 191.245 ;
        RECT -49.805 189.555 -49.475 189.885 ;
        RECT -49.805 188.195 -49.475 188.525 ;
        RECT -49.805 186.835 -49.475 187.165 ;
        RECT -49.805 185.475 -49.475 185.805 ;
        RECT -49.805 184.115 -49.475 184.445 ;
        RECT -49.805 182.755 -49.475 183.085 ;
        RECT -49.805 181.395 -49.475 181.725 ;
        RECT -49.805 180.035 -49.475 180.365 ;
        RECT -49.805 178.675 -49.475 179.005 ;
        RECT -49.805 177.315 -49.475 177.645 ;
        RECT -49.805 175.955 -49.475 176.285 ;
        RECT -49.805 174.595 -49.475 174.925 ;
        RECT -49.805 173.235 -49.475 173.565 ;
        RECT -49.805 171.875 -49.475 172.205 ;
        RECT -49.805 170.515 -49.475 170.845 ;
        RECT -49.805 169.155 -49.475 169.485 ;
        RECT -49.805 167.795 -49.475 168.125 ;
        RECT -49.805 166.435 -49.475 166.765 ;
        RECT -49.805 165.075 -49.475 165.405 ;
        RECT -49.805 163.715 -49.475 164.045 ;
        RECT -49.805 162.355 -49.475 162.685 ;
        RECT -49.805 160.995 -49.475 161.325 ;
        RECT -49.805 159.635 -49.475 159.965 ;
        RECT -49.805 158.275 -49.475 158.605 ;
        RECT -49.805 156.915 -49.475 157.245 ;
        RECT -49.805 155.555 -49.475 155.885 ;
        RECT -49.805 154.195 -49.475 154.525 ;
        RECT -49.805 152.835 -49.475 153.165 ;
        RECT -49.805 151.475 -49.475 151.805 ;
        RECT -49.805 150.115 -49.475 150.445 ;
        RECT -49.805 148.755 -49.475 149.085 ;
        RECT -49.805 147.395 -49.475 147.725 ;
        RECT -49.805 146.035 -49.475 146.365 ;
        RECT -49.805 144.675 -49.475 145.005 ;
        RECT -49.805 143.315 -49.475 143.645 ;
        RECT -49.805 141.955 -49.475 142.285 ;
        RECT -49.805 140.595 -49.475 140.925 ;
        RECT -49.805 139.235 -49.475 139.565 ;
        RECT -49.8 138.56 -49.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 97.075 -49.475 97.405 ;
        RECT -49.805 95.715 -49.475 96.045 ;
        RECT -49.805 94.355 -49.475 94.685 ;
        RECT -49.805 92.995 -49.475 93.325 ;
        RECT -49.805 88.915 -49.475 89.245 ;
        RECT -49.805 84.835 -49.475 85.165 ;
        RECT -49.805 83.475 -49.475 83.805 ;
        RECT -49.805 82.115 -49.475 82.445 ;
        RECT -49.805 80.755 -49.475 81.085 ;
        RECT -49.805 79.395 -49.475 79.725 ;
        RECT -49.805 78.035 -49.475 78.365 ;
        RECT -49.805 76.675 -49.475 77.005 ;
        RECT -49.805 75.315 -49.475 75.645 ;
        RECT -49.805 73.955 -49.475 74.285 ;
        RECT -49.805 72.595 -49.475 72.925 ;
        RECT -49.805 71.235 -49.475 71.565 ;
        RECT -49.805 69.875 -49.475 70.205 ;
        RECT -49.805 68.515 -49.475 68.845 ;
        RECT -49.805 67.155 -49.475 67.485 ;
        RECT -49.805 65.795 -49.475 66.125 ;
        RECT -49.805 64.435 -49.475 64.765 ;
        RECT -49.805 63.075 -49.475 63.405 ;
        RECT -49.805 61.715 -49.475 62.045 ;
        RECT -49.805 60.355 -49.475 60.685 ;
        RECT -49.805 58.995 -49.475 59.325 ;
        RECT -49.805 57.635 -49.475 57.965 ;
        RECT -49.805 56.275 -49.475 56.605 ;
        RECT -49.805 54.915 -49.475 55.245 ;
        RECT -49.805 53.555 -49.475 53.885 ;
        RECT -49.805 52.195 -49.475 52.525 ;
        RECT -49.805 50.835 -49.475 51.165 ;
        RECT -49.805 49.475 -49.475 49.805 ;
        RECT -49.805 48.115 -49.475 48.445 ;
        RECT -49.805 46.755 -49.475 47.085 ;
        RECT -49.805 45.395 -49.475 45.725 ;
        RECT -49.805 44.035 -49.475 44.365 ;
        RECT -49.805 42.675 -49.475 43.005 ;
        RECT -49.805 41.315 -49.475 41.645 ;
        RECT -49.805 39.955 -49.475 40.285 ;
        RECT -49.805 38.595 -49.475 38.925 ;
        RECT -49.805 37.235 -49.475 37.565 ;
        RECT -49.805 35.875 -49.475 36.205 ;
        RECT -49.805 34.515 -49.475 34.845 ;
        RECT -49.805 33.155 -49.475 33.485 ;
        RECT -49.805 31.795 -49.475 32.125 ;
        RECT -49.805 30.435 -49.475 30.765 ;
        RECT -49.805 29.075 -49.475 29.405 ;
        RECT -49.805 27.715 -49.475 28.045 ;
        RECT -49.805 26.355 -49.475 26.685 ;
        RECT -49.805 24.995 -49.475 25.325 ;
        RECT -49.805 23.635 -49.475 23.965 ;
        RECT -49.805 22.275 -49.475 22.605 ;
        RECT -49.805 20.915 -49.475 21.245 ;
        RECT -49.805 19.555 -49.475 19.885 ;
        RECT -49.805 18.195 -49.475 18.525 ;
        RECT -49.805 16.835 -49.475 17.165 ;
        RECT -49.805 15.475 -49.475 15.805 ;
        RECT -49.805 14.115 -49.475 14.445 ;
        RECT -49.805 12.755 -49.475 13.085 ;
        RECT -49.805 11.395 -49.475 11.725 ;
        RECT -49.805 10.035 -49.475 10.365 ;
        RECT -49.805 8.675 -49.475 9.005 ;
        RECT -49.805 7.315 -49.475 7.645 ;
        RECT -49.805 5.955 -49.475 6.285 ;
        RECT -49.805 4.595 -49.475 4.925 ;
        RECT -49.805 3.235 -49.475 3.565 ;
        RECT -49.805 1.875 -49.475 2.205 ;
        RECT -49.805 0.515 -49.475 0.845 ;
        RECT -49.805 -0.845 -49.475 -0.515 ;
        RECT -49.805 -2.205 -49.475 -1.875 ;
        RECT -49.805 -3.565 -49.475 -3.235 ;
        RECT -49.805 -4.925 -49.475 -4.595 ;
        RECT -49.805 -6.285 -49.475 -5.955 ;
        RECT -49.805 -7.645 -49.475 -7.315 ;
        RECT -49.805 -9.005 -49.475 -8.675 ;
        RECT -49.805 -10.365 -49.475 -10.035 ;
        RECT -49.805 -11.725 -49.475 -11.395 ;
        RECT -49.805 -13.085 -49.475 -12.755 ;
        RECT -49.805 -14.445 -49.475 -14.115 ;
        RECT -49.805 -15.805 -49.475 -15.475 ;
        RECT -49.805 -17.165 -49.475 -16.835 ;
        RECT -49.805 -18.525 -49.475 -18.195 ;
        RECT -49.805 -19.885 -49.475 -19.555 ;
        RECT -49.805 -21.245 -49.475 -20.915 ;
        RECT -49.805 -22.605 -49.475 -22.275 ;
        RECT -49.805 -23.965 -49.475 -23.635 ;
        RECT -49.805 -25.325 -49.475 -24.995 ;
        RECT -49.805 -26.685 -49.475 -26.355 ;
        RECT -49.805 -28.045 -49.475 -27.715 ;
        RECT -49.805 -29.405 -49.475 -29.075 ;
        RECT -49.805 -32.125 -49.475 -31.795 ;
        RECT -49.805 -33.485 -49.475 -33.155 ;
        RECT -49.805 -36.205 -49.475 -35.875 ;
        RECT -49.805 -38.925 -49.475 -38.595 ;
        RECT -49.805 -48.445 -49.475 -48.115 ;
        RECT -49.805 -49.805 -49.475 -49.475 ;
        RECT -49.805 -51.165 -49.475 -50.835 ;
        RECT -49.805 -53.885 -49.475 -53.555 ;
        RECT -49.805 -57.965 -49.475 -57.635 ;
        RECT -49.805 -62.045 -49.475 -61.715 ;
        RECT -49.805 -63.405 -49.475 -63.075 ;
        RECT -49.805 -64.765 -49.475 -64.435 ;
        RECT -49.805 -66.125 -49.475 -65.795 ;
        RECT -49.805 -67.485 -49.475 -67.155 ;
        RECT -49.805 -68.845 -49.475 -68.515 ;
        RECT -49.805 -70.205 -49.475 -69.875 ;
        RECT -49.805 -71.565 -49.475 -71.235 ;
        RECT -49.805 -72.925 -49.475 -72.595 ;
        RECT -49.805 -74.285 -49.475 -73.955 ;
        RECT -49.805 -75.645 -49.475 -75.315 ;
        RECT -49.805 -77.005 -49.475 -76.675 ;
        RECT -49.805 -78.365 -49.475 -78.035 ;
        RECT -49.805 -79.725 -49.475 -79.395 ;
        RECT -49.805 -81.085 -49.475 -80.755 ;
        RECT -49.805 -82.445 -49.475 -82.115 ;
        RECT -49.805 -83.805 -49.475 -83.475 ;
        RECT -49.805 -85.165 -49.475 -84.835 ;
        RECT -49.805 -86.525 -49.475 -86.195 ;
        RECT -49.805 -87.885 -49.475 -87.555 ;
        RECT -49.805 -89.245 -49.475 -88.915 ;
        RECT -49.805 -90.605 -49.475 -90.275 ;
        RECT -49.805 -91.965 -49.475 -91.635 ;
        RECT -49.805 -93.325 -49.475 -92.995 ;
        RECT -49.805 -94.685 -49.475 -94.355 ;
        RECT -49.805 -96.045 -49.475 -95.715 ;
        RECT -49.805 -97.405 -49.475 -97.075 ;
        RECT -49.805 -98.765 -49.475 -98.435 ;
        RECT -49.805 -100.125 -49.475 -99.795 ;
        RECT -49.805 -101.485 -49.475 -101.155 ;
        RECT -49.805 -102.845 -49.475 -102.515 ;
        RECT -49.805 -104.205 -49.475 -103.875 ;
        RECT -49.805 -105.565 -49.475 -105.235 ;
        RECT -49.805 -106.925 -49.475 -106.595 ;
        RECT -49.805 -108.285 -49.475 -107.955 ;
        RECT -49.805 -109.645 -49.475 -109.315 ;
        RECT -49.805 -111.005 -49.475 -110.675 ;
        RECT -49.805 -112.365 -49.475 -112.035 ;
        RECT -49.805 -113.725 -49.475 -113.395 ;
        RECT -49.805 -115.085 -49.475 -114.755 ;
        RECT -49.805 -116.445 -49.475 -116.115 ;
        RECT -49.805 -117.805 -49.475 -117.475 ;
        RECT -49.805 -119.165 -49.475 -118.835 ;
        RECT -49.805 -120.525 -49.475 -120.195 ;
        RECT -49.805 -121.885 -49.475 -121.555 ;
        RECT -49.805 -128.685 -49.475 -128.355 ;
        RECT -49.805 -130.045 -49.475 -129.715 ;
        RECT -49.805 -132.765 -49.475 -132.435 ;
        RECT -49.805 -134.125 -49.475 -133.795 ;
        RECT -49.805 -135.485 -49.475 -135.155 ;
        RECT -49.805 -136.845 -49.475 -136.515 ;
        RECT -49.805 -138.205 -49.475 -137.875 ;
        RECT -49.805 -139.39 -49.475 -139.06 ;
        RECT -49.805 -140.925 -49.475 -140.595 ;
        RECT -49.805 -142.285 -49.475 -141.955 ;
        RECT -49.805 -145.005 -49.475 -144.675 ;
        RECT -49.805 -146.365 -49.475 -146.035 ;
        RECT -49.805 -148.03 -49.475 -147.7 ;
        RECT -49.805 -149.085 -49.475 -148.755 ;
        RECT -49.805 -150.445 -49.475 -150.115 ;
        RECT -49.805 -153.165 -49.475 -152.835 ;
        RECT -49.805 -154.525 -49.475 -154.195 ;
        RECT -49.805 -155.885 -49.475 -155.555 ;
        RECT -49.805 -157.245 -49.475 -156.915 ;
        RECT -49.805 -158.605 -49.475 -158.275 ;
        RECT -49.805 -159.965 -49.475 -159.635 ;
        RECT -49.805 -162.685 -49.475 -162.355 ;
        RECT -49.805 -164.045 -49.475 -163.715 ;
        RECT -49.805 -165.405 -49.475 -165.075 ;
        RECT -49.805 -166.765 -49.475 -166.435 ;
        RECT -49.805 -168.125 -49.475 -167.795 ;
        RECT -49.805 -169.485 -49.475 -169.155 ;
        RECT -49.805 -170.845 -49.475 -170.515 ;
        RECT -49.805 -172.205 -49.475 -171.875 ;
        RECT -49.805 -173.565 -49.475 -173.235 ;
        RECT -49.805 -174.925 -49.475 -174.595 ;
        RECT -49.805 -176.285 -49.475 -175.955 ;
        RECT -49.805 -177.645 -49.475 -177.315 ;
        RECT -49.805 -179.005 -49.475 -178.675 ;
        RECT -49.805 -180.365 -49.475 -180.035 ;
        RECT -49.805 -181.725 -49.475 -181.395 ;
        RECT -49.805 -183.085 -49.475 -182.755 ;
        RECT -49.805 -184.445 -49.475 -184.115 ;
        RECT -49.805 -185.805 -49.475 -185.475 ;
        RECT -49.805 -187.165 -49.475 -186.835 ;
        RECT -49.805 -188.525 -49.475 -188.195 ;
        RECT -49.805 -189.885 -49.475 -189.555 ;
        RECT -49.805 -191.245 -49.475 -190.915 ;
        RECT -49.805 -192.605 -49.475 -192.275 ;
        RECT -49.805 -193.965 -49.475 -193.635 ;
        RECT -49.805 -195.325 -49.475 -194.995 ;
        RECT -49.805 -196.685 -49.475 -196.355 ;
        RECT -49.805 -198.045 -49.475 -197.715 ;
        RECT -49.805 -199.405 -49.475 -199.075 ;
        RECT -49.805 -200.765 -49.475 -200.435 ;
        RECT -49.805 -202.125 -49.475 -201.795 ;
        RECT -49.805 -203.485 -49.475 -203.155 ;
        RECT -49.805 -204.845 -49.475 -204.515 ;
        RECT -49.805 -206.205 -49.475 -205.875 ;
        RECT -49.805 -207.565 -49.475 -207.235 ;
        RECT -49.805 -208.925 -49.475 -208.595 ;
        RECT -49.805 -210.285 -49.475 -209.955 ;
        RECT -49.805 -211.645 -49.475 -211.315 ;
        RECT -49.805 -213.005 -49.475 -212.675 ;
        RECT -49.805 -214.365 -49.475 -214.035 ;
        RECT -49.805 -215.725 -49.475 -215.395 ;
        RECT -49.805 -217.085 -49.475 -216.755 ;
        RECT -49.805 -218.445 -49.475 -218.115 ;
        RECT -49.805 -219.805 -49.475 -219.475 ;
        RECT -49.805 -221.165 -49.475 -220.835 ;
        RECT -49.805 -222.525 -49.475 -222.195 ;
        RECT -49.805 -223.885 -49.475 -223.555 ;
        RECT -49.805 -225.245 -49.475 -224.915 ;
        RECT -49.805 -227.965 -49.475 -227.635 ;
        RECT -49.805 -230.685 -49.475 -230.355 ;
        RECT -49.805 -232.045 -49.475 -231.715 ;
        RECT -49.805 -233.225 -49.475 -232.895 ;
        RECT -49.805 -234.765 -49.475 -234.435 ;
        RECT -49.805 -236.125 -49.475 -235.795 ;
        RECT -49.805 -237.485 -49.475 -237.155 ;
        RECT -49.805 -238.845 -49.475 -238.515 ;
        RECT -49.805 -241.09 -49.475 -239.96 ;
        RECT -49.8 -241.205 -49.48 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 244.04 -48.115 245.17 ;
        RECT -48.445 242.595 -48.115 242.925 ;
        RECT -48.445 241.235 -48.115 241.565 ;
        RECT -48.445 239.875 -48.115 240.205 ;
        RECT -48.445 238.515 -48.115 238.845 ;
        RECT -48.445 237.155 -48.115 237.485 ;
        RECT -48.445 235.795 -48.115 236.125 ;
        RECT -48.445 234.435 -48.115 234.765 ;
        RECT -48.445 233.075 -48.115 233.405 ;
        RECT -48.445 231.715 -48.115 232.045 ;
        RECT -48.445 230.355 -48.115 230.685 ;
        RECT -48.445 228.995 -48.115 229.325 ;
        RECT -48.445 227.635 -48.115 227.965 ;
        RECT -48.445 226.275 -48.115 226.605 ;
        RECT -48.445 224.915 -48.115 225.245 ;
        RECT -48.445 223.555 -48.115 223.885 ;
        RECT -48.445 222.195 -48.115 222.525 ;
        RECT -48.445 220.835 -48.115 221.165 ;
        RECT -48.445 219.475 -48.115 219.805 ;
        RECT -48.445 218.115 -48.115 218.445 ;
        RECT -48.445 216.755 -48.115 217.085 ;
        RECT -48.445 215.395 -48.115 215.725 ;
        RECT -48.445 214.035 -48.115 214.365 ;
        RECT -48.445 212.675 -48.115 213.005 ;
        RECT -48.445 211.315 -48.115 211.645 ;
        RECT -48.445 209.955 -48.115 210.285 ;
        RECT -48.445 208.595 -48.115 208.925 ;
        RECT -48.445 207.235 -48.115 207.565 ;
        RECT -48.445 205.875 -48.115 206.205 ;
        RECT -48.445 204.515 -48.115 204.845 ;
        RECT -48.445 203.155 -48.115 203.485 ;
        RECT -48.445 201.795 -48.115 202.125 ;
        RECT -48.445 200.435 -48.115 200.765 ;
        RECT -48.445 199.075 -48.115 199.405 ;
        RECT -48.445 197.715 -48.115 198.045 ;
        RECT -48.445 196.355 -48.115 196.685 ;
        RECT -48.445 194.995 -48.115 195.325 ;
        RECT -48.445 193.635 -48.115 193.965 ;
        RECT -48.445 192.275 -48.115 192.605 ;
        RECT -48.445 190.915 -48.115 191.245 ;
        RECT -48.445 189.555 -48.115 189.885 ;
        RECT -48.445 188.195 -48.115 188.525 ;
        RECT -48.445 186.835 -48.115 187.165 ;
        RECT -48.445 185.475 -48.115 185.805 ;
        RECT -48.445 184.115 -48.115 184.445 ;
        RECT -48.445 182.755 -48.115 183.085 ;
        RECT -48.445 181.395 -48.115 181.725 ;
        RECT -48.445 180.035 -48.115 180.365 ;
        RECT -48.445 178.675 -48.115 179.005 ;
        RECT -48.445 177.315 -48.115 177.645 ;
        RECT -48.445 175.955 -48.115 176.285 ;
        RECT -48.445 174.595 -48.115 174.925 ;
        RECT -48.445 173.235 -48.115 173.565 ;
        RECT -48.445 171.875 -48.115 172.205 ;
        RECT -48.445 170.515 -48.115 170.845 ;
        RECT -48.445 169.155 -48.115 169.485 ;
        RECT -48.445 167.795 -48.115 168.125 ;
        RECT -48.445 166.435 -48.115 166.765 ;
        RECT -48.445 165.075 -48.115 165.405 ;
        RECT -48.445 163.715 -48.115 164.045 ;
        RECT -48.445 162.355 -48.115 162.685 ;
        RECT -48.445 160.995 -48.115 161.325 ;
        RECT -48.445 159.635 -48.115 159.965 ;
        RECT -48.445 158.275 -48.115 158.605 ;
        RECT -48.445 156.915 -48.115 157.245 ;
        RECT -48.445 155.555 -48.115 155.885 ;
        RECT -48.445 154.195 -48.115 154.525 ;
        RECT -48.445 152.835 -48.115 153.165 ;
        RECT -48.445 151.475 -48.115 151.805 ;
        RECT -48.445 150.115 -48.115 150.445 ;
        RECT -48.445 148.755 -48.115 149.085 ;
        RECT -48.445 147.395 -48.115 147.725 ;
        RECT -48.445 146.035 -48.115 146.365 ;
        RECT -48.445 144.675 -48.115 145.005 ;
        RECT -48.445 143.315 -48.115 143.645 ;
        RECT -48.445 141.955 -48.115 142.285 ;
        RECT -48.445 140.595 -48.115 140.925 ;
        RECT -48.445 139.235 -48.115 139.565 ;
        RECT -48.445 137.225 -48.115 137.555 ;
        RECT -48.445 135.175 -48.115 135.505 ;
        RECT -48.445 132.815 -48.115 133.145 ;
        RECT -48.445 131.665 -48.115 131.995 ;
        RECT -48.445 129.655 -48.115 129.985 ;
        RECT -48.445 128.505 -48.115 128.835 ;
        RECT -48.445 126.495 -48.115 126.825 ;
        RECT -48.445 125.345 -48.115 125.675 ;
        RECT -48.445 123.335 -48.115 123.665 ;
        RECT -48.445 122.185 -48.115 122.515 ;
        RECT -48.445 120.175 -48.115 120.505 ;
        RECT -48.445 119.025 -48.115 119.355 ;
        RECT -48.445 117.185 -48.115 117.515 ;
        RECT -48.445 115.865 -48.115 116.195 ;
        RECT -48.445 113.855 -48.115 114.185 ;
        RECT -48.445 112.705 -48.115 113.035 ;
        RECT -48.445 110.695 -48.115 111.025 ;
        RECT -48.445 109.545 -48.115 109.875 ;
        RECT -48.445 107.535 -48.115 107.865 ;
        RECT -48.445 106.385 -48.115 106.715 ;
        RECT -48.445 104.375 -48.115 104.705 ;
        RECT -48.445 103.225 -48.115 103.555 ;
        RECT -48.445 100.865 -48.115 101.195 ;
        RECT -48.445 98.81 -48.115 99.14 ;
        RECT -48.445 97.075 -48.115 97.405 ;
        RECT -48.445 95.715 -48.115 96.045 ;
        RECT -48.445 94.355 -48.115 94.685 ;
        RECT -48.445 92.995 -48.115 93.325 ;
        RECT -48.445 91.635 -48.115 91.965 ;
        RECT -48.445 90.275 -48.115 90.605 ;
        RECT -48.445 88.915 -48.115 89.245 ;
        RECT -48.445 87.555 -48.115 87.885 ;
        RECT -48.445 86.195 -48.115 86.525 ;
        RECT -48.445 84.835 -48.115 85.165 ;
        RECT -48.445 83.475 -48.115 83.805 ;
        RECT -48.445 82.115 -48.115 82.445 ;
        RECT -48.445 80.755 -48.115 81.085 ;
        RECT -48.445 79.395 -48.115 79.725 ;
        RECT -48.445 78.035 -48.115 78.365 ;
        RECT -48.445 76.675 -48.115 77.005 ;
        RECT -48.445 75.315 -48.115 75.645 ;
        RECT -48.445 73.955 -48.115 74.285 ;
        RECT -48.445 72.595 -48.115 72.925 ;
        RECT -48.445 71.235 -48.115 71.565 ;
        RECT -48.445 69.875 -48.115 70.205 ;
        RECT -48.445 68.515 -48.115 68.845 ;
        RECT -48.445 67.155 -48.115 67.485 ;
        RECT -48.445 65.795 -48.115 66.125 ;
        RECT -48.445 64.435 -48.115 64.765 ;
        RECT -48.445 63.075 -48.115 63.405 ;
        RECT -48.445 61.715 -48.115 62.045 ;
        RECT -48.445 60.355 -48.115 60.685 ;
        RECT -48.445 58.995 -48.115 59.325 ;
        RECT -48.445 57.635 -48.115 57.965 ;
        RECT -48.445 56.275 -48.115 56.605 ;
        RECT -48.445 54.915 -48.115 55.245 ;
        RECT -48.445 53.555 -48.115 53.885 ;
        RECT -48.445 52.195 -48.115 52.525 ;
        RECT -48.445 50.835 -48.115 51.165 ;
        RECT -48.445 49.475 -48.115 49.805 ;
        RECT -48.445 48.115 -48.115 48.445 ;
        RECT -48.445 46.755 -48.115 47.085 ;
        RECT -48.445 45.395 -48.115 45.725 ;
        RECT -48.445 44.035 -48.115 44.365 ;
        RECT -48.445 42.675 -48.115 43.005 ;
        RECT -48.445 41.315 -48.115 41.645 ;
        RECT -48.445 39.955 -48.115 40.285 ;
        RECT -48.445 38.595 -48.115 38.925 ;
        RECT -48.445 37.235 -48.115 37.565 ;
        RECT -48.445 35.875 -48.115 36.205 ;
        RECT -48.445 34.515 -48.115 34.845 ;
        RECT -48.445 33.155 -48.115 33.485 ;
        RECT -48.445 31.795 -48.115 32.125 ;
        RECT -48.445 30.435 -48.115 30.765 ;
        RECT -48.445 29.075 -48.115 29.405 ;
        RECT -48.445 27.715 -48.115 28.045 ;
        RECT -48.445 26.355 -48.115 26.685 ;
        RECT -48.445 24.995 -48.115 25.325 ;
        RECT -48.445 23.635 -48.115 23.965 ;
        RECT -48.445 22.275 -48.115 22.605 ;
        RECT -48.445 20.915 -48.115 21.245 ;
        RECT -48.445 19.555 -48.115 19.885 ;
        RECT -48.445 18.195 -48.115 18.525 ;
        RECT -48.445 16.835 -48.115 17.165 ;
        RECT -48.445 15.475 -48.115 15.805 ;
        RECT -48.445 14.115 -48.115 14.445 ;
        RECT -48.445 12.755 -48.115 13.085 ;
        RECT -48.445 11.395 -48.115 11.725 ;
        RECT -48.445 10.035 -48.115 10.365 ;
        RECT -48.445 8.675 -48.115 9.005 ;
        RECT -48.445 7.315 -48.115 7.645 ;
        RECT -48.445 5.955 -48.115 6.285 ;
        RECT -48.445 4.595 -48.115 4.925 ;
        RECT -48.445 3.235 -48.115 3.565 ;
        RECT -48.445 1.875 -48.115 2.205 ;
        RECT -48.445 0.515 -48.115 0.845 ;
        RECT -48.445 -0.845 -48.115 -0.515 ;
        RECT -48.445 -2.205 -48.115 -1.875 ;
        RECT -48.445 -3.565 -48.115 -3.235 ;
        RECT -48.445 -4.925 -48.115 -4.595 ;
        RECT -48.445 -6.285 -48.115 -5.955 ;
        RECT -48.445 -7.645 -48.115 -7.315 ;
        RECT -48.445 -9.005 -48.115 -8.675 ;
        RECT -48.445 -10.365 -48.115 -10.035 ;
        RECT -48.445 -11.725 -48.115 -11.395 ;
        RECT -48.445 -13.085 -48.115 -12.755 ;
        RECT -48.445 -14.445 -48.115 -14.115 ;
        RECT -48.445 -15.805 -48.115 -15.475 ;
        RECT -48.445 -17.165 -48.115 -16.835 ;
        RECT -48.445 -18.525 -48.115 -18.195 ;
        RECT -48.445 -19.885 -48.115 -19.555 ;
        RECT -48.445 -21.245 -48.115 -20.915 ;
        RECT -48.445 -22.605 -48.115 -22.275 ;
        RECT -48.445 -23.965 -48.115 -23.635 ;
        RECT -48.445 -25.325 -48.115 -24.995 ;
        RECT -48.445 -26.685 -48.115 -26.355 ;
        RECT -48.445 -28.045 -48.115 -27.715 ;
        RECT -48.445 -29.405 -48.115 -29.075 ;
        RECT -48.445 -32.125 -48.115 -31.795 ;
        RECT -48.445 -33.485 -48.115 -33.155 ;
        RECT -48.445 -34.88 -48.115 -34.55 ;
        RECT -48.445 -36.205 -48.115 -35.875 ;
        RECT -48.445 -38.925 -48.115 -38.595 ;
        RECT -48.445 -39.97 -48.115 -39.64 ;
        RECT -48.445 -48.445 -48.115 -48.115 ;
        RECT -48.445 -49.805 -48.115 -49.475 ;
        RECT -48.445 -51.165 -48.115 -50.835 ;
        RECT -48.445 -53.885 -48.115 -53.555 ;
        RECT -48.445 -57.965 -48.115 -57.635 ;
        RECT -48.445 -62.045 -48.115 -61.715 ;
        RECT -48.445 -63.405 -48.115 -63.075 ;
        RECT -48.445 -64.765 -48.115 -64.435 ;
        RECT -48.445 -66.125 -48.115 -65.795 ;
        RECT -48.445 -67.485 -48.115 -67.155 ;
        RECT -48.445 -68.845 -48.115 -68.515 ;
        RECT -48.445 -70.205 -48.115 -69.875 ;
        RECT -48.445 -71.565 -48.115 -71.235 ;
        RECT -48.445 -72.925 -48.115 -72.595 ;
        RECT -48.445 -74.285 -48.115 -73.955 ;
        RECT -48.445 -75.645 -48.115 -75.315 ;
        RECT -48.445 -77.005 -48.115 -76.675 ;
        RECT -48.445 -78.365 -48.115 -78.035 ;
        RECT -48.445 -79.725 -48.115 -79.395 ;
        RECT -48.445 -81.085 -48.115 -80.755 ;
        RECT -48.445 -82.445 -48.115 -82.115 ;
        RECT -48.445 -83.805 -48.115 -83.475 ;
        RECT -48.445 -85.165 -48.115 -84.835 ;
        RECT -48.445 -86.525 -48.115 -86.195 ;
        RECT -48.445 -87.885 -48.115 -87.555 ;
        RECT -48.445 -89.245 -48.115 -88.915 ;
        RECT -48.445 -90.605 -48.115 -90.275 ;
        RECT -48.445 -91.965 -48.115 -91.635 ;
        RECT -48.445 -93.325 -48.115 -92.995 ;
        RECT -48.445 -94.685 -48.115 -94.355 ;
        RECT -48.445 -96.045 -48.115 -95.715 ;
        RECT -48.445 -97.405 -48.115 -97.075 ;
        RECT -48.445 -98.765 -48.115 -98.435 ;
        RECT -48.445 -100.125 -48.115 -99.795 ;
        RECT -48.445 -101.485 -48.115 -101.155 ;
        RECT -48.445 -102.845 -48.115 -102.515 ;
        RECT -48.445 -104.205 -48.115 -103.875 ;
        RECT -48.445 -105.565 -48.115 -105.235 ;
        RECT -48.445 -106.925 -48.115 -106.595 ;
        RECT -48.445 -108.285 -48.115 -107.955 ;
        RECT -48.445 -109.645 -48.115 -109.315 ;
        RECT -48.445 -111.005 -48.115 -110.675 ;
        RECT -48.445 -112.365 -48.115 -112.035 ;
        RECT -48.445 -113.725 -48.115 -113.395 ;
        RECT -48.445 -115.085 -48.115 -114.755 ;
        RECT -48.445 -116.445 -48.115 -116.115 ;
        RECT -48.445 -117.805 -48.115 -117.475 ;
        RECT -48.445 -119.165 -48.115 -118.835 ;
        RECT -48.445 -120.525 -48.115 -120.195 ;
        RECT -48.445 -128.685 -48.115 -128.355 ;
        RECT -48.445 -130.045 -48.115 -129.715 ;
        RECT -48.445 -132.765 -48.115 -132.435 ;
        RECT -48.445 -134.125 -48.115 -133.795 ;
        RECT -48.445 -135.485 -48.115 -135.155 ;
        RECT -48.445 -136.845 -48.115 -136.515 ;
        RECT -48.445 -138.205 -48.115 -137.875 ;
        RECT -48.445 -139.39 -48.115 -139.06 ;
        RECT -48.445 -140.925 -48.115 -140.595 ;
        RECT -48.445 -142.285 -48.115 -141.955 ;
        RECT -48.445 -145.005 -48.115 -144.675 ;
        RECT -48.445 -146.365 -48.115 -146.035 ;
        RECT -48.445 -148.03 -48.115 -147.7 ;
        RECT -48.445 -149.085 -48.115 -148.755 ;
        RECT -48.44 -149.76 -48.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 -232.045 -48.115 -231.715 ;
        RECT -48.445 -233.225 -48.115 -232.895 ;
        RECT -48.445 -234.765 -48.115 -234.435 ;
        RECT -48.445 -236.125 -48.115 -235.795 ;
        RECT -48.445 -237.485 -48.115 -237.155 ;
        RECT -48.445 -238.845 -48.115 -238.515 ;
        RECT -48.445 -241.09 -48.115 -239.96 ;
        RECT -48.44 -241.205 -48.12 -231.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 132.815 -46.755 133.145 ;
        RECT -47.085 131.665 -46.755 131.995 ;
        RECT -47.085 129.655 -46.755 129.985 ;
        RECT -47.085 128.505 -46.755 128.835 ;
        RECT -47.085 126.495 -46.755 126.825 ;
        RECT -47.085 125.345 -46.755 125.675 ;
        RECT -47.085 123.335 -46.755 123.665 ;
        RECT -47.085 122.185 -46.755 122.515 ;
        RECT -47.085 120.175 -46.755 120.505 ;
        RECT -47.085 119.025 -46.755 119.355 ;
        RECT -47.085 117.185 -46.755 117.515 ;
        RECT -47.085 115.865 -46.755 116.195 ;
        RECT -47.085 113.855 -46.755 114.185 ;
        RECT -47.085 112.705 -46.755 113.035 ;
        RECT -47.085 110.695 -46.755 111.025 ;
        RECT -47.085 109.545 -46.755 109.875 ;
        RECT -47.085 107.535 -46.755 107.865 ;
        RECT -47.085 106.385 -46.755 106.715 ;
        RECT -47.085 104.375 -46.755 104.705 ;
        RECT -47.085 103.225 -46.755 103.555 ;
        RECT -47.085 100.865 -46.755 101.195 ;
        RECT -47.085 98.81 -46.755 99.14 ;
        RECT -47.085 97.075 -46.755 97.405 ;
        RECT -47.085 95.715 -46.755 96.045 ;
        RECT -47.085 94.355 -46.755 94.685 ;
        RECT -47.085 92.995 -46.755 93.325 ;
        RECT -47.085 91.635 -46.755 91.965 ;
        RECT -47.085 90.275 -46.755 90.605 ;
        RECT -47.085 88.915 -46.755 89.245 ;
        RECT -47.085 87.555 -46.755 87.885 ;
        RECT -47.085 86.195 -46.755 86.525 ;
        RECT -47.085 84.835 -46.755 85.165 ;
        RECT -47.085 83.475 -46.755 83.805 ;
        RECT -47.085 82.115 -46.755 82.445 ;
        RECT -47.085 80.755 -46.755 81.085 ;
        RECT -47.085 79.395 -46.755 79.725 ;
        RECT -47.085 78.035 -46.755 78.365 ;
        RECT -47.085 76.675 -46.755 77.005 ;
        RECT -47.085 75.315 -46.755 75.645 ;
        RECT -47.085 73.955 -46.755 74.285 ;
        RECT -47.085 72.595 -46.755 72.925 ;
        RECT -47.085 71.235 -46.755 71.565 ;
        RECT -47.085 69.875 -46.755 70.205 ;
        RECT -47.085 68.515 -46.755 68.845 ;
        RECT -47.085 67.155 -46.755 67.485 ;
        RECT -47.085 65.795 -46.755 66.125 ;
        RECT -47.085 64.435 -46.755 64.765 ;
        RECT -47.085 63.075 -46.755 63.405 ;
        RECT -47.085 61.715 -46.755 62.045 ;
        RECT -47.085 60.355 -46.755 60.685 ;
        RECT -47.085 58.995 -46.755 59.325 ;
        RECT -47.085 57.635 -46.755 57.965 ;
        RECT -47.085 56.275 -46.755 56.605 ;
        RECT -47.085 54.915 -46.755 55.245 ;
        RECT -47.085 53.555 -46.755 53.885 ;
        RECT -47.085 52.195 -46.755 52.525 ;
        RECT -47.085 50.835 -46.755 51.165 ;
        RECT -47.085 49.475 -46.755 49.805 ;
        RECT -47.085 48.115 -46.755 48.445 ;
        RECT -47.085 46.755 -46.755 47.085 ;
        RECT -47.085 45.395 -46.755 45.725 ;
        RECT -47.085 44.035 -46.755 44.365 ;
        RECT -47.085 42.675 -46.755 43.005 ;
        RECT -47.085 41.315 -46.755 41.645 ;
        RECT -47.085 39.955 -46.755 40.285 ;
        RECT -47.085 38.595 -46.755 38.925 ;
        RECT -47.085 37.235 -46.755 37.565 ;
        RECT -47.085 35.875 -46.755 36.205 ;
        RECT -47.085 34.515 -46.755 34.845 ;
        RECT -47.085 33.155 -46.755 33.485 ;
        RECT -47.085 31.795 -46.755 32.125 ;
        RECT -47.085 30.435 -46.755 30.765 ;
        RECT -47.085 29.075 -46.755 29.405 ;
        RECT -47.085 27.715 -46.755 28.045 ;
        RECT -47.085 26.355 -46.755 26.685 ;
        RECT -47.085 24.995 -46.755 25.325 ;
        RECT -47.085 23.635 -46.755 23.965 ;
        RECT -47.085 22.275 -46.755 22.605 ;
        RECT -47.085 20.915 -46.755 21.245 ;
        RECT -47.085 19.555 -46.755 19.885 ;
        RECT -47.085 18.195 -46.755 18.525 ;
        RECT -47.085 16.835 -46.755 17.165 ;
        RECT -47.085 15.475 -46.755 15.805 ;
        RECT -47.085 14.115 -46.755 14.445 ;
        RECT -47.085 12.755 -46.755 13.085 ;
        RECT -47.085 11.395 -46.755 11.725 ;
        RECT -47.085 10.035 -46.755 10.365 ;
        RECT -47.085 8.675 -46.755 9.005 ;
        RECT -47.085 7.315 -46.755 7.645 ;
        RECT -47.085 5.955 -46.755 6.285 ;
        RECT -47.085 4.595 -46.755 4.925 ;
        RECT -47.085 3.235 -46.755 3.565 ;
        RECT -47.085 1.875 -46.755 2.205 ;
        RECT -47.085 0.515 -46.755 0.845 ;
        RECT -47.085 -0.845 -46.755 -0.515 ;
        RECT -47.08 -1.52 -46.76 245.285 ;
        RECT -47.085 244.04 -46.755 245.17 ;
        RECT -47.085 242.595 -46.755 242.925 ;
        RECT -47.085 241.235 -46.755 241.565 ;
        RECT -47.085 239.875 -46.755 240.205 ;
        RECT -47.085 238.515 -46.755 238.845 ;
        RECT -47.085 237.155 -46.755 237.485 ;
        RECT -47.085 235.795 -46.755 236.125 ;
        RECT -47.085 234.435 -46.755 234.765 ;
        RECT -47.085 233.075 -46.755 233.405 ;
        RECT -47.085 231.715 -46.755 232.045 ;
        RECT -47.085 230.355 -46.755 230.685 ;
        RECT -47.085 228.995 -46.755 229.325 ;
        RECT -47.085 227.635 -46.755 227.965 ;
        RECT -47.085 226.275 -46.755 226.605 ;
        RECT -47.085 224.915 -46.755 225.245 ;
        RECT -47.085 223.555 -46.755 223.885 ;
        RECT -47.085 222.195 -46.755 222.525 ;
        RECT -47.085 220.835 -46.755 221.165 ;
        RECT -47.085 219.475 -46.755 219.805 ;
        RECT -47.085 218.115 -46.755 218.445 ;
        RECT -47.085 216.755 -46.755 217.085 ;
        RECT -47.085 215.395 -46.755 215.725 ;
        RECT -47.085 214.035 -46.755 214.365 ;
        RECT -47.085 212.675 -46.755 213.005 ;
        RECT -47.085 211.315 -46.755 211.645 ;
        RECT -47.085 209.955 -46.755 210.285 ;
        RECT -47.085 208.595 -46.755 208.925 ;
        RECT -47.085 207.235 -46.755 207.565 ;
        RECT -47.085 205.875 -46.755 206.205 ;
        RECT -47.085 204.515 -46.755 204.845 ;
        RECT -47.085 203.155 -46.755 203.485 ;
        RECT -47.085 201.795 -46.755 202.125 ;
        RECT -47.085 200.435 -46.755 200.765 ;
        RECT -47.085 199.075 -46.755 199.405 ;
        RECT -47.085 197.715 -46.755 198.045 ;
        RECT -47.085 196.355 -46.755 196.685 ;
        RECT -47.085 194.995 -46.755 195.325 ;
        RECT -47.085 193.635 -46.755 193.965 ;
        RECT -47.085 192.275 -46.755 192.605 ;
        RECT -47.085 190.915 -46.755 191.245 ;
        RECT -47.085 189.555 -46.755 189.885 ;
        RECT -47.085 188.195 -46.755 188.525 ;
        RECT -47.085 186.835 -46.755 187.165 ;
        RECT -47.085 185.475 -46.755 185.805 ;
        RECT -47.085 184.115 -46.755 184.445 ;
        RECT -47.085 182.755 -46.755 183.085 ;
        RECT -47.085 181.395 -46.755 181.725 ;
        RECT -47.085 180.035 -46.755 180.365 ;
        RECT -47.085 178.675 -46.755 179.005 ;
        RECT -47.085 177.315 -46.755 177.645 ;
        RECT -47.085 175.955 -46.755 176.285 ;
        RECT -47.085 174.595 -46.755 174.925 ;
        RECT -47.085 173.235 -46.755 173.565 ;
        RECT -47.085 171.875 -46.755 172.205 ;
        RECT -47.085 170.515 -46.755 170.845 ;
        RECT -47.085 169.155 -46.755 169.485 ;
        RECT -47.085 167.795 -46.755 168.125 ;
        RECT -47.085 166.435 -46.755 166.765 ;
        RECT -47.085 165.075 -46.755 165.405 ;
        RECT -47.085 163.715 -46.755 164.045 ;
        RECT -47.085 162.355 -46.755 162.685 ;
        RECT -47.085 160.995 -46.755 161.325 ;
        RECT -47.085 159.635 -46.755 159.965 ;
        RECT -47.085 158.275 -46.755 158.605 ;
        RECT -47.085 156.915 -46.755 157.245 ;
        RECT -47.085 155.555 -46.755 155.885 ;
        RECT -47.085 154.195 -46.755 154.525 ;
        RECT -47.085 152.835 -46.755 153.165 ;
        RECT -47.085 151.475 -46.755 151.805 ;
        RECT -47.085 150.115 -46.755 150.445 ;
        RECT -47.085 148.755 -46.755 149.085 ;
        RECT -47.085 147.395 -46.755 147.725 ;
        RECT -47.085 146.035 -46.755 146.365 ;
        RECT -47.085 144.675 -46.755 145.005 ;
        RECT -47.085 143.315 -46.755 143.645 ;
        RECT -47.085 141.955 -46.755 142.285 ;
        RECT -47.085 140.595 -46.755 140.925 ;
        RECT -47.085 139.235 -46.755 139.565 ;
        RECT -47.085 137.225 -46.755 137.555 ;
        RECT -47.085 135.175 -46.755 135.505 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 -162.685 -56.275 -162.355 ;
        RECT -56.605 -164.045 -56.275 -163.715 ;
        RECT -56.605 -165.405 -56.275 -165.075 ;
        RECT -56.605 -166.765 -56.275 -166.435 ;
        RECT -56.605 -168.125 -56.275 -167.795 ;
        RECT -56.605 -169.485 -56.275 -169.155 ;
        RECT -56.605 -170.845 -56.275 -170.515 ;
        RECT -56.605 -172.205 -56.275 -171.875 ;
        RECT -56.605 -173.565 -56.275 -173.235 ;
        RECT -56.605 -174.925 -56.275 -174.595 ;
        RECT -56.605 -176.285 -56.275 -175.955 ;
        RECT -56.605 -177.645 -56.275 -177.315 ;
        RECT -56.605 -179.005 -56.275 -178.675 ;
        RECT -56.605 -180.365 -56.275 -180.035 ;
        RECT -56.605 -181.725 -56.275 -181.395 ;
        RECT -56.605 -183.085 -56.275 -182.755 ;
        RECT -56.605 -184.445 -56.275 -184.115 ;
        RECT -56.605 -185.805 -56.275 -185.475 ;
        RECT -56.605 -187.165 -56.275 -186.835 ;
        RECT -56.605 -188.525 -56.275 -188.195 ;
        RECT -56.605 -189.885 -56.275 -189.555 ;
        RECT -56.605 -191.245 -56.275 -190.915 ;
        RECT -56.605 -192.605 -56.275 -192.275 ;
        RECT -56.605 -193.965 -56.275 -193.635 ;
        RECT -56.605 -195.325 -56.275 -194.995 ;
        RECT -56.605 -196.685 -56.275 -196.355 ;
        RECT -56.605 -198.045 -56.275 -197.715 ;
        RECT -56.605 -199.405 -56.275 -199.075 ;
        RECT -56.605 -200.765 -56.275 -200.435 ;
        RECT -56.605 -202.125 -56.275 -201.795 ;
        RECT -56.605 -203.485 -56.275 -203.155 ;
        RECT -56.605 -204.845 -56.275 -204.515 ;
        RECT -56.605 -206.205 -56.275 -205.875 ;
        RECT -56.605 -207.565 -56.275 -207.235 ;
        RECT -56.605 -208.925 -56.275 -208.595 ;
        RECT -56.605 -210.285 -56.275 -209.955 ;
        RECT -56.605 -211.645 -56.275 -211.315 ;
        RECT -56.605 -213.005 -56.275 -212.675 ;
        RECT -56.605 -214.365 -56.275 -214.035 ;
        RECT -56.605 -215.725 -56.275 -215.395 ;
        RECT -56.605 -217.085 -56.275 -216.755 ;
        RECT -56.605 -218.445 -56.275 -218.115 ;
        RECT -56.605 -219.805 -56.275 -219.475 ;
        RECT -56.605 -221.165 -56.275 -220.835 ;
        RECT -56.605 -222.525 -56.275 -222.195 ;
        RECT -56.605 -223.885 -56.275 -223.555 ;
        RECT -56.605 -225.245 -56.275 -224.915 ;
        RECT -56.605 -227.965 -56.275 -227.635 ;
        RECT -56.605 -230.685 -56.275 -230.355 ;
        RECT -56.605 -232.045 -56.275 -231.715 ;
        RECT -56.605 -233.225 -56.275 -232.895 ;
        RECT -56.605 -234.765 -56.275 -234.435 ;
        RECT -56.605 -236.125 -56.275 -235.795 ;
        RECT -56.605 -237.485 -56.275 -237.155 ;
        RECT -56.605 -238.845 -56.275 -238.515 ;
        RECT -56.605 -241.09 -56.275 -239.96 ;
        RECT -56.6 -241.205 -56.28 -161.68 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 244.04 -54.915 245.17 ;
        RECT -55.245 242.595 -54.915 242.925 ;
        RECT -55.245 241.235 -54.915 241.565 ;
        RECT -55.245 239.875 -54.915 240.205 ;
        RECT -55.245 238.515 -54.915 238.845 ;
        RECT -55.245 237.155 -54.915 237.485 ;
        RECT -55.245 235.795 -54.915 236.125 ;
        RECT -55.245 234.435 -54.915 234.765 ;
        RECT -55.245 233.075 -54.915 233.405 ;
        RECT -55.245 231.715 -54.915 232.045 ;
        RECT -55.245 230.355 -54.915 230.685 ;
        RECT -55.245 228.995 -54.915 229.325 ;
        RECT -55.245 227.635 -54.915 227.965 ;
        RECT -55.245 226.275 -54.915 226.605 ;
        RECT -55.245 224.915 -54.915 225.245 ;
        RECT -55.245 223.555 -54.915 223.885 ;
        RECT -55.245 222.195 -54.915 222.525 ;
        RECT -55.245 220.835 -54.915 221.165 ;
        RECT -55.245 219.475 -54.915 219.805 ;
        RECT -55.245 218.115 -54.915 218.445 ;
        RECT -55.245 216.755 -54.915 217.085 ;
        RECT -55.245 215.395 -54.915 215.725 ;
        RECT -55.245 214.035 -54.915 214.365 ;
        RECT -55.245 212.675 -54.915 213.005 ;
        RECT -55.245 211.315 -54.915 211.645 ;
        RECT -55.245 209.955 -54.915 210.285 ;
        RECT -55.245 208.595 -54.915 208.925 ;
        RECT -55.245 207.235 -54.915 207.565 ;
        RECT -55.245 205.875 -54.915 206.205 ;
        RECT -55.245 204.515 -54.915 204.845 ;
        RECT -55.245 203.155 -54.915 203.485 ;
        RECT -55.245 201.795 -54.915 202.125 ;
        RECT -55.245 200.435 -54.915 200.765 ;
        RECT -55.245 199.075 -54.915 199.405 ;
        RECT -55.245 197.715 -54.915 198.045 ;
        RECT -55.245 196.355 -54.915 196.685 ;
        RECT -55.245 194.995 -54.915 195.325 ;
        RECT -55.245 193.635 -54.915 193.965 ;
        RECT -55.245 192.275 -54.915 192.605 ;
        RECT -55.245 190.915 -54.915 191.245 ;
        RECT -55.245 189.555 -54.915 189.885 ;
        RECT -55.245 188.195 -54.915 188.525 ;
        RECT -55.245 186.835 -54.915 187.165 ;
        RECT -55.245 185.475 -54.915 185.805 ;
        RECT -55.245 184.115 -54.915 184.445 ;
        RECT -55.245 182.755 -54.915 183.085 ;
        RECT -55.245 181.395 -54.915 181.725 ;
        RECT -55.245 180.035 -54.915 180.365 ;
        RECT -55.245 178.675 -54.915 179.005 ;
        RECT -55.245 177.315 -54.915 177.645 ;
        RECT -55.245 175.955 -54.915 176.285 ;
        RECT -55.245 174.595 -54.915 174.925 ;
        RECT -55.245 173.235 -54.915 173.565 ;
        RECT -55.245 171.875 -54.915 172.205 ;
        RECT -55.245 170.515 -54.915 170.845 ;
        RECT -55.245 169.155 -54.915 169.485 ;
        RECT -55.245 167.795 -54.915 168.125 ;
        RECT -55.245 166.435 -54.915 166.765 ;
        RECT -55.245 165.075 -54.915 165.405 ;
        RECT -55.245 163.715 -54.915 164.045 ;
        RECT -55.245 162.355 -54.915 162.685 ;
        RECT -55.245 160.995 -54.915 161.325 ;
        RECT -55.245 159.635 -54.915 159.965 ;
        RECT -55.245 158.275 -54.915 158.605 ;
        RECT -55.245 156.915 -54.915 157.245 ;
        RECT -55.245 155.555 -54.915 155.885 ;
        RECT -55.245 154.195 -54.915 154.525 ;
        RECT -55.245 152.835 -54.915 153.165 ;
        RECT -55.245 151.475 -54.915 151.805 ;
        RECT -55.245 150.115 -54.915 150.445 ;
        RECT -55.245 148.755 -54.915 149.085 ;
        RECT -55.245 147.395 -54.915 147.725 ;
        RECT -55.245 146.035 -54.915 146.365 ;
        RECT -55.245 144.675 -54.915 145.005 ;
        RECT -55.245 143.315 -54.915 143.645 ;
        RECT -55.245 141.955 -54.915 142.285 ;
        RECT -55.245 140.595 -54.915 140.925 ;
        RECT -55.245 139.235 -54.915 139.565 ;
        RECT -55.24 138.56 -54.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 97.075 -54.915 97.405 ;
        RECT -55.245 95.715 -54.915 96.045 ;
        RECT -55.245 94.355 -54.915 94.685 ;
        RECT -55.245 92.995 -54.915 93.325 ;
        RECT -55.245 88.915 -54.915 89.245 ;
        RECT -55.245 84.835 -54.915 85.165 ;
        RECT -55.245 83.475 -54.915 83.805 ;
        RECT -55.245 82.115 -54.915 82.445 ;
        RECT -55.245 80.755 -54.915 81.085 ;
        RECT -55.245 79.395 -54.915 79.725 ;
        RECT -55.245 78.035 -54.915 78.365 ;
        RECT -55.245 76.675 -54.915 77.005 ;
        RECT -55.245 75.315 -54.915 75.645 ;
        RECT -55.245 73.955 -54.915 74.285 ;
        RECT -55.245 72.595 -54.915 72.925 ;
        RECT -55.245 71.235 -54.915 71.565 ;
        RECT -55.245 69.875 -54.915 70.205 ;
        RECT -55.245 68.515 -54.915 68.845 ;
        RECT -55.245 67.155 -54.915 67.485 ;
        RECT -55.245 65.795 -54.915 66.125 ;
        RECT -55.245 64.435 -54.915 64.765 ;
        RECT -55.245 63.075 -54.915 63.405 ;
        RECT -55.245 61.715 -54.915 62.045 ;
        RECT -55.245 60.355 -54.915 60.685 ;
        RECT -55.245 58.995 -54.915 59.325 ;
        RECT -55.245 57.635 -54.915 57.965 ;
        RECT -55.245 56.275 -54.915 56.605 ;
        RECT -55.245 54.915 -54.915 55.245 ;
        RECT -55.245 53.555 -54.915 53.885 ;
        RECT -55.245 52.195 -54.915 52.525 ;
        RECT -55.245 50.835 -54.915 51.165 ;
        RECT -55.245 49.475 -54.915 49.805 ;
        RECT -55.245 48.115 -54.915 48.445 ;
        RECT -55.245 46.755 -54.915 47.085 ;
        RECT -55.245 45.395 -54.915 45.725 ;
        RECT -55.245 44.035 -54.915 44.365 ;
        RECT -55.245 42.675 -54.915 43.005 ;
        RECT -55.245 41.315 -54.915 41.645 ;
        RECT -55.245 39.955 -54.915 40.285 ;
        RECT -55.245 38.595 -54.915 38.925 ;
        RECT -55.245 37.235 -54.915 37.565 ;
        RECT -55.245 35.875 -54.915 36.205 ;
        RECT -55.245 34.515 -54.915 34.845 ;
        RECT -55.245 33.155 -54.915 33.485 ;
        RECT -55.245 31.795 -54.915 32.125 ;
        RECT -55.245 30.435 -54.915 30.765 ;
        RECT -55.245 29.075 -54.915 29.405 ;
        RECT -55.245 27.715 -54.915 28.045 ;
        RECT -55.245 26.355 -54.915 26.685 ;
        RECT -55.245 24.995 -54.915 25.325 ;
        RECT -55.245 23.635 -54.915 23.965 ;
        RECT -55.245 22.275 -54.915 22.605 ;
        RECT -55.245 20.915 -54.915 21.245 ;
        RECT -55.245 19.555 -54.915 19.885 ;
        RECT -55.245 18.195 -54.915 18.525 ;
        RECT -55.245 16.835 -54.915 17.165 ;
        RECT -55.245 15.475 -54.915 15.805 ;
        RECT -55.245 14.115 -54.915 14.445 ;
        RECT -55.245 12.755 -54.915 13.085 ;
        RECT -55.245 11.395 -54.915 11.725 ;
        RECT -55.245 10.035 -54.915 10.365 ;
        RECT -55.245 8.675 -54.915 9.005 ;
        RECT -55.245 7.315 -54.915 7.645 ;
        RECT -55.245 5.955 -54.915 6.285 ;
        RECT -55.245 4.595 -54.915 4.925 ;
        RECT -55.245 3.235 -54.915 3.565 ;
        RECT -55.245 1.875 -54.915 2.205 ;
        RECT -55.245 0.515 -54.915 0.845 ;
        RECT -55.245 -0.845 -54.915 -0.515 ;
        RECT -55.245 -2.205 -54.915 -1.875 ;
        RECT -55.245 -3.565 -54.915 -3.235 ;
        RECT -55.245 -4.925 -54.915 -4.595 ;
        RECT -55.245 -6.285 -54.915 -5.955 ;
        RECT -55.245 -7.645 -54.915 -7.315 ;
        RECT -55.245 -9.005 -54.915 -8.675 ;
        RECT -55.245 -10.365 -54.915 -10.035 ;
        RECT -55.245 -11.725 -54.915 -11.395 ;
        RECT -55.245 -13.085 -54.915 -12.755 ;
        RECT -55.245 -14.445 -54.915 -14.115 ;
        RECT -55.245 -15.805 -54.915 -15.475 ;
        RECT -55.245 -17.165 -54.915 -16.835 ;
        RECT -55.245 -18.525 -54.915 -18.195 ;
        RECT -55.245 -19.885 -54.915 -19.555 ;
        RECT -55.245 -21.245 -54.915 -20.915 ;
        RECT -55.245 -22.605 -54.915 -22.275 ;
        RECT -55.245 -23.965 -54.915 -23.635 ;
        RECT -55.245 -25.325 -54.915 -24.995 ;
        RECT -55.245 -26.685 -54.915 -26.355 ;
        RECT -55.245 -28.045 -54.915 -27.715 ;
        RECT -55.245 -29.405 -54.915 -29.075 ;
        RECT -55.245 -30.765 -54.915 -30.435 ;
        RECT -55.245 -32.125 -54.915 -31.795 ;
        RECT -55.245 -33.485 -54.915 -33.155 ;
        RECT -55.245 -34.845 -54.915 -34.515 ;
        RECT -55.245 -36.205 -54.915 -35.875 ;
        RECT -55.245 -37.565 -54.915 -37.235 ;
        RECT -55.245 -38.925 -54.915 -38.595 ;
        RECT -55.245 -40.285 -54.915 -39.955 ;
        RECT -55.245 -41.645 -54.915 -41.315 ;
        RECT -55.245 -43.005 -54.915 -42.675 ;
        RECT -55.245 -44.365 -54.915 -44.035 ;
        RECT -55.245 -45.725 -54.915 -45.395 ;
        RECT -55.245 -47.085 -54.915 -46.755 ;
        RECT -55.245 -48.445 -54.915 -48.115 ;
        RECT -55.245 -49.805 -54.915 -49.475 ;
        RECT -55.245 -51.165 -54.915 -50.835 ;
        RECT -55.245 -52.525 -54.915 -52.195 ;
        RECT -55.245 -53.885 -54.915 -53.555 ;
        RECT -55.245 -55.245 -54.915 -54.915 ;
        RECT -55.245 -56.605 -54.915 -56.275 ;
        RECT -55.245 -57.965 -54.915 -57.635 ;
        RECT -55.245 -59.325 -54.915 -58.995 ;
        RECT -55.245 -60.685 -54.915 -60.355 ;
        RECT -55.245 -62.045 -54.915 -61.715 ;
        RECT -55.245 -63.405 -54.915 -63.075 ;
        RECT -55.245 -64.765 -54.915 -64.435 ;
        RECT -55.245 -66.125 -54.915 -65.795 ;
        RECT -55.245 -67.485 -54.915 -67.155 ;
        RECT -55.245 -68.845 -54.915 -68.515 ;
        RECT -55.245 -70.205 -54.915 -69.875 ;
        RECT -55.245 -71.565 -54.915 -71.235 ;
        RECT -55.245 -72.925 -54.915 -72.595 ;
        RECT -55.245 -74.285 -54.915 -73.955 ;
        RECT -55.245 -75.645 -54.915 -75.315 ;
        RECT -55.245 -77.005 -54.915 -76.675 ;
        RECT -55.245 -78.365 -54.915 -78.035 ;
        RECT -55.245 -79.725 -54.915 -79.395 ;
        RECT -55.245 -81.085 -54.915 -80.755 ;
        RECT -55.245 -82.445 -54.915 -82.115 ;
        RECT -55.245 -83.805 -54.915 -83.475 ;
        RECT -55.245 -85.165 -54.915 -84.835 ;
        RECT -55.245 -86.525 -54.915 -86.195 ;
        RECT -55.245 -87.885 -54.915 -87.555 ;
        RECT -55.245 -89.245 -54.915 -88.915 ;
        RECT -55.245 -90.605 -54.915 -90.275 ;
        RECT -55.245 -91.965 -54.915 -91.635 ;
        RECT -55.245 -93.325 -54.915 -92.995 ;
        RECT -55.245 -94.685 -54.915 -94.355 ;
        RECT -55.245 -96.045 -54.915 -95.715 ;
        RECT -55.245 -97.405 -54.915 -97.075 ;
        RECT -55.245 -98.765 -54.915 -98.435 ;
        RECT -55.245 -100.125 -54.915 -99.795 ;
        RECT -55.245 -101.485 -54.915 -101.155 ;
        RECT -55.245 -102.845 -54.915 -102.515 ;
        RECT -55.245 -104.205 -54.915 -103.875 ;
        RECT -55.245 -105.565 -54.915 -105.235 ;
        RECT -55.245 -106.925 -54.915 -106.595 ;
        RECT -55.245 -108.285 -54.915 -107.955 ;
        RECT -55.245 -109.645 -54.915 -109.315 ;
        RECT -55.245 -111.005 -54.915 -110.675 ;
        RECT -55.245 -112.365 -54.915 -112.035 ;
        RECT -55.245 -113.725 -54.915 -113.395 ;
        RECT -55.245 -115.085 -54.915 -114.755 ;
        RECT -55.245 -116.445 -54.915 -116.115 ;
        RECT -55.245 -117.805 -54.915 -117.475 ;
        RECT -55.245 -119.165 -54.915 -118.835 ;
        RECT -55.245 -120.525 -54.915 -120.195 ;
        RECT -55.245 -121.885 -54.915 -121.555 ;
        RECT -55.245 -124.605 -54.915 -124.275 ;
        RECT -55.245 -128.685 -54.915 -128.355 ;
        RECT -55.245 -130.045 -54.915 -129.715 ;
        RECT -55.245 -132.765 -54.915 -132.435 ;
        RECT -55.245 -134.125 -54.915 -133.795 ;
        RECT -55.245 -135.485 -54.915 -135.155 ;
        RECT -55.245 -136.845 -54.915 -136.515 ;
        RECT -55.245 -138.205 -54.915 -137.875 ;
        RECT -55.245 -139.39 -54.915 -139.06 ;
        RECT -55.245 -140.925 -54.915 -140.595 ;
        RECT -55.245 -142.285 -54.915 -141.955 ;
        RECT -55.245 -145.005 -54.915 -144.675 ;
        RECT -55.245 -146.365 -54.915 -146.035 ;
        RECT -55.245 -148.03 -54.915 -147.7 ;
        RECT -55.245 -149.085 -54.915 -148.755 ;
        RECT -55.245 -150.445 -54.915 -150.115 ;
        RECT -55.245 -153.165 -54.915 -152.835 ;
        RECT -55.245 -154.525 -54.915 -154.195 ;
        RECT -55.245 -155.885 -54.915 -155.555 ;
        RECT -55.245 -157.245 -54.915 -156.915 ;
        RECT -55.245 -158.605 -54.915 -158.275 ;
        RECT -55.245 -159.965 -54.915 -159.635 ;
        RECT -55.245 -162.685 -54.915 -162.355 ;
        RECT -55.245 -164.045 -54.915 -163.715 ;
        RECT -55.245 -165.405 -54.915 -165.075 ;
        RECT -55.245 -166.765 -54.915 -166.435 ;
        RECT -55.245 -168.125 -54.915 -167.795 ;
        RECT -55.245 -169.485 -54.915 -169.155 ;
        RECT -55.245 -170.845 -54.915 -170.515 ;
        RECT -55.245 -172.205 -54.915 -171.875 ;
        RECT -55.245 -173.565 -54.915 -173.235 ;
        RECT -55.245 -174.925 -54.915 -174.595 ;
        RECT -55.245 -176.285 -54.915 -175.955 ;
        RECT -55.245 -177.645 -54.915 -177.315 ;
        RECT -55.245 -179.005 -54.915 -178.675 ;
        RECT -55.245 -180.365 -54.915 -180.035 ;
        RECT -55.245 -181.725 -54.915 -181.395 ;
        RECT -55.245 -183.085 -54.915 -182.755 ;
        RECT -55.245 -184.445 -54.915 -184.115 ;
        RECT -55.245 -185.805 -54.915 -185.475 ;
        RECT -55.245 -187.165 -54.915 -186.835 ;
        RECT -55.245 -188.525 -54.915 -188.195 ;
        RECT -55.245 -189.885 -54.915 -189.555 ;
        RECT -55.245 -191.245 -54.915 -190.915 ;
        RECT -55.245 -192.605 -54.915 -192.275 ;
        RECT -55.245 -193.965 -54.915 -193.635 ;
        RECT -55.245 -195.325 -54.915 -194.995 ;
        RECT -55.245 -196.685 -54.915 -196.355 ;
        RECT -55.245 -198.045 -54.915 -197.715 ;
        RECT -55.245 -199.405 -54.915 -199.075 ;
        RECT -55.245 -200.765 -54.915 -200.435 ;
        RECT -55.245 -202.125 -54.915 -201.795 ;
        RECT -55.245 -203.485 -54.915 -203.155 ;
        RECT -55.245 -204.845 -54.915 -204.515 ;
        RECT -55.245 -206.205 -54.915 -205.875 ;
        RECT -55.245 -207.565 -54.915 -207.235 ;
        RECT -55.245 -208.925 -54.915 -208.595 ;
        RECT -55.245 -210.285 -54.915 -209.955 ;
        RECT -55.245 -211.645 -54.915 -211.315 ;
        RECT -55.245 -213.005 -54.915 -212.675 ;
        RECT -55.245 -214.365 -54.915 -214.035 ;
        RECT -55.245 -215.725 -54.915 -215.395 ;
        RECT -55.245 -217.085 -54.915 -216.755 ;
        RECT -55.245 -218.445 -54.915 -218.115 ;
        RECT -55.245 -219.805 -54.915 -219.475 ;
        RECT -55.245 -221.165 -54.915 -220.835 ;
        RECT -55.245 -222.525 -54.915 -222.195 ;
        RECT -55.245 -223.885 -54.915 -223.555 ;
        RECT -55.245 -225.245 -54.915 -224.915 ;
        RECT -55.245 -227.965 -54.915 -227.635 ;
        RECT -55.245 -232.045 -54.915 -231.715 ;
        RECT -55.245 -233.225 -54.915 -232.895 ;
        RECT -55.245 -234.765 -54.915 -234.435 ;
        RECT -55.245 -236.125 -54.915 -235.795 ;
        RECT -55.245 -237.485 -54.915 -237.155 ;
        RECT -55.245 -238.845 -54.915 -238.515 ;
        RECT -55.245 -241.09 -54.915 -239.96 ;
        RECT -55.24 -241.205 -54.92 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 244.04 -53.555 245.17 ;
        RECT -53.885 242.595 -53.555 242.925 ;
        RECT -53.885 241.235 -53.555 241.565 ;
        RECT -53.885 239.875 -53.555 240.205 ;
        RECT -53.885 238.515 -53.555 238.845 ;
        RECT -53.885 237.155 -53.555 237.485 ;
        RECT -53.885 235.795 -53.555 236.125 ;
        RECT -53.885 234.435 -53.555 234.765 ;
        RECT -53.885 233.075 -53.555 233.405 ;
        RECT -53.885 231.715 -53.555 232.045 ;
        RECT -53.885 230.355 -53.555 230.685 ;
        RECT -53.885 228.995 -53.555 229.325 ;
        RECT -53.885 227.635 -53.555 227.965 ;
        RECT -53.885 226.275 -53.555 226.605 ;
        RECT -53.885 224.915 -53.555 225.245 ;
        RECT -53.885 223.555 -53.555 223.885 ;
        RECT -53.885 222.195 -53.555 222.525 ;
        RECT -53.885 220.835 -53.555 221.165 ;
        RECT -53.885 219.475 -53.555 219.805 ;
        RECT -53.885 218.115 -53.555 218.445 ;
        RECT -53.885 216.755 -53.555 217.085 ;
        RECT -53.885 215.395 -53.555 215.725 ;
        RECT -53.885 214.035 -53.555 214.365 ;
        RECT -53.885 212.675 -53.555 213.005 ;
        RECT -53.885 211.315 -53.555 211.645 ;
        RECT -53.885 209.955 -53.555 210.285 ;
        RECT -53.885 208.595 -53.555 208.925 ;
        RECT -53.885 207.235 -53.555 207.565 ;
        RECT -53.885 205.875 -53.555 206.205 ;
        RECT -53.885 204.515 -53.555 204.845 ;
        RECT -53.885 203.155 -53.555 203.485 ;
        RECT -53.885 201.795 -53.555 202.125 ;
        RECT -53.885 200.435 -53.555 200.765 ;
        RECT -53.885 199.075 -53.555 199.405 ;
        RECT -53.885 197.715 -53.555 198.045 ;
        RECT -53.885 196.355 -53.555 196.685 ;
        RECT -53.885 194.995 -53.555 195.325 ;
        RECT -53.885 193.635 -53.555 193.965 ;
        RECT -53.885 192.275 -53.555 192.605 ;
        RECT -53.885 190.915 -53.555 191.245 ;
        RECT -53.885 189.555 -53.555 189.885 ;
        RECT -53.885 188.195 -53.555 188.525 ;
        RECT -53.885 186.835 -53.555 187.165 ;
        RECT -53.885 185.475 -53.555 185.805 ;
        RECT -53.885 184.115 -53.555 184.445 ;
        RECT -53.885 182.755 -53.555 183.085 ;
        RECT -53.885 181.395 -53.555 181.725 ;
        RECT -53.885 180.035 -53.555 180.365 ;
        RECT -53.885 178.675 -53.555 179.005 ;
        RECT -53.885 177.315 -53.555 177.645 ;
        RECT -53.885 175.955 -53.555 176.285 ;
        RECT -53.885 174.595 -53.555 174.925 ;
        RECT -53.885 173.235 -53.555 173.565 ;
        RECT -53.885 171.875 -53.555 172.205 ;
        RECT -53.885 170.515 -53.555 170.845 ;
        RECT -53.885 169.155 -53.555 169.485 ;
        RECT -53.885 167.795 -53.555 168.125 ;
        RECT -53.885 166.435 -53.555 166.765 ;
        RECT -53.885 165.075 -53.555 165.405 ;
        RECT -53.885 163.715 -53.555 164.045 ;
        RECT -53.885 162.355 -53.555 162.685 ;
        RECT -53.885 160.995 -53.555 161.325 ;
        RECT -53.885 159.635 -53.555 159.965 ;
        RECT -53.885 158.275 -53.555 158.605 ;
        RECT -53.885 156.915 -53.555 157.245 ;
        RECT -53.885 155.555 -53.555 155.885 ;
        RECT -53.885 154.195 -53.555 154.525 ;
        RECT -53.885 152.835 -53.555 153.165 ;
        RECT -53.885 151.475 -53.555 151.805 ;
        RECT -53.885 150.115 -53.555 150.445 ;
        RECT -53.885 148.755 -53.555 149.085 ;
        RECT -53.885 147.395 -53.555 147.725 ;
        RECT -53.885 146.035 -53.555 146.365 ;
        RECT -53.885 144.675 -53.555 145.005 ;
        RECT -53.885 143.315 -53.555 143.645 ;
        RECT -53.885 141.955 -53.555 142.285 ;
        RECT -53.885 140.595 -53.555 140.925 ;
        RECT -53.885 139.235 -53.555 139.565 ;
        RECT -53.88 138.56 -53.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 97.075 -53.555 97.405 ;
        RECT -53.885 95.715 -53.555 96.045 ;
        RECT -53.885 94.355 -53.555 94.685 ;
        RECT -53.885 92.995 -53.555 93.325 ;
        RECT -53.885 88.915 -53.555 89.245 ;
        RECT -53.885 84.835 -53.555 85.165 ;
        RECT -53.885 83.475 -53.555 83.805 ;
        RECT -53.885 82.115 -53.555 82.445 ;
        RECT -53.885 80.755 -53.555 81.085 ;
        RECT -53.885 79.395 -53.555 79.725 ;
        RECT -53.885 78.035 -53.555 78.365 ;
        RECT -53.885 76.675 -53.555 77.005 ;
        RECT -53.885 75.315 -53.555 75.645 ;
        RECT -53.885 73.955 -53.555 74.285 ;
        RECT -53.885 72.595 -53.555 72.925 ;
        RECT -53.885 71.235 -53.555 71.565 ;
        RECT -53.885 69.875 -53.555 70.205 ;
        RECT -53.885 68.515 -53.555 68.845 ;
        RECT -53.885 67.155 -53.555 67.485 ;
        RECT -53.885 65.795 -53.555 66.125 ;
        RECT -53.885 64.435 -53.555 64.765 ;
        RECT -53.885 63.075 -53.555 63.405 ;
        RECT -53.885 61.715 -53.555 62.045 ;
        RECT -53.885 60.355 -53.555 60.685 ;
        RECT -53.885 58.995 -53.555 59.325 ;
        RECT -53.885 57.635 -53.555 57.965 ;
        RECT -53.885 56.275 -53.555 56.605 ;
        RECT -53.885 54.915 -53.555 55.245 ;
        RECT -53.885 53.555 -53.555 53.885 ;
        RECT -53.885 52.195 -53.555 52.525 ;
        RECT -53.885 50.835 -53.555 51.165 ;
        RECT -53.885 49.475 -53.555 49.805 ;
        RECT -53.885 48.115 -53.555 48.445 ;
        RECT -53.885 46.755 -53.555 47.085 ;
        RECT -53.885 45.395 -53.555 45.725 ;
        RECT -53.885 44.035 -53.555 44.365 ;
        RECT -53.885 42.675 -53.555 43.005 ;
        RECT -53.885 41.315 -53.555 41.645 ;
        RECT -53.885 39.955 -53.555 40.285 ;
        RECT -53.885 38.595 -53.555 38.925 ;
        RECT -53.885 37.235 -53.555 37.565 ;
        RECT -53.885 35.875 -53.555 36.205 ;
        RECT -53.885 34.515 -53.555 34.845 ;
        RECT -53.885 33.155 -53.555 33.485 ;
        RECT -53.885 31.795 -53.555 32.125 ;
        RECT -53.885 30.435 -53.555 30.765 ;
        RECT -53.885 29.075 -53.555 29.405 ;
        RECT -53.885 27.715 -53.555 28.045 ;
        RECT -53.885 26.355 -53.555 26.685 ;
        RECT -53.885 24.995 -53.555 25.325 ;
        RECT -53.885 23.635 -53.555 23.965 ;
        RECT -53.885 22.275 -53.555 22.605 ;
        RECT -53.885 20.915 -53.555 21.245 ;
        RECT -53.885 19.555 -53.555 19.885 ;
        RECT -53.885 18.195 -53.555 18.525 ;
        RECT -53.885 16.835 -53.555 17.165 ;
        RECT -53.885 15.475 -53.555 15.805 ;
        RECT -53.885 14.115 -53.555 14.445 ;
        RECT -53.885 12.755 -53.555 13.085 ;
        RECT -53.885 11.395 -53.555 11.725 ;
        RECT -53.885 10.035 -53.555 10.365 ;
        RECT -53.885 8.675 -53.555 9.005 ;
        RECT -53.885 7.315 -53.555 7.645 ;
        RECT -53.885 5.955 -53.555 6.285 ;
        RECT -53.885 4.595 -53.555 4.925 ;
        RECT -53.885 3.235 -53.555 3.565 ;
        RECT -53.885 1.875 -53.555 2.205 ;
        RECT -53.885 0.515 -53.555 0.845 ;
        RECT -53.885 -0.845 -53.555 -0.515 ;
        RECT -53.885 -2.205 -53.555 -1.875 ;
        RECT -53.885 -3.565 -53.555 -3.235 ;
        RECT -53.885 -4.925 -53.555 -4.595 ;
        RECT -53.885 -6.285 -53.555 -5.955 ;
        RECT -53.885 -7.645 -53.555 -7.315 ;
        RECT -53.885 -9.005 -53.555 -8.675 ;
        RECT -53.885 -10.365 -53.555 -10.035 ;
        RECT -53.885 -11.725 -53.555 -11.395 ;
        RECT -53.885 -13.085 -53.555 -12.755 ;
        RECT -53.885 -14.445 -53.555 -14.115 ;
        RECT -53.885 -15.805 -53.555 -15.475 ;
        RECT -53.885 -17.165 -53.555 -16.835 ;
        RECT -53.885 -18.525 -53.555 -18.195 ;
        RECT -53.885 -19.885 -53.555 -19.555 ;
        RECT -53.885 -21.245 -53.555 -20.915 ;
        RECT -53.885 -22.605 -53.555 -22.275 ;
        RECT -53.885 -23.965 -53.555 -23.635 ;
        RECT -53.885 -25.325 -53.555 -24.995 ;
        RECT -53.885 -26.685 -53.555 -26.355 ;
        RECT -53.885 -28.045 -53.555 -27.715 ;
        RECT -53.885 -29.405 -53.555 -29.075 ;
        RECT -53.885 -30.765 -53.555 -30.435 ;
        RECT -53.885 -32.125 -53.555 -31.795 ;
        RECT -53.885 -33.485 -53.555 -33.155 ;
        RECT -53.885 -34.845 -53.555 -34.515 ;
        RECT -53.885 -36.205 -53.555 -35.875 ;
        RECT -53.885 -37.565 -53.555 -37.235 ;
        RECT -53.885 -38.925 -53.555 -38.595 ;
        RECT -53.885 -40.285 -53.555 -39.955 ;
        RECT -53.885 -41.645 -53.555 -41.315 ;
        RECT -53.885 -43.005 -53.555 -42.675 ;
        RECT -53.885 -44.365 -53.555 -44.035 ;
        RECT -53.885 -45.725 -53.555 -45.395 ;
        RECT -53.885 -47.085 -53.555 -46.755 ;
        RECT -53.885 -48.445 -53.555 -48.115 ;
        RECT -53.885 -49.805 -53.555 -49.475 ;
        RECT -53.885 -51.165 -53.555 -50.835 ;
        RECT -53.885 -52.525 -53.555 -52.195 ;
        RECT -53.885 -53.885 -53.555 -53.555 ;
        RECT -53.885 -55.245 -53.555 -54.915 ;
        RECT -53.885 -56.605 -53.555 -56.275 ;
        RECT -53.885 -57.965 -53.555 -57.635 ;
        RECT -53.885 -59.325 -53.555 -58.995 ;
        RECT -53.885 -60.685 -53.555 -60.355 ;
        RECT -53.885 -62.045 -53.555 -61.715 ;
        RECT -53.885 -63.405 -53.555 -63.075 ;
        RECT -53.885 -64.765 -53.555 -64.435 ;
        RECT -53.885 -66.125 -53.555 -65.795 ;
        RECT -53.885 -67.485 -53.555 -67.155 ;
        RECT -53.885 -68.845 -53.555 -68.515 ;
        RECT -53.885 -70.205 -53.555 -69.875 ;
        RECT -53.885 -71.565 -53.555 -71.235 ;
        RECT -53.885 -72.925 -53.555 -72.595 ;
        RECT -53.885 -74.285 -53.555 -73.955 ;
        RECT -53.885 -75.645 -53.555 -75.315 ;
        RECT -53.885 -77.005 -53.555 -76.675 ;
        RECT -53.885 -78.365 -53.555 -78.035 ;
        RECT -53.885 -79.725 -53.555 -79.395 ;
        RECT -53.885 -81.085 -53.555 -80.755 ;
        RECT -53.885 -82.445 -53.555 -82.115 ;
        RECT -53.885 -83.805 -53.555 -83.475 ;
        RECT -53.885 -85.165 -53.555 -84.835 ;
        RECT -53.885 -86.525 -53.555 -86.195 ;
        RECT -53.885 -87.885 -53.555 -87.555 ;
        RECT -53.885 -89.245 -53.555 -88.915 ;
        RECT -53.885 -90.605 -53.555 -90.275 ;
        RECT -53.885 -91.965 -53.555 -91.635 ;
        RECT -53.885 -93.325 -53.555 -92.995 ;
        RECT -53.885 -94.685 -53.555 -94.355 ;
        RECT -53.885 -96.045 -53.555 -95.715 ;
        RECT -53.885 -97.405 -53.555 -97.075 ;
        RECT -53.885 -98.765 -53.555 -98.435 ;
        RECT -53.885 -100.125 -53.555 -99.795 ;
        RECT -53.885 -101.485 -53.555 -101.155 ;
        RECT -53.885 -102.845 -53.555 -102.515 ;
        RECT -53.885 -104.205 -53.555 -103.875 ;
        RECT -53.885 -105.565 -53.555 -105.235 ;
        RECT -53.885 -106.925 -53.555 -106.595 ;
        RECT -53.885 -108.285 -53.555 -107.955 ;
        RECT -53.885 -109.645 -53.555 -109.315 ;
        RECT -53.885 -111.005 -53.555 -110.675 ;
        RECT -53.885 -112.365 -53.555 -112.035 ;
        RECT -53.885 -113.725 -53.555 -113.395 ;
        RECT -53.885 -115.085 -53.555 -114.755 ;
        RECT -53.885 -116.445 -53.555 -116.115 ;
        RECT -53.885 -117.805 -53.555 -117.475 ;
        RECT -53.885 -119.165 -53.555 -118.835 ;
        RECT -53.885 -120.525 -53.555 -120.195 ;
        RECT -53.885 -121.885 -53.555 -121.555 ;
        RECT -53.885 -128.685 -53.555 -128.355 ;
        RECT -53.885 -130.045 -53.555 -129.715 ;
        RECT -53.885 -132.765 -53.555 -132.435 ;
        RECT -53.885 -134.125 -53.555 -133.795 ;
        RECT -53.885 -135.485 -53.555 -135.155 ;
        RECT -53.885 -136.845 -53.555 -136.515 ;
        RECT -53.885 -138.205 -53.555 -137.875 ;
        RECT -53.885 -139.39 -53.555 -139.06 ;
        RECT -53.885 -140.925 -53.555 -140.595 ;
        RECT -53.885 -142.285 -53.555 -141.955 ;
        RECT -53.885 -145.005 -53.555 -144.675 ;
        RECT -53.885 -146.365 -53.555 -146.035 ;
        RECT -53.885 -148.03 -53.555 -147.7 ;
        RECT -53.885 -149.085 -53.555 -148.755 ;
        RECT -53.885 -150.445 -53.555 -150.115 ;
        RECT -53.885 -153.165 -53.555 -152.835 ;
        RECT -53.885 -154.525 -53.555 -154.195 ;
        RECT -53.885 -155.885 -53.555 -155.555 ;
        RECT -53.885 -157.245 -53.555 -156.915 ;
        RECT -53.885 -158.605 -53.555 -158.275 ;
        RECT -53.885 -159.965 -53.555 -159.635 ;
        RECT -53.885 -162.685 -53.555 -162.355 ;
        RECT -53.885 -164.045 -53.555 -163.715 ;
        RECT -53.885 -165.405 -53.555 -165.075 ;
        RECT -53.885 -166.765 -53.555 -166.435 ;
        RECT -53.885 -168.125 -53.555 -167.795 ;
        RECT -53.885 -169.485 -53.555 -169.155 ;
        RECT -53.885 -170.845 -53.555 -170.515 ;
        RECT -53.885 -172.205 -53.555 -171.875 ;
        RECT -53.885 -173.565 -53.555 -173.235 ;
        RECT -53.885 -174.925 -53.555 -174.595 ;
        RECT -53.885 -176.285 -53.555 -175.955 ;
        RECT -53.885 -177.645 -53.555 -177.315 ;
        RECT -53.885 -179.005 -53.555 -178.675 ;
        RECT -53.885 -180.365 -53.555 -180.035 ;
        RECT -53.885 -181.725 -53.555 -181.395 ;
        RECT -53.885 -183.085 -53.555 -182.755 ;
        RECT -53.885 -184.445 -53.555 -184.115 ;
        RECT -53.885 -185.805 -53.555 -185.475 ;
        RECT -53.885 -187.165 -53.555 -186.835 ;
        RECT -53.885 -188.525 -53.555 -188.195 ;
        RECT -53.885 -189.885 -53.555 -189.555 ;
        RECT -53.885 -191.245 -53.555 -190.915 ;
        RECT -53.885 -192.605 -53.555 -192.275 ;
        RECT -53.885 -193.965 -53.555 -193.635 ;
        RECT -53.885 -195.325 -53.555 -194.995 ;
        RECT -53.885 -196.685 -53.555 -196.355 ;
        RECT -53.885 -198.045 -53.555 -197.715 ;
        RECT -53.885 -199.405 -53.555 -199.075 ;
        RECT -53.885 -200.765 -53.555 -200.435 ;
        RECT -53.885 -202.125 -53.555 -201.795 ;
        RECT -53.885 -203.485 -53.555 -203.155 ;
        RECT -53.885 -204.845 -53.555 -204.515 ;
        RECT -53.885 -206.205 -53.555 -205.875 ;
        RECT -53.885 -207.565 -53.555 -207.235 ;
        RECT -53.885 -208.925 -53.555 -208.595 ;
        RECT -53.885 -210.285 -53.555 -209.955 ;
        RECT -53.885 -211.645 -53.555 -211.315 ;
        RECT -53.885 -213.005 -53.555 -212.675 ;
        RECT -53.885 -214.365 -53.555 -214.035 ;
        RECT -53.885 -215.725 -53.555 -215.395 ;
        RECT -53.885 -217.085 -53.555 -216.755 ;
        RECT -53.885 -218.445 -53.555 -218.115 ;
        RECT -53.885 -219.805 -53.555 -219.475 ;
        RECT -53.885 -221.165 -53.555 -220.835 ;
        RECT -53.885 -222.525 -53.555 -222.195 ;
        RECT -53.885 -223.885 -53.555 -223.555 ;
        RECT -53.885 -225.245 -53.555 -224.915 ;
        RECT -53.885 -227.965 -53.555 -227.635 ;
        RECT -53.885 -232.045 -53.555 -231.715 ;
        RECT -53.885 -234.765 -53.555 -234.435 ;
        RECT -53.885 -236.125 -53.555 -235.795 ;
        RECT -53.885 -237.485 -53.555 -237.155 ;
        RECT -53.885 -238.845 -53.555 -238.515 ;
        RECT -53.885 -241.09 -53.555 -239.96 ;
        RECT -53.88 -241.205 -53.56 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 244.04 -52.195 245.17 ;
        RECT -52.525 242.595 -52.195 242.925 ;
        RECT -52.525 241.235 -52.195 241.565 ;
        RECT -52.525 239.875 -52.195 240.205 ;
        RECT -52.525 238.515 -52.195 238.845 ;
        RECT -52.525 237.155 -52.195 237.485 ;
        RECT -52.525 235.795 -52.195 236.125 ;
        RECT -52.525 234.435 -52.195 234.765 ;
        RECT -52.525 233.075 -52.195 233.405 ;
        RECT -52.525 231.715 -52.195 232.045 ;
        RECT -52.525 230.355 -52.195 230.685 ;
        RECT -52.525 228.995 -52.195 229.325 ;
        RECT -52.525 227.635 -52.195 227.965 ;
        RECT -52.525 226.275 -52.195 226.605 ;
        RECT -52.525 224.915 -52.195 225.245 ;
        RECT -52.525 223.555 -52.195 223.885 ;
        RECT -52.525 222.195 -52.195 222.525 ;
        RECT -52.525 220.835 -52.195 221.165 ;
        RECT -52.525 219.475 -52.195 219.805 ;
        RECT -52.525 218.115 -52.195 218.445 ;
        RECT -52.525 216.755 -52.195 217.085 ;
        RECT -52.525 215.395 -52.195 215.725 ;
        RECT -52.525 214.035 -52.195 214.365 ;
        RECT -52.525 212.675 -52.195 213.005 ;
        RECT -52.525 211.315 -52.195 211.645 ;
        RECT -52.525 209.955 -52.195 210.285 ;
        RECT -52.525 208.595 -52.195 208.925 ;
        RECT -52.525 207.235 -52.195 207.565 ;
        RECT -52.525 205.875 -52.195 206.205 ;
        RECT -52.525 204.515 -52.195 204.845 ;
        RECT -52.525 203.155 -52.195 203.485 ;
        RECT -52.525 201.795 -52.195 202.125 ;
        RECT -52.525 200.435 -52.195 200.765 ;
        RECT -52.525 199.075 -52.195 199.405 ;
        RECT -52.525 197.715 -52.195 198.045 ;
        RECT -52.525 196.355 -52.195 196.685 ;
        RECT -52.525 194.995 -52.195 195.325 ;
        RECT -52.525 193.635 -52.195 193.965 ;
        RECT -52.525 192.275 -52.195 192.605 ;
        RECT -52.525 190.915 -52.195 191.245 ;
        RECT -52.525 189.555 -52.195 189.885 ;
        RECT -52.525 188.195 -52.195 188.525 ;
        RECT -52.525 186.835 -52.195 187.165 ;
        RECT -52.525 185.475 -52.195 185.805 ;
        RECT -52.525 184.115 -52.195 184.445 ;
        RECT -52.525 182.755 -52.195 183.085 ;
        RECT -52.525 181.395 -52.195 181.725 ;
        RECT -52.525 180.035 -52.195 180.365 ;
        RECT -52.525 178.675 -52.195 179.005 ;
        RECT -52.525 177.315 -52.195 177.645 ;
        RECT -52.525 175.955 -52.195 176.285 ;
        RECT -52.525 174.595 -52.195 174.925 ;
        RECT -52.525 173.235 -52.195 173.565 ;
        RECT -52.525 171.875 -52.195 172.205 ;
        RECT -52.525 170.515 -52.195 170.845 ;
        RECT -52.525 169.155 -52.195 169.485 ;
        RECT -52.525 167.795 -52.195 168.125 ;
        RECT -52.525 166.435 -52.195 166.765 ;
        RECT -52.525 165.075 -52.195 165.405 ;
        RECT -52.525 163.715 -52.195 164.045 ;
        RECT -52.525 162.355 -52.195 162.685 ;
        RECT -52.525 160.995 -52.195 161.325 ;
        RECT -52.525 159.635 -52.195 159.965 ;
        RECT -52.525 158.275 -52.195 158.605 ;
        RECT -52.525 156.915 -52.195 157.245 ;
        RECT -52.525 155.555 -52.195 155.885 ;
        RECT -52.525 154.195 -52.195 154.525 ;
        RECT -52.525 152.835 -52.195 153.165 ;
        RECT -52.525 151.475 -52.195 151.805 ;
        RECT -52.525 150.115 -52.195 150.445 ;
        RECT -52.525 148.755 -52.195 149.085 ;
        RECT -52.525 147.395 -52.195 147.725 ;
        RECT -52.525 146.035 -52.195 146.365 ;
        RECT -52.525 144.675 -52.195 145.005 ;
        RECT -52.525 143.315 -52.195 143.645 ;
        RECT -52.525 141.955 -52.195 142.285 ;
        RECT -52.525 140.595 -52.195 140.925 ;
        RECT -52.525 139.235 -52.195 139.565 ;
        RECT -52.52 138.56 -52.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 72.595 -52.195 72.925 ;
        RECT -52.525 71.235 -52.195 71.565 ;
        RECT -52.525 69.875 -52.195 70.205 ;
        RECT -52.525 68.515 -52.195 68.845 ;
        RECT -52.525 67.155 -52.195 67.485 ;
        RECT -52.525 65.795 -52.195 66.125 ;
        RECT -52.525 64.435 -52.195 64.765 ;
        RECT -52.525 63.075 -52.195 63.405 ;
        RECT -52.525 61.715 -52.195 62.045 ;
        RECT -52.525 60.355 -52.195 60.685 ;
        RECT -52.525 58.995 -52.195 59.325 ;
        RECT -52.525 57.635 -52.195 57.965 ;
        RECT -52.525 56.275 -52.195 56.605 ;
        RECT -52.525 54.915 -52.195 55.245 ;
        RECT -52.525 53.555 -52.195 53.885 ;
        RECT -52.525 52.195 -52.195 52.525 ;
        RECT -52.525 50.835 -52.195 51.165 ;
        RECT -52.525 49.475 -52.195 49.805 ;
        RECT -52.525 48.115 -52.195 48.445 ;
        RECT -52.525 46.755 -52.195 47.085 ;
        RECT -52.525 45.395 -52.195 45.725 ;
        RECT -52.525 44.035 -52.195 44.365 ;
        RECT -52.525 42.675 -52.195 43.005 ;
        RECT -52.525 41.315 -52.195 41.645 ;
        RECT -52.525 39.955 -52.195 40.285 ;
        RECT -52.525 38.595 -52.195 38.925 ;
        RECT -52.525 37.235 -52.195 37.565 ;
        RECT -52.525 35.875 -52.195 36.205 ;
        RECT -52.525 34.515 -52.195 34.845 ;
        RECT -52.525 33.155 -52.195 33.485 ;
        RECT -52.525 31.795 -52.195 32.125 ;
        RECT -52.525 30.435 -52.195 30.765 ;
        RECT -52.525 29.075 -52.195 29.405 ;
        RECT -52.525 27.715 -52.195 28.045 ;
        RECT -52.525 26.355 -52.195 26.685 ;
        RECT -52.525 24.995 -52.195 25.325 ;
        RECT -52.525 23.635 -52.195 23.965 ;
        RECT -52.525 22.275 -52.195 22.605 ;
        RECT -52.525 20.915 -52.195 21.245 ;
        RECT -52.525 19.555 -52.195 19.885 ;
        RECT -52.525 18.195 -52.195 18.525 ;
        RECT -52.525 16.835 -52.195 17.165 ;
        RECT -52.525 15.475 -52.195 15.805 ;
        RECT -52.525 14.115 -52.195 14.445 ;
        RECT -52.525 12.755 -52.195 13.085 ;
        RECT -52.525 11.395 -52.195 11.725 ;
        RECT -52.525 10.035 -52.195 10.365 ;
        RECT -52.525 8.675 -52.195 9.005 ;
        RECT -52.525 7.315 -52.195 7.645 ;
        RECT -52.525 5.955 -52.195 6.285 ;
        RECT -52.525 4.595 -52.195 4.925 ;
        RECT -52.525 3.235 -52.195 3.565 ;
        RECT -52.525 1.875 -52.195 2.205 ;
        RECT -52.525 0.515 -52.195 0.845 ;
        RECT -52.525 -0.845 -52.195 -0.515 ;
        RECT -52.525 -2.205 -52.195 -1.875 ;
        RECT -52.525 -3.565 -52.195 -3.235 ;
        RECT -52.525 -4.925 -52.195 -4.595 ;
        RECT -52.525 -6.285 -52.195 -5.955 ;
        RECT -52.525 -7.645 -52.195 -7.315 ;
        RECT -52.525 -9.005 -52.195 -8.675 ;
        RECT -52.525 -10.365 -52.195 -10.035 ;
        RECT -52.525 -11.725 -52.195 -11.395 ;
        RECT -52.525 -13.085 -52.195 -12.755 ;
        RECT -52.525 -14.445 -52.195 -14.115 ;
        RECT -52.525 -15.805 -52.195 -15.475 ;
        RECT -52.525 -17.165 -52.195 -16.835 ;
        RECT -52.525 -18.525 -52.195 -18.195 ;
        RECT -52.525 -19.885 -52.195 -19.555 ;
        RECT -52.525 -21.245 -52.195 -20.915 ;
        RECT -52.525 -22.605 -52.195 -22.275 ;
        RECT -52.525 -23.965 -52.195 -23.635 ;
        RECT -52.525 -25.325 -52.195 -24.995 ;
        RECT -52.525 -26.685 -52.195 -26.355 ;
        RECT -52.525 -28.045 -52.195 -27.715 ;
        RECT -52.525 -29.405 -52.195 -29.075 ;
        RECT -52.525 -30.765 -52.195 -30.435 ;
        RECT -52.525 -32.125 -52.195 -31.795 ;
        RECT -52.525 -33.485 -52.195 -33.155 ;
        RECT -52.525 -34.845 -52.195 -34.515 ;
        RECT -52.525 -36.205 -52.195 -35.875 ;
        RECT -52.525 -37.565 -52.195 -37.235 ;
        RECT -52.525 -38.925 -52.195 -38.595 ;
        RECT -52.525 -40.285 -52.195 -39.955 ;
        RECT -52.525 -41.645 -52.195 -41.315 ;
        RECT -52.525 -43.005 -52.195 -42.675 ;
        RECT -52.525 -44.365 -52.195 -44.035 ;
        RECT -52.525 -45.725 -52.195 -45.395 ;
        RECT -52.525 -47.085 -52.195 -46.755 ;
        RECT -52.525 -48.445 -52.195 -48.115 ;
        RECT -52.525 -49.805 -52.195 -49.475 ;
        RECT -52.525 -51.165 -52.195 -50.835 ;
        RECT -52.525 -52.525 -52.195 -52.195 ;
        RECT -52.525 -53.885 -52.195 -53.555 ;
        RECT -52.525 -55.245 -52.195 -54.915 ;
        RECT -52.525 -56.605 -52.195 -56.275 ;
        RECT -52.525 -57.965 -52.195 -57.635 ;
        RECT -52.525 -59.325 -52.195 -58.995 ;
        RECT -52.525 -60.685 -52.195 -60.355 ;
        RECT -52.525 -62.045 -52.195 -61.715 ;
        RECT -52.525 -63.405 -52.195 -63.075 ;
        RECT -52.525 -64.765 -52.195 -64.435 ;
        RECT -52.525 -66.125 -52.195 -65.795 ;
        RECT -52.525 -67.485 -52.195 -67.155 ;
        RECT -52.525 -68.845 -52.195 -68.515 ;
        RECT -52.525 -70.205 -52.195 -69.875 ;
        RECT -52.525 -71.565 -52.195 -71.235 ;
        RECT -52.525 -72.925 -52.195 -72.595 ;
        RECT -52.525 -74.285 -52.195 -73.955 ;
        RECT -52.525 -75.645 -52.195 -75.315 ;
        RECT -52.525 -77.005 -52.195 -76.675 ;
        RECT -52.525 -78.365 -52.195 -78.035 ;
        RECT -52.525 -79.725 -52.195 -79.395 ;
        RECT -52.525 -81.085 -52.195 -80.755 ;
        RECT -52.525 -82.445 -52.195 -82.115 ;
        RECT -52.525 -83.805 -52.195 -83.475 ;
        RECT -52.525 -85.165 -52.195 -84.835 ;
        RECT -52.525 -86.525 -52.195 -86.195 ;
        RECT -52.525 -87.885 -52.195 -87.555 ;
        RECT -52.525 -89.245 -52.195 -88.915 ;
        RECT -52.525 -90.605 -52.195 -90.275 ;
        RECT -52.525 -91.965 -52.195 -91.635 ;
        RECT -52.525 -93.325 -52.195 -92.995 ;
        RECT -52.525 -94.685 -52.195 -94.355 ;
        RECT -52.525 -96.045 -52.195 -95.715 ;
        RECT -52.525 -97.405 -52.195 -97.075 ;
        RECT -52.525 -98.765 -52.195 -98.435 ;
        RECT -52.525 -100.125 -52.195 -99.795 ;
        RECT -52.525 -101.485 -52.195 -101.155 ;
        RECT -52.525 -102.845 -52.195 -102.515 ;
        RECT -52.525 -104.205 -52.195 -103.875 ;
        RECT -52.525 -105.565 -52.195 -105.235 ;
        RECT -52.525 -106.925 -52.195 -106.595 ;
        RECT -52.525 -108.285 -52.195 -107.955 ;
        RECT -52.525 -109.645 -52.195 -109.315 ;
        RECT -52.525 -111.005 -52.195 -110.675 ;
        RECT -52.525 -112.365 -52.195 -112.035 ;
        RECT -52.525 -113.725 -52.195 -113.395 ;
        RECT -52.525 -115.085 -52.195 -114.755 ;
        RECT -52.525 -116.445 -52.195 -116.115 ;
        RECT -52.525 -117.805 -52.195 -117.475 ;
        RECT -52.525 -119.165 -52.195 -118.835 ;
        RECT -52.525 -120.525 -52.195 -120.195 ;
        RECT -52.525 -121.885 -52.195 -121.555 ;
        RECT -52.525 -128.685 -52.195 -128.355 ;
        RECT -52.525 -130.045 -52.195 -129.715 ;
        RECT -52.525 -132.765 -52.195 -132.435 ;
        RECT -52.525 -134.125 -52.195 -133.795 ;
        RECT -52.525 -135.485 -52.195 -135.155 ;
        RECT -52.525 -136.845 -52.195 -136.515 ;
        RECT -52.525 -138.205 -52.195 -137.875 ;
        RECT -52.525 -139.39 -52.195 -139.06 ;
        RECT -52.525 -140.925 -52.195 -140.595 ;
        RECT -52.525 -142.285 -52.195 -141.955 ;
        RECT -52.525 -145.005 -52.195 -144.675 ;
        RECT -52.525 -146.365 -52.195 -146.035 ;
        RECT -52.525 -148.03 -52.195 -147.7 ;
        RECT -52.525 -149.085 -52.195 -148.755 ;
        RECT -52.525 -150.445 -52.195 -150.115 ;
        RECT -52.525 -153.165 -52.195 -152.835 ;
        RECT -52.525 -154.525 -52.195 -154.195 ;
        RECT -52.525 -155.885 -52.195 -155.555 ;
        RECT -52.525 -157.245 -52.195 -156.915 ;
        RECT -52.525 -158.605 -52.195 -158.275 ;
        RECT -52.525 -159.965 -52.195 -159.635 ;
        RECT -52.525 -162.685 -52.195 -162.355 ;
        RECT -52.525 -164.045 -52.195 -163.715 ;
        RECT -52.525 -165.405 -52.195 -165.075 ;
        RECT -52.525 -166.765 -52.195 -166.435 ;
        RECT -52.525 -168.125 -52.195 -167.795 ;
        RECT -52.525 -169.485 -52.195 -169.155 ;
        RECT -52.525 -170.845 -52.195 -170.515 ;
        RECT -52.525 -172.205 -52.195 -171.875 ;
        RECT -52.525 -173.565 -52.195 -173.235 ;
        RECT -52.525 -174.925 -52.195 -174.595 ;
        RECT -52.525 -176.285 -52.195 -175.955 ;
        RECT -52.525 -177.645 -52.195 -177.315 ;
        RECT -52.525 -179.005 -52.195 -178.675 ;
        RECT -52.525 -180.365 -52.195 -180.035 ;
        RECT -52.525 -181.725 -52.195 -181.395 ;
        RECT -52.525 -183.085 -52.195 -182.755 ;
        RECT -52.525 -184.445 -52.195 -184.115 ;
        RECT -52.525 -185.805 -52.195 -185.475 ;
        RECT -52.525 -187.165 -52.195 -186.835 ;
        RECT -52.525 -188.525 -52.195 -188.195 ;
        RECT -52.525 -189.885 -52.195 -189.555 ;
        RECT -52.525 -191.245 -52.195 -190.915 ;
        RECT -52.525 -192.605 -52.195 -192.275 ;
        RECT -52.525 -193.965 -52.195 -193.635 ;
        RECT -52.525 -195.325 -52.195 -194.995 ;
        RECT -52.525 -196.685 -52.195 -196.355 ;
        RECT -52.525 -198.045 -52.195 -197.715 ;
        RECT -52.525 -199.405 -52.195 -199.075 ;
        RECT -52.525 -200.765 -52.195 -200.435 ;
        RECT -52.525 -202.125 -52.195 -201.795 ;
        RECT -52.525 -203.485 -52.195 -203.155 ;
        RECT -52.525 -204.845 -52.195 -204.515 ;
        RECT -52.525 -206.205 -52.195 -205.875 ;
        RECT -52.525 -207.565 -52.195 -207.235 ;
        RECT -52.525 -208.925 -52.195 -208.595 ;
        RECT -52.525 -210.285 -52.195 -209.955 ;
        RECT -52.525 -211.645 -52.195 -211.315 ;
        RECT -52.525 -213.005 -52.195 -212.675 ;
        RECT -52.525 -214.365 -52.195 -214.035 ;
        RECT -52.525 -215.725 -52.195 -215.395 ;
        RECT -52.525 -217.085 -52.195 -216.755 ;
        RECT -52.525 -218.445 -52.195 -218.115 ;
        RECT -52.525 -219.805 -52.195 -219.475 ;
        RECT -52.525 -221.165 -52.195 -220.835 ;
        RECT -52.525 -222.525 -52.195 -222.195 ;
        RECT -52.525 -223.885 -52.195 -223.555 ;
        RECT -52.525 -225.245 -52.195 -224.915 ;
        RECT -52.525 -227.965 -52.195 -227.635 ;
        RECT -52.52 -229.32 -52.2 98.08 ;
        RECT -52.525 97.075 -52.195 97.405 ;
        RECT -52.525 95.715 -52.195 96.045 ;
        RECT -52.525 94.355 -52.195 94.685 ;
        RECT -52.525 92.995 -52.195 93.325 ;
        RECT -52.525 88.915 -52.195 89.245 ;
        RECT -52.525 84.835 -52.195 85.165 ;
        RECT -52.525 83.475 -52.195 83.805 ;
        RECT -52.525 82.115 -52.195 82.445 ;
        RECT -52.525 80.755 -52.195 81.085 ;
        RECT -52.525 79.395 -52.195 79.725 ;
        RECT -52.525 78.035 -52.195 78.365 ;
        RECT -52.525 76.675 -52.195 77.005 ;
        RECT -52.525 75.315 -52.195 75.645 ;
        RECT -52.525 73.955 -52.195 74.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 -232.045 -60.355 -231.715 ;
        RECT -60.685 -233.225 -60.355 -232.895 ;
        RECT -60.685 -234.765 -60.355 -234.435 ;
        RECT -60.685 -236.125 -60.355 -235.795 ;
        RECT -60.685 -237.485 -60.355 -237.155 ;
        RECT -60.685 -238.845 -60.355 -238.515 ;
        RECT -60.685 -241.09 -60.355 -239.96 ;
        RECT -60.68 -241.205 -60.36 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.325 244.04 -58.995 245.17 ;
        RECT -59.325 242.595 -58.995 242.925 ;
        RECT -59.325 241.235 -58.995 241.565 ;
        RECT -59.325 239.875 -58.995 240.205 ;
        RECT -59.325 238.515 -58.995 238.845 ;
        RECT -59.325 237.155 -58.995 237.485 ;
        RECT -59.325 235.795 -58.995 236.125 ;
        RECT -59.325 234.435 -58.995 234.765 ;
        RECT -59.325 233.075 -58.995 233.405 ;
        RECT -59.325 231.715 -58.995 232.045 ;
        RECT -59.325 230.355 -58.995 230.685 ;
        RECT -59.325 228.995 -58.995 229.325 ;
        RECT -59.325 227.635 -58.995 227.965 ;
        RECT -59.325 226.275 -58.995 226.605 ;
        RECT -59.325 224.915 -58.995 225.245 ;
        RECT -59.325 223.555 -58.995 223.885 ;
        RECT -59.325 222.195 -58.995 222.525 ;
        RECT -59.325 220.835 -58.995 221.165 ;
        RECT -59.325 219.475 -58.995 219.805 ;
        RECT -59.325 218.115 -58.995 218.445 ;
        RECT -59.325 216.755 -58.995 217.085 ;
        RECT -59.325 215.395 -58.995 215.725 ;
        RECT -59.325 214.035 -58.995 214.365 ;
        RECT -59.325 212.675 -58.995 213.005 ;
        RECT -59.325 211.315 -58.995 211.645 ;
        RECT -59.325 209.955 -58.995 210.285 ;
        RECT -59.325 208.595 -58.995 208.925 ;
        RECT -59.325 207.235 -58.995 207.565 ;
        RECT -59.325 205.875 -58.995 206.205 ;
        RECT -59.325 204.515 -58.995 204.845 ;
        RECT -59.325 203.155 -58.995 203.485 ;
        RECT -59.325 201.795 -58.995 202.125 ;
        RECT -59.325 200.435 -58.995 200.765 ;
        RECT -59.325 199.075 -58.995 199.405 ;
        RECT -59.325 197.715 -58.995 198.045 ;
        RECT -59.325 196.355 -58.995 196.685 ;
        RECT -59.325 194.995 -58.995 195.325 ;
        RECT -59.325 193.635 -58.995 193.965 ;
        RECT -59.325 192.275 -58.995 192.605 ;
        RECT -59.325 190.915 -58.995 191.245 ;
        RECT -59.325 189.555 -58.995 189.885 ;
        RECT -59.325 188.195 -58.995 188.525 ;
        RECT -59.325 186.835 -58.995 187.165 ;
        RECT -59.325 185.475 -58.995 185.805 ;
        RECT -59.325 184.115 -58.995 184.445 ;
        RECT -59.325 182.755 -58.995 183.085 ;
        RECT -59.325 181.395 -58.995 181.725 ;
        RECT -59.325 180.035 -58.995 180.365 ;
        RECT -59.325 178.675 -58.995 179.005 ;
        RECT -59.325 177.315 -58.995 177.645 ;
        RECT -59.325 175.955 -58.995 176.285 ;
        RECT -59.325 174.595 -58.995 174.925 ;
        RECT -59.325 173.235 -58.995 173.565 ;
        RECT -59.325 171.875 -58.995 172.205 ;
        RECT -59.325 170.515 -58.995 170.845 ;
        RECT -59.325 169.155 -58.995 169.485 ;
        RECT -59.325 167.795 -58.995 168.125 ;
        RECT -59.325 166.435 -58.995 166.765 ;
        RECT -59.325 165.075 -58.995 165.405 ;
        RECT -59.325 163.715 -58.995 164.045 ;
        RECT -59.325 162.355 -58.995 162.685 ;
        RECT -59.325 160.995 -58.995 161.325 ;
        RECT -59.325 159.635 -58.995 159.965 ;
        RECT -59.325 158.275 -58.995 158.605 ;
        RECT -59.325 156.915 -58.995 157.245 ;
        RECT -59.325 155.555 -58.995 155.885 ;
        RECT -59.325 154.195 -58.995 154.525 ;
        RECT -59.325 152.835 -58.995 153.165 ;
        RECT -59.325 151.475 -58.995 151.805 ;
        RECT -59.325 150.115 -58.995 150.445 ;
        RECT -59.325 148.755 -58.995 149.085 ;
        RECT -59.325 147.395 -58.995 147.725 ;
        RECT -59.325 146.035 -58.995 146.365 ;
        RECT -59.325 144.675 -58.995 145.005 ;
        RECT -59.325 143.315 -58.995 143.645 ;
        RECT -59.325 141.955 -58.995 142.285 ;
        RECT -59.325 140.595 -58.995 140.925 ;
        RECT -59.325 139.235 -58.995 139.565 ;
        RECT -59.325 137.225 -58.995 137.555 ;
        RECT -59.325 135.175 -58.995 135.505 ;
        RECT -59.325 132.815 -58.995 133.145 ;
        RECT -59.325 131.665 -58.995 131.995 ;
        RECT -59.325 129.655 -58.995 129.985 ;
        RECT -59.325 128.505 -58.995 128.835 ;
        RECT -59.325 126.495 -58.995 126.825 ;
        RECT -59.325 125.345 -58.995 125.675 ;
        RECT -59.325 123.335 -58.995 123.665 ;
        RECT -59.325 122.185 -58.995 122.515 ;
        RECT -59.325 120.175 -58.995 120.505 ;
        RECT -59.325 119.025 -58.995 119.355 ;
        RECT -59.325 117.185 -58.995 117.515 ;
        RECT -59.325 115.865 -58.995 116.195 ;
        RECT -59.325 113.855 -58.995 114.185 ;
        RECT -59.325 112.705 -58.995 113.035 ;
        RECT -59.325 110.695 -58.995 111.025 ;
        RECT -59.325 109.545 -58.995 109.875 ;
        RECT -59.325 107.535 -58.995 107.865 ;
        RECT -59.325 106.385 -58.995 106.715 ;
        RECT -59.325 104.375 -58.995 104.705 ;
        RECT -59.325 103.225 -58.995 103.555 ;
        RECT -59.325 100.865 -58.995 101.195 ;
        RECT -59.325 98.81 -58.995 99.14 ;
        RECT -59.325 97.075 -58.995 97.405 ;
        RECT -59.325 95.715 -58.995 96.045 ;
        RECT -59.325 94.355 -58.995 94.685 ;
        RECT -59.325 92.995 -58.995 93.325 ;
        RECT -59.325 91.635 -58.995 91.965 ;
        RECT -59.325 90.275 -58.995 90.605 ;
        RECT -59.325 88.915 -58.995 89.245 ;
        RECT -59.325 87.555 -58.995 87.885 ;
        RECT -59.325 86.195 -58.995 86.525 ;
        RECT -59.325 84.835 -58.995 85.165 ;
        RECT -59.325 83.475 -58.995 83.805 ;
        RECT -59.325 82.115 -58.995 82.445 ;
        RECT -59.325 80.755 -58.995 81.085 ;
        RECT -59.325 79.395 -58.995 79.725 ;
        RECT -59.325 78.035 -58.995 78.365 ;
        RECT -59.325 76.675 -58.995 77.005 ;
        RECT -59.325 75.315 -58.995 75.645 ;
        RECT -59.325 73.955 -58.995 74.285 ;
        RECT -59.325 72.595 -58.995 72.925 ;
        RECT -59.325 71.235 -58.995 71.565 ;
        RECT -59.325 69.875 -58.995 70.205 ;
        RECT -59.325 68.515 -58.995 68.845 ;
        RECT -59.325 67.155 -58.995 67.485 ;
        RECT -59.325 65.795 -58.995 66.125 ;
        RECT -59.325 64.435 -58.995 64.765 ;
        RECT -59.325 63.075 -58.995 63.405 ;
        RECT -59.325 61.715 -58.995 62.045 ;
        RECT -59.325 60.355 -58.995 60.685 ;
        RECT -59.325 58.995 -58.995 59.325 ;
        RECT -59.325 57.635 -58.995 57.965 ;
        RECT -59.325 56.275 -58.995 56.605 ;
        RECT -59.325 54.915 -58.995 55.245 ;
        RECT -59.325 53.555 -58.995 53.885 ;
        RECT -59.325 52.195 -58.995 52.525 ;
        RECT -59.325 50.835 -58.995 51.165 ;
        RECT -59.325 49.475 -58.995 49.805 ;
        RECT -59.325 48.115 -58.995 48.445 ;
        RECT -59.325 46.755 -58.995 47.085 ;
        RECT -59.325 45.395 -58.995 45.725 ;
        RECT -59.325 44.035 -58.995 44.365 ;
        RECT -59.325 42.675 -58.995 43.005 ;
        RECT -59.325 41.315 -58.995 41.645 ;
        RECT -59.325 39.955 -58.995 40.285 ;
        RECT -59.325 38.595 -58.995 38.925 ;
        RECT -59.325 37.235 -58.995 37.565 ;
        RECT -59.325 35.875 -58.995 36.205 ;
        RECT -59.325 34.515 -58.995 34.845 ;
        RECT -59.325 33.155 -58.995 33.485 ;
        RECT -59.325 31.795 -58.995 32.125 ;
        RECT -59.325 30.435 -58.995 30.765 ;
        RECT -59.325 29.075 -58.995 29.405 ;
        RECT -59.325 27.715 -58.995 28.045 ;
        RECT -59.325 26.355 -58.995 26.685 ;
        RECT -59.325 24.995 -58.995 25.325 ;
        RECT -59.325 23.635 -58.995 23.965 ;
        RECT -59.325 22.275 -58.995 22.605 ;
        RECT -59.325 20.915 -58.995 21.245 ;
        RECT -59.325 19.555 -58.995 19.885 ;
        RECT -59.325 18.195 -58.995 18.525 ;
        RECT -59.325 16.835 -58.995 17.165 ;
        RECT -59.325 15.475 -58.995 15.805 ;
        RECT -59.325 14.115 -58.995 14.445 ;
        RECT -59.325 12.755 -58.995 13.085 ;
        RECT -59.325 11.395 -58.995 11.725 ;
        RECT -59.325 10.035 -58.995 10.365 ;
        RECT -59.325 8.675 -58.995 9.005 ;
        RECT -59.325 7.315 -58.995 7.645 ;
        RECT -59.325 5.955 -58.995 6.285 ;
        RECT -59.325 4.595 -58.995 4.925 ;
        RECT -59.325 3.235 -58.995 3.565 ;
        RECT -59.325 1.875 -58.995 2.205 ;
        RECT -59.325 0.515 -58.995 0.845 ;
        RECT -59.325 -0.845 -58.995 -0.515 ;
        RECT -59.325 -2.205 -58.995 -1.875 ;
        RECT -59.325 -3.565 -58.995 -3.235 ;
        RECT -59.325 -4.925 -58.995 -4.595 ;
        RECT -59.325 -6.285 -58.995 -5.955 ;
        RECT -59.325 -7.645 -58.995 -7.315 ;
        RECT -59.325 -9.005 -58.995 -8.675 ;
        RECT -59.325 -10.365 -58.995 -10.035 ;
        RECT -59.325 -11.725 -58.995 -11.395 ;
        RECT -59.325 -13.085 -58.995 -12.755 ;
        RECT -59.325 -14.445 -58.995 -14.115 ;
        RECT -59.325 -15.805 -58.995 -15.475 ;
        RECT -59.325 -17.165 -58.995 -16.835 ;
        RECT -59.325 -18.525 -58.995 -18.195 ;
        RECT -59.325 -19.885 -58.995 -19.555 ;
        RECT -59.325 -21.245 -58.995 -20.915 ;
        RECT -59.325 -22.605 -58.995 -22.275 ;
        RECT -59.325 -23.965 -58.995 -23.635 ;
        RECT -59.325 -25.325 -58.995 -24.995 ;
        RECT -59.325 -26.685 -58.995 -26.355 ;
        RECT -59.325 -28.045 -58.995 -27.715 ;
        RECT -59.325 -29.405 -58.995 -29.075 ;
        RECT -59.325 -30.765 -58.995 -30.435 ;
        RECT -59.325 -32.125 -58.995 -31.795 ;
        RECT -59.325 -33.485 -58.995 -33.155 ;
        RECT -59.325 -34.845 -58.995 -34.515 ;
        RECT -59.325 -36.205 -58.995 -35.875 ;
        RECT -59.325 -37.565 -58.995 -37.235 ;
        RECT -59.325 -38.925 -58.995 -38.595 ;
        RECT -59.325 -40.285 -58.995 -39.955 ;
        RECT -59.325 -41.645 -58.995 -41.315 ;
        RECT -59.325 -43.005 -58.995 -42.675 ;
        RECT -59.325 -44.365 -58.995 -44.035 ;
        RECT -59.325 -45.725 -58.995 -45.395 ;
        RECT -59.325 -47.085 -58.995 -46.755 ;
        RECT -59.325 -48.445 -58.995 -48.115 ;
        RECT -59.325 -49.805 -58.995 -49.475 ;
        RECT -59.325 -51.165 -58.995 -50.835 ;
        RECT -59.325 -52.525 -58.995 -52.195 ;
        RECT -59.325 -53.885 -58.995 -53.555 ;
        RECT -59.325 -55.245 -58.995 -54.915 ;
        RECT -59.325 -56.605 -58.995 -56.275 ;
        RECT -59.325 -57.965 -58.995 -57.635 ;
        RECT -59.325 -59.325 -58.995 -58.995 ;
        RECT -59.325 -60.685 -58.995 -60.355 ;
        RECT -59.325 -62.045 -58.995 -61.715 ;
        RECT -59.325 -63.405 -58.995 -63.075 ;
        RECT -59.325 -64.765 -58.995 -64.435 ;
        RECT -59.325 -66.125 -58.995 -65.795 ;
        RECT -59.325 -67.485 -58.995 -67.155 ;
        RECT -59.325 -68.845 -58.995 -68.515 ;
        RECT -59.325 -70.205 -58.995 -69.875 ;
        RECT -59.325 -71.565 -58.995 -71.235 ;
        RECT -59.325 -72.925 -58.995 -72.595 ;
        RECT -59.325 -74.285 -58.995 -73.955 ;
        RECT -59.325 -75.645 -58.995 -75.315 ;
        RECT -59.325 -77.005 -58.995 -76.675 ;
        RECT -59.325 -78.365 -58.995 -78.035 ;
        RECT -59.325 -79.725 -58.995 -79.395 ;
        RECT -59.325 -81.085 -58.995 -80.755 ;
        RECT -59.325 -82.445 -58.995 -82.115 ;
        RECT -59.325 -83.805 -58.995 -83.475 ;
        RECT -59.325 -85.165 -58.995 -84.835 ;
        RECT -59.325 -86.525 -58.995 -86.195 ;
        RECT -59.325 -87.885 -58.995 -87.555 ;
        RECT -59.325 -89.245 -58.995 -88.915 ;
        RECT -59.325 -90.605 -58.995 -90.275 ;
        RECT -59.325 -91.965 -58.995 -91.635 ;
        RECT -59.325 -93.325 -58.995 -92.995 ;
        RECT -59.325 -94.685 -58.995 -94.355 ;
        RECT -59.325 -96.045 -58.995 -95.715 ;
        RECT -59.325 -97.405 -58.995 -97.075 ;
        RECT -59.325 -98.765 -58.995 -98.435 ;
        RECT -59.325 -100.125 -58.995 -99.795 ;
        RECT -59.325 -101.485 -58.995 -101.155 ;
        RECT -59.325 -102.845 -58.995 -102.515 ;
        RECT -59.325 -104.205 -58.995 -103.875 ;
        RECT -59.325 -105.565 -58.995 -105.235 ;
        RECT -59.325 -106.925 -58.995 -106.595 ;
        RECT -59.325 -108.285 -58.995 -107.955 ;
        RECT -59.325 -109.645 -58.995 -109.315 ;
        RECT -59.325 -111.005 -58.995 -110.675 ;
        RECT -59.325 -112.365 -58.995 -112.035 ;
        RECT -59.325 -113.725 -58.995 -113.395 ;
        RECT -59.325 -115.085 -58.995 -114.755 ;
        RECT -59.325 -116.445 -58.995 -116.115 ;
        RECT -59.325 -117.805 -58.995 -117.475 ;
        RECT -59.325 -119.165 -58.995 -118.835 ;
        RECT -59.325 -120.525 -58.995 -120.195 ;
        RECT -59.325 -121.885 -58.995 -121.555 ;
        RECT -59.325 -123.245 -58.995 -122.915 ;
        RECT -59.325 -124.605 -58.995 -124.275 ;
        RECT -59.325 -128.685 -58.995 -128.355 ;
        RECT -59.325 -130.045 -58.995 -129.715 ;
        RECT -59.325 -132.765 -58.995 -132.435 ;
        RECT -59.325 -134.125 -58.995 -133.795 ;
        RECT -59.325 -135.485 -58.995 -135.155 ;
        RECT -59.325 -136.845 -58.995 -136.515 ;
        RECT -59.325 -138.205 -58.995 -137.875 ;
        RECT -59.325 -139.39 -58.995 -139.06 ;
        RECT -59.325 -140.925 -58.995 -140.595 ;
        RECT -59.325 -142.285 -58.995 -141.955 ;
        RECT -59.325 -145.005 -58.995 -144.675 ;
        RECT -59.325 -146.365 -58.995 -146.035 ;
        RECT -59.325 -148.03 -58.995 -147.7 ;
        RECT -59.325 -149.085 -58.995 -148.755 ;
        RECT -59.325 -150.445 -58.995 -150.115 ;
        RECT -59.325 -153.165 -58.995 -152.835 ;
        RECT -59.325 -154.525 -58.995 -154.195 ;
        RECT -59.325 -155.885 -58.995 -155.555 ;
        RECT -59.325 -157.245 -58.995 -156.915 ;
        RECT -59.325 -158.605 -58.995 -158.275 ;
        RECT -59.325 -159.965 -58.995 -159.635 ;
        RECT -59.325 -161.325 -58.995 -160.995 ;
        RECT -59.325 -162.685 -58.995 -162.355 ;
        RECT -59.325 -164.045 -58.995 -163.715 ;
        RECT -59.325 -165.405 -58.995 -165.075 ;
        RECT -59.325 -166.765 -58.995 -166.435 ;
        RECT -59.325 -168.125 -58.995 -167.795 ;
        RECT -59.325 -169.485 -58.995 -169.155 ;
        RECT -59.325 -170.845 -58.995 -170.515 ;
        RECT -59.325 -172.205 -58.995 -171.875 ;
        RECT -59.325 -173.565 -58.995 -173.235 ;
        RECT -59.325 -174.925 -58.995 -174.595 ;
        RECT -59.325 -176.285 -58.995 -175.955 ;
        RECT -59.325 -177.645 -58.995 -177.315 ;
        RECT -59.325 -179.005 -58.995 -178.675 ;
        RECT -59.325 -180.365 -58.995 -180.035 ;
        RECT -59.325 -181.725 -58.995 -181.395 ;
        RECT -59.325 -183.085 -58.995 -182.755 ;
        RECT -59.325 -184.445 -58.995 -184.115 ;
        RECT -59.325 -185.805 -58.995 -185.475 ;
        RECT -59.325 -187.165 -58.995 -186.835 ;
        RECT -59.325 -188.525 -58.995 -188.195 ;
        RECT -59.325 -189.885 -58.995 -189.555 ;
        RECT -59.325 -191.245 -58.995 -190.915 ;
        RECT -59.325 -192.605 -58.995 -192.275 ;
        RECT -59.325 -193.965 -58.995 -193.635 ;
        RECT -59.325 -195.325 -58.995 -194.995 ;
        RECT -59.325 -196.685 -58.995 -196.355 ;
        RECT -59.325 -198.045 -58.995 -197.715 ;
        RECT -59.325 -199.405 -58.995 -199.075 ;
        RECT -59.325 -200.765 -58.995 -200.435 ;
        RECT -59.325 -202.125 -58.995 -201.795 ;
        RECT -59.325 -203.485 -58.995 -203.155 ;
        RECT -59.325 -204.845 -58.995 -204.515 ;
        RECT -59.325 -206.205 -58.995 -205.875 ;
        RECT -59.325 -207.565 -58.995 -207.235 ;
        RECT -59.325 -208.925 -58.995 -208.595 ;
        RECT -59.325 -210.285 -58.995 -209.955 ;
        RECT -59.325 -211.645 -58.995 -211.315 ;
        RECT -59.325 -213.005 -58.995 -212.675 ;
        RECT -59.325 -214.365 -58.995 -214.035 ;
        RECT -59.325 -215.725 -58.995 -215.395 ;
        RECT -59.325 -217.085 -58.995 -216.755 ;
        RECT -59.325 -218.445 -58.995 -218.115 ;
        RECT -59.325 -219.805 -58.995 -219.475 ;
        RECT -59.325 -221.165 -58.995 -220.835 ;
        RECT -59.325 -222.525 -58.995 -222.195 ;
        RECT -59.325 -223.885 -58.995 -223.555 ;
        RECT -59.325 -225.245 -58.995 -224.915 ;
        RECT -59.325 -227.965 -58.995 -227.635 ;
        RECT -59.325 -232.045 -58.995 -231.715 ;
        RECT -59.325 -233.225 -58.995 -232.895 ;
        RECT -59.325 -234.765 -58.995 -234.435 ;
        RECT -59.325 -236.125 -58.995 -235.795 ;
        RECT -59.325 -237.485 -58.995 -237.155 ;
        RECT -59.325 -238.845 -58.995 -238.515 ;
        RECT -59.325 -241.09 -58.995 -239.96 ;
        RECT -59.32 -241.205 -59 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.965 244.04 -57.635 245.17 ;
        RECT -57.965 242.595 -57.635 242.925 ;
        RECT -57.965 241.235 -57.635 241.565 ;
        RECT -57.965 239.875 -57.635 240.205 ;
        RECT -57.965 238.515 -57.635 238.845 ;
        RECT -57.965 237.155 -57.635 237.485 ;
        RECT -57.965 235.795 -57.635 236.125 ;
        RECT -57.965 234.435 -57.635 234.765 ;
        RECT -57.965 233.075 -57.635 233.405 ;
        RECT -57.965 231.715 -57.635 232.045 ;
        RECT -57.965 230.355 -57.635 230.685 ;
        RECT -57.965 228.995 -57.635 229.325 ;
        RECT -57.965 227.635 -57.635 227.965 ;
        RECT -57.965 226.275 -57.635 226.605 ;
        RECT -57.965 224.915 -57.635 225.245 ;
        RECT -57.965 223.555 -57.635 223.885 ;
        RECT -57.965 222.195 -57.635 222.525 ;
        RECT -57.965 220.835 -57.635 221.165 ;
        RECT -57.965 219.475 -57.635 219.805 ;
        RECT -57.965 218.115 -57.635 218.445 ;
        RECT -57.965 216.755 -57.635 217.085 ;
        RECT -57.965 215.395 -57.635 215.725 ;
        RECT -57.965 214.035 -57.635 214.365 ;
        RECT -57.965 212.675 -57.635 213.005 ;
        RECT -57.965 211.315 -57.635 211.645 ;
        RECT -57.965 209.955 -57.635 210.285 ;
        RECT -57.965 208.595 -57.635 208.925 ;
        RECT -57.965 207.235 -57.635 207.565 ;
        RECT -57.965 205.875 -57.635 206.205 ;
        RECT -57.965 204.515 -57.635 204.845 ;
        RECT -57.965 203.155 -57.635 203.485 ;
        RECT -57.965 201.795 -57.635 202.125 ;
        RECT -57.965 200.435 -57.635 200.765 ;
        RECT -57.965 199.075 -57.635 199.405 ;
        RECT -57.965 197.715 -57.635 198.045 ;
        RECT -57.965 196.355 -57.635 196.685 ;
        RECT -57.965 194.995 -57.635 195.325 ;
        RECT -57.965 193.635 -57.635 193.965 ;
        RECT -57.965 192.275 -57.635 192.605 ;
        RECT -57.965 190.915 -57.635 191.245 ;
        RECT -57.965 189.555 -57.635 189.885 ;
        RECT -57.965 188.195 -57.635 188.525 ;
        RECT -57.965 186.835 -57.635 187.165 ;
        RECT -57.965 185.475 -57.635 185.805 ;
        RECT -57.965 184.115 -57.635 184.445 ;
        RECT -57.965 182.755 -57.635 183.085 ;
        RECT -57.965 181.395 -57.635 181.725 ;
        RECT -57.965 180.035 -57.635 180.365 ;
        RECT -57.965 178.675 -57.635 179.005 ;
        RECT -57.965 177.315 -57.635 177.645 ;
        RECT -57.965 175.955 -57.635 176.285 ;
        RECT -57.965 174.595 -57.635 174.925 ;
        RECT -57.965 173.235 -57.635 173.565 ;
        RECT -57.965 171.875 -57.635 172.205 ;
        RECT -57.965 170.515 -57.635 170.845 ;
        RECT -57.965 169.155 -57.635 169.485 ;
        RECT -57.965 167.795 -57.635 168.125 ;
        RECT -57.965 166.435 -57.635 166.765 ;
        RECT -57.965 165.075 -57.635 165.405 ;
        RECT -57.965 163.715 -57.635 164.045 ;
        RECT -57.965 162.355 -57.635 162.685 ;
        RECT -57.965 160.995 -57.635 161.325 ;
        RECT -57.965 159.635 -57.635 159.965 ;
        RECT -57.965 158.275 -57.635 158.605 ;
        RECT -57.965 156.915 -57.635 157.245 ;
        RECT -57.965 155.555 -57.635 155.885 ;
        RECT -57.965 154.195 -57.635 154.525 ;
        RECT -57.965 152.835 -57.635 153.165 ;
        RECT -57.965 151.475 -57.635 151.805 ;
        RECT -57.965 150.115 -57.635 150.445 ;
        RECT -57.965 148.755 -57.635 149.085 ;
        RECT -57.965 147.395 -57.635 147.725 ;
        RECT -57.965 146.035 -57.635 146.365 ;
        RECT -57.965 144.675 -57.635 145.005 ;
        RECT -57.965 143.315 -57.635 143.645 ;
        RECT -57.965 141.955 -57.635 142.285 ;
        RECT -57.965 140.595 -57.635 140.925 ;
        RECT -57.965 139.235 -57.635 139.565 ;
        RECT -57.965 137.225 -57.635 137.555 ;
        RECT -57.965 135.175 -57.635 135.505 ;
        RECT -57.965 132.815 -57.635 133.145 ;
        RECT -57.965 131.665 -57.635 131.995 ;
        RECT -57.965 129.655 -57.635 129.985 ;
        RECT -57.965 128.505 -57.635 128.835 ;
        RECT -57.965 126.495 -57.635 126.825 ;
        RECT -57.965 125.345 -57.635 125.675 ;
        RECT -57.965 123.335 -57.635 123.665 ;
        RECT -57.965 122.185 -57.635 122.515 ;
        RECT -57.965 120.175 -57.635 120.505 ;
        RECT -57.965 119.025 -57.635 119.355 ;
        RECT -57.965 117.185 -57.635 117.515 ;
        RECT -57.965 115.865 -57.635 116.195 ;
        RECT -57.965 113.855 -57.635 114.185 ;
        RECT -57.965 112.705 -57.635 113.035 ;
        RECT -57.965 110.695 -57.635 111.025 ;
        RECT -57.965 109.545 -57.635 109.875 ;
        RECT -57.965 107.535 -57.635 107.865 ;
        RECT -57.965 106.385 -57.635 106.715 ;
        RECT -57.965 104.375 -57.635 104.705 ;
        RECT -57.965 103.225 -57.635 103.555 ;
        RECT -57.965 100.865 -57.635 101.195 ;
        RECT -57.965 98.81 -57.635 99.14 ;
        RECT -57.965 97.075 -57.635 97.405 ;
        RECT -57.965 95.715 -57.635 96.045 ;
        RECT -57.965 94.355 -57.635 94.685 ;
        RECT -57.965 92.995 -57.635 93.325 ;
        RECT -57.965 91.635 -57.635 91.965 ;
        RECT -57.965 90.275 -57.635 90.605 ;
        RECT -57.965 88.915 -57.635 89.245 ;
        RECT -57.965 87.555 -57.635 87.885 ;
        RECT -57.965 86.195 -57.635 86.525 ;
        RECT -57.965 84.835 -57.635 85.165 ;
        RECT -57.965 83.475 -57.635 83.805 ;
        RECT -57.965 82.115 -57.635 82.445 ;
        RECT -57.965 80.755 -57.635 81.085 ;
        RECT -57.965 79.395 -57.635 79.725 ;
        RECT -57.965 78.035 -57.635 78.365 ;
        RECT -57.965 76.675 -57.635 77.005 ;
        RECT -57.965 75.315 -57.635 75.645 ;
        RECT -57.965 73.955 -57.635 74.285 ;
        RECT -57.965 72.595 -57.635 72.925 ;
        RECT -57.965 71.235 -57.635 71.565 ;
        RECT -57.965 69.875 -57.635 70.205 ;
        RECT -57.965 68.515 -57.635 68.845 ;
        RECT -57.965 67.155 -57.635 67.485 ;
        RECT -57.965 65.795 -57.635 66.125 ;
        RECT -57.965 64.435 -57.635 64.765 ;
        RECT -57.965 63.075 -57.635 63.405 ;
        RECT -57.965 61.715 -57.635 62.045 ;
        RECT -57.965 60.355 -57.635 60.685 ;
        RECT -57.965 58.995 -57.635 59.325 ;
        RECT -57.965 57.635 -57.635 57.965 ;
        RECT -57.965 56.275 -57.635 56.605 ;
        RECT -57.965 54.915 -57.635 55.245 ;
        RECT -57.965 53.555 -57.635 53.885 ;
        RECT -57.965 52.195 -57.635 52.525 ;
        RECT -57.965 50.835 -57.635 51.165 ;
        RECT -57.965 49.475 -57.635 49.805 ;
        RECT -57.965 48.115 -57.635 48.445 ;
        RECT -57.965 46.755 -57.635 47.085 ;
        RECT -57.965 45.395 -57.635 45.725 ;
        RECT -57.965 44.035 -57.635 44.365 ;
        RECT -57.965 42.675 -57.635 43.005 ;
        RECT -57.965 41.315 -57.635 41.645 ;
        RECT -57.965 39.955 -57.635 40.285 ;
        RECT -57.965 38.595 -57.635 38.925 ;
        RECT -57.965 37.235 -57.635 37.565 ;
        RECT -57.965 35.875 -57.635 36.205 ;
        RECT -57.965 34.515 -57.635 34.845 ;
        RECT -57.965 33.155 -57.635 33.485 ;
        RECT -57.965 31.795 -57.635 32.125 ;
        RECT -57.965 30.435 -57.635 30.765 ;
        RECT -57.965 29.075 -57.635 29.405 ;
        RECT -57.965 27.715 -57.635 28.045 ;
        RECT -57.965 26.355 -57.635 26.685 ;
        RECT -57.965 24.995 -57.635 25.325 ;
        RECT -57.965 23.635 -57.635 23.965 ;
        RECT -57.965 22.275 -57.635 22.605 ;
        RECT -57.965 20.915 -57.635 21.245 ;
        RECT -57.965 19.555 -57.635 19.885 ;
        RECT -57.965 18.195 -57.635 18.525 ;
        RECT -57.965 16.835 -57.635 17.165 ;
        RECT -57.965 15.475 -57.635 15.805 ;
        RECT -57.965 14.115 -57.635 14.445 ;
        RECT -57.965 12.755 -57.635 13.085 ;
        RECT -57.965 11.395 -57.635 11.725 ;
        RECT -57.965 10.035 -57.635 10.365 ;
        RECT -57.965 8.675 -57.635 9.005 ;
        RECT -57.965 7.315 -57.635 7.645 ;
        RECT -57.965 5.955 -57.635 6.285 ;
        RECT -57.965 4.595 -57.635 4.925 ;
        RECT -57.965 3.235 -57.635 3.565 ;
        RECT -57.965 1.875 -57.635 2.205 ;
        RECT -57.965 0.515 -57.635 0.845 ;
        RECT -57.965 -0.845 -57.635 -0.515 ;
        RECT -57.965 -2.205 -57.635 -1.875 ;
        RECT -57.965 -3.565 -57.635 -3.235 ;
        RECT -57.965 -4.925 -57.635 -4.595 ;
        RECT -57.965 -6.285 -57.635 -5.955 ;
        RECT -57.965 -7.645 -57.635 -7.315 ;
        RECT -57.965 -9.005 -57.635 -8.675 ;
        RECT -57.965 -10.365 -57.635 -10.035 ;
        RECT -57.965 -11.725 -57.635 -11.395 ;
        RECT -57.965 -13.085 -57.635 -12.755 ;
        RECT -57.965 -14.445 -57.635 -14.115 ;
        RECT -57.965 -15.805 -57.635 -15.475 ;
        RECT -57.965 -17.165 -57.635 -16.835 ;
        RECT -57.965 -18.525 -57.635 -18.195 ;
        RECT -57.965 -19.885 -57.635 -19.555 ;
        RECT -57.965 -21.245 -57.635 -20.915 ;
        RECT -57.965 -22.605 -57.635 -22.275 ;
        RECT -57.965 -23.965 -57.635 -23.635 ;
        RECT -57.965 -25.325 -57.635 -24.995 ;
        RECT -57.965 -26.685 -57.635 -26.355 ;
        RECT -57.965 -28.045 -57.635 -27.715 ;
        RECT -57.965 -29.405 -57.635 -29.075 ;
        RECT -57.965 -30.765 -57.635 -30.435 ;
        RECT -57.965 -32.125 -57.635 -31.795 ;
        RECT -57.965 -33.485 -57.635 -33.155 ;
        RECT -57.965 -34.845 -57.635 -34.515 ;
        RECT -57.965 -36.205 -57.635 -35.875 ;
        RECT -57.965 -37.565 -57.635 -37.235 ;
        RECT -57.965 -38.925 -57.635 -38.595 ;
        RECT -57.965 -40.285 -57.635 -39.955 ;
        RECT -57.965 -41.645 -57.635 -41.315 ;
        RECT -57.965 -43.005 -57.635 -42.675 ;
        RECT -57.965 -44.365 -57.635 -44.035 ;
        RECT -57.965 -45.725 -57.635 -45.395 ;
        RECT -57.965 -47.085 -57.635 -46.755 ;
        RECT -57.965 -48.445 -57.635 -48.115 ;
        RECT -57.965 -49.805 -57.635 -49.475 ;
        RECT -57.965 -51.165 -57.635 -50.835 ;
        RECT -57.965 -52.525 -57.635 -52.195 ;
        RECT -57.965 -53.885 -57.635 -53.555 ;
        RECT -57.965 -55.245 -57.635 -54.915 ;
        RECT -57.965 -56.605 -57.635 -56.275 ;
        RECT -57.965 -57.965 -57.635 -57.635 ;
        RECT -57.965 -59.325 -57.635 -58.995 ;
        RECT -57.965 -60.685 -57.635 -60.355 ;
        RECT -57.965 -62.045 -57.635 -61.715 ;
        RECT -57.965 -63.405 -57.635 -63.075 ;
        RECT -57.965 -64.765 -57.635 -64.435 ;
        RECT -57.965 -66.125 -57.635 -65.795 ;
        RECT -57.965 -67.485 -57.635 -67.155 ;
        RECT -57.965 -68.845 -57.635 -68.515 ;
        RECT -57.965 -70.205 -57.635 -69.875 ;
        RECT -57.965 -71.565 -57.635 -71.235 ;
        RECT -57.965 -72.925 -57.635 -72.595 ;
        RECT -57.965 -74.285 -57.635 -73.955 ;
        RECT -57.965 -75.645 -57.635 -75.315 ;
        RECT -57.965 -77.005 -57.635 -76.675 ;
        RECT -57.965 -78.365 -57.635 -78.035 ;
        RECT -57.965 -79.725 -57.635 -79.395 ;
        RECT -57.965 -81.085 -57.635 -80.755 ;
        RECT -57.965 -82.445 -57.635 -82.115 ;
        RECT -57.965 -83.805 -57.635 -83.475 ;
        RECT -57.965 -85.165 -57.635 -84.835 ;
        RECT -57.965 -86.525 -57.635 -86.195 ;
        RECT -57.965 -87.885 -57.635 -87.555 ;
        RECT -57.965 -89.245 -57.635 -88.915 ;
        RECT -57.965 -90.605 -57.635 -90.275 ;
        RECT -57.965 -91.965 -57.635 -91.635 ;
        RECT -57.965 -93.325 -57.635 -92.995 ;
        RECT -57.965 -94.685 -57.635 -94.355 ;
        RECT -57.965 -96.045 -57.635 -95.715 ;
        RECT -57.965 -97.405 -57.635 -97.075 ;
        RECT -57.965 -98.765 -57.635 -98.435 ;
        RECT -57.965 -100.125 -57.635 -99.795 ;
        RECT -57.965 -101.485 -57.635 -101.155 ;
        RECT -57.965 -102.845 -57.635 -102.515 ;
        RECT -57.965 -104.205 -57.635 -103.875 ;
        RECT -57.965 -105.565 -57.635 -105.235 ;
        RECT -57.965 -106.925 -57.635 -106.595 ;
        RECT -57.965 -108.285 -57.635 -107.955 ;
        RECT -57.965 -109.645 -57.635 -109.315 ;
        RECT -57.965 -111.005 -57.635 -110.675 ;
        RECT -57.965 -112.365 -57.635 -112.035 ;
        RECT -57.965 -113.725 -57.635 -113.395 ;
        RECT -57.965 -115.085 -57.635 -114.755 ;
        RECT -57.965 -116.445 -57.635 -116.115 ;
        RECT -57.965 -117.805 -57.635 -117.475 ;
        RECT -57.965 -119.165 -57.635 -118.835 ;
        RECT -57.965 -120.525 -57.635 -120.195 ;
        RECT -57.965 -121.885 -57.635 -121.555 ;
        RECT -57.965 -124.605 -57.635 -124.275 ;
        RECT -57.965 -128.685 -57.635 -128.355 ;
        RECT -57.965 -130.045 -57.635 -129.715 ;
        RECT -57.965 -132.765 -57.635 -132.435 ;
        RECT -57.965 -134.125 -57.635 -133.795 ;
        RECT -57.965 -135.485 -57.635 -135.155 ;
        RECT -57.965 -136.845 -57.635 -136.515 ;
        RECT -57.965 -138.205 -57.635 -137.875 ;
        RECT -57.965 -139.39 -57.635 -139.06 ;
        RECT -57.965 -140.925 -57.635 -140.595 ;
        RECT -57.965 -142.285 -57.635 -141.955 ;
        RECT -57.965 -145.005 -57.635 -144.675 ;
        RECT -57.965 -146.365 -57.635 -146.035 ;
        RECT -57.965 -148.03 -57.635 -147.7 ;
        RECT -57.965 -149.085 -57.635 -148.755 ;
        RECT -57.96 -149.76 -57.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.965 -232.045 -57.635 -231.715 ;
        RECT -57.965 -233.225 -57.635 -232.895 ;
        RECT -57.965 -234.765 -57.635 -234.435 ;
        RECT -57.965 -236.125 -57.635 -235.795 ;
        RECT -57.965 -237.485 -57.635 -237.155 ;
        RECT -57.965 -238.845 -57.635 -238.515 ;
        RECT -57.965 -241.09 -57.635 -239.96 ;
        RECT -57.96 -241.205 -57.64 -231.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 214.035 -56.275 214.365 ;
        RECT -56.605 212.675 -56.275 213.005 ;
        RECT -56.605 211.315 -56.275 211.645 ;
        RECT -56.605 209.955 -56.275 210.285 ;
        RECT -56.605 208.595 -56.275 208.925 ;
        RECT -56.605 207.235 -56.275 207.565 ;
        RECT -56.605 205.875 -56.275 206.205 ;
        RECT -56.605 204.515 -56.275 204.845 ;
        RECT -56.605 203.155 -56.275 203.485 ;
        RECT -56.605 201.795 -56.275 202.125 ;
        RECT -56.605 200.435 -56.275 200.765 ;
        RECT -56.605 199.075 -56.275 199.405 ;
        RECT -56.605 197.715 -56.275 198.045 ;
        RECT -56.605 196.355 -56.275 196.685 ;
        RECT -56.605 194.995 -56.275 195.325 ;
        RECT -56.605 193.635 -56.275 193.965 ;
        RECT -56.605 192.275 -56.275 192.605 ;
        RECT -56.605 190.915 -56.275 191.245 ;
        RECT -56.605 189.555 -56.275 189.885 ;
        RECT -56.605 188.195 -56.275 188.525 ;
        RECT -56.605 186.835 -56.275 187.165 ;
        RECT -56.605 185.475 -56.275 185.805 ;
        RECT -56.605 184.115 -56.275 184.445 ;
        RECT -56.605 182.755 -56.275 183.085 ;
        RECT -56.605 181.395 -56.275 181.725 ;
        RECT -56.605 180.035 -56.275 180.365 ;
        RECT -56.605 178.675 -56.275 179.005 ;
        RECT -56.605 177.315 -56.275 177.645 ;
        RECT -56.605 175.955 -56.275 176.285 ;
        RECT -56.605 174.595 -56.275 174.925 ;
        RECT -56.605 173.235 -56.275 173.565 ;
        RECT -56.605 171.875 -56.275 172.205 ;
        RECT -56.605 170.515 -56.275 170.845 ;
        RECT -56.605 169.155 -56.275 169.485 ;
        RECT -56.605 167.795 -56.275 168.125 ;
        RECT -56.605 166.435 -56.275 166.765 ;
        RECT -56.605 165.075 -56.275 165.405 ;
        RECT -56.605 163.715 -56.275 164.045 ;
        RECT -56.605 162.355 -56.275 162.685 ;
        RECT -56.605 160.995 -56.275 161.325 ;
        RECT -56.605 159.635 -56.275 159.965 ;
        RECT -56.605 158.275 -56.275 158.605 ;
        RECT -56.605 156.915 -56.275 157.245 ;
        RECT -56.605 155.555 -56.275 155.885 ;
        RECT -56.605 154.195 -56.275 154.525 ;
        RECT -56.605 152.835 -56.275 153.165 ;
        RECT -56.605 151.475 -56.275 151.805 ;
        RECT -56.605 150.115 -56.275 150.445 ;
        RECT -56.605 148.755 -56.275 149.085 ;
        RECT -56.605 147.395 -56.275 147.725 ;
        RECT -56.605 146.035 -56.275 146.365 ;
        RECT -56.605 144.675 -56.275 145.005 ;
        RECT -56.605 143.315 -56.275 143.645 ;
        RECT -56.605 141.955 -56.275 142.285 ;
        RECT -56.605 140.595 -56.275 140.925 ;
        RECT -56.605 139.235 -56.275 139.565 ;
        RECT -56.605 137.225 -56.275 137.555 ;
        RECT -56.605 135.175 -56.275 135.505 ;
        RECT -56.605 132.815 -56.275 133.145 ;
        RECT -56.605 131.665 -56.275 131.995 ;
        RECT -56.605 129.655 -56.275 129.985 ;
        RECT -56.605 128.505 -56.275 128.835 ;
        RECT -56.605 126.495 -56.275 126.825 ;
        RECT -56.605 125.345 -56.275 125.675 ;
        RECT -56.605 123.335 -56.275 123.665 ;
        RECT -56.605 122.185 -56.275 122.515 ;
        RECT -56.605 120.175 -56.275 120.505 ;
        RECT -56.605 119.025 -56.275 119.355 ;
        RECT -56.605 117.185 -56.275 117.515 ;
        RECT -56.605 115.865 -56.275 116.195 ;
        RECT -56.605 113.855 -56.275 114.185 ;
        RECT -56.605 112.705 -56.275 113.035 ;
        RECT -56.605 110.695 -56.275 111.025 ;
        RECT -56.605 109.545 -56.275 109.875 ;
        RECT -56.605 107.535 -56.275 107.865 ;
        RECT -56.605 106.385 -56.275 106.715 ;
        RECT -56.605 104.375 -56.275 104.705 ;
        RECT -56.605 103.225 -56.275 103.555 ;
        RECT -56.605 100.865 -56.275 101.195 ;
        RECT -56.605 98.81 -56.275 99.14 ;
        RECT -56.605 97.075 -56.275 97.405 ;
        RECT -56.605 95.715 -56.275 96.045 ;
        RECT -56.605 94.355 -56.275 94.685 ;
        RECT -56.605 92.995 -56.275 93.325 ;
        RECT -56.605 91.635 -56.275 91.965 ;
        RECT -56.605 90.275 -56.275 90.605 ;
        RECT -56.605 88.915 -56.275 89.245 ;
        RECT -56.6 86.88 -56.28 245.285 ;
        RECT -56.605 244.04 -56.275 245.17 ;
        RECT -56.605 242.595 -56.275 242.925 ;
        RECT -56.605 241.235 -56.275 241.565 ;
        RECT -56.605 239.875 -56.275 240.205 ;
        RECT -56.605 238.515 -56.275 238.845 ;
        RECT -56.605 237.155 -56.275 237.485 ;
        RECT -56.605 235.795 -56.275 236.125 ;
        RECT -56.605 234.435 -56.275 234.765 ;
        RECT -56.605 233.075 -56.275 233.405 ;
        RECT -56.605 231.715 -56.275 232.045 ;
        RECT -56.605 230.355 -56.275 230.685 ;
        RECT -56.605 228.995 -56.275 229.325 ;
        RECT -56.605 227.635 -56.275 227.965 ;
        RECT -56.605 226.275 -56.275 226.605 ;
        RECT -56.605 224.915 -56.275 225.245 ;
        RECT -56.605 223.555 -56.275 223.885 ;
        RECT -56.605 222.195 -56.275 222.525 ;
        RECT -56.605 220.835 -56.275 221.165 ;
        RECT -56.605 219.475 -56.275 219.805 ;
        RECT -56.605 218.115 -56.275 218.445 ;
        RECT -56.605 216.755 -56.275 217.085 ;
        RECT -56.605 215.395 -56.275 215.725 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.405 244.04 -63.075 245.17 ;
        RECT -63.405 242.595 -63.075 242.925 ;
        RECT -63.405 241.235 -63.075 241.565 ;
        RECT -63.405 239.875 -63.075 240.205 ;
        RECT -63.405 238.515 -63.075 238.845 ;
        RECT -63.405 237.155 -63.075 237.485 ;
        RECT -63.405 235.795 -63.075 236.125 ;
        RECT -63.405 234.435 -63.075 234.765 ;
        RECT -63.405 233.075 -63.075 233.405 ;
        RECT -63.405 231.715 -63.075 232.045 ;
        RECT -63.405 230.355 -63.075 230.685 ;
        RECT -63.405 228.995 -63.075 229.325 ;
        RECT -63.405 227.635 -63.075 227.965 ;
        RECT -63.405 226.275 -63.075 226.605 ;
        RECT -63.405 224.915 -63.075 225.245 ;
        RECT -63.405 223.555 -63.075 223.885 ;
        RECT -63.405 222.195 -63.075 222.525 ;
        RECT -63.405 220.835 -63.075 221.165 ;
        RECT -63.405 219.475 -63.075 219.805 ;
        RECT -63.405 218.115 -63.075 218.445 ;
        RECT -63.405 216.755 -63.075 217.085 ;
        RECT -63.405 215.395 -63.075 215.725 ;
        RECT -63.405 214.035 -63.075 214.365 ;
        RECT -63.405 212.675 -63.075 213.005 ;
        RECT -63.405 211.315 -63.075 211.645 ;
        RECT -63.405 209.955 -63.075 210.285 ;
        RECT -63.405 208.595 -63.075 208.925 ;
        RECT -63.405 207.235 -63.075 207.565 ;
        RECT -63.405 205.875 -63.075 206.205 ;
        RECT -63.405 204.515 -63.075 204.845 ;
        RECT -63.405 203.155 -63.075 203.485 ;
        RECT -63.405 201.795 -63.075 202.125 ;
        RECT -63.405 200.435 -63.075 200.765 ;
        RECT -63.405 199.075 -63.075 199.405 ;
        RECT -63.405 197.715 -63.075 198.045 ;
        RECT -63.405 196.355 -63.075 196.685 ;
        RECT -63.405 194.995 -63.075 195.325 ;
        RECT -63.405 193.635 -63.075 193.965 ;
        RECT -63.405 192.275 -63.075 192.605 ;
        RECT -63.405 190.915 -63.075 191.245 ;
        RECT -63.405 189.555 -63.075 189.885 ;
        RECT -63.405 188.195 -63.075 188.525 ;
        RECT -63.405 186.835 -63.075 187.165 ;
        RECT -63.405 185.475 -63.075 185.805 ;
        RECT -63.405 184.115 -63.075 184.445 ;
        RECT -63.405 182.755 -63.075 183.085 ;
        RECT -63.405 181.395 -63.075 181.725 ;
        RECT -63.405 180.035 -63.075 180.365 ;
        RECT -63.405 178.675 -63.075 179.005 ;
        RECT -63.405 177.315 -63.075 177.645 ;
        RECT -63.405 175.955 -63.075 176.285 ;
        RECT -63.405 174.595 -63.075 174.925 ;
        RECT -63.405 173.235 -63.075 173.565 ;
        RECT -63.405 171.875 -63.075 172.205 ;
        RECT -63.405 170.515 -63.075 170.845 ;
        RECT -63.405 169.155 -63.075 169.485 ;
        RECT -63.405 167.795 -63.075 168.125 ;
        RECT -63.405 166.435 -63.075 166.765 ;
        RECT -63.405 165.075 -63.075 165.405 ;
        RECT -63.405 163.715 -63.075 164.045 ;
        RECT -63.405 162.355 -63.075 162.685 ;
        RECT -63.405 160.995 -63.075 161.325 ;
        RECT -63.405 159.635 -63.075 159.965 ;
        RECT -63.405 158.275 -63.075 158.605 ;
        RECT -63.405 156.915 -63.075 157.245 ;
        RECT -63.405 155.555 -63.075 155.885 ;
        RECT -63.405 154.195 -63.075 154.525 ;
        RECT -63.405 152.835 -63.075 153.165 ;
        RECT -63.405 151.475 -63.075 151.805 ;
        RECT -63.405 150.115 -63.075 150.445 ;
        RECT -63.405 148.755 -63.075 149.085 ;
        RECT -63.405 147.395 -63.075 147.725 ;
        RECT -63.405 146.035 -63.075 146.365 ;
        RECT -63.405 144.675 -63.075 145.005 ;
        RECT -63.405 143.315 -63.075 143.645 ;
        RECT -63.405 141.955 -63.075 142.285 ;
        RECT -63.405 140.595 -63.075 140.925 ;
        RECT -63.405 139.235 -63.075 139.565 ;
        RECT -63.405 137.875 -63.075 138.205 ;
        RECT -63.405 136.515 -63.075 136.845 ;
        RECT -63.405 135.155 -63.075 135.485 ;
        RECT -63.405 133.795 -63.075 134.125 ;
        RECT -63.405 132.435 -63.075 132.765 ;
        RECT -63.405 131.075 -63.075 131.405 ;
        RECT -63.405 129.715 -63.075 130.045 ;
        RECT -63.405 128.355 -63.075 128.685 ;
        RECT -63.405 126.995 -63.075 127.325 ;
        RECT -63.405 125.635 -63.075 125.965 ;
        RECT -63.405 124.275 -63.075 124.605 ;
        RECT -63.405 122.915 -63.075 123.245 ;
        RECT -63.405 121.555 -63.075 121.885 ;
        RECT -63.405 120.195 -63.075 120.525 ;
        RECT -63.405 118.835 -63.075 119.165 ;
        RECT -63.405 117.475 -63.075 117.805 ;
        RECT -63.405 116.115 -63.075 116.445 ;
        RECT -63.405 114.755 -63.075 115.085 ;
        RECT -63.405 113.395 -63.075 113.725 ;
        RECT -63.405 112.035 -63.075 112.365 ;
        RECT -63.405 110.675 -63.075 111.005 ;
        RECT -63.405 109.315 -63.075 109.645 ;
        RECT -63.405 107.955 -63.075 108.285 ;
        RECT -63.405 106.595 -63.075 106.925 ;
        RECT -63.405 105.235 -63.075 105.565 ;
        RECT -63.405 103.875 -63.075 104.205 ;
        RECT -63.405 102.515 -63.075 102.845 ;
        RECT -63.405 101.155 -63.075 101.485 ;
        RECT -63.405 99.795 -63.075 100.125 ;
        RECT -63.405 98.435 -63.075 98.765 ;
        RECT -63.405 97.075 -63.075 97.405 ;
        RECT -63.405 95.715 -63.075 96.045 ;
        RECT -63.405 94.355 -63.075 94.685 ;
        RECT -63.405 92.995 -63.075 93.325 ;
        RECT -63.405 91.635 -63.075 91.965 ;
        RECT -63.405 90.275 -63.075 90.605 ;
        RECT -63.405 88.915 -63.075 89.245 ;
        RECT -63.405 87.555 -63.075 87.885 ;
        RECT -63.405 86.195 -63.075 86.525 ;
        RECT -63.405 84.835 -63.075 85.165 ;
        RECT -63.405 83.475 -63.075 83.805 ;
        RECT -63.405 82.115 -63.075 82.445 ;
        RECT -63.405 80.755 -63.075 81.085 ;
        RECT -63.405 79.395 -63.075 79.725 ;
        RECT -63.405 78.035 -63.075 78.365 ;
        RECT -63.405 76.675 -63.075 77.005 ;
        RECT -63.405 75.315 -63.075 75.645 ;
        RECT -63.405 73.955 -63.075 74.285 ;
        RECT -63.405 72.595 -63.075 72.925 ;
        RECT -63.405 71.235 -63.075 71.565 ;
        RECT -63.405 69.875 -63.075 70.205 ;
        RECT -63.405 68.515 -63.075 68.845 ;
        RECT -63.405 67.155 -63.075 67.485 ;
        RECT -63.405 65.795 -63.075 66.125 ;
        RECT -63.405 64.435 -63.075 64.765 ;
        RECT -63.405 63.075 -63.075 63.405 ;
        RECT -63.405 61.715 -63.075 62.045 ;
        RECT -63.405 60.355 -63.075 60.685 ;
        RECT -63.405 58.995 -63.075 59.325 ;
        RECT -63.405 57.635 -63.075 57.965 ;
        RECT -63.405 56.275 -63.075 56.605 ;
        RECT -63.405 54.915 -63.075 55.245 ;
        RECT -63.405 53.555 -63.075 53.885 ;
        RECT -63.405 52.195 -63.075 52.525 ;
        RECT -63.405 50.835 -63.075 51.165 ;
        RECT -63.405 49.475 -63.075 49.805 ;
        RECT -63.405 48.115 -63.075 48.445 ;
        RECT -63.405 46.755 -63.075 47.085 ;
        RECT -63.405 45.395 -63.075 45.725 ;
        RECT -63.405 44.035 -63.075 44.365 ;
        RECT -63.405 42.675 -63.075 43.005 ;
        RECT -63.405 41.315 -63.075 41.645 ;
        RECT -63.405 39.955 -63.075 40.285 ;
        RECT -63.405 38.595 -63.075 38.925 ;
        RECT -63.405 37.235 -63.075 37.565 ;
        RECT -63.405 35.875 -63.075 36.205 ;
        RECT -63.405 34.515 -63.075 34.845 ;
        RECT -63.405 33.155 -63.075 33.485 ;
        RECT -63.405 31.795 -63.075 32.125 ;
        RECT -63.405 30.435 -63.075 30.765 ;
        RECT -63.405 29.075 -63.075 29.405 ;
        RECT -63.405 27.715 -63.075 28.045 ;
        RECT -63.405 26.355 -63.075 26.685 ;
        RECT -63.405 24.995 -63.075 25.325 ;
        RECT -63.405 23.635 -63.075 23.965 ;
        RECT -63.405 22.275 -63.075 22.605 ;
        RECT -63.405 20.915 -63.075 21.245 ;
        RECT -63.405 19.555 -63.075 19.885 ;
        RECT -63.405 18.195 -63.075 18.525 ;
        RECT -63.405 16.835 -63.075 17.165 ;
        RECT -63.405 15.475 -63.075 15.805 ;
        RECT -63.405 14.115 -63.075 14.445 ;
        RECT -63.405 12.755 -63.075 13.085 ;
        RECT -63.405 11.395 -63.075 11.725 ;
        RECT -63.405 10.035 -63.075 10.365 ;
        RECT -63.405 8.675 -63.075 9.005 ;
        RECT -63.405 7.315 -63.075 7.645 ;
        RECT -63.405 5.955 -63.075 6.285 ;
        RECT -63.405 4.595 -63.075 4.925 ;
        RECT -63.405 3.235 -63.075 3.565 ;
        RECT -63.405 1.875 -63.075 2.205 ;
        RECT -63.405 0.515 -63.075 0.845 ;
        RECT -63.405 -0.845 -63.075 -0.515 ;
        RECT -63.405 -2.205 -63.075 -1.875 ;
        RECT -63.405 -3.565 -63.075 -3.235 ;
        RECT -63.405 -4.925 -63.075 -4.595 ;
        RECT -63.405 -6.285 -63.075 -5.955 ;
        RECT -63.405 -7.645 -63.075 -7.315 ;
        RECT -63.405 -9.005 -63.075 -8.675 ;
        RECT -63.405 -10.365 -63.075 -10.035 ;
        RECT -63.405 -11.725 -63.075 -11.395 ;
        RECT -63.405 -13.085 -63.075 -12.755 ;
        RECT -63.405 -14.445 -63.075 -14.115 ;
        RECT -63.405 -15.805 -63.075 -15.475 ;
        RECT -63.405 -17.165 -63.075 -16.835 ;
        RECT -63.405 -18.525 -63.075 -18.195 ;
        RECT -63.405 -19.885 -63.075 -19.555 ;
        RECT -63.405 -21.245 -63.075 -20.915 ;
        RECT -63.405 -22.605 -63.075 -22.275 ;
        RECT -63.405 -23.965 -63.075 -23.635 ;
        RECT -63.405 -25.325 -63.075 -24.995 ;
        RECT -63.405 -26.685 -63.075 -26.355 ;
        RECT -63.405 -28.045 -63.075 -27.715 ;
        RECT -63.405 -29.405 -63.075 -29.075 ;
        RECT -63.405 -30.765 -63.075 -30.435 ;
        RECT -63.405 -32.125 -63.075 -31.795 ;
        RECT -63.405 -33.485 -63.075 -33.155 ;
        RECT -63.405 -34.845 -63.075 -34.515 ;
        RECT -63.405 -36.205 -63.075 -35.875 ;
        RECT -63.405 -37.565 -63.075 -37.235 ;
        RECT -63.405 -38.925 -63.075 -38.595 ;
        RECT -63.405 -40.285 -63.075 -39.955 ;
        RECT -63.405 -41.645 -63.075 -41.315 ;
        RECT -63.405 -43.005 -63.075 -42.675 ;
        RECT -63.405 -44.365 -63.075 -44.035 ;
        RECT -63.405 -45.725 -63.075 -45.395 ;
        RECT -63.405 -47.085 -63.075 -46.755 ;
        RECT -63.405 -48.445 -63.075 -48.115 ;
        RECT -63.405 -49.805 -63.075 -49.475 ;
        RECT -63.405 -51.165 -63.075 -50.835 ;
        RECT -63.405 -52.525 -63.075 -52.195 ;
        RECT -63.405 -53.885 -63.075 -53.555 ;
        RECT -63.405 -55.245 -63.075 -54.915 ;
        RECT -63.405 -56.605 -63.075 -56.275 ;
        RECT -63.405 -57.965 -63.075 -57.635 ;
        RECT -63.405 -59.325 -63.075 -58.995 ;
        RECT -63.405 -60.685 -63.075 -60.355 ;
        RECT -63.405 -62.045 -63.075 -61.715 ;
        RECT -63.405 -63.405 -63.075 -63.075 ;
        RECT -63.405 -64.765 -63.075 -64.435 ;
        RECT -63.405 -66.125 -63.075 -65.795 ;
        RECT -63.405 -67.485 -63.075 -67.155 ;
        RECT -63.405 -68.845 -63.075 -68.515 ;
        RECT -63.405 -70.205 -63.075 -69.875 ;
        RECT -63.405 -71.565 -63.075 -71.235 ;
        RECT -63.405 -72.925 -63.075 -72.595 ;
        RECT -63.405 -74.285 -63.075 -73.955 ;
        RECT -63.405 -75.645 -63.075 -75.315 ;
        RECT -63.405 -77.005 -63.075 -76.675 ;
        RECT -63.405 -78.365 -63.075 -78.035 ;
        RECT -63.405 -79.725 -63.075 -79.395 ;
        RECT -63.405 -81.085 -63.075 -80.755 ;
        RECT -63.405 -82.445 -63.075 -82.115 ;
        RECT -63.405 -83.805 -63.075 -83.475 ;
        RECT -63.405 -85.165 -63.075 -84.835 ;
        RECT -63.405 -86.525 -63.075 -86.195 ;
        RECT -63.405 -87.885 -63.075 -87.555 ;
        RECT -63.405 -89.245 -63.075 -88.915 ;
        RECT -63.405 -90.605 -63.075 -90.275 ;
        RECT -63.405 -91.965 -63.075 -91.635 ;
        RECT -63.405 -93.325 -63.075 -92.995 ;
        RECT -63.405 -94.685 -63.075 -94.355 ;
        RECT -63.405 -96.045 -63.075 -95.715 ;
        RECT -63.405 -97.405 -63.075 -97.075 ;
        RECT -63.405 -98.765 -63.075 -98.435 ;
        RECT -63.405 -100.125 -63.075 -99.795 ;
        RECT -63.405 -101.485 -63.075 -101.155 ;
        RECT -63.405 -102.845 -63.075 -102.515 ;
        RECT -63.405 -104.205 -63.075 -103.875 ;
        RECT -63.405 -105.565 -63.075 -105.235 ;
        RECT -63.405 -106.925 -63.075 -106.595 ;
        RECT -63.405 -108.285 -63.075 -107.955 ;
        RECT -63.405 -109.645 -63.075 -109.315 ;
        RECT -63.405 -111.005 -63.075 -110.675 ;
        RECT -63.405 -112.365 -63.075 -112.035 ;
        RECT -63.405 -113.725 -63.075 -113.395 ;
        RECT -63.405 -115.085 -63.075 -114.755 ;
        RECT -63.405 -116.445 -63.075 -116.115 ;
        RECT -63.405 -117.805 -63.075 -117.475 ;
        RECT -63.405 -119.165 -63.075 -118.835 ;
        RECT -63.405 -120.525 -63.075 -120.195 ;
        RECT -63.405 -121.885 -63.075 -121.555 ;
        RECT -63.405 -123.245 -63.075 -122.915 ;
        RECT -63.405 -124.605 -63.075 -124.275 ;
        RECT -63.405 -125.965 -63.075 -125.635 ;
        RECT -63.405 -128.685 -63.075 -128.355 ;
        RECT -63.405 -130.045 -63.075 -129.715 ;
        RECT -63.405 -132.765 -63.075 -132.435 ;
        RECT -63.405 -134.125 -63.075 -133.795 ;
        RECT -63.405 -135.485 -63.075 -135.155 ;
        RECT -63.405 -136.845 -63.075 -136.515 ;
        RECT -63.405 -138.205 -63.075 -137.875 ;
        RECT -63.405 -139.39 -63.075 -139.06 ;
        RECT -63.405 -140.925 -63.075 -140.595 ;
        RECT -63.405 -142.285 -63.075 -141.955 ;
        RECT -63.405 -145.005 -63.075 -144.675 ;
        RECT -63.405 -146.365 -63.075 -146.035 ;
        RECT -63.405 -148.03 -63.075 -147.7 ;
        RECT -63.405 -149.085 -63.075 -148.755 ;
        RECT -63.405 -150.445 -63.075 -150.115 ;
        RECT -63.4 -151.8 -63.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.405 -232.045 -63.075 -231.715 ;
        RECT -63.405 -233.225 -63.075 -232.895 ;
        RECT -63.405 -234.765 -63.075 -234.435 ;
        RECT -63.405 -236.125 -63.075 -235.795 ;
        RECT -63.405 -237.485 -63.075 -237.155 ;
        RECT -63.405 -238.845 -63.075 -238.515 ;
        RECT -63.405 -241.09 -63.075 -239.96 ;
        RECT -63.4 -241.205 -63.08 -231.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.045 244.04 -61.715 245.17 ;
        RECT -62.045 242.595 -61.715 242.925 ;
        RECT -62.045 241.235 -61.715 241.565 ;
        RECT -62.045 239.875 -61.715 240.205 ;
        RECT -62.045 238.515 -61.715 238.845 ;
        RECT -62.045 237.155 -61.715 237.485 ;
        RECT -62.045 235.795 -61.715 236.125 ;
        RECT -62.045 234.435 -61.715 234.765 ;
        RECT -62.045 233.075 -61.715 233.405 ;
        RECT -62.045 231.715 -61.715 232.045 ;
        RECT -62.045 230.355 -61.715 230.685 ;
        RECT -62.045 228.995 -61.715 229.325 ;
        RECT -62.045 227.635 -61.715 227.965 ;
        RECT -62.045 226.275 -61.715 226.605 ;
        RECT -62.045 224.915 -61.715 225.245 ;
        RECT -62.045 223.555 -61.715 223.885 ;
        RECT -62.045 222.195 -61.715 222.525 ;
        RECT -62.045 220.835 -61.715 221.165 ;
        RECT -62.045 219.475 -61.715 219.805 ;
        RECT -62.045 218.115 -61.715 218.445 ;
        RECT -62.045 216.755 -61.715 217.085 ;
        RECT -62.045 215.395 -61.715 215.725 ;
        RECT -62.045 214.035 -61.715 214.365 ;
        RECT -62.045 212.675 -61.715 213.005 ;
        RECT -62.045 211.315 -61.715 211.645 ;
        RECT -62.045 209.955 -61.715 210.285 ;
        RECT -62.045 208.595 -61.715 208.925 ;
        RECT -62.045 207.235 -61.715 207.565 ;
        RECT -62.045 205.875 -61.715 206.205 ;
        RECT -62.045 204.515 -61.715 204.845 ;
        RECT -62.045 203.155 -61.715 203.485 ;
        RECT -62.045 201.795 -61.715 202.125 ;
        RECT -62.045 200.435 -61.715 200.765 ;
        RECT -62.045 199.075 -61.715 199.405 ;
        RECT -62.045 197.715 -61.715 198.045 ;
        RECT -62.045 196.355 -61.715 196.685 ;
        RECT -62.045 194.995 -61.715 195.325 ;
        RECT -62.045 193.635 -61.715 193.965 ;
        RECT -62.045 192.275 -61.715 192.605 ;
        RECT -62.045 190.915 -61.715 191.245 ;
        RECT -62.045 189.555 -61.715 189.885 ;
        RECT -62.045 188.195 -61.715 188.525 ;
        RECT -62.045 186.835 -61.715 187.165 ;
        RECT -62.045 185.475 -61.715 185.805 ;
        RECT -62.045 184.115 -61.715 184.445 ;
        RECT -62.045 182.755 -61.715 183.085 ;
        RECT -62.045 181.395 -61.715 181.725 ;
        RECT -62.045 180.035 -61.715 180.365 ;
        RECT -62.045 178.675 -61.715 179.005 ;
        RECT -62.045 177.315 -61.715 177.645 ;
        RECT -62.045 175.955 -61.715 176.285 ;
        RECT -62.045 174.595 -61.715 174.925 ;
        RECT -62.045 173.235 -61.715 173.565 ;
        RECT -62.045 171.875 -61.715 172.205 ;
        RECT -62.045 170.515 -61.715 170.845 ;
        RECT -62.045 169.155 -61.715 169.485 ;
        RECT -62.045 167.795 -61.715 168.125 ;
        RECT -62.045 166.435 -61.715 166.765 ;
        RECT -62.045 165.075 -61.715 165.405 ;
        RECT -62.045 163.715 -61.715 164.045 ;
        RECT -62.045 162.355 -61.715 162.685 ;
        RECT -62.045 160.995 -61.715 161.325 ;
        RECT -62.045 159.635 -61.715 159.965 ;
        RECT -62.045 158.275 -61.715 158.605 ;
        RECT -62.045 156.915 -61.715 157.245 ;
        RECT -62.045 155.555 -61.715 155.885 ;
        RECT -62.045 154.195 -61.715 154.525 ;
        RECT -62.045 152.835 -61.715 153.165 ;
        RECT -62.045 151.475 -61.715 151.805 ;
        RECT -62.045 150.115 -61.715 150.445 ;
        RECT -62.045 148.755 -61.715 149.085 ;
        RECT -62.045 147.395 -61.715 147.725 ;
        RECT -62.045 146.035 -61.715 146.365 ;
        RECT -62.045 144.675 -61.715 145.005 ;
        RECT -62.045 143.315 -61.715 143.645 ;
        RECT -62.045 141.955 -61.715 142.285 ;
        RECT -62.045 140.595 -61.715 140.925 ;
        RECT -62.045 139.235 -61.715 139.565 ;
        RECT -62.045 137.875 -61.715 138.205 ;
        RECT -62.045 136.515 -61.715 136.845 ;
        RECT -62.045 135.155 -61.715 135.485 ;
        RECT -62.045 133.795 -61.715 134.125 ;
        RECT -62.045 132.435 -61.715 132.765 ;
        RECT -62.045 131.075 -61.715 131.405 ;
        RECT -62.045 129.715 -61.715 130.045 ;
        RECT -62.045 128.355 -61.715 128.685 ;
        RECT -62.045 126.995 -61.715 127.325 ;
        RECT -62.045 125.635 -61.715 125.965 ;
        RECT -62.045 124.275 -61.715 124.605 ;
        RECT -62.045 122.915 -61.715 123.245 ;
        RECT -62.045 121.555 -61.715 121.885 ;
        RECT -62.045 120.195 -61.715 120.525 ;
        RECT -62.045 118.835 -61.715 119.165 ;
        RECT -62.045 117.475 -61.715 117.805 ;
        RECT -62.045 116.115 -61.715 116.445 ;
        RECT -62.045 114.755 -61.715 115.085 ;
        RECT -62.045 113.395 -61.715 113.725 ;
        RECT -62.045 112.035 -61.715 112.365 ;
        RECT -62.045 110.675 -61.715 111.005 ;
        RECT -62.045 109.315 -61.715 109.645 ;
        RECT -62.045 107.955 -61.715 108.285 ;
        RECT -62.045 106.595 -61.715 106.925 ;
        RECT -62.045 105.235 -61.715 105.565 ;
        RECT -62.045 103.875 -61.715 104.205 ;
        RECT -62.045 102.515 -61.715 102.845 ;
        RECT -62.045 101.155 -61.715 101.485 ;
        RECT -62.045 99.795 -61.715 100.125 ;
        RECT -62.045 98.435 -61.715 98.765 ;
        RECT -62.045 97.075 -61.715 97.405 ;
        RECT -62.045 95.715 -61.715 96.045 ;
        RECT -62.045 94.355 -61.715 94.685 ;
        RECT -62.045 92.995 -61.715 93.325 ;
        RECT -62.045 91.635 -61.715 91.965 ;
        RECT -62.045 90.275 -61.715 90.605 ;
        RECT -62.045 88.915 -61.715 89.245 ;
        RECT -62.045 87.555 -61.715 87.885 ;
        RECT -62.045 86.195 -61.715 86.525 ;
        RECT -62.045 84.835 -61.715 85.165 ;
        RECT -62.045 83.475 -61.715 83.805 ;
        RECT -62.045 82.115 -61.715 82.445 ;
        RECT -62.045 80.755 -61.715 81.085 ;
        RECT -62.045 79.395 -61.715 79.725 ;
        RECT -62.045 78.035 -61.715 78.365 ;
        RECT -62.045 76.675 -61.715 77.005 ;
        RECT -62.045 75.315 -61.715 75.645 ;
        RECT -62.045 73.955 -61.715 74.285 ;
        RECT -62.045 72.595 -61.715 72.925 ;
        RECT -62.045 71.235 -61.715 71.565 ;
        RECT -62.045 69.875 -61.715 70.205 ;
        RECT -62.045 68.515 -61.715 68.845 ;
        RECT -62.045 67.155 -61.715 67.485 ;
        RECT -62.045 65.795 -61.715 66.125 ;
        RECT -62.045 64.435 -61.715 64.765 ;
        RECT -62.045 63.075 -61.715 63.405 ;
        RECT -62.045 61.715 -61.715 62.045 ;
        RECT -62.045 60.355 -61.715 60.685 ;
        RECT -62.045 58.995 -61.715 59.325 ;
        RECT -62.045 57.635 -61.715 57.965 ;
        RECT -62.045 56.275 -61.715 56.605 ;
        RECT -62.045 54.915 -61.715 55.245 ;
        RECT -62.045 53.555 -61.715 53.885 ;
        RECT -62.045 52.195 -61.715 52.525 ;
        RECT -62.045 50.835 -61.715 51.165 ;
        RECT -62.045 49.475 -61.715 49.805 ;
        RECT -62.045 48.115 -61.715 48.445 ;
        RECT -62.045 46.755 -61.715 47.085 ;
        RECT -62.045 45.395 -61.715 45.725 ;
        RECT -62.045 44.035 -61.715 44.365 ;
        RECT -62.045 42.675 -61.715 43.005 ;
        RECT -62.045 41.315 -61.715 41.645 ;
        RECT -62.045 39.955 -61.715 40.285 ;
        RECT -62.045 38.595 -61.715 38.925 ;
        RECT -62.045 37.235 -61.715 37.565 ;
        RECT -62.045 35.875 -61.715 36.205 ;
        RECT -62.045 34.515 -61.715 34.845 ;
        RECT -62.045 33.155 -61.715 33.485 ;
        RECT -62.045 31.795 -61.715 32.125 ;
        RECT -62.045 30.435 -61.715 30.765 ;
        RECT -62.045 29.075 -61.715 29.405 ;
        RECT -62.045 27.715 -61.715 28.045 ;
        RECT -62.045 26.355 -61.715 26.685 ;
        RECT -62.045 24.995 -61.715 25.325 ;
        RECT -62.045 23.635 -61.715 23.965 ;
        RECT -62.045 22.275 -61.715 22.605 ;
        RECT -62.045 20.915 -61.715 21.245 ;
        RECT -62.045 19.555 -61.715 19.885 ;
        RECT -62.045 18.195 -61.715 18.525 ;
        RECT -62.045 16.835 -61.715 17.165 ;
        RECT -62.045 15.475 -61.715 15.805 ;
        RECT -62.045 14.115 -61.715 14.445 ;
        RECT -62.045 12.755 -61.715 13.085 ;
        RECT -62.045 11.395 -61.715 11.725 ;
        RECT -62.045 10.035 -61.715 10.365 ;
        RECT -62.045 8.675 -61.715 9.005 ;
        RECT -62.045 7.315 -61.715 7.645 ;
        RECT -62.045 5.955 -61.715 6.285 ;
        RECT -62.045 4.595 -61.715 4.925 ;
        RECT -62.045 3.235 -61.715 3.565 ;
        RECT -62.045 1.875 -61.715 2.205 ;
        RECT -62.045 0.515 -61.715 0.845 ;
        RECT -62.045 -0.845 -61.715 -0.515 ;
        RECT -62.045 -2.205 -61.715 -1.875 ;
        RECT -62.045 -3.565 -61.715 -3.235 ;
        RECT -62.045 -4.925 -61.715 -4.595 ;
        RECT -62.045 -6.285 -61.715 -5.955 ;
        RECT -62.045 -7.645 -61.715 -7.315 ;
        RECT -62.045 -9.005 -61.715 -8.675 ;
        RECT -62.045 -10.365 -61.715 -10.035 ;
        RECT -62.045 -11.725 -61.715 -11.395 ;
        RECT -62.045 -13.085 -61.715 -12.755 ;
        RECT -62.045 -14.445 -61.715 -14.115 ;
        RECT -62.045 -15.805 -61.715 -15.475 ;
        RECT -62.045 -17.165 -61.715 -16.835 ;
        RECT -62.045 -18.525 -61.715 -18.195 ;
        RECT -62.045 -19.885 -61.715 -19.555 ;
        RECT -62.045 -21.245 -61.715 -20.915 ;
        RECT -62.045 -22.605 -61.715 -22.275 ;
        RECT -62.045 -23.965 -61.715 -23.635 ;
        RECT -62.045 -25.325 -61.715 -24.995 ;
        RECT -62.045 -26.685 -61.715 -26.355 ;
        RECT -62.045 -28.045 -61.715 -27.715 ;
        RECT -62.045 -29.405 -61.715 -29.075 ;
        RECT -62.045 -30.765 -61.715 -30.435 ;
        RECT -62.045 -32.125 -61.715 -31.795 ;
        RECT -62.045 -33.485 -61.715 -33.155 ;
        RECT -62.045 -34.845 -61.715 -34.515 ;
        RECT -62.045 -36.205 -61.715 -35.875 ;
        RECT -62.045 -37.565 -61.715 -37.235 ;
        RECT -62.045 -38.925 -61.715 -38.595 ;
        RECT -62.045 -40.285 -61.715 -39.955 ;
        RECT -62.045 -41.645 -61.715 -41.315 ;
        RECT -62.045 -43.005 -61.715 -42.675 ;
        RECT -62.045 -44.365 -61.715 -44.035 ;
        RECT -62.045 -45.725 -61.715 -45.395 ;
        RECT -62.045 -47.085 -61.715 -46.755 ;
        RECT -62.045 -48.445 -61.715 -48.115 ;
        RECT -62.045 -49.805 -61.715 -49.475 ;
        RECT -62.045 -51.165 -61.715 -50.835 ;
        RECT -62.045 -52.525 -61.715 -52.195 ;
        RECT -62.045 -53.885 -61.715 -53.555 ;
        RECT -62.045 -55.245 -61.715 -54.915 ;
        RECT -62.045 -56.605 -61.715 -56.275 ;
        RECT -62.045 -57.965 -61.715 -57.635 ;
        RECT -62.045 -59.325 -61.715 -58.995 ;
        RECT -62.045 -60.685 -61.715 -60.355 ;
        RECT -62.045 -62.045 -61.715 -61.715 ;
        RECT -62.045 -63.405 -61.715 -63.075 ;
        RECT -62.045 -64.765 -61.715 -64.435 ;
        RECT -62.045 -66.125 -61.715 -65.795 ;
        RECT -62.045 -67.485 -61.715 -67.155 ;
        RECT -62.045 -68.845 -61.715 -68.515 ;
        RECT -62.045 -70.205 -61.715 -69.875 ;
        RECT -62.045 -71.565 -61.715 -71.235 ;
        RECT -62.045 -72.925 -61.715 -72.595 ;
        RECT -62.045 -74.285 -61.715 -73.955 ;
        RECT -62.045 -75.645 -61.715 -75.315 ;
        RECT -62.045 -77.005 -61.715 -76.675 ;
        RECT -62.045 -78.365 -61.715 -78.035 ;
        RECT -62.045 -79.725 -61.715 -79.395 ;
        RECT -62.045 -81.085 -61.715 -80.755 ;
        RECT -62.045 -82.445 -61.715 -82.115 ;
        RECT -62.045 -83.805 -61.715 -83.475 ;
        RECT -62.045 -85.165 -61.715 -84.835 ;
        RECT -62.045 -86.525 -61.715 -86.195 ;
        RECT -62.045 -87.885 -61.715 -87.555 ;
        RECT -62.045 -89.245 -61.715 -88.915 ;
        RECT -62.045 -90.605 -61.715 -90.275 ;
        RECT -62.045 -91.965 -61.715 -91.635 ;
        RECT -62.045 -93.325 -61.715 -92.995 ;
        RECT -62.045 -94.685 -61.715 -94.355 ;
        RECT -62.045 -96.045 -61.715 -95.715 ;
        RECT -62.045 -97.405 -61.715 -97.075 ;
        RECT -62.045 -98.765 -61.715 -98.435 ;
        RECT -62.045 -100.125 -61.715 -99.795 ;
        RECT -62.045 -101.485 -61.715 -101.155 ;
        RECT -62.045 -102.845 -61.715 -102.515 ;
        RECT -62.045 -104.205 -61.715 -103.875 ;
        RECT -62.045 -105.565 -61.715 -105.235 ;
        RECT -62.045 -106.925 -61.715 -106.595 ;
        RECT -62.045 -108.285 -61.715 -107.955 ;
        RECT -62.045 -109.645 -61.715 -109.315 ;
        RECT -62.045 -111.005 -61.715 -110.675 ;
        RECT -62.045 -112.365 -61.715 -112.035 ;
        RECT -62.045 -113.725 -61.715 -113.395 ;
        RECT -62.045 -115.085 -61.715 -114.755 ;
        RECT -62.045 -116.445 -61.715 -116.115 ;
        RECT -62.045 -117.805 -61.715 -117.475 ;
        RECT -62.045 -119.165 -61.715 -118.835 ;
        RECT -62.045 -120.525 -61.715 -120.195 ;
        RECT -62.045 -121.885 -61.715 -121.555 ;
        RECT -62.045 -123.245 -61.715 -122.915 ;
        RECT -62.045 -124.605 -61.715 -124.275 ;
        RECT -62.045 -128.685 -61.715 -128.355 ;
        RECT -62.045 -130.045 -61.715 -129.715 ;
        RECT -62.045 -132.765 -61.715 -132.435 ;
        RECT -62.045 -134.125 -61.715 -133.795 ;
        RECT -62.045 -135.485 -61.715 -135.155 ;
        RECT -62.045 -136.845 -61.715 -136.515 ;
        RECT -62.045 -138.205 -61.715 -137.875 ;
        RECT -62.045 -139.39 -61.715 -139.06 ;
        RECT -62.045 -140.925 -61.715 -140.595 ;
        RECT -62.045 -142.285 -61.715 -141.955 ;
        RECT -62.045 -145.005 -61.715 -144.675 ;
        RECT -62.045 -146.365 -61.715 -146.035 ;
        RECT -62.045 -148.03 -61.715 -147.7 ;
        RECT -62.045 -149.085 -61.715 -148.755 ;
        RECT -62.045 -150.445 -61.715 -150.115 ;
        RECT -62.045 -153.165 -61.715 -152.835 ;
        RECT -62.045 -154.525 -61.715 -154.195 ;
        RECT -62.045 -155.885 -61.715 -155.555 ;
        RECT -62.045 -157.245 -61.715 -156.915 ;
        RECT -62.045 -158.605 -61.715 -158.275 ;
        RECT -62.045 -159.965 -61.715 -159.635 ;
        RECT -62.045 -161.325 -61.715 -160.995 ;
        RECT -62.045 -162.685 -61.715 -162.355 ;
        RECT -62.045 -164.045 -61.715 -163.715 ;
        RECT -62.045 -165.405 -61.715 -165.075 ;
        RECT -62.045 -166.765 -61.715 -166.435 ;
        RECT -62.045 -168.125 -61.715 -167.795 ;
        RECT -62.045 -169.485 -61.715 -169.155 ;
        RECT -62.045 -170.845 -61.715 -170.515 ;
        RECT -62.045 -172.205 -61.715 -171.875 ;
        RECT -62.045 -173.565 -61.715 -173.235 ;
        RECT -62.045 -174.925 -61.715 -174.595 ;
        RECT -62.045 -176.285 -61.715 -175.955 ;
        RECT -62.045 -177.645 -61.715 -177.315 ;
        RECT -62.045 -179.005 -61.715 -178.675 ;
        RECT -62.045 -180.365 -61.715 -180.035 ;
        RECT -62.045 -181.725 -61.715 -181.395 ;
        RECT -62.045 -183.085 -61.715 -182.755 ;
        RECT -62.045 -184.445 -61.715 -184.115 ;
        RECT -62.045 -185.805 -61.715 -185.475 ;
        RECT -62.045 -187.165 -61.715 -186.835 ;
        RECT -62.045 -188.525 -61.715 -188.195 ;
        RECT -62.045 -189.885 -61.715 -189.555 ;
        RECT -62.045 -191.245 -61.715 -190.915 ;
        RECT -62.045 -192.605 -61.715 -192.275 ;
        RECT -62.045 -193.965 -61.715 -193.635 ;
        RECT -62.045 -195.325 -61.715 -194.995 ;
        RECT -62.045 -196.685 -61.715 -196.355 ;
        RECT -62.045 -198.045 -61.715 -197.715 ;
        RECT -62.045 -199.405 -61.715 -199.075 ;
        RECT -62.045 -200.765 -61.715 -200.435 ;
        RECT -62.045 -202.125 -61.715 -201.795 ;
        RECT -62.045 -203.485 -61.715 -203.155 ;
        RECT -62.045 -204.845 -61.715 -204.515 ;
        RECT -62.045 -206.205 -61.715 -205.875 ;
        RECT -62.045 -207.565 -61.715 -207.235 ;
        RECT -62.045 -208.925 -61.715 -208.595 ;
        RECT -62.045 -210.285 -61.715 -209.955 ;
        RECT -62.045 -211.645 -61.715 -211.315 ;
        RECT -62.045 -213.005 -61.715 -212.675 ;
        RECT -62.045 -214.365 -61.715 -214.035 ;
        RECT -62.045 -215.725 -61.715 -215.395 ;
        RECT -62.045 -217.085 -61.715 -216.755 ;
        RECT -62.045 -218.445 -61.715 -218.115 ;
        RECT -62.045 -219.805 -61.715 -219.475 ;
        RECT -62.045 -221.165 -61.715 -220.835 ;
        RECT -62.045 -222.525 -61.715 -222.195 ;
        RECT -62.045 -223.885 -61.715 -223.555 ;
        RECT -62.045 -225.245 -61.715 -224.915 ;
        RECT -62.045 -227.965 -61.715 -227.635 ;
        RECT -62.045 -230.685 -61.715 -230.355 ;
        RECT -62.045 -232.045 -61.715 -231.715 ;
        RECT -62.045 -233.225 -61.715 -232.895 ;
        RECT -62.045 -234.765 -61.715 -234.435 ;
        RECT -62.045 -236.125 -61.715 -235.795 ;
        RECT -62.045 -237.485 -61.715 -237.155 ;
        RECT -62.045 -238.845 -61.715 -238.515 ;
        RECT -62.045 -241.09 -61.715 -239.96 ;
        RECT -62.04 -241.205 -61.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 -138.205 -60.355 -137.875 ;
        RECT -60.685 -139.39 -60.355 -139.06 ;
        RECT -60.685 -140.925 -60.355 -140.595 ;
        RECT -60.685 -142.285 -60.355 -141.955 ;
        RECT -60.685 -145.005 -60.355 -144.675 ;
        RECT -60.685 -146.365 -60.355 -146.035 ;
        RECT -60.685 -148.03 -60.355 -147.7 ;
        RECT -60.685 -149.085 -60.355 -148.755 ;
        RECT -60.685 -150.445 -60.355 -150.115 ;
        RECT -60.68 -151.8 -60.36 245.285 ;
        RECT -60.685 244.04 -60.355 245.17 ;
        RECT -60.685 242.595 -60.355 242.925 ;
        RECT -60.685 241.235 -60.355 241.565 ;
        RECT -60.685 239.875 -60.355 240.205 ;
        RECT -60.685 238.515 -60.355 238.845 ;
        RECT -60.685 237.155 -60.355 237.485 ;
        RECT -60.685 235.795 -60.355 236.125 ;
        RECT -60.685 234.435 -60.355 234.765 ;
        RECT -60.685 233.075 -60.355 233.405 ;
        RECT -60.685 231.715 -60.355 232.045 ;
        RECT -60.685 230.355 -60.355 230.685 ;
        RECT -60.685 228.995 -60.355 229.325 ;
        RECT -60.685 227.635 -60.355 227.965 ;
        RECT -60.685 226.275 -60.355 226.605 ;
        RECT -60.685 224.915 -60.355 225.245 ;
        RECT -60.685 223.555 -60.355 223.885 ;
        RECT -60.685 222.195 -60.355 222.525 ;
        RECT -60.685 220.835 -60.355 221.165 ;
        RECT -60.685 219.475 -60.355 219.805 ;
        RECT -60.685 218.115 -60.355 218.445 ;
        RECT -60.685 216.755 -60.355 217.085 ;
        RECT -60.685 215.395 -60.355 215.725 ;
        RECT -60.685 214.035 -60.355 214.365 ;
        RECT -60.685 212.675 -60.355 213.005 ;
        RECT -60.685 211.315 -60.355 211.645 ;
        RECT -60.685 209.955 -60.355 210.285 ;
        RECT -60.685 208.595 -60.355 208.925 ;
        RECT -60.685 207.235 -60.355 207.565 ;
        RECT -60.685 205.875 -60.355 206.205 ;
        RECT -60.685 204.515 -60.355 204.845 ;
        RECT -60.685 203.155 -60.355 203.485 ;
        RECT -60.685 201.795 -60.355 202.125 ;
        RECT -60.685 200.435 -60.355 200.765 ;
        RECT -60.685 199.075 -60.355 199.405 ;
        RECT -60.685 197.715 -60.355 198.045 ;
        RECT -60.685 196.355 -60.355 196.685 ;
        RECT -60.685 194.995 -60.355 195.325 ;
        RECT -60.685 193.635 -60.355 193.965 ;
        RECT -60.685 192.275 -60.355 192.605 ;
        RECT -60.685 190.915 -60.355 191.245 ;
        RECT -60.685 189.555 -60.355 189.885 ;
        RECT -60.685 188.195 -60.355 188.525 ;
        RECT -60.685 186.835 -60.355 187.165 ;
        RECT -60.685 185.475 -60.355 185.805 ;
        RECT -60.685 184.115 -60.355 184.445 ;
        RECT -60.685 182.755 -60.355 183.085 ;
        RECT -60.685 181.395 -60.355 181.725 ;
        RECT -60.685 180.035 -60.355 180.365 ;
        RECT -60.685 178.675 -60.355 179.005 ;
        RECT -60.685 177.315 -60.355 177.645 ;
        RECT -60.685 175.955 -60.355 176.285 ;
        RECT -60.685 174.595 -60.355 174.925 ;
        RECT -60.685 173.235 -60.355 173.565 ;
        RECT -60.685 171.875 -60.355 172.205 ;
        RECT -60.685 170.515 -60.355 170.845 ;
        RECT -60.685 169.155 -60.355 169.485 ;
        RECT -60.685 167.795 -60.355 168.125 ;
        RECT -60.685 166.435 -60.355 166.765 ;
        RECT -60.685 165.075 -60.355 165.405 ;
        RECT -60.685 163.715 -60.355 164.045 ;
        RECT -60.685 162.355 -60.355 162.685 ;
        RECT -60.685 160.995 -60.355 161.325 ;
        RECT -60.685 159.635 -60.355 159.965 ;
        RECT -60.685 158.275 -60.355 158.605 ;
        RECT -60.685 156.915 -60.355 157.245 ;
        RECT -60.685 155.555 -60.355 155.885 ;
        RECT -60.685 154.195 -60.355 154.525 ;
        RECT -60.685 152.835 -60.355 153.165 ;
        RECT -60.685 151.475 -60.355 151.805 ;
        RECT -60.685 150.115 -60.355 150.445 ;
        RECT -60.685 148.755 -60.355 149.085 ;
        RECT -60.685 147.395 -60.355 147.725 ;
        RECT -60.685 146.035 -60.355 146.365 ;
        RECT -60.685 144.675 -60.355 145.005 ;
        RECT -60.685 143.315 -60.355 143.645 ;
        RECT -60.685 141.955 -60.355 142.285 ;
        RECT -60.685 140.595 -60.355 140.925 ;
        RECT -60.685 139.235 -60.355 139.565 ;
        RECT -60.685 137.225 -60.355 137.555 ;
        RECT -60.685 135.175 -60.355 135.505 ;
        RECT -60.685 132.815 -60.355 133.145 ;
        RECT -60.685 131.665 -60.355 131.995 ;
        RECT -60.685 129.655 -60.355 129.985 ;
        RECT -60.685 128.505 -60.355 128.835 ;
        RECT -60.685 126.495 -60.355 126.825 ;
        RECT -60.685 125.345 -60.355 125.675 ;
        RECT -60.685 123.335 -60.355 123.665 ;
        RECT -60.685 122.185 -60.355 122.515 ;
        RECT -60.685 120.175 -60.355 120.505 ;
        RECT -60.685 119.025 -60.355 119.355 ;
        RECT -60.685 117.185 -60.355 117.515 ;
        RECT -60.685 115.865 -60.355 116.195 ;
        RECT -60.685 113.855 -60.355 114.185 ;
        RECT -60.685 112.705 -60.355 113.035 ;
        RECT -60.685 110.695 -60.355 111.025 ;
        RECT -60.685 109.545 -60.355 109.875 ;
        RECT -60.685 107.535 -60.355 107.865 ;
        RECT -60.685 106.385 -60.355 106.715 ;
        RECT -60.685 104.375 -60.355 104.705 ;
        RECT -60.685 103.225 -60.355 103.555 ;
        RECT -60.685 100.865 -60.355 101.195 ;
        RECT -60.685 98.81 -60.355 99.14 ;
        RECT -60.685 97.075 -60.355 97.405 ;
        RECT -60.685 95.715 -60.355 96.045 ;
        RECT -60.685 94.355 -60.355 94.685 ;
        RECT -60.685 92.995 -60.355 93.325 ;
        RECT -60.685 91.635 -60.355 91.965 ;
        RECT -60.685 90.275 -60.355 90.605 ;
        RECT -60.685 88.915 -60.355 89.245 ;
        RECT -60.685 87.555 -60.355 87.885 ;
        RECT -60.685 86.195 -60.355 86.525 ;
        RECT -60.685 84.835 -60.355 85.165 ;
        RECT -60.685 83.475 -60.355 83.805 ;
        RECT -60.685 82.115 -60.355 82.445 ;
        RECT -60.685 80.755 -60.355 81.085 ;
        RECT -60.685 79.395 -60.355 79.725 ;
        RECT -60.685 78.035 -60.355 78.365 ;
        RECT -60.685 76.675 -60.355 77.005 ;
        RECT -60.685 75.315 -60.355 75.645 ;
        RECT -60.685 73.955 -60.355 74.285 ;
        RECT -60.685 72.595 -60.355 72.925 ;
        RECT -60.685 71.235 -60.355 71.565 ;
        RECT -60.685 69.875 -60.355 70.205 ;
        RECT -60.685 68.515 -60.355 68.845 ;
        RECT -60.685 67.155 -60.355 67.485 ;
        RECT -60.685 65.795 -60.355 66.125 ;
        RECT -60.685 64.435 -60.355 64.765 ;
        RECT -60.685 63.075 -60.355 63.405 ;
        RECT -60.685 61.715 -60.355 62.045 ;
        RECT -60.685 60.355 -60.355 60.685 ;
        RECT -60.685 58.995 -60.355 59.325 ;
        RECT -60.685 57.635 -60.355 57.965 ;
        RECT -60.685 56.275 -60.355 56.605 ;
        RECT -60.685 54.915 -60.355 55.245 ;
        RECT -60.685 53.555 -60.355 53.885 ;
        RECT -60.685 52.195 -60.355 52.525 ;
        RECT -60.685 50.835 -60.355 51.165 ;
        RECT -60.685 49.475 -60.355 49.805 ;
        RECT -60.685 48.115 -60.355 48.445 ;
        RECT -60.685 46.755 -60.355 47.085 ;
        RECT -60.685 45.395 -60.355 45.725 ;
        RECT -60.685 44.035 -60.355 44.365 ;
        RECT -60.685 42.675 -60.355 43.005 ;
        RECT -60.685 41.315 -60.355 41.645 ;
        RECT -60.685 39.955 -60.355 40.285 ;
        RECT -60.685 38.595 -60.355 38.925 ;
        RECT -60.685 37.235 -60.355 37.565 ;
        RECT -60.685 35.875 -60.355 36.205 ;
        RECT -60.685 34.515 -60.355 34.845 ;
        RECT -60.685 33.155 -60.355 33.485 ;
        RECT -60.685 31.795 -60.355 32.125 ;
        RECT -60.685 30.435 -60.355 30.765 ;
        RECT -60.685 29.075 -60.355 29.405 ;
        RECT -60.685 27.715 -60.355 28.045 ;
        RECT -60.685 26.355 -60.355 26.685 ;
        RECT -60.685 24.995 -60.355 25.325 ;
        RECT -60.685 23.635 -60.355 23.965 ;
        RECT -60.685 22.275 -60.355 22.605 ;
        RECT -60.685 20.915 -60.355 21.245 ;
        RECT -60.685 19.555 -60.355 19.885 ;
        RECT -60.685 18.195 -60.355 18.525 ;
        RECT -60.685 16.835 -60.355 17.165 ;
        RECT -60.685 15.475 -60.355 15.805 ;
        RECT -60.685 14.115 -60.355 14.445 ;
        RECT -60.685 12.755 -60.355 13.085 ;
        RECT -60.685 11.395 -60.355 11.725 ;
        RECT -60.685 10.035 -60.355 10.365 ;
        RECT -60.685 8.675 -60.355 9.005 ;
        RECT -60.685 7.315 -60.355 7.645 ;
        RECT -60.685 5.955 -60.355 6.285 ;
        RECT -60.685 4.595 -60.355 4.925 ;
        RECT -60.685 3.235 -60.355 3.565 ;
        RECT -60.685 1.875 -60.355 2.205 ;
        RECT -60.685 0.515 -60.355 0.845 ;
        RECT -60.685 -0.845 -60.355 -0.515 ;
        RECT -60.685 -2.205 -60.355 -1.875 ;
        RECT -60.685 -3.565 -60.355 -3.235 ;
        RECT -60.685 -4.925 -60.355 -4.595 ;
        RECT -60.685 -6.285 -60.355 -5.955 ;
        RECT -60.685 -7.645 -60.355 -7.315 ;
        RECT -60.685 -9.005 -60.355 -8.675 ;
        RECT -60.685 -10.365 -60.355 -10.035 ;
        RECT -60.685 -11.725 -60.355 -11.395 ;
        RECT -60.685 -13.085 -60.355 -12.755 ;
        RECT -60.685 -14.445 -60.355 -14.115 ;
        RECT -60.685 -15.805 -60.355 -15.475 ;
        RECT -60.685 -17.165 -60.355 -16.835 ;
        RECT -60.685 -18.525 -60.355 -18.195 ;
        RECT -60.685 -19.885 -60.355 -19.555 ;
        RECT -60.685 -21.245 -60.355 -20.915 ;
        RECT -60.685 -22.605 -60.355 -22.275 ;
        RECT -60.685 -23.965 -60.355 -23.635 ;
        RECT -60.685 -25.325 -60.355 -24.995 ;
        RECT -60.685 -26.685 -60.355 -26.355 ;
        RECT -60.685 -28.045 -60.355 -27.715 ;
        RECT -60.685 -29.405 -60.355 -29.075 ;
        RECT -60.685 -30.765 -60.355 -30.435 ;
        RECT -60.685 -32.125 -60.355 -31.795 ;
        RECT -60.685 -33.485 -60.355 -33.155 ;
        RECT -60.685 -34.845 -60.355 -34.515 ;
        RECT -60.685 -36.205 -60.355 -35.875 ;
        RECT -60.685 -37.565 -60.355 -37.235 ;
        RECT -60.685 -38.925 -60.355 -38.595 ;
        RECT -60.685 -40.285 -60.355 -39.955 ;
        RECT -60.685 -41.645 -60.355 -41.315 ;
        RECT -60.685 -43.005 -60.355 -42.675 ;
        RECT -60.685 -44.365 -60.355 -44.035 ;
        RECT -60.685 -45.725 -60.355 -45.395 ;
        RECT -60.685 -47.085 -60.355 -46.755 ;
        RECT -60.685 -48.445 -60.355 -48.115 ;
        RECT -60.685 -49.805 -60.355 -49.475 ;
        RECT -60.685 -51.165 -60.355 -50.835 ;
        RECT -60.685 -52.525 -60.355 -52.195 ;
        RECT -60.685 -53.885 -60.355 -53.555 ;
        RECT -60.685 -55.245 -60.355 -54.915 ;
        RECT -60.685 -56.605 -60.355 -56.275 ;
        RECT -60.685 -57.965 -60.355 -57.635 ;
        RECT -60.685 -59.325 -60.355 -58.995 ;
        RECT -60.685 -60.685 -60.355 -60.355 ;
        RECT -60.685 -62.045 -60.355 -61.715 ;
        RECT -60.685 -63.405 -60.355 -63.075 ;
        RECT -60.685 -64.765 -60.355 -64.435 ;
        RECT -60.685 -66.125 -60.355 -65.795 ;
        RECT -60.685 -67.485 -60.355 -67.155 ;
        RECT -60.685 -68.845 -60.355 -68.515 ;
        RECT -60.685 -70.205 -60.355 -69.875 ;
        RECT -60.685 -71.565 -60.355 -71.235 ;
        RECT -60.685 -72.925 -60.355 -72.595 ;
        RECT -60.685 -74.285 -60.355 -73.955 ;
        RECT -60.685 -75.645 -60.355 -75.315 ;
        RECT -60.685 -77.005 -60.355 -76.675 ;
        RECT -60.685 -78.365 -60.355 -78.035 ;
        RECT -60.685 -79.725 -60.355 -79.395 ;
        RECT -60.685 -81.085 -60.355 -80.755 ;
        RECT -60.685 -82.445 -60.355 -82.115 ;
        RECT -60.685 -83.805 -60.355 -83.475 ;
        RECT -60.685 -85.165 -60.355 -84.835 ;
        RECT -60.685 -86.525 -60.355 -86.195 ;
        RECT -60.685 -87.885 -60.355 -87.555 ;
        RECT -60.685 -89.245 -60.355 -88.915 ;
        RECT -60.685 -90.605 -60.355 -90.275 ;
        RECT -60.685 -91.965 -60.355 -91.635 ;
        RECT -60.685 -93.325 -60.355 -92.995 ;
        RECT -60.685 -94.685 -60.355 -94.355 ;
        RECT -60.685 -96.045 -60.355 -95.715 ;
        RECT -60.685 -97.405 -60.355 -97.075 ;
        RECT -60.685 -98.765 -60.355 -98.435 ;
        RECT -60.685 -100.125 -60.355 -99.795 ;
        RECT -60.685 -101.485 -60.355 -101.155 ;
        RECT -60.685 -102.845 -60.355 -102.515 ;
        RECT -60.685 -104.205 -60.355 -103.875 ;
        RECT -60.685 -105.565 -60.355 -105.235 ;
        RECT -60.685 -106.925 -60.355 -106.595 ;
        RECT -60.685 -108.285 -60.355 -107.955 ;
        RECT -60.685 -109.645 -60.355 -109.315 ;
        RECT -60.685 -111.005 -60.355 -110.675 ;
        RECT -60.685 -112.365 -60.355 -112.035 ;
        RECT -60.685 -113.725 -60.355 -113.395 ;
        RECT -60.685 -115.085 -60.355 -114.755 ;
        RECT -60.685 -116.445 -60.355 -116.115 ;
        RECT -60.685 -117.805 -60.355 -117.475 ;
        RECT -60.685 -119.165 -60.355 -118.835 ;
        RECT -60.685 -120.525 -60.355 -120.195 ;
        RECT -60.685 -121.885 -60.355 -121.555 ;
        RECT -60.685 -123.245 -60.355 -122.915 ;
        RECT -60.685 -124.605 -60.355 -124.275 ;
        RECT -60.685 -128.685 -60.355 -128.355 ;
        RECT -60.685 -130.045 -60.355 -129.715 ;
        RECT -60.685 -132.765 -60.355 -132.435 ;
        RECT -60.685 -134.125 -60.355 -133.795 ;
        RECT -60.685 -135.485 -60.355 -135.155 ;
        RECT -60.685 -136.845 -60.355 -136.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.485 244.04 -67.155 245.17 ;
        RECT -67.485 242.595 -67.155 242.925 ;
        RECT -67.485 241.235 -67.155 241.565 ;
        RECT -67.485 239.875 -67.155 240.205 ;
        RECT -67.485 238.515 -67.155 238.845 ;
        RECT -67.485 237.155 -67.155 237.485 ;
        RECT -67.485 235.795 -67.155 236.125 ;
        RECT -67.485 234.435 -67.155 234.765 ;
        RECT -67.485 233.075 -67.155 233.405 ;
        RECT -67.485 231.715 -67.155 232.045 ;
        RECT -67.485 230.355 -67.155 230.685 ;
        RECT -67.485 228.995 -67.155 229.325 ;
        RECT -67.485 227.635 -67.155 227.965 ;
        RECT -67.485 226.275 -67.155 226.605 ;
        RECT -67.485 224.915 -67.155 225.245 ;
        RECT -67.485 223.555 -67.155 223.885 ;
        RECT -67.485 222.195 -67.155 222.525 ;
        RECT -67.485 220.835 -67.155 221.165 ;
        RECT -67.485 219.475 -67.155 219.805 ;
        RECT -67.485 218.115 -67.155 218.445 ;
        RECT -67.485 216.755 -67.155 217.085 ;
        RECT -67.485 215.395 -67.155 215.725 ;
        RECT -67.485 214.035 -67.155 214.365 ;
        RECT -67.485 212.675 -67.155 213.005 ;
        RECT -67.485 211.315 -67.155 211.645 ;
        RECT -67.485 209.955 -67.155 210.285 ;
        RECT -67.485 208.595 -67.155 208.925 ;
        RECT -67.485 207.235 -67.155 207.565 ;
        RECT -67.485 205.875 -67.155 206.205 ;
        RECT -67.485 204.515 -67.155 204.845 ;
        RECT -67.485 203.155 -67.155 203.485 ;
        RECT -67.485 201.795 -67.155 202.125 ;
        RECT -67.485 200.435 -67.155 200.765 ;
        RECT -67.485 199.075 -67.155 199.405 ;
        RECT -67.485 197.715 -67.155 198.045 ;
        RECT -67.485 196.355 -67.155 196.685 ;
        RECT -67.485 194.995 -67.155 195.325 ;
        RECT -67.485 193.635 -67.155 193.965 ;
        RECT -67.485 192.275 -67.155 192.605 ;
        RECT -67.485 190.915 -67.155 191.245 ;
        RECT -67.485 189.555 -67.155 189.885 ;
        RECT -67.485 188.195 -67.155 188.525 ;
        RECT -67.485 186.835 -67.155 187.165 ;
        RECT -67.485 185.475 -67.155 185.805 ;
        RECT -67.485 184.115 -67.155 184.445 ;
        RECT -67.485 182.755 -67.155 183.085 ;
        RECT -67.485 181.395 -67.155 181.725 ;
        RECT -67.485 180.035 -67.155 180.365 ;
        RECT -67.485 178.675 -67.155 179.005 ;
        RECT -67.485 177.315 -67.155 177.645 ;
        RECT -67.485 175.955 -67.155 176.285 ;
        RECT -67.485 174.595 -67.155 174.925 ;
        RECT -67.485 173.235 -67.155 173.565 ;
        RECT -67.485 171.875 -67.155 172.205 ;
        RECT -67.485 170.515 -67.155 170.845 ;
        RECT -67.485 169.155 -67.155 169.485 ;
        RECT -67.485 167.795 -67.155 168.125 ;
        RECT -67.485 166.435 -67.155 166.765 ;
        RECT -67.485 165.075 -67.155 165.405 ;
        RECT -67.485 163.715 -67.155 164.045 ;
        RECT -67.485 162.355 -67.155 162.685 ;
        RECT -67.485 160.995 -67.155 161.325 ;
        RECT -67.485 159.635 -67.155 159.965 ;
        RECT -67.485 158.275 -67.155 158.605 ;
        RECT -67.485 156.915 -67.155 157.245 ;
        RECT -67.485 155.555 -67.155 155.885 ;
        RECT -67.485 154.195 -67.155 154.525 ;
        RECT -67.485 152.835 -67.155 153.165 ;
        RECT -67.485 151.475 -67.155 151.805 ;
        RECT -67.485 150.115 -67.155 150.445 ;
        RECT -67.485 148.755 -67.155 149.085 ;
        RECT -67.485 147.395 -67.155 147.725 ;
        RECT -67.485 146.035 -67.155 146.365 ;
        RECT -67.485 144.675 -67.155 145.005 ;
        RECT -67.485 143.315 -67.155 143.645 ;
        RECT -67.485 141.955 -67.155 142.285 ;
        RECT -67.485 140.595 -67.155 140.925 ;
        RECT -67.485 139.235 -67.155 139.565 ;
        RECT -67.485 137.875 -67.155 138.205 ;
        RECT -67.485 136.515 -67.155 136.845 ;
        RECT -67.485 135.155 -67.155 135.485 ;
        RECT -67.485 133.795 -67.155 134.125 ;
        RECT -67.485 132.435 -67.155 132.765 ;
        RECT -67.485 131.075 -67.155 131.405 ;
        RECT -67.485 129.715 -67.155 130.045 ;
        RECT -67.485 128.355 -67.155 128.685 ;
        RECT -67.485 126.995 -67.155 127.325 ;
        RECT -67.485 125.635 -67.155 125.965 ;
        RECT -67.485 124.275 -67.155 124.605 ;
        RECT -67.485 122.915 -67.155 123.245 ;
        RECT -67.485 121.555 -67.155 121.885 ;
        RECT -67.485 120.195 -67.155 120.525 ;
        RECT -67.485 118.835 -67.155 119.165 ;
        RECT -67.485 117.475 -67.155 117.805 ;
        RECT -67.485 116.115 -67.155 116.445 ;
        RECT -67.485 114.755 -67.155 115.085 ;
        RECT -67.485 113.395 -67.155 113.725 ;
        RECT -67.485 112.035 -67.155 112.365 ;
        RECT -67.485 110.675 -67.155 111.005 ;
        RECT -67.485 109.315 -67.155 109.645 ;
        RECT -67.485 107.955 -67.155 108.285 ;
        RECT -67.485 106.595 -67.155 106.925 ;
        RECT -67.485 105.235 -67.155 105.565 ;
        RECT -67.485 103.875 -67.155 104.205 ;
        RECT -67.485 102.515 -67.155 102.845 ;
        RECT -67.485 101.155 -67.155 101.485 ;
        RECT -67.485 99.795 -67.155 100.125 ;
        RECT -67.485 98.435 -67.155 98.765 ;
        RECT -67.485 97.075 -67.155 97.405 ;
        RECT -67.485 95.715 -67.155 96.045 ;
        RECT -67.485 94.355 -67.155 94.685 ;
        RECT -67.485 92.995 -67.155 93.325 ;
        RECT -67.485 91.635 -67.155 91.965 ;
        RECT -67.485 90.275 -67.155 90.605 ;
        RECT -67.485 88.915 -67.155 89.245 ;
        RECT -67.485 87.555 -67.155 87.885 ;
        RECT -67.485 86.195 -67.155 86.525 ;
        RECT -67.485 84.835 -67.155 85.165 ;
        RECT -67.485 83.475 -67.155 83.805 ;
        RECT -67.485 82.115 -67.155 82.445 ;
        RECT -67.485 80.755 -67.155 81.085 ;
        RECT -67.485 79.395 -67.155 79.725 ;
        RECT -67.485 78.035 -67.155 78.365 ;
        RECT -67.485 76.675 -67.155 77.005 ;
        RECT -67.485 75.315 -67.155 75.645 ;
        RECT -67.485 73.955 -67.155 74.285 ;
        RECT -67.485 72.595 -67.155 72.925 ;
        RECT -67.485 71.235 -67.155 71.565 ;
        RECT -67.485 69.875 -67.155 70.205 ;
        RECT -67.485 68.515 -67.155 68.845 ;
        RECT -67.485 67.155 -67.155 67.485 ;
        RECT -67.485 65.795 -67.155 66.125 ;
        RECT -67.485 64.435 -67.155 64.765 ;
        RECT -67.485 63.075 -67.155 63.405 ;
        RECT -67.485 61.715 -67.155 62.045 ;
        RECT -67.485 60.355 -67.155 60.685 ;
        RECT -67.485 58.995 -67.155 59.325 ;
        RECT -67.485 57.635 -67.155 57.965 ;
        RECT -67.485 56.275 -67.155 56.605 ;
        RECT -67.485 54.915 -67.155 55.245 ;
        RECT -67.485 53.555 -67.155 53.885 ;
        RECT -67.485 52.195 -67.155 52.525 ;
        RECT -67.485 50.835 -67.155 51.165 ;
        RECT -67.485 49.475 -67.155 49.805 ;
        RECT -67.485 48.115 -67.155 48.445 ;
        RECT -67.485 46.755 -67.155 47.085 ;
        RECT -67.485 45.395 -67.155 45.725 ;
        RECT -67.485 44.035 -67.155 44.365 ;
        RECT -67.485 42.675 -67.155 43.005 ;
        RECT -67.485 41.315 -67.155 41.645 ;
        RECT -67.485 39.955 -67.155 40.285 ;
        RECT -67.485 38.595 -67.155 38.925 ;
        RECT -67.485 37.235 -67.155 37.565 ;
        RECT -67.485 35.875 -67.155 36.205 ;
        RECT -67.485 34.515 -67.155 34.845 ;
        RECT -67.485 33.155 -67.155 33.485 ;
        RECT -67.485 31.795 -67.155 32.125 ;
        RECT -67.485 30.435 -67.155 30.765 ;
        RECT -67.485 29.075 -67.155 29.405 ;
        RECT -67.485 27.715 -67.155 28.045 ;
        RECT -67.485 26.355 -67.155 26.685 ;
        RECT -67.485 24.995 -67.155 25.325 ;
        RECT -67.485 23.635 -67.155 23.965 ;
        RECT -67.485 22.275 -67.155 22.605 ;
        RECT -67.485 20.915 -67.155 21.245 ;
        RECT -67.485 19.555 -67.155 19.885 ;
        RECT -67.485 18.195 -67.155 18.525 ;
        RECT -67.485 16.835 -67.155 17.165 ;
        RECT -67.485 15.475 -67.155 15.805 ;
        RECT -67.485 14.115 -67.155 14.445 ;
        RECT -67.485 12.755 -67.155 13.085 ;
        RECT -67.485 11.395 -67.155 11.725 ;
        RECT -67.485 10.035 -67.155 10.365 ;
        RECT -67.485 8.675 -67.155 9.005 ;
        RECT -67.485 7.315 -67.155 7.645 ;
        RECT -67.485 5.955 -67.155 6.285 ;
        RECT -67.485 4.595 -67.155 4.925 ;
        RECT -67.485 3.235 -67.155 3.565 ;
        RECT -67.485 1.875 -67.155 2.205 ;
        RECT -67.485 0.515 -67.155 0.845 ;
        RECT -67.485 -0.845 -67.155 -0.515 ;
        RECT -67.485 -2.205 -67.155 -1.875 ;
        RECT -67.485 -3.565 -67.155 -3.235 ;
        RECT -67.485 -4.925 -67.155 -4.595 ;
        RECT -67.485 -6.285 -67.155 -5.955 ;
        RECT -67.485 -7.645 -67.155 -7.315 ;
        RECT -67.485 -9.005 -67.155 -8.675 ;
        RECT -67.485 -10.365 -67.155 -10.035 ;
        RECT -67.485 -11.725 -67.155 -11.395 ;
        RECT -67.485 -13.085 -67.155 -12.755 ;
        RECT -67.485 -14.445 -67.155 -14.115 ;
        RECT -67.485 -15.805 -67.155 -15.475 ;
        RECT -67.485 -17.165 -67.155 -16.835 ;
        RECT -67.485 -18.525 -67.155 -18.195 ;
        RECT -67.485 -19.885 -67.155 -19.555 ;
        RECT -67.485 -21.245 -67.155 -20.915 ;
        RECT -67.485 -22.605 -67.155 -22.275 ;
        RECT -67.485 -23.965 -67.155 -23.635 ;
        RECT -67.485 -25.325 -67.155 -24.995 ;
        RECT -67.485 -26.685 -67.155 -26.355 ;
        RECT -67.485 -28.045 -67.155 -27.715 ;
        RECT -67.485 -29.405 -67.155 -29.075 ;
        RECT -67.485 -30.765 -67.155 -30.435 ;
        RECT -67.485 -32.125 -67.155 -31.795 ;
        RECT -67.485 -33.485 -67.155 -33.155 ;
        RECT -67.485 -34.845 -67.155 -34.515 ;
        RECT -67.485 -36.205 -67.155 -35.875 ;
        RECT -67.485 -37.565 -67.155 -37.235 ;
        RECT -67.485 -38.925 -67.155 -38.595 ;
        RECT -67.485 -40.285 -67.155 -39.955 ;
        RECT -67.485 -41.645 -67.155 -41.315 ;
        RECT -67.485 -43.005 -67.155 -42.675 ;
        RECT -67.485 -44.365 -67.155 -44.035 ;
        RECT -67.485 -45.725 -67.155 -45.395 ;
        RECT -67.485 -47.085 -67.155 -46.755 ;
        RECT -67.485 -48.445 -67.155 -48.115 ;
        RECT -67.485 -49.805 -67.155 -49.475 ;
        RECT -67.485 -51.165 -67.155 -50.835 ;
        RECT -67.485 -52.525 -67.155 -52.195 ;
        RECT -67.485 -53.885 -67.155 -53.555 ;
        RECT -67.485 -55.245 -67.155 -54.915 ;
        RECT -67.485 -56.605 -67.155 -56.275 ;
        RECT -67.485 -57.965 -67.155 -57.635 ;
        RECT -67.485 -59.325 -67.155 -58.995 ;
        RECT -67.485 -60.685 -67.155 -60.355 ;
        RECT -67.485 -62.045 -67.155 -61.715 ;
        RECT -67.485 -63.405 -67.155 -63.075 ;
        RECT -67.485 -64.765 -67.155 -64.435 ;
        RECT -67.485 -66.125 -67.155 -65.795 ;
        RECT -67.485 -67.485 -67.155 -67.155 ;
        RECT -67.485 -68.845 -67.155 -68.515 ;
        RECT -67.485 -70.205 -67.155 -69.875 ;
        RECT -67.485 -71.565 -67.155 -71.235 ;
        RECT -67.485 -72.925 -67.155 -72.595 ;
        RECT -67.485 -74.285 -67.155 -73.955 ;
        RECT -67.485 -75.645 -67.155 -75.315 ;
        RECT -67.485 -77.005 -67.155 -76.675 ;
        RECT -67.485 -78.365 -67.155 -78.035 ;
        RECT -67.485 -79.725 -67.155 -79.395 ;
        RECT -67.485 -81.085 -67.155 -80.755 ;
        RECT -67.485 -82.445 -67.155 -82.115 ;
        RECT -67.485 -83.805 -67.155 -83.475 ;
        RECT -67.485 -85.165 -67.155 -84.835 ;
        RECT -67.485 -86.525 -67.155 -86.195 ;
        RECT -67.485 -87.885 -67.155 -87.555 ;
        RECT -67.485 -89.245 -67.155 -88.915 ;
        RECT -67.485 -90.605 -67.155 -90.275 ;
        RECT -67.485 -91.965 -67.155 -91.635 ;
        RECT -67.485 -93.325 -67.155 -92.995 ;
        RECT -67.485 -94.685 -67.155 -94.355 ;
        RECT -67.485 -96.045 -67.155 -95.715 ;
        RECT -67.485 -97.405 -67.155 -97.075 ;
        RECT -67.485 -98.765 -67.155 -98.435 ;
        RECT -67.485 -100.125 -67.155 -99.795 ;
        RECT -67.485 -101.485 -67.155 -101.155 ;
        RECT -67.485 -102.845 -67.155 -102.515 ;
        RECT -67.485 -104.205 -67.155 -103.875 ;
        RECT -67.485 -105.565 -67.155 -105.235 ;
        RECT -67.485 -106.925 -67.155 -106.595 ;
        RECT -67.485 -108.285 -67.155 -107.955 ;
        RECT -67.485 -109.645 -67.155 -109.315 ;
        RECT -67.485 -111.005 -67.155 -110.675 ;
        RECT -67.485 -112.365 -67.155 -112.035 ;
        RECT -67.485 -113.725 -67.155 -113.395 ;
        RECT -67.485 -115.085 -67.155 -114.755 ;
        RECT -67.485 -116.445 -67.155 -116.115 ;
        RECT -67.485 -117.805 -67.155 -117.475 ;
        RECT -67.485 -119.165 -67.155 -118.835 ;
        RECT -67.485 -120.525 -67.155 -120.195 ;
        RECT -67.485 -121.885 -67.155 -121.555 ;
        RECT -67.485 -123.245 -67.155 -122.915 ;
        RECT -67.485 -124.605 -67.155 -124.275 ;
        RECT -67.485 -125.965 -67.155 -125.635 ;
        RECT -67.485 -128.685 -67.155 -128.355 ;
        RECT -67.485 -130.045 -67.155 -129.715 ;
        RECT -67.485 -132.765 -67.155 -132.435 ;
        RECT -67.485 -134.125 -67.155 -133.795 ;
        RECT -67.485 -135.485 -67.155 -135.155 ;
        RECT -67.485 -136.845 -67.155 -136.515 ;
        RECT -67.485 -138.205 -67.155 -137.875 ;
        RECT -67.485 -139.39 -67.155 -139.06 ;
        RECT -67.485 -140.925 -67.155 -140.595 ;
        RECT -67.485 -142.285 -67.155 -141.955 ;
        RECT -67.485 -145.005 -67.155 -144.675 ;
        RECT -67.485 -146.365 -67.155 -146.035 ;
        RECT -67.485 -148.03 -67.155 -147.7 ;
        RECT -67.485 -149.085 -67.155 -148.755 ;
        RECT -67.485 -150.445 -67.155 -150.115 ;
        RECT -67.485 -153.165 -67.155 -152.835 ;
        RECT -67.485 -154.525 -67.155 -154.195 ;
        RECT -67.485 -155.885 -67.155 -155.555 ;
        RECT -67.485 -157.245 -67.155 -156.915 ;
        RECT -67.485 -158.605 -67.155 -158.275 ;
        RECT -67.485 -159.965 -67.155 -159.635 ;
        RECT -67.485 -161.325 -67.155 -160.995 ;
        RECT -67.485 -162.685 -67.155 -162.355 ;
        RECT -67.485 -164.045 -67.155 -163.715 ;
        RECT -67.485 -165.405 -67.155 -165.075 ;
        RECT -67.485 -166.765 -67.155 -166.435 ;
        RECT -67.485 -168.125 -67.155 -167.795 ;
        RECT -67.485 -169.485 -67.155 -169.155 ;
        RECT -67.485 -170.845 -67.155 -170.515 ;
        RECT -67.485 -172.205 -67.155 -171.875 ;
        RECT -67.485 -173.565 -67.155 -173.235 ;
        RECT -67.485 -174.925 -67.155 -174.595 ;
        RECT -67.485 -176.285 -67.155 -175.955 ;
        RECT -67.485 -177.645 -67.155 -177.315 ;
        RECT -67.485 -179.005 -67.155 -178.675 ;
        RECT -67.485 -180.365 -67.155 -180.035 ;
        RECT -67.485 -181.725 -67.155 -181.395 ;
        RECT -67.485 -183.085 -67.155 -182.755 ;
        RECT -67.485 -184.445 -67.155 -184.115 ;
        RECT -67.485 -185.805 -67.155 -185.475 ;
        RECT -67.485 -187.165 -67.155 -186.835 ;
        RECT -67.485 -188.525 -67.155 -188.195 ;
        RECT -67.485 -189.885 -67.155 -189.555 ;
        RECT -67.485 -191.245 -67.155 -190.915 ;
        RECT -67.485 -192.605 -67.155 -192.275 ;
        RECT -67.485 -193.965 -67.155 -193.635 ;
        RECT -67.485 -195.325 -67.155 -194.995 ;
        RECT -67.485 -196.685 -67.155 -196.355 ;
        RECT -67.485 -198.045 -67.155 -197.715 ;
        RECT -67.485 -199.405 -67.155 -199.075 ;
        RECT -67.485 -200.765 -67.155 -200.435 ;
        RECT -67.485 -202.125 -67.155 -201.795 ;
        RECT -67.485 -203.485 -67.155 -203.155 ;
        RECT -67.485 -204.845 -67.155 -204.515 ;
        RECT -67.485 -206.205 -67.155 -205.875 ;
        RECT -67.485 -207.565 -67.155 -207.235 ;
        RECT -67.485 -208.925 -67.155 -208.595 ;
        RECT -67.485 -210.285 -67.155 -209.955 ;
        RECT -67.485 -211.645 -67.155 -211.315 ;
        RECT -67.485 -213.005 -67.155 -212.675 ;
        RECT -67.485 -214.365 -67.155 -214.035 ;
        RECT -67.485 -215.725 -67.155 -215.395 ;
        RECT -67.485 -217.085 -67.155 -216.755 ;
        RECT -67.485 -218.445 -67.155 -218.115 ;
        RECT -67.485 -219.805 -67.155 -219.475 ;
        RECT -67.485 -221.165 -67.155 -220.835 ;
        RECT -67.485 -222.525 -67.155 -222.195 ;
        RECT -67.485 -223.885 -67.155 -223.555 ;
        RECT -67.485 -225.245 -67.155 -224.915 ;
        RECT -67.485 -227.965 -67.155 -227.635 ;
        RECT -67.485 -232.045 -67.155 -231.715 ;
        RECT -67.485 -233.225 -67.155 -232.895 ;
        RECT -67.485 -234.765 -67.155 -234.435 ;
        RECT -67.485 -236.125 -67.155 -235.795 ;
        RECT -67.485 -237.485 -67.155 -237.155 ;
        RECT -67.485 -238.845 -67.155 -238.515 ;
        RECT -67.485 -241.09 -67.155 -239.96 ;
        RECT -67.48 -241.205 -67.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.125 244.04 -65.795 245.17 ;
        RECT -66.125 242.595 -65.795 242.925 ;
        RECT -66.125 241.235 -65.795 241.565 ;
        RECT -66.125 239.875 -65.795 240.205 ;
        RECT -66.125 238.515 -65.795 238.845 ;
        RECT -66.125 237.155 -65.795 237.485 ;
        RECT -66.125 235.795 -65.795 236.125 ;
        RECT -66.125 234.435 -65.795 234.765 ;
        RECT -66.125 233.075 -65.795 233.405 ;
        RECT -66.125 231.715 -65.795 232.045 ;
        RECT -66.125 230.355 -65.795 230.685 ;
        RECT -66.125 228.995 -65.795 229.325 ;
        RECT -66.125 227.635 -65.795 227.965 ;
        RECT -66.125 226.275 -65.795 226.605 ;
        RECT -66.125 224.915 -65.795 225.245 ;
        RECT -66.125 223.555 -65.795 223.885 ;
        RECT -66.125 222.195 -65.795 222.525 ;
        RECT -66.125 220.835 -65.795 221.165 ;
        RECT -66.125 219.475 -65.795 219.805 ;
        RECT -66.125 218.115 -65.795 218.445 ;
        RECT -66.125 216.755 -65.795 217.085 ;
        RECT -66.125 215.395 -65.795 215.725 ;
        RECT -66.125 214.035 -65.795 214.365 ;
        RECT -66.125 212.675 -65.795 213.005 ;
        RECT -66.125 211.315 -65.795 211.645 ;
        RECT -66.125 209.955 -65.795 210.285 ;
        RECT -66.125 208.595 -65.795 208.925 ;
        RECT -66.125 207.235 -65.795 207.565 ;
        RECT -66.125 205.875 -65.795 206.205 ;
        RECT -66.125 204.515 -65.795 204.845 ;
        RECT -66.125 203.155 -65.795 203.485 ;
        RECT -66.125 201.795 -65.795 202.125 ;
        RECT -66.125 200.435 -65.795 200.765 ;
        RECT -66.125 199.075 -65.795 199.405 ;
        RECT -66.125 197.715 -65.795 198.045 ;
        RECT -66.125 196.355 -65.795 196.685 ;
        RECT -66.125 194.995 -65.795 195.325 ;
        RECT -66.125 193.635 -65.795 193.965 ;
        RECT -66.125 192.275 -65.795 192.605 ;
        RECT -66.125 190.915 -65.795 191.245 ;
        RECT -66.125 189.555 -65.795 189.885 ;
        RECT -66.125 188.195 -65.795 188.525 ;
        RECT -66.125 186.835 -65.795 187.165 ;
        RECT -66.125 185.475 -65.795 185.805 ;
        RECT -66.125 184.115 -65.795 184.445 ;
        RECT -66.125 182.755 -65.795 183.085 ;
        RECT -66.125 181.395 -65.795 181.725 ;
        RECT -66.125 180.035 -65.795 180.365 ;
        RECT -66.125 178.675 -65.795 179.005 ;
        RECT -66.125 177.315 -65.795 177.645 ;
        RECT -66.125 175.955 -65.795 176.285 ;
        RECT -66.125 174.595 -65.795 174.925 ;
        RECT -66.125 173.235 -65.795 173.565 ;
        RECT -66.125 171.875 -65.795 172.205 ;
        RECT -66.125 170.515 -65.795 170.845 ;
        RECT -66.125 169.155 -65.795 169.485 ;
        RECT -66.125 167.795 -65.795 168.125 ;
        RECT -66.125 166.435 -65.795 166.765 ;
        RECT -66.125 165.075 -65.795 165.405 ;
        RECT -66.125 163.715 -65.795 164.045 ;
        RECT -66.125 162.355 -65.795 162.685 ;
        RECT -66.125 160.995 -65.795 161.325 ;
        RECT -66.125 159.635 -65.795 159.965 ;
        RECT -66.125 158.275 -65.795 158.605 ;
        RECT -66.125 156.915 -65.795 157.245 ;
        RECT -66.125 155.555 -65.795 155.885 ;
        RECT -66.125 154.195 -65.795 154.525 ;
        RECT -66.125 152.835 -65.795 153.165 ;
        RECT -66.125 151.475 -65.795 151.805 ;
        RECT -66.125 150.115 -65.795 150.445 ;
        RECT -66.125 148.755 -65.795 149.085 ;
        RECT -66.125 147.395 -65.795 147.725 ;
        RECT -66.125 146.035 -65.795 146.365 ;
        RECT -66.125 144.675 -65.795 145.005 ;
        RECT -66.125 143.315 -65.795 143.645 ;
        RECT -66.125 141.955 -65.795 142.285 ;
        RECT -66.125 140.595 -65.795 140.925 ;
        RECT -66.125 139.235 -65.795 139.565 ;
        RECT -66.125 137.875 -65.795 138.205 ;
        RECT -66.125 136.515 -65.795 136.845 ;
        RECT -66.125 135.155 -65.795 135.485 ;
        RECT -66.125 133.795 -65.795 134.125 ;
        RECT -66.125 132.435 -65.795 132.765 ;
        RECT -66.125 131.075 -65.795 131.405 ;
        RECT -66.125 129.715 -65.795 130.045 ;
        RECT -66.125 128.355 -65.795 128.685 ;
        RECT -66.125 126.995 -65.795 127.325 ;
        RECT -66.125 125.635 -65.795 125.965 ;
        RECT -66.125 124.275 -65.795 124.605 ;
        RECT -66.125 122.915 -65.795 123.245 ;
        RECT -66.125 121.555 -65.795 121.885 ;
        RECT -66.125 120.195 -65.795 120.525 ;
        RECT -66.125 118.835 -65.795 119.165 ;
        RECT -66.125 117.475 -65.795 117.805 ;
        RECT -66.125 116.115 -65.795 116.445 ;
        RECT -66.125 114.755 -65.795 115.085 ;
        RECT -66.125 113.395 -65.795 113.725 ;
        RECT -66.125 112.035 -65.795 112.365 ;
        RECT -66.125 110.675 -65.795 111.005 ;
        RECT -66.125 109.315 -65.795 109.645 ;
        RECT -66.125 107.955 -65.795 108.285 ;
        RECT -66.125 106.595 -65.795 106.925 ;
        RECT -66.125 105.235 -65.795 105.565 ;
        RECT -66.125 103.875 -65.795 104.205 ;
        RECT -66.125 102.515 -65.795 102.845 ;
        RECT -66.125 101.155 -65.795 101.485 ;
        RECT -66.125 99.795 -65.795 100.125 ;
        RECT -66.125 98.435 -65.795 98.765 ;
        RECT -66.125 97.075 -65.795 97.405 ;
        RECT -66.125 95.715 -65.795 96.045 ;
        RECT -66.125 94.355 -65.795 94.685 ;
        RECT -66.125 92.995 -65.795 93.325 ;
        RECT -66.125 91.635 -65.795 91.965 ;
        RECT -66.125 90.275 -65.795 90.605 ;
        RECT -66.125 88.915 -65.795 89.245 ;
        RECT -66.125 87.555 -65.795 87.885 ;
        RECT -66.125 86.195 -65.795 86.525 ;
        RECT -66.125 84.835 -65.795 85.165 ;
        RECT -66.125 83.475 -65.795 83.805 ;
        RECT -66.125 82.115 -65.795 82.445 ;
        RECT -66.125 80.755 -65.795 81.085 ;
        RECT -66.125 79.395 -65.795 79.725 ;
        RECT -66.125 78.035 -65.795 78.365 ;
        RECT -66.125 76.675 -65.795 77.005 ;
        RECT -66.125 75.315 -65.795 75.645 ;
        RECT -66.125 73.955 -65.795 74.285 ;
        RECT -66.125 72.595 -65.795 72.925 ;
        RECT -66.125 71.235 -65.795 71.565 ;
        RECT -66.125 69.875 -65.795 70.205 ;
        RECT -66.125 68.515 -65.795 68.845 ;
        RECT -66.125 67.155 -65.795 67.485 ;
        RECT -66.125 65.795 -65.795 66.125 ;
        RECT -66.125 64.435 -65.795 64.765 ;
        RECT -66.125 63.075 -65.795 63.405 ;
        RECT -66.125 61.715 -65.795 62.045 ;
        RECT -66.125 60.355 -65.795 60.685 ;
        RECT -66.125 58.995 -65.795 59.325 ;
        RECT -66.125 57.635 -65.795 57.965 ;
        RECT -66.125 56.275 -65.795 56.605 ;
        RECT -66.125 54.915 -65.795 55.245 ;
        RECT -66.125 53.555 -65.795 53.885 ;
        RECT -66.125 52.195 -65.795 52.525 ;
        RECT -66.125 50.835 -65.795 51.165 ;
        RECT -66.125 49.475 -65.795 49.805 ;
        RECT -66.125 48.115 -65.795 48.445 ;
        RECT -66.125 46.755 -65.795 47.085 ;
        RECT -66.125 45.395 -65.795 45.725 ;
        RECT -66.125 44.035 -65.795 44.365 ;
        RECT -66.125 42.675 -65.795 43.005 ;
        RECT -66.125 41.315 -65.795 41.645 ;
        RECT -66.125 39.955 -65.795 40.285 ;
        RECT -66.125 38.595 -65.795 38.925 ;
        RECT -66.125 37.235 -65.795 37.565 ;
        RECT -66.125 35.875 -65.795 36.205 ;
        RECT -66.125 34.515 -65.795 34.845 ;
        RECT -66.125 33.155 -65.795 33.485 ;
        RECT -66.125 31.795 -65.795 32.125 ;
        RECT -66.125 30.435 -65.795 30.765 ;
        RECT -66.125 29.075 -65.795 29.405 ;
        RECT -66.125 27.715 -65.795 28.045 ;
        RECT -66.125 26.355 -65.795 26.685 ;
        RECT -66.125 24.995 -65.795 25.325 ;
        RECT -66.125 23.635 -65.795 23.965 ;
        RECT -66.125 22.275 -65.795 22.605 ;
        RECT -66.125 20.915 -65.795 21.245 ;
        RECT -66.125 19.555 -65.795 19.885 ;
        RECT -66.125 18.195 -65.795 18.525 ;
        RECT -66.125 16.835 -65.795 17.165 ;
        RECT -66.125 15.475 -65.795 15.805 ;
        RECT -66.125 14.115 -65.795 14.445 ;
        RECT -66.125 12.755 -65.795 13.085 ;
        RECT -66.125 11.395 -65.795 11.725 ;
        RECT -66.125 10.035 -65.795 10.365 ;
        RECT -66.125 8.675 -65.795 9.005 ;
        RECT -66.125 7.315 -65.795 7.645 ;
        RECT -66.125 5.955 -65.795 6.285 ;
        RECT -66.125 4.595 -65.795 4.925 ;
        RECT -66.125 3.235 -65.795 3.565 ;
        RECT -66.125 1.875 -65.795 2.205 ;
        RECT -66.125 0.515 -65.795 0.845 ;
        RECT -66.125 -0.845 -65.795 -0.515 ;
        RECT -66.125 -2.205 -65.795 -1.875 ;
        RECT -66.125 -3.565 -65.795 -3.235 ;
        RECT -66.125 -4.925 -65.795 -4.595 ;
        RECT -66.125 -6.285 -65.795 -5.955 ;
        RECT -66.125 -7.645 -65.795 -7.315 ;
        RECT -66.125 -9.005 -65.795 -8.675 ;
        RECT -66.125 -10.365 -65.795 -10.035 ;
        RECT -66.125 -11.725 -65.795 -11.395 ;
        RECT -66.125 -13.085 -65.795 -12.755 ;
        RECT -66.125 -14.445 -65.795 -14.115 ;
        RECT -66.125 -15.805 -65.795 -15.475 ;
        RECT -66.125 -17.165 -65.795 -16.835 ;
        RECT -66.125 -18.525 -65.795 -18.195 ;
        RECT -66.125 -19.885 -65.795 -19.555 ;
        RECT -66.125 -21.245 -65.795 -20.915 ;
        RECT -66.125 -22.605 -65.795 -22.275 ;
        RECT -66.125 -23.965 -65.795 -23.635 ;
        RECT -66.125 -25.325 -65.795 -24.995 ;
        RECT -66.125 -26.685 -65.795 -26.355 ;
        RECT -66.125 -28.045 -65.795 -27.715 ;
        RECT -66.125 -29.405 -65.795 -29.075 ;
        RECT -66.125 -30.765 -65.795 -30.435 ;
        RECT -66.125 -32.125 -65.795 -31.795 ;
        RECT -66.125 -33.485 -65.795 -33.155 ;
        RECT -66.125 -34.845 -65.795 -34.515 ;
        RECT -66.125 -36.205 -65.795 -35.875 ;
        RECT -66.125 -37.565 -65.795 -37.235 ;
        RECT -66.125 -38.925 -65.795 -38.595 ;
        RECT -66.125 -40.285 -65.795 -39.955 ;
        RECT -66.125 -41.645 -65.795 -41.315 ;
        RECT -66.125 -43.005 -65.795 -42.675 ;
        RECT -66.125 -44.365 -65.795 -44.035 ;
        RECT -66.125 -45.725 -65.795 -45.395 ;
        RECT -66.125 -47.085 -65.795 -46.755 ;
        RECT -66.125 -48.445 -65.795 -48.115 ;
        RECT -66.125 -49.805 -65.795 -49.475 ;
        RECT -66.125 -51.165 -65.795 -50.835 ;
        RECT -66.125 -52.525 -65.795 -52.195 ;
        RECT -66.125 -53.885 -65.795 -53.555 ;
        RECT -66.125 -55.245 -65.795 -54.915 ;
        RECT -66.125 -56.605 -65.795 -56.275 ;
        RECT -66.125 -57.965 -65.795 -57.635 ;
        RECT -66.125 -59.325 -65.795 -58.995 ;
        RECT -66.125 -60.685 -65.795 -60.355 ;
        RECT -66.125 -62.045 -65.795 -61.715 ;
        RECT -66.125 -63.405 -65.795 -63.075 ;
        RECT -66.125 -64.765 -65.795 -64.435 ;
        RECT -66.125 -66.125 -65.795 -65.795 ;
        RECT -66.125 -67.485 -65.795 -67.155 ;
        RECT -66.125 -68.845 -65.795 -68.515 ;
        RECT -66.125 -70.205 -65.795 -69.875 ;
        RECT -66.125 -71.565 -65.795 -71.235 ;
        RECT -66.125 -72.925 -65.795 -72.595 ;
        RECT -66.125 -74.285 -65.795 -73.955 ;
        RECT -66.125 -75.645 -65.795 -75.315 ;
        RECT -66.125 -77.005 -65.795 -76.675 ;
        RECT -66.125 -78.365 -65.795 -78.035 ;
        RECT -66.125 -79.725 -65.795 -79.395 ;
        RECT -66.125 -81.085 -65.795 -80.755 ;
        RECT -66.125 -82.445 -65.795 -82.115 ;
        RECT -66.125 -83.805 -65.795 -83.475 ;
        RECT -66.125 -85.165 -65.795 -84.835 ;
        RECT -66.125 -86.525 -65.795 -86.195 ;
        RECT -66.125 -87.885 -65.795 -87.555 ;
        RECT -66.125 -89.245 -65.795 -88.915 ;
        RECT -66.125 -90.605 -65.795 -90.275 ;
        RECT -66.125 -91.965 -65.795 -91.635 ;
        RECT -66.125 -93.325 -65.795 -92.995 ;
        RECT -66.125 -94.685 -65.795 -94.355 ;
        RECT -66.125 -96.045 -65.795 -95.715 ;
        RECT -66.125 -97.405 -65.795 -97.075 ;
        RECT -66.125 -98.765 -65.795 -98.435 ;
        RECT -66.125 -100.125 -65.795 -99.795 ;
        RECT -66.125 -101.485 -65.795 -101.155 ;
        RECT -66.125 -102.845 -65.795 -102.515 ;
        RECT -66.125 -104.205 -65.795 -103.875 ;
        RECT -66.125 -105.565 -65.795 -105.235 ;
        RECT -66.125 -106.925 -65.795 -106.595 ;
        RECT -66.125 -108.285 -65.795 -107.955 ;
        RECT -66.125 -109.645 -65.795 -109.315 ;
        RECT -66.125 -111.005 -65.795 -110.675 ;
        RECT -66.125 -112.365 -65.795 -112.035 ;
        RECT -66.125 -113.725 -65.795 -113.395 ;
        RECT -66.125 -115.085 -65.795 -114.755 ;
        RECT -66.125 -116.445 -65.795 -116.115 ;
        RECT -66.125 -117.805 -65.795 -117.475 ;
        RECT -66.125 -119.165 -65.795 -118.835 ;
        RECT -66.125 -120.525 -65.795 -120.195 ;
        RECT -66.125 -121.885 -65.795 -121.555 ;
        RECT -66.125 -123.245 -65.795 -122.915 ;
        RECT -66.125 -124.605 -65.795 -124.275 ;
        RECT -66.125 -125.965 -65.795 -125.635 ;
        RECT -66.125 -128.685 -65.795 -128.355 ;
        RECT -66.125 -130.045 -65.795 -129.715 ;
        RECT -66.125 -132.765 -65.795 -132.435 ;
        RECT -66.125 -134.125 -65.795 -133.795 ;
        RECT -66.125 -135.485 -65.795 -135.155 ;
        RECT -66.125 -136.845 -65.795 -136.515 ;
        RECT -66.125 -138.205 -65.795 -137.875 ;
        RECT -66.125 -139.39 -65.795 -139.06 ;
        RECT -66.125 -140.925 -65.795 -140.595 ;
        RECT -66.125 -142.285 -65.795 -141.955 ;
        RECT -66.125 -145.005 -65.795 -144.675 ;
        RECT -66.125 -146.365 -65.795 -146.035 ;
        RECT -66.125 -148.03 -65.795 -147.7 ;
        RECT -66.125 -149.085 -65.795 -148.755 ;
        RECT -66.125 -153.165 -65.795 -152.835 ;
        RECT -66.125 -154.525 -65.795 -154.195 ;
        RECT -66.125 -155.885 -65.795 -155.555 ;
        RECT -66.125 -157.245 -65.795 -156.915 ;
        RECT -66.125 -158.605 -65.795 -158.275 ;
        RECT -66.125 -159.965 -65.795 -159.635 ;
        RECT -66.125 -161.325 -65.795 -160.995 ;
        RECT -66.125 -162.685 -65.795 -162.355 ;
        RECT -66.125 -164.045 -65.795 -163.715 ;
        RECT -66.125 -165.405 -65.795 -165.075 ;
        RECT -66.125 -166.765 -65.795 -166.435 ;
        RECT -66.125 -168.125 -65.795 -167.795 ;
        RECT -66.125 -169.485 -65.795 -169.155 ;
        RECT -66.125 -170.845 -65.795 -170.515 ;
        RECT -66.125 -172.205 -65.795 -171.875 ;
        RECT -66.125 -173.565 -65.795 -173.235 ;
        RECT -66.125 -174.925 -65.795 -174.595 ;
        RECT -66.125 -176.285 -65.795 -175.955 ;
        RECT -66.125 -177.645 -65.795 -177.315 ;
        RECT -66.125 -179.005 -65.795 -178.675 ;
        RECT -66.125 -180.365 -65.795 -180.035 ;
        RECT -66.125 -181.725 -65.795 -181.395 ;
        RECT -66.125 -183.085 -65.795 -182.755 ;
        RECT -66.125 -184.445 -65.795 -184.115 ;
        RECT -66.125 -185.805 -65.795 -185.475 ;
        RECT -66.125 -187.165 -65.795 -186.835 ;
        RECT -66.125 -188.525 -65.795 -188.195 ;
        RECT -66.125 -189.885 -65.795 -189.555 ;
        RECT -66.125 -191.245 -65.795 -190.915 ;
        RECT -66.125 -192.605 -65.795 -192.275 ;
        RECT -66.125 -193.965 -65.795 -193.635 ;
        RECT -66.125 -195.325 -65.795 -194.995 ;
        RECT -66.125 -196.685 -65.795 -196.355 ;
        RECT -66.125 -198.045 -65.795 -197.715 ;
        RECT -66.125 -199.405 -65.795 -199.075 ;
        RECT -66.125 -200.765 -65.795 -200.435 ;
        RECT -66.125 -202.125 -65.795 -201.795 ;
        RECT -66.125 -203.485 -65.795 -203.155 ;
        RECT -66.125 -204.845 -65.795 -204.515 ;
        RECT -66.125 -206.205 -65.795 -205.875 ;
        RECT -66.125 -207.565 -65.795 -207.235 ;
        RECT -66.125 -208.925 -65.795 -208.595 ;
        RECT -66.125 -210.285 -65.795 -209.955 ;
        RECT -66.125 -211.645 -65.795 -211.315 ;
        RECT -66.125 -213.005 -65.795 -212.675 ;
        RECT -66.125 -214.365 -65.795 -214.035 ;
        RECT -66.125 -215.725 -65.795 -215.395 ;
        RECT -66.125 -217.085 -65.795 -216.755 ;
        RECT -66.125 -218.445 -65.795 -218.115 ;
        RECT -66.125 -219.805 -65.795 -219.475 ;
        RECT -66.125 -221.165 -65.795 -220.835 ;
        RECT -66.125 -222.525 -65.795 -222.195 ;
        RECT -66.125 -223.885 -65.795 -223.555 ;
        RECT -66.125 -225.245 -65.795 -224.915 ;
        RECT -66.125 -227.965 -65.795 -227.635 ;
        RECT -66.125 -232.045 -65.795 -231.715 ;
        RECT -66.125 -234.765 -65.795 -234.435 ;
        RECT -66.125 -236.125 -65.795 -235.795 ;
        RECT -66.125 -237.485 -65.795 -237.155 ;
        RECT -66.125 -238.845 -65.795 -238.515 ;
        RECT -66.125 -241.09 -65.795 -239.96 ;
        RECT -66.12 -241.205 -65.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.765 -232.045 -64.435 -231.715 ;
        RECT -64.765 -233.225 -64.435 -232.895 ;
        RECT -64.765 -234.765 -64.435 -234.435 ;
        RECT -64.765 -236.125 -64.435 -235.795 ;
        RECT -64.765 -237.485 -64.435 -237.155 ;
        RECT -64.765 -238.845 -64.435 -238.515 ;
        RECT -64.765 -241.09 -64.435 -239.96 ;
        RECT -64.76 -241.205 -64.44 245.285 ;
        RECT -64.765 244.04 -64.435 245.17 ;
        RECT -64.765 242.595 -64.435 242.925 ;
        RECT -64.765 241.235 -64.435 241.565 ;
        RECT -64.765 239.875 -64.435 240.205 ;
        RECT -64.765 238.515 -64.435 238.845 ;
        RECT -64.765 237.155 -64.435 237.485 ;
        RECT -64.765 235.795 -64.435 236.125 ;
        RECT -64.765 234.435 -64.435 234.765 ;
        RECT -64.765 233.075 -64.435 233.405 ;
        RECT -64.765 231.715 -64.435 232.045 ;
        RECT -64.765 230.355 -64.435 230.685 ;
        RECT -64.765 228.995 -64.435 229.325 ;
        RECT -64.765 227.635 -64.435 227.965 ;
        RECT -64.765 226.275 -64.435 226.605 ;
        RECT -64.765 224.915 -64.435 225.245 ;
        RECT -64.765 223.555 -64.435 223.885 ;
        RECT -64.765 222.195 -64.435 222.525 ;
        RECT -64.765 220.835 -64.435 221.165 ;
        RECT -64.765 219.475 -64.435 219.805 ;
        RECT -64.765 218.115 -64.435 218.445 ;
        RECT -64.765 216.755 -64.435 217.085 ;
        RECT -64.765 215.395 -64.435 215.725 ;
        RECT -64.765 214.035 -64.435 214.365 ;
        RECT -64.765 212.675 -64.435 213.005 ;
        RECT -64.765 211.315 -64.435 211.645 ;
        RECT -64.765 209.955 -64.435 210.285 ;
        RECT -64.765 208.595 -64.435 208.925 ;
        RECT -64.765 207.235 -64.435 207.565 ;
        RECT -64.765 205.875 -64.435 206.205 ;
        RECT -64.765 204.515 -64.435 204.845 ;
        RECT -64.765 203.155 -64.435 203.485 ;
        RECT -64.765 201.795 -64.435 202.125 ;
        RECT -64.765 200.435 -64.435 200.765 ;
        RECT -64.765 199.075 -64.435 199.405 ;
        RECT -64.765 197.715 -64.435 198.045 ;
        RECT -64.765 196.355 -64.435 196.685 ;
        RECT -64.765 194.995 -64.435 195.325 ;
        RECT -64.765 193.635 -64.435 193.965 ;
        RECT -64.765 192.275 -64.435 192.605 ;
        RECT -64.765 190.915 -64.435 191.245 ;
        RECT -64.765 189.555 -64.435 189.885 ;
        RECT -64.765 188.195 -64.435 188.525 ;
        RECT -64.765 186.835 -64.435 187.165 ;
        RECT -64.765 185.475 -64.435 185.805 ;
        RECT -64.765 184.115 -64.435 184.445 ;
        RECT -64.765 182.755 -64.435 183.085 ;
        RECT -64.765 181.395 -64.435 181.725 ;
        RECT -64.765 180.035 -64.435 180.365 ;
        RECT -64.765 178.675 -64.435 179.005 ;
        RECT -64.765 177.315 -64.435 177.645 ;
        RECT -64.765 175.955 -64.435 176.285 ;
        RECT -64.765 174.595 -64.435 174.925 ;
        RECT -64.765 173.235 -64.435 173.565 ;
        RECT -64.765 171.875 -64.435 172.205 ;
        RECT -64.765 170.515 -64.435 170.845 ;
        RECT -64.765 169.155 -64.435 169.485 ;
        RECT -64.765 167.795 -64.435 168.125 ;
        RECT -64.765 166.435 -64.435 166.765 ;
        RECT -64.765 165.075 -64.435 165.405 ;
        RECT -64.765 163.715 -64.435 164.045 ;
        RECT -64.765 162.355 -64.435 162.685 ;
        RECT -64.765 160.995 -64.435 161.325 ;
        RECT -64.765 159.635 -64.435 159.965 ;
        RECT -64.765 158.275 -64.435 158.605 ;
        RECT -64.765 156.915 -64.435 157.245 ;
        RECT -64.765 155.555 -64.435 155.885 ;
        RECT -64.765 154.195 -64.435 154.525 ;
        RECT -64.765 152.835 -64.435 153.165 ;
        RECT -64.765 151.475 -64.435 151.805 ;
        RECT -64.765 150.115 -64.435 150.445 ;
        RECT -64.765 148.755 -64.435 149.085 ;
        RECT -64.765 147.395 -64.435 147.725 ;
        RECT -64.765 146.035 -64.435 146.365 ;
        RECT -64.765 144.675 -64.435 145.005 ;
        RECT -64.765 143.315 -64.435 143.645 ;
        RECT -64.765 141.955 -64.435 142.285 ;
        RECT -64.765 140.595 -64.435 140.925 ;
        RECT -64.765 139.235 -64.435 139.565 ;
        RECT -64.765 137.875 -64.435 138.205 ;
        RECT -64.765 136.515 -64.435 136.845 ;
        RECT -64.765 135.155 -64.435 135.485 ;
        RECT -64.765 133.795 -64.435 134.125 ;
        RECT -64.765 132.435 -64.435 132.765 ;
        RECT -64.765 131.075 -64.435 131.405 ;
        RECT -64.765 129.715 -64.435 130.045 ;
        RECT -64.765 128.355 -64.435 128.685 ;
        RECT -64.765 126.995 -64.435 127.325 ;
        RECT -64.765 125.635 -64.435 125.965 ;
        RECT -64.765 124.275 -64.435 124.605 ;
        RECT -64.765 122.915 -64.435 123.245 ;
        RECT -64.765 121.555 -64.435 121.885 ;
        RECT -64.765 120.195 -64.435 120.525 ;
        RECT -64.765 118.835 -64.435 119.165 ;
        RECT -64.765 117.475 -64.435 117.805 ;
        RECT -64.765 116.115 -64.435 116.445 ;
        RECT -64.765 114.755 -64.435 115.085 ;
        RECT -64.765 113.395 -64.435 113.725 ;
        RECT -64.765 112.035 -64.435 112.365 ;
        RECT -64.765 110.675 -64.435 111.005 ;
        RECT -64.765 109.315 -64.435 109.645 ;
        RECT -64.765 107.955 -64.435 108.285 ;
        RECT -64.765 106.595 -64.435 106.925 ;
        RECT -64.765 105.235 -64.435 105.565 ;
        RECT -64.765 103.875 -64.435 104.205 ;
        RECT -64.765 102.515 -64.435 102.845 ;
        RECT -64.765 101.155 -64.435 101.485 ;
        RECT -64.765 99.795 -64.435 100.125 ;
        RECT -64.765 98.435 -64.435 98.765 ;
        RECT -64.765 97.075 -64.435 97.405 ;
        RECT -64.765 95.715 -64.435 96.045 ;
        RECT -64.765 94.355 -64.435 94.685 ;
        RECT -64.765 92.995 -64.435 93.325 ;
        RECT -64.765 91.635 -64.435 91.965 ;
        RECT -64.765 90.275 -64.435 90.605 ;
        RECT -64.765 88.915 -64.435 89.245 ;
        RECT -64.765 87.555 -64.435 87.885 ;
        RECT -64.765 86.195 -64.435 86.525 ;
        RECT -64.765 84.835 -64.435 85.165 ;
        RECT -64.765 83.475 -64.435 83.805 ;
        RECT -64.765 82.115 -64.435 82.445 ;
        RECT -64.765 80.755 -64.435 81.085 ;
        RECT -64.765 79.395 -64.435 79.725 ;
        RECT -64.765 78.035 -64.435 78.365 ;
        RECT -64.765 76.675 -64.435 77.005 ;
        RECT -64.765 75.315 -64.435 75.645 ;
        RECT -64.765 73.955 -64.435 74.285 ;
        RECT -64.765 72.595 -64.435 72.925 ;
        RECT -64.765 71.235 -64.435 71.565 ;
        RECT -64.765 69.875 -64.435 70.205 ;
        RECT -64.765 68.515 -64.435 68.845 ;
        RECT -64.765 67.155 -64.435 67.485 ;
        RECT -64.765 65.795 -64.435 66.125 ;
        RECT -64.765 64.435 -64.435 64.765 ;
        RECT -64.765 63.075 -64.435 63.405 ;
        RECT -64.765 61.715 -64.435 62.045 ;
        RECT -64.765 60.355 -64.435 60.685 ;
        RECT -64.765 58.995 -64.435 59.325 ;
        RECT -64.765 57.635 -64.435 57.965 ;
        RECT -64.765 56.275 -64.435 56.605 ;
        RECT -64.765 54.915 -64.435 55.245 ;
        RECT -64.765 53.555 -64.435 53.885 ;
        RECT -64.765 52.195 -64.435 52.525 ;
        RECT -64.765 50.835 -64.435 51.165 ;
        RECT -64.765 49.475 -64.435 49.805 ;
        RECT -64.765 48.115 -64.435 48.445 ;
        RECT -64.765 46.755 -64.435 47.085 ;
        RECT -64.765 45.395 -64.435 45.725 ;
        RECT -64.765 44.035 -64.435 44.365 ;
        RECT -64.765 42.675 -64.435 43.005 ;
        RECT -64.765 41.315 -64.435 41.645 ;
        RECT -64.765 39.955 -64.435 40.285 ;
        RECT -64.765 38.595 -64.435 38.925 ;
        RECT -64.765 37.235 -64.435 37.565 ;
        RECT -64.765 35.875 -64.435 36.205 ;
        RECT -64.765 34.515 -64.435 34.845 ;
        RECT -64.765 33.155 -64.435 33.485 ;
        RECT -64.765 31.795 -64.435 32.125 ;
        RECT -64.765 30.435 -64.435 30.765 ;
        RECT -64.765 29.075 -64.435 29.405 ;
        RECT -64.765 27.715 -64.435 28.045 ;
        RECT -64.765 26.355 -64.435 26.685 ;
        RECT -64.765 24.995 -64.435 25.325 ;
        RECT -64.765 23.635 -64.435 23.965 ;
        RECT -64.765 22.275 -64.435 22.605 ;
        RECT -64.765 20.915 -64.435 21.245 ;
        RECT -64.765 19.555 -64.435 19.885 ;
        RECT -64.765 18.195 -64.435 18.525 ;
        RECT -64.765 16.835 -64.435 17.165 ;
        RECT -64.765 15.475 -64.435 15.805 ;
        RECT -64.765 14.115 -64.435 14.445 ;
        RECT -64.765 12.755 -64.435 13.085 ;
        RECT -64.765 11.395 -64.435 11.725 ;
        RECT -64.765 10.035 -64.435 10.365 ;
        RECT -64.765 8.675 -64.435 9.005 ;
        RECT -64.765 7.315 -64.435 7.645 ;
        RECT -64.765 5.955 -64.435 6.285 ;
        RECT -64.765 4.595 -64.435 4.925 ;
        RECT -64.765 3.235 -64.435 3.565 ;
        RECT -64.765 1.875 -64.435 2.205 ;
        RECT -64.765 0.515 -64.435 0.845 ;
        RECT -64.765 -0.845 -64.435 -0.515 ;
        RECT -64.765 -2.205 -64.435 -1.875 ;
        RECT -64.765 -3.565 -64.435 -3.235 ;
        RECT -64.765 -4.925 -64.435 -4.595 ;
        RECT -64.765 -6.285 -64.435 -5.955 ;
        RECT -64.765 -7.645 -64.435 -7.315 ;
        RECT -64.765 -9.005 -64.435 -8.675 ;
        RECT -64.765 -10.365 -64.435 -10.035 ;
        RECT -64.765 -11.725 -64.435 -11.395 ;
        RECT -64.765 -13.085 -64.435 -12.755 ;
        RECT -64.765 -14.445 -64.435 -14.115 ;
        RECT -64.765 -15.805 -64.435 -15.475 ;
        RECT -64.765 -17.165 -64.435 -16.835 ;
        RECT -64.765 -18.525 -64.435 -18.195 ;
        RECT -64.765 -19.885 -64.435 -19.555 ;
        RECT -64.765 -21.245 -64.435 -20.915 ;
        RECT -64.765 -22.605 -64.435 -22.275 ;
        RECT -64.765 -23.965 -64.435 -23.635 ;
        RECT -64.765 -25.325 -64.435 -24.995 ;
        RECT -64.765 -26.685 -64.435 -26.355 ;
        RECT -64.765 -28.045 -64.435 -27.715 ;
        RECT -64.765 -29.405 -64.435 -29.075 ;
        RECT -64.765 -30.765 -64.435 -30.435 ;
        RECT -64.765 -32.125 -64.435 -31.795 ;
        RECT -64.765 -33.485 -64.435 -33.155 ;
        RECT -64.765 -34.845 -64.435 -34.515 ;
        RECT -64.765 -36.205 -64.435 -35.875 ;
        RECT -64.765 -37.565 -64.435 -37.235 ;
        RECT -64.765 -38.925 -64.435 -38.595 ;
        RECT -64.765 -40.285 -64.435 -39.955 ;
        RECT -64.765 -41.645 -64.435 -41.315 ;
        RECT -64.765 -43.005 -64.435 -42.675 ;
        RECT -64.765 -44.365 -64.435 -44.035 ;
        RECT -64.765 -45.725 -64.435 -45.395 ;
        RECT -64.765 -47.085 -64.435 -46.755 ;
        RECT -64.765 -48.445 -64.435 -48.115 ;
        RECT -64.765 -49.805 -64.435 -49.475 ;
        RECT -64.765 -51.165 -64.435 -50.835 ;
        RECT -64.765 -52.525 -64.435 -52.195 ;
        RECT -64.765 -53.885 -64.435 -53.555 ;
        RECT -64.765 -55.245 -64.435 -54.915 ;
        RECT -64.765 -56.605 -64.435 -56.275 ;
        RECT -64.765 -57.965 -64.435 -57.635 ;
        RECT -64.765 -59.325 -64.435 -58.995 ;
        RECT -64.765 -60.685 -64.435 -60.355 ;
        RECT -64.765 -62.045 -64.435 -61.715 ;
        RECT -64.765 -63.405 -64.435 -63.075 ;
        RECT -64.765 -64.765 -64.435 -64.435 ;
        RECT -64.765 -66.125 -64.435 -65.795 ;
        RECT -64.765 -67.485 -64.435 -67.155 ;
        RECT -64.765 -68.845 -64.435 -68.515 ;
        RECT -64.765 -70.205 -64.435 -69.875 ;
        RECT -64.765 -71.565 -64.435 -71.235 ;
        RECT -64.765 -72.925 -64.435 -72.595 ;
        RECT -64.765 -74.285 -64.435 -73.955 ;
        RECT -64.765 -75.645 -64.435 -75.315 ;
        RECT -64.765 -77.005 -64.435 -76.675 ;
        RECT -64.765 -78.365 -64.435 -78.035 ;
        RECT -64.765 -79.725 -64.435 -79.395 ;
        RECT -64.765 -81.085 -64.435 -80.755 ;
        RECT -64.765 -82.445 -64.435 -82.115 ;
        RECT -64.765 -83.805 -64.435 -83.475 ;
        RECT -64.765 -85.165 -64.435 -84.835 ;
        RECT -64.765 -86.525 -64.435 -86.195 ;
        RECT -64.765 -87.885 -64.435 -87.555 ;
        RECT -64.765 -89.245 -64.435 -88.915 ;
        RECT -64.765 -90.605 -64.435 -90.275 ;
        RECT -64.765 -91.965 -64.435 -91.635 ;
        RECT -64.765 -93.325 -64.435 -92.995 ;
        RECT -64.765 -94.685 -64.435 -94.355 ;
        RECT -64.765 -96.045 -64.435 -95.715 ;
        RECT -64.765 -97.405 -64.435 -97.075 ;
        RECT -64.765 -98.765 -64.435 -98.435 ;
        RECT -64.765 -100.125 -64.435 -99.795 ;
        RECT -64.765 -101.485 -64.435 -101.155 ;
        RECT -64.765 -102.845 -64.435 -102.515 ;
        RECT -64.765 -104.205 -64.435 -103.875 ;
        RECT -64.765 -105.565 -64.435 -105.235 ;
        RECT -64.765 -106.925 -64.435 -106.595 ;
        RECT -64.765 -108.285 -64.435 -107.955 ;
        RECT -64.765 -109.645 -64.435 -109.315 ;
        RECT -64.765 -111.005 -64.435 -110.675 ;
        RECT -64.765 -112.365 -64.435 -112.035 ;
        RECT -64.765 -113.725 -64.435 -113.395 ;
        RECT -64.765 -115.085 -64.435 -114.755 ;
        RECT -64.765 -116.445 -64.435 -116.115 ;
        RECT -64.765 -117.805 -64.435 -117.475 ;
        RECT -64.765 -119.165 -64.435 -118.835 ;
        RECT -64.765 -120.525 -64.435 -120.195 ;
        RECT -64.765 -121.885 -64.435 -121.555 ;
        RECT -64.765 -123.245 -64.435 -122.915 ;
        RECT -64.765 -124.605 -64.435 -124.275 ;
        RECT -64.765 -125.965 -64.435 -125.635 ;
        RECT -64.765 -128.685 -64.435 -128.355 ;
        RECT -64.765 -130.045 -64.435 -129.715 ;
        RECT -64.765 -132.765 -64.435 -132.435 ;
        RECT -64.765 -134.125 -64.435 -133.795 ;
        RECT -64.765 -135.485 -64.435 -135.155 ;
        RECT -64.765 -136.845 -64.435 -136.515 ;
        RECT -64.765 -138.205 -64.435 -137.875 ;
        RECT -64.765 -139.39 -64.435 -139.06 ;
        RECT -64.765 -140.925 -64.435 -140.595 ;
        RECT -64.765 -142.285 -64.435 -141.955 ;
        RECT -64.765 -145.005 -64.435 -144.675 ;
        RECT -64.765 -146.365 -64.435 -146.035 ;
        RECT -64.765 -148.03 -64.435 -147.7 ;
        RECT -64.765 -149.085 -64.435 -148.755 ;
        RECT -64.765 -153.165 -64.435 -152.835 ;
        RECT -64.765 -154.525 -64.435 -154.195 ;
        RECT -64.765 -155.885 -64.435 -155.555 ;
        RECT -64.765 -157.245 -64.435 -156.915 ;
        RECT -64.765 -158.605 -64.435 -158.275 ;
        RECT -64.765 -159.965 -64.435 -159.635 ;
        RECT -64.765 -161.325 -64.435 -160.995 ;
        RECT -64.765 -162.685 -64.435 -162.355 ;
        RECT -64.765 -164.045 -64.435 -163.715 ;
        RECT -64.765 -165.405 -64.435 -165.075 ;
        RECT -64.765 -166.765 -64.435 -166.435 ;
        RECT -64.765 -168.125 -64.435 -167.795 ;
        RECT -64.765 -169.485 -64.435 -169.155 ;
        RECT -64.765 -170.845 -64.435 -170.515 ;
        RECT -64.765 -172.205 -64.435 -171.875 ;
        RECT -64.765 -173.565 -64.435 -173.235 ;
        RECT -64.765 -174.925 -64.435 -174.595 ;
        RECT -64.765 -176.285 -64.435 -175.955 ;
        RECT -64.765 -177.645 -64.435 -177.315 ;
        RECT -64.765 -179.005 -64.435 -178.675 ;
        RECT -64.765 -180.365 -64.435 -180.035 ;
        RECT -64.765 -181.725 -64.435 -181.395 ;
        RECT -64.765 -183.085 -64.435 -182.755 ;
        RECT -64.765 -184.445 -64.435 -184.115 ;
        RECT -64.765 -185.805 -64.435 -185.475 ;
        RECT -64.765 -187.165 -64.435 -186.835 ;
        RECT -64.765 -188.525 -64.435 -188.195 ;
        RECT -64.765 -189.885 -64.435 -189.555 ;
        RECT -64.765 -191.245 -64.435 -190.915 ;
        RECT -64.765 -192.605 -64.435 -192.275 ;
        RECT -64.765 -193.965 -64.435 -193.635 ;
        RECT -64.765 -195.325 -64.435 -194.995 ;
        RECT -64.765 -196.685 -64.435 -196.355 ;
        RECT -64.765 -198.045 -64.435 -197.715 ;
        RECT -64.765 -199.405 -64.435 -199.075 ;
        RECT -64.765 -200.765 -64.435 -200.435 ;
        RECT -64.765 -202.125 -64.435 -201.795 ;
        RECT -64.765 -203.485 -64.435 -203.155 ;
        RECT -64.765 -204.845 -64.435 -204.515 ;
        RECT -64.765 -206.205 -64.435 -205.875 ;
        RECT -64.765 -207.565 -64.435 -207.235 ;
        RECT -64.765 -208.925 -64.435 -208.595 ;
        RECT -64.765 -210.285 -64.435 -209.955 ;
        RECT -64.765 -211.645 -64.435 -211.315 ;
        RECT -64.765 -213.005 -64.435 -212.675 ;
        RECT -64.765 -214.365 -64.435 -214.035 ;
        RECT -64.765 -215.725 -64.435 -215.395 ;
        RECT -64.765 -217.085 -64.435 -216.755 ;
        RECT -64.765 -218.445 -64.435 -218.115 ;
        RECT -64.765 -219.805 -64.435 -219.475 ;
        RECT -64.765 -221.165 -64.435 -220.835 ;
        RECT -64.765 -222.525 -64.435 -222.195 ;
        RECT -64.765 -223.885 -64.435 -223.555 ;
        RECT -64.765 -225.245 -64.435 -224.915 ;
        RECT -64.765 -227.965 -64.435 -227.635 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.925 -232.045 -72.595 -231.715 ;
        RECT -72.925 -233.225 -72.595 -232.895 ;
        RECT -72.925 -234.765 -72.595 -234.435 ;
        RECT -72.925 -236.125 -72.595 -235.795 ;
        RECT -72.925 -237.485 -72.595 -237.155 ;
        RECT -72.925 -238.845 -72.595 -238.515 ;
        RECT -72.925 -241.09 -72.595 -239.96 ;
        RECT -72.92 -241.205 -72.6 -230.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.565 244.04 -71.235 245.17 ;
        RECT -71.565 242.595 -71.235 242.925 ;
        RECT -71.565 241.235 -71.235 241.565 ;
        RECT -71.565 239.875 -71.235 240.205 ;
        RECT -71.565 238.515 -71.235 238.845 ;
        RECT -71.565 237.155 -71.235 237.485 ;
        RECT -71.565 235.795 -71.235 236.125 ;
        RECT -71.565 234.435 -71.235 234.765 ;
        RECT -71.565 233.075 -71.235 233.405 ;
        RECT -71.565 231.715 -71.235 232.045 ;
        RECT -71.565 230.355 -71.235 230.685 ;
        RECT -71.565 228.995 -71.235 229.325 ;
        RECT -71.565 227.635 -71.235 227.965 ;
        RECT -71.565 226.275 -71.235 226.605 ;
        RECT -71.565 224.915 -71.235 225.245 ;
        RECT -71.565 223.555 -71.235 223.885 ;
        RECT -71.565 222.195 -71.235 222.525 ;
        RECT -71.565 220.835 -71.235 221.165 ;
        RECT -71.565 219.475 -71.235 219.805 ;
        RECT -71.565 218.115 -71.235 218.445 ;
        RECT -71.565 216.755 -71.235 217.085 ;
        RECT -71.565 215.395 -71.235 215.725 ;
        RECT -71.565 214.035 -71.235 214.365 ;
        RECT -71.565 212.675 -71.235 213.005 ;
        RECT -71.565 211.315 -71.235 211.645 ;
        RECT -71.565 209.955 -71.235 210.285 ;
        RECT -71.565 208.595 -71.235 208.925 ;
        RECT -71.565 207.235 -71.235 207.565 ;
        RECT -71.565 205.875 -71.235 206.205 ;
        RECT -71.565 204.515 -71.235 204.845 ;
        RECT -71.565 203.155 -71.235 203.485 ;
        RECT -71.565 201.795 -71.235 202.125 ;
        RECT -71.565 200.435 -71.235 200.765 ;
        RECT -71.565 199.075 -71.235 199.405 ;
        RECT -71.565 197.715 -71.235 198.045 ;
        RECT -71.565 196.355 -71.235 196.685 ;
        RECT -71.565 194.995 -71.235 195.325 ;
        RECT -71.565 193.635 -71.235 193.965 ;
        RECT -71.565 192.275 -71.235 192.605 ;
        RECT -71.565 190.915 -71.235 191.245 ;
        RECT -71.565 189.555 -71.235 189.885 ;
        RECT -71.565 188.195 -71.235 188.525 ;
        RECT -71.565 186.835 -71.235 187.165 ;
        RECT -71.565 185.475 -71.235 185.805 ;
        RECT -71.565 184.115 -71.235 184.445 ;
        RECT -71.565 182.755 -71.235 183.085 ;
        RECT -71.565 181.395 -71.235 181.725 ;
        RECT -71.565 180.035 -71.235 180.365 ;
        RECT -71.565 178.675 -71.235 179.005 ;
        RECT -71.565 177.315 -71.235 177.645 ;
        RECT -71.565 175.955 -71.235 176.285 ;
        RECT -71.565 174.595 -71.235 174.925 ;
        RECT -71.565 173.235 -71.235 173.565 ;
        RECT -71.565 171.875 -71.235 172.205 ;
        RECT -71.565 170.515 -71.235 170.845 ;
        RECT -71.565 169.155 -71.235 169.485 ;
        RECT -71.565 167.795 -71.235 168.125 ;
        RECT -71.565 166.435 -71.235 166.765 ;
        RECT -71.565 165.075 -71.235 165.405 ;
        RECT -71.565 163.715 -71.235 164.045 ;
        RECT -71.565 162.355 -71.235 162.685 ;
        RECT -71.565 160.995 -71.235 161.325 ;
        RECT -71.565 159.635 -71.235 159.965 ;
        RECT -71.565 158.275 -71.235 158.605 ;
        RECT -71.565 156.915 -71.235 157.245 ;
        RECT -71.565 155.555 -71.235 155.885 ;
        RECT -71.565 154.195 -71.235 154.525 ;
        RECT -71.565 152.835 -71.235 153.165 ;
        RECT -71.565 151.475 -71.235 151.805 ;
        RECT -71.565 150.115 -71.235 150.445 ;
        RECT -71.565 148.755 -71.235 149.085 ;
        RECT -71.565 147.395 -71.235 147.725 ;
        RECT -71.565 146.035 -71.235 146.365 ;
        RECT -71.565 144.675 -71.235 145.005 ;
        RECT -71.565 143.315 -71.235 143.645 ;
        RECT -71.565 141.955 -71.235 142.285 ;
        RECT -71.565 140.595 -71.235 140.925 ;
        RECT -71.565 139.235 -71.235 139.565 ;
        RECT -71.565 137.875 -71.235 138.205 ;
        RECT -71.565 136.515 -71.235 136.845 ;
        RECT -71.565 135.155 -71.235 135.485 ;
        RECT -71.565 133.795 -71.235 134.125 ;
        RECT -71.565 132.435 -71.235 132.765 ;
        RECT -71.565 131.075 -71.235 131.405 ;
        RECT -71.565 129.715 -71.235 130.045 ;
        RECT -71.565 128.355 -71.235 128.685 ;
        RECT -71.565 126.995 -71.235 127.325 ;
        RECT -71.565 125.635 -71.235 125.965 ;
        RECT -71.565 124.275 -71.235 124.605 ;
        RECT -71.565 122.915 -71.235 123.245 ;
        RECT -71.565 121.555 -71.235 121.885 ;
        RECT -71.565 120.195 -71.235 120.525 ;
        RECT -71.565 118.835 -71.235 119.165 ;
        RECT -71.565 117.475 -71.235 117.805 ;
        RECT -71.565 116.115 -71.235 116.445 ;
        RECT -71.565 114.755 -71.235 115.085 ;
        RECT -71.565 113.395 -71.235 113.725 ;
        RECT -71.565 112.035 -71.235 112.365 ;
        RECT -71.565 110.675 -71.235 111.005 ;
        RECT -71.565 109.315 -71.235 109.645 ;
        RECT -71.565 107.955 -71.235 108.285 ;
        RECT -71.565 106.595 -71.235 106.925 ;
        RECT -71.565 105.235 -71.235 105.565 ;
        RECT -71.565 103.875 -71.235 104.205 ;
        RECT -71.565 102.515 -71.235 102.845 ;
        RECT -71.565 101.155 -71.235 101.485 ;
        RECT -71.565 99.795 -71.235 100.125 ;
        RECT -71.565 98.435 -71.235 98.765 ;
        RECT -71.565 97.075 -71.235 97.405 ;
        RECT -71.565 95.715 -71.235 96.045 ;
        RECT -71.565 94.355 -71.235 94.685 ;
        RECT -71.565 92.995 -71.235 93.325 ;
        RECT -71.565 91.635 -71.235 91.965 ;
        RECT -71.565 90.275 -71.235 90.605 ;
        RECT -71.565 88.915 -71.235 89.245 ;
        RECT -71.565 87.555 -71.235 87.885 ;
        RECT -71.565 86.195 -71.235 86.525 ;
        RECT -71.565 84.835 -71.235 85.165 ;
        RECT -71.565 83.475 -71.235 83.805 ;
        RECT -71.565 82.115 -71.235 82.445 ;
        RECT -71.565 80.755 -71.235 81.085 ;
        RECT -71.565 79.395 -71.235 79.725 ;
        RECT -71.565 78.035 -71.235 78.365 ;
        RECT -71.565 76.675 -71.235 77.005 ;
        RECT -71.565 75.315 -71.235 75.645 ;
        RECT -71.565 73.955 -71.235 74.285 ;
        RECT -71.565 72.595 -71.235 72.925 ;
        RECT -71.565 71.235 -71.235 71.565 ;
        RECT -71.565 69.875 -71.235 70.205 ;
        RECT -71.565 68.515 -71.235 68.845 ;
        RECT -71.565 67.155 -71.235 67.485 ;
        RECT -71.565 65.795 -71.235 66.125 ;
        RECT -71.565 64.435 -71.235 64.765 ;
        RECT -71.565 63.075 -71.235 63.405 ;
        RECT -71.565 61.715 -71.235 62.045 ;
        RECT -71.565 60.355 -71.235 60.685 ;
        RECT -71.565 58.995 -71.235 59.325 ;
        RECT -71.565 57.635 -71.235 57.965 ;
        RECT -71.565 56.275 -71.235 56.605 ;
        RECT -71.565 54.915 -71.235 55.245 ;
        RECT -71.565 53.555 -71.235 53.885 ;
        RECT -71.565 52.195 -71.235 52.525 ;
        RECT -71.565 50.835 -71.235 51.165 ;
        RECT -71.565 49.475 -71.235 49.805 ;
        RECT -71.565 48.115 -71.235 48.445 ;
        RECT -71.565 46.755 -71.235 47.085 ;
        RECT -71.565 45.395 -71.235 45.725 ;
        RECT -71.565 44.035 -71.235 44.365 ;
        RECT -71.565 42.675 -71.235 43.005 ;
        RECT -71.565 41.315 -71.235 41.645 ;
        RECT -71.565 39.955 -71.235 40.285 ;
        RECT -71.565 38.595 -71.235 38.925 ;
        RECT -71.565 37.235 -71.235 37.565 ;
        RECT -71.565 35.875 -71.235 36.205 ;
        RECT -71.565 34.515 -71.235 34.845 ;
        RECT -71.565 33.155 -71.235 33.485 ;
        RECT -71.565 31.795 -71.235 32.125 ;
        RECT -71.565 30.435 -71.235 30.765 ;
        RECT -71.565 29.075 -71.235 29.405 ;
        RECT -71.565 27.715 -71.235 28.045 ;
        RECT -71.565 26.355 -71.235 26.685 ;
        RECT -71.565 24.995 -71.235 25.325 ;
        RECT -71.565 23.635 -71.235 23.965 ;
        RECT -71.565 22.275 -71.235 22.605 ;
        RECT -71.565 20.915 -71.235 21.245 ;
        RECT -71.565 19.555 -71.235 19.885 ;
        RECT -71.565 18.195 -71.235 18.525 ;
        RECT -71.565 16.835 -71.235 17.165 ;
        RECT -71.565 15.475 -71.235 15.805 ;
        RECT -71.565 14.115 -71.235 14.445 ;
        RECT -71.565 12.755 -71.235 13.085 ;
        RECT -71.565 11.395 -71.235 11.725 ;
        RECT -71.565 10.035 -71.235 10.365 ;
        RECT -71.565 8.675 -71.235 9.005 ;
        RECT -71.565 7.315 -71.235 7.645 ;
        RECT -71.565 5.955 -71.235 6.285 ;
        RECT -71.565 4.595 -71.235 4.925 ;
        RECT -71.565 3.235 -71.235 3.565 ;
        RECT -71.565 1.875 -71.235 2.205 ;
        RECT -71.565 0.515 -71.235 0.845 ;
        RECT -71.565 -0.845 -71.235 -0.515 ;
        RECT -71.565 -2.205 -71.235 -1.875 ;
        RECT -71.565 -3.565 -71.235 -3.235 ;
        RECT -71.565 -4.925 -71.235 -4.595 ;
        RECT -71.565 -6.285 -71.235 -5.955 ;
        RECT -71.565 -7.645 -71.235 -7.315 ;
        RECT -71.565 -9.005 -71.235 -8.675 ;
        RECT -71.565 -10.365 -71.235 -10.035 ;
        RECT -71.565 -11.725 -71.235 -11.395 ;
        RECT -71.565 -13.085 -71.235 -12.755 ;
        RECT -71.565 -14.445 -71.235 -14.115 ;
        RECT -71.565 -15.805 -71.235 -15.475 ;
        RECT -71.565 -17.165 -71.235 -16.835 ;
        RECT -71.565 -18.525 -71.235 -18.195 ;
        RECT -71.565 -19.885 -71.235 -19.555 ;
        RECT -71.565 -21.245 -71.235 -20.915 ;
        RECT -71.565 -22.605 -71.235 -22.275 ;
        RECT -71.565 -23.965 -71.235 -23.635 ;
        RECT -71.565 -25.325 -71.235 -24.995 ;
        RECT -71.565 -26.685 -71.235 -26.355 ;
        RECT -71.565 -28.045 -71.235 -27.715 ;
        RECT -71.565 -29.405 -71.235 -29.075 ;
        RECT -71.565 -30.765 -71.235 -30.435 ;
        RECT -71.565 -32.125 -71.235 -31.795 ;
        RECT -71.565 -33.485 -71.235 -33.155 ;
        RECT -71.565 -34.845 -71.235 -34.515 ;
        RECT -71.565 -36.205 -71.235 -35.875 ;
        RECT -71.565 -37.565 -71.235 -37.235 ;
        RECT -71.565 -38.925 -71.235 -38.595 ;
        RECT -71.565 -40.285 -71.235 -39.955 ;
        RECT -71.565 -41.645 -71.235 -41.315 ;
        RECT -71.565 -43.005 -71.235 -42.675 ;
        RECT -71.565 -44.365 -71.235 -44.035 ;
        RECT -71.565 -45.725 -71.235 -45.395 ;
        RECT -71.565 -47.085 -71.235 -46.755 ;
        RECT -71.565 -48.445 -71.235 -48.115 ;
        RECT -71.565 -49.805 -71.235 -49.475 ;
        RECT -71.565 -51.165 -71.235 -50.835 ;
        RECT -71.565 -52.525 -71.235 -52.195 ;
        RECT -71.565 -53.885 -71.235 -53.555 ;
        RECT -71.565 -55.245 -71.235 -54.915 ;
        RECT -71.565 -56.605 -71.235 -56.275 ;
        RECT -71.565 -57.965 -71.235 -57.635 ;
        RECT -71.565 -59.325 -71.235 -58.995 ;
        RECT -71.565 -60.685 -71.235 -60.355 ;
        RECT -71.565 -62.045 -71.235 -61.715 ;
        RECT -71.565 -63.405 -71.235 -63.075 ;
        RECT -71.565 -64.765 -71.235 -64.435 ;
        RECT -71.565 -66.125 -71.235 -65.795 ;
        RECT -71.565 -67.485 -71.235 -67.155 ;
        RECT -71.565 -68.845 -71.235 -68.515 ;
        RECT -71.565 -70.205 -71.235 -69.875 ;
        RECT -71.565 -71.565 -71.235 -71.235 ;
        RECT -71.565 -72.925 -71.235 -72.595 ;
        RECT -71.565 -74.285 -71.235 -73.955 ;
        RECT -71.565 -75.645 -71.235 -75.315 ;
        RECT -71.565 -77.005 -71.235 -76.675 ;
        RECT -71.565 -78.365 -71.235 -78.035 ;
        RECT -71.565 -79.725 -71.235 -79.395 ;
        RECT -71.565 -81.085 -71.235 -80.755 ;
        RECT -71.565 -82.445 -71.235 -82.115 ;
        RECT -71.565 -83.805 -71.235 -83.475 ;
        RECT -71.565 -85.165 -71.235 -84.835 ;
        RECT -71.565 -86.525 -71.235 -86.195 ;
        RECT -71.565 -87.885 -71.235 -87.555 ;
        RECT -71.565 -89.245 -71.235 -88.915 ;
        RECT -71.565 -90.605 -71.235 -90.275 ;
        RECT -71.565 -91.965 -71.235 -91.635 ;
        RECT -71.565 -93.325 -71.235 -92.995 ;
        RECT -71.565 -94.685 -71.235 -94.355 ;
        RECT -71.565 -96.045 -71.235 -95.715 ;
        RECT -71.565 -97.405 -71.235 -97.075 ;
        RECT -71.565 -98.765 -71.235 -98.435 ;
        RECT -71.565 -100.125 -71.235 -99.795 ;
        RECT -71.565 -101.485 -71.235 -101.155 ;
        RECT -71.565 -102.845 -71.235 -102.515 ;
        RECT -71.565 -104.205 -71.235 -103.875 ;
        RECT -71.565 -105.565 -71.235 -105.235 ;
        RECT -71.565 -106.925 -71.235 -106.595 ;
        RECT -71.565 -108.285 -71.235 -107.955 ;
        RECT -71.565 -109.645 -71.235 -109.315 ;
        RECT -71.565 -111.005 -71.235 -110.675 ;
        RECT -71.565 -112.365 -71.235 -112.035 ;
        RECT -71.565 -113.725 -71.235 -113.395 ;
        RECT -71.565 -115.085 -71.235 -114.755 ;
        RECT -71.565 -116.445 -71.235 -116.115 ;
        RECT -71.565 -117.805 -71.235 -117.475 ;
        RECT -71.565 -119.165 -71.235 -118.835 ;
        RECT -71.565 -120.525 -71.235 -120.195 ;
        RECT -71.565 -121.885 -71.235 -121.555 ;
        RECT -71.565 -123.245 -71.235 -122.915 ;
        RECT -71.565 -124.605 -71.235 -124.275 ;
        RECT -71.565 -125.965 -71.235 -125.635 ;
        RECT -71.565 -127.325 -71.235 -126.995 ;
        RECT -71.565 -128.685 -71.235 -128.355 ;
        RECT -71.565 -130.045 -71.235 -129.715 ;
        RECT -71.565 -131.405 -71.235 -131.075 ;
        RECT -71.565 -132.765 -71.235 -132.435 ;
        RECT -71.565 -134.125 -71.235 -133.795 ;
        RECT -71.565 -135.485 -71.235 -135.155 ;
        RECT -71.565 -136.845 -71.235 -136.515 ;
        RECT -71.565 -138.205 -71.235 -137.875 ;
        RECT -71.565 -139.565 -71.235 -139.235 ;
        RECT -71.565 -140.925 -71.235 -140.595 ;
        RECT -71.565 -142.285 -71.235 -141.955 ;
        RECT -71.565 -143.645 -71.235 -143.315 ;
        RECT -71.565 -145.005 -71.235 -144.675 ;
        RECT -71.565 -146.365 -71.235 -146.035 ;
        RECT -71.565 -147.725 -71.235 -147.395 ;
        RECT -71.565 -149.085 -71.235 -148.755 ;
        RECT -71.56 -151.12 -71.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.565 -161.325 -71.235 -160.995 ;
        RECT -71.565 -162.685 -71.235 -162.355 ;
        RECT -71.565 -164.045 -71.235 -163.715 ;
        RECT -71.565 -165.405 -71.235 -165.075 ;
        RECT -71.565 -166.765 -71.235 -166.435 ;
        RECT -71.565 -168.125 -71.235 -167.795 ;
        RECT -71.565 -169.485 -71.235 -169.155 ;
        RECT -71.565 -170.845 -71.235 -170.515 ;
        RECT -71.565 -172.205 -71.235 -171.875 ;
        RECT -71.565 -173.565 -71.235 -173.235 ;
        RECT -71.565 -174.925 -71.235 -174.595 ;
        RECT -71.565 -176.285 -71.235 -175.955 ;
        RECT -71.565 -177.645 -71.235 -177.315 ;
        RECT -71.565 -179.005 -71.235 -178.675 ;
        RECT -71.565 -180.365 -71.235 -180.035 ;
        RECT -71.565 -181.725 -71.235 -181.395 ;
        RECT -71.565 -183.085 -71.235 -182.755 ;
        RECT -71.565 -184.445 -71.235 -184.115 ;
        RECT -71.565 -185.805 -71.235 -185.475 ;
        RECT -71.565 -187.165 -71.235 -186.835 ;
        RECT -71.565 -188.525 -71.235 -188.195 ;
        RECT -71.565 -189.885 -71.235 -189.555 ;
        RECT -71.565 -191.245 -71.235 -190.915 ;
        RECT -71.565 -192.605 -71.235 -192.275 ;
        RECT -71.565 -193.965 -71.235 -193.635 ;
        RECT -71.565 -195.325 -71.235 -194.995 ;
        RECT -71.565 -196.685 -71.235 -196.355 ;
        RECT -71.565 -198.045 -71.235 -197.715 ;
        RECT -71.565 -199.405 -71.235 -199.075 ;
        RECT -71.565 -200.765 -71.235 -200.435 ;
        RECT -71.565 -202.125 -71.235 -201.795 ;
        RECT -71.565 -203.485 -71.235 -203.155 ;
        RECT -71.565 -204.845 -71.235 -204.515 ;
        RECT -71.565 -206.205 -71.235 -205.875 ;
        RECT -71.565 -207.565 -71.235 -207.235 ;
        RECT -71.565 -208.925 -71.235 -208.595 ;
        RECT -71.565 -210.285 -71.235 -209.955 ;
        RECT -71.565 -211.645 -71.235 -211.315 ;
        RECT -71.565 -213.005 -71.235 -212.675 ;
        RECT -71.565 -214.365 -71.235 -214.035 ;
        RECT -71.565 -215.725 -71.235 -215.395 ;
        RECT -71.565 -217.085 -71.235 -216.755 ;
        RECT -71.565 -218.445 -71.235 -218.115 ;
        RECT -71.565 -219.805 -71.235 -219.475 ;
        RECT -71.565 -221.165 -71.235 -220.835 ;
        RECT -71.565 -222.525 -71.235 -222.195 ;
        RECT -71.565 -223.885 -71.235 -223.555 ;
        RECT -71.565 -225.245 -71.235 -224.915 ;
        RECT -71.565 -227.965 -71.235 -227.635 ;
        RECT -71.56 -229.32 -71.24 -160.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.205 244.04 -69.875 245.17 ;
        RECT -70.205 242.595 -69.875 242.925 ;
        RECT -70.205 241.235 -69.875 241.565 ;
        RECT -70.205 239.875 -69.875 240.205 ;
        RECT -70.205 238.515 -69.875 238.845 ;
        RECT -70.205 237.155 -69.875 237.485 ;
        RECT -70.205 235.795 -69.875 236.125 ;
        RECT -70.205 234.435 -69.875 234.765 ;
        RECT -70.205 233.075 -69.875 233.405 ;
        RECT -70.205 231.715 -69.875 232.045 ;
        RECT -70.205 230.355 -69.875 230.685 ;
        RECT -70.205 228.995 -69.875 229.325 ;
        RECT -70.205 227.635 -69.875 227.965 ;
        RECT -70.205 226.275 -69.875 226.605 ;
        RECT -70.205 224.915 -69.875 225.245 ;
        RECT -70.205 223.555 -69.875 223.885 ;
        RECT -70.205 222.195 -69.875 222.525 ;
        RECT -70.205 220.835 -69.875 221.165 ;
        RECT -70.205 219.475 -69.875 219.805 ;
        RECT -70.205 218.115 -69.875 218.445 ;
        RECT -70.205 216.755 -69.875 217.085 ;
        RECT -70.205 215.395 -69.875 215.725 ;
        RECT -70.205 214.035 -69.875 214.365 ;
        RECT -70.205 212.675 -69.875 213.005 ;
        RECT -70.205 211.315 -69.875 211.645 ;
        RECT -70.205 209.955 -69.875 210.285 ;
        RECT -70.205 208.595 -69.875 208.925 ;
        RECT -70.205 207.235 -69.875 207.565 ;
        RECT -70.205 205.875 -69.875 206.205 ;
        RECT -70.205 204.515 -69.875 204.845 ;
        RECT -70.205 203.155 -69.875 203.485 ;
        RECT -70.205 201.795 -69.875 202.125 ;
        RECT -70.205 200.435 -69.875 200.765 ;
        RECT -70.205 199.075 -69.875 199.405 ;
        RECT -70.205 197.715 -69.875 198.045 ;
        RECT -70.205 196.355 -69.875 196.685 ;
        RECT -70.205 194.995 -69.875 195.325 ;
        RECT -70.205 193.635 -69.875 193.965 ;
        RECT -70.205 192.275 -69.875 192.605 ;
        RECT -70.205 190.915 -69.875 191.245 ;
        RECT -70.205 189.555 -69.875 189.885 ;
        RECT -70.205 188.195 -69.875 188.525 ;
        RECT -70.205 186.835 -69.875 187.165 ;
        RECT -70.205 185.475 -69.875 185.805 ;
        RECT -70.205 184.115 -69.875 184.445 ;
        RECT -70.205 182.755 -69.875 183.085 ;
        RECT -70.205 181.395 -69.875 181.725 ;
        RECT -70.205 180.035 -69.875 180.365 ;
        RECT -70.205 178.675 -69.875 179.005 ;
        RECT -70.205 177.315 -69.875 177.645 ;
        RECT -70.205 175.955 -69.875 176.285 ;
        RECT -70.205 174.595 -69.875 174.925 ;
        RECT -70.205 173.235 -69.875 173.565 ;
        RECT -70.205 171.875 -69.875 172.205 ;
        RECT -70.205 170.515 -69.875 170.845 ;
        RECT -70.205 169.155 -69.875 169.485 ;
        RECT -70.205 167.795 -69.875 168.125 ;
        RECT -70.205 166.435 -69.875 166.765 ;
        RECT -70.205 165.075 -69.875 165.405 ;
        RECT -70.205 163.715 -69.875 164.045 ;
        RECT -70.205 162.355 -69.875 162.685 ;
        RECT -70.205 160.995 -69.875 161.325 ;
        RECT -70.205 159.635 -69.875 159.965 ;
        RECT -70.205 158.275 -69.875 158.605 ;
        RECT -70.205 156.915 -69.875 157.245 ;
        RECT -70.205 155.555 -69.875 155.885 ;
        RECT -70.205 154.195 -69.875 154.525 ;
        RECT -70.205 152.835 -69.875 153.165 ;
        RECT -70.205 151.475 -69.875 151.805 ;
        RECT -70.205 150.115 -69.875 150.445 ;
        RECT -70.205 148.755 -69.875 149.085 ;
        RECT -70.205 147.395 -69.875 147.725 ;
        RECT -70.205 146.035 -69.875 146.365 ;
        RECT -70.205 144.675 -69.875 145.005 ;
        RECT -70.205 143.315 -69.875 143.645 ;
        RECT -70.205 141.955 -69.875 142.285 ;
        RECT -70.205 140.595 -69.875 140.925 ;
        RECT -70.205 139.235 -69.875 139.565 ;
        RECT -70.205 137.875 -69.875 138.205 ;
        RECT -70.205 136.515 -69.875 136.845 ;
        RECT -70.205 135.155 -69.875 135.485 ;
        RECT -70.205 133.795 -69.875 134.125 ;
        RECT -70.205 132.435 -69.875 132.765 ;
        RECT -70.205 131.075 -69.875 131.405 ;
        RECT -70.205 129.715 -69.875 130.045 ;
        RECT -70.205 128.355 -69.875 128.685 ;
        RECT -70.205 126.995 -69.875 127.325 ;
        RECT -70.205 125.635 -69.875 125.965 ;
        RECT -70.205 124.275 -69.875 124.605 ;
        RECT -70.205 122.915 -69.875 123.245 ;
        RECT -70.205 121.555 -69.875 121.885 ;
        RECT -70.205 120.195 -69.875 120.525 ;
        RECT -70.205 118.835 -69.875 119.165 ;
        RECT -70.205 117.475 -69.875 117.805 ;
        RECT -70.205 116.115 -69.875 116.445 ;
        RECT -70.205 114.755 -69.875 115.085 ;
        RECT -70.205 113.395 -69.875 113.725 ;
        RECT -70.205 112.035 -69.875 112.365 ;
        RECT -70.205 110.675 -69.875 111.005 ;
        RECT -70.205 109.315 -69.875 109.645 ;
        RECT -70.205 107.955 -69.875 108.285 ;
        RECT -70.205 106.595 -69.875 106.925 ;
        RECT -70.205 105.235 -69.875 105.565 ;
        RECT -70.205 103.875 -69.875 104.205 ;
        RECT -70.205 102.515 -69.875 102.845 ;
        RECT -70.205 101.155 -69.875 101.485 ;
        RECT -70.205 99.795 -69.875 100.125 ;
        RECT -70.205 98.435 -69.875 98.765 ;
        RECT -70.205 97.075 -69.875 97.405 ;
        RECT -70.205 95.715 -69.875 96.045 ;
        RECT -70.205 94.355 -69.875 94.685 ;
        RECT -70.205 92.995 -69.875 93.325 ;
        RECT -70.205 91.635 -69.875 91.965 ;
        RECT -70.205 90.275 -69.875 90.605 ;
        RECT -70.205 88.915 -69.875 89.245 ;
        RECT -70.205 87.555 -69.875 87.885 ;
        RECT -70.205 86.195 -69.875 86.525 ;
        RECT -70.205 84.835 -69.875 85.165 ;
        RECT -70.205 83.475 -69.875 83.805 ;
        RECT -70.205 82.115 -69.875 82.445 ;
        RECT -70.205 80.755 -69.875 81.085 ;
        RECT -70.205 79.395 -69.875 79.725 ;
        RECT -70.205 78.035 -69.875 78.365 ;
        RECT -70.205 76.675 -69.875 77.005 ;
        RECT -70.205 75.315 -69.875 75.645 ;
        RECT -70.205 73.955 -69.875 74.285 ;
        RECT -70.205 72.595 -69.875 72.925 ;
        RECT -70.205 71.235 -69.875 71.565 ;
        RECT -70.205 69.875 -69.875 70.205 ;
        RECT -70.205 68.515 -69.875 68.845 ;
        RECT -70.205 67.155 -69.875 67.485 ;
        RECT -70.205 65.795 -69.875 66.125 ;
        RECT -70.205 64.435 -69.875 64.765 ;
        RECT -70.205 63.075 -69.875 63.405 ;
        RECT -70.205 61.715 -69.875 62.045 ;
        RECT -70.205 60.355 -69.875 60.685 ;
        RECT -70.205 58.995 -69.875 59.325 ;
        RECT -70.205 57.635 -69.875 57.965 ;
        RECT -70.205 56.275 -69.875 56.605 ;
        RECT -70.205 54.915 -69.875 55.245 ;
        RECT -70.205 53.555 -69.875 53.885 ;
        RECT -70.205 52.195 -69.875 52.525 ;
        RECT -70.205 50.835 -69.875 51.165 ;
        RECT -70.205 49.475 -69.875 49.805 ;
        RECT -70.205 48.115 -69.875 48.445 ;
        RECT -70.205 46.755 -69.875 47.085 ;
        RECT -70.205 45.395 -69.875 45.725 ;
        RECT -70.205 44.035 -69.875 44.365 ;
        RECT -70.205 42.675 -69.875 43.005 ;
        RECT -70.205 41.315 -69.875 41.645 ;
        RECT -70.205 39.955 -69.875 40.285 ;
        RECT -70.205 38.595 -69.875 38.925 ;
        RECT -70.205 37.235 -69.875 37.565 ;
        RECT -70.205 35.875 -69.875 36.205 ;
        RECT -70.205 34.515 -69.875 34.845 ;
        RECT -70.205 33.155 -69.875 33.485 ;
        RECT -70.205 31.795 -69.875 32.125 ;
        RECT -70.205 30.435 -69.875 30.765 ;
        RECT -70.205 29.075 -69.875 29.405 ;
        RECT -70.205 27.715 -69.875 28.045 ;
        RECT -70.205 26.355 -69.875 26.685 ;
        RECT -70.205 24.995 -69.875 25.325 ;
        RECT -70.205 23.635 -69.875 23.965 ;
        RECT -70.205 22.275 -69.875 22.605 ;
        RECT -70.205 20.915 -69.875 21.245 ;
        RECT -70.205 19.555 -69.875 19.885 ;
        RECT -70.205 18.195 -69.875 18.525 ;
        RECT -70.205 16.835 -69.875 17.165 ;
        RECT -70.205 15.475 -69.875 15.805 ;
        RECT -70.205 14.115 -69.875 14.445 ;
        RECT -70.205 12.755 -69.875 13.085 ;
        RECT -70.205 11.395 -69.875 11.725 ;
        RECT -70.205 10.035 -69.875 10.365 ;
        RECT -70.205 8.675 -69.875 9.005 ;
        RECT -70.205 7.315 -69.875 7.645 ;
        RECT -70.205 5.955 -69.875 6.285 ;
        RECT -70.205 4.595 -69.875 4.925 ;
        RECT -70.205 3.235 -69.875 3.565 ;
        RECT -70.205 1.875 -69.875 2.205 ;
        RECT -70.205 0.515 -69.875 0.845 ;
        RECT -70.205 -0.845 -69.875 -0.515 ;
        RECT -70.205 -2.205 -69.875 -1.875 ;
        RECT -70.205 -3.565 -69.875 -3.235 ;
        RECT -70.205 -4.925 -69.875 -4.595 ;
        RECT -70.205 -6.285 -69.875 -5.955 ;
        RECT -70.205 -7.645 -69.875 -7.315 ;
        RECT -70.205 -9.005 -69.875 -8.675 ;
        RECT -70.205 -10.365 -69.875 -10.035 ;
        RECT -70.205 -11.725 -69.875 -11.395 ;
        RECT -70.205 -13.085 -69.875 -12.755 ;
        RECT -70.205 -14.445 -69.875 -14.115 ;
        RECT -70.205 -15.805 -69.875 -15.475 ;
        RECT -70.205 -17.165 -69.875 -16.835 ;
        RECT -70.205 -18.525 -69.875 -18.195 ;
        RECT -70.205 -19.885 -69.875 -19.555 ;
        RECT -70.205 -21.245 -69.875 -20.915 ;
        RECT -70.205 -22.605 -69.875 -22.275 ;
        RECT -70.205 -23.965 -69.875 -23.635 ;
        RECT -70.205 -25.325 -69.875 -24.995 ;
        RECT -70.205 -26.685 -69.875 -26.355 ;
        RECT -70.205 -28.045 -69.875 -27.715 ;
        RECT -70.205 -29.405 -69.875 -29.075 ;
        RECT -70.205 -30.765 -69.875 -30.435 ;
        RECT -70.205 -32.125 -69.875 -31.795 ;
        RECT -70.205 -33.485 -69.875 -33.155 ;
        RECT -70.205 -34.845 -69.875 -34.515 ;
        RECT -70.205 -36.205 -69.875 -35.875 ;
        RECT -70.205 -37.565 -69.875 -37.235 ;
        RECT -70.205 -38.925 -69.875 -38.595 ;
        RECT -70.205 -40.285 -69.875 -39.955 ;
        RECT -70.205 -41.645 -69.875 -41.315 ;
        RECT -70.205 -43.005 -69.875 -42.675 ;
        RECT -70.205 -44.365 -69.875 -44.035 ;
        RECT -70.205 -45.725 -69.875 -45.395 ;
        RECT -70.205 -47.085 -69.875 -46.755 ;
        RECT -70.205 -48.445 -69.875 -48.115 ;
        RECT -70.205 -49.805 -69.875 -49.475 ;
        RECT -70.205 -51.165 -69.875 -50.835 ;
        RECT -70.205 -52.525 -69.875 -52.195 ;
        RECT -70.205 -53.885 -69.875 -53.555 ;
        RECT -70.205 -55.245 -69.875 -54.915 ;
        RECT -70.205 -56.605 -69.875 -56.275 ;
        RECT -70.205 -57.965 -69.875 -57.635 ;
        RECT -70.205 -59.325 -69.875 -58.995 ;
        RECT -70.205 -60.685 -69.875 -60.355 ;
        RECT -70.205 -62.045 -69.875 -61.715 ;
        RECT -70.205 -63.405 -69.875 -63.075 ;
        RECT -70.205 -64.765 -69.875 -64.435 ;
        RECT -70.205 -66.125 -69.875 -65.795 ;
        RECT -70.205 -67.485 -69.875 -67.155 ;
        RECT -70.205 -68.845 -69.875 -68.515 ;
        RECT -70.205 -70.205 -69.875 -69.875 ;
        RECT -70.205 -71.565 -69.875 -71.235 ;
        RECT -70.205 -72.925 -69.875 -72.595 ;
        RECT -70.205 -74.285 -69.875 -73.955 ;
        RECT -70.205 -75.645 -69.875 -75.315 ;
        RECT -70.205 -77.005 -69.875 -76.675 ;
        RECT -70.205 -78.365 -69.875 -78.035 ;
        RECT -70.205 -79.725 -69.875 -79.395 ;
        RECT -70.205 -81.085 -69.875 -80.755 ;
        RECT -70.205 -82.445 -69.875 -82.115 ;
        RECT -70.205 -83.805 -69.875 -83.475 ;
        RECT -70.205 -85.165 -69.875 -84.835 ;
        RECT -70.205 -86.525 -69.875 -86.195 ;
        RECT -70.205 -87.885 -69.875 -87.555 ;
        RECT -70.205 -89.245 -69.875 -88.915 ;
        RECT -70.205 -90.605 -69.875 -90.275 ;
        RECT -70.205 -91.965 -69.875 -91.635 ;
        RECT -70.205 -93.325 -69.875 -92.995 ;
        RECT -70.205 -94.685 -69.875 -94.355 ;
        RECT -70.205 -96.045 -69.875 -95.715 ;
        RECT -70.205 -97.405 -69.875 -97.075 ;
        RECT -70.205 -98.765 -69.875 -98.435 ;
        RECT -70.205 -100.125 -69.875 -99.795 ;
        RECT -70.205 -101.485 -69.875 -101.155 ;
        RECT -70.205 -102.845 -69.875 -102.515 ;
        RECT -70.205 -104.205 -69.875 -103.875 ;
        RECT -70.205 -105.565 -69.875 -105.235 ;
        RECT -70.205 -106.925 -69.875 -106.595 ;
        RECT -70.205 -108.285 -69.875 -107.955 ;
        RECT -70.205 -109.645 -69.875 -109.315 ;
        RECT -70.205 -111.005 -69.875 -110.675 ;
        RECT -70.205 -112.365 -69.875 -112.035 ;
        RECT -70.205 -113.725 -69.875 -113.395 ;
        RECT -70.205 -115.085 -69.875 -114.755 ;
        RECT -70.205 -116.445 -69.875 -116.115 ;
        RECT -70.205 -117.805 -69.875 -117.475 ;
        RECT -70.205 -119.165 -69.875 -118.835 ;
        RECT -70.205 -120.525 -69.875 -120.195 ;
        RECT -70.205 -121.885 -69.875 -121.555 ;
        RECT -70.205 -123.245 -69.875 -122.915 ;
        RECT -70.205 -124.605 -69.875 -124.275 ;
        RECT -70.205 -125.965 -69.875 -125.635 ;
        RECT -70.205 -127.325 -69.875 -126.995 ;
        RECT -70.205 -128.685 -69.875 -128.355 ;
        RECT -70.205 -130.045 -69.875 -129.715 ;
        RECT -70.205 -132.765 -69.875 -132.435 ;
        RECT -70.205 -134.125 -69.875 -133.795 ;
        RECT -70.205 -135.485 -69.875 -135.155 ;
        RECT -70.205 -136.845 -69.875 -136.515 ;
        RECT -70.205 -138.205 -69.875 -137.875 ;
        RECT -70.205 -139.39 -69.875 -139.06 ;
        RECT -70.205 -140.925 -69.875 -140.595 ;
        RECT -70.205 -142.285 -69.875 -141.955 ;
        RECT -70.205 -145.005 -69.875 -144.675 ;
        RECT -70.205 -146.365 -69.875 -146.035 ;
        RECT -70.205 -148.03 -69.875 -147.7 ;
        RECT -70.205 -149.085 -69.875 -148.755 ;
        RECT -70.205 -153.165 -69.875 -152.835 ;
        RECT -70.205 -154.525 -69.875 -154.195 ;
        RECT -70.205 -155.885 -69.875 -155.555 ;
        RECT -70.205 -157.245 -69.875 -156.915 ;
        RECT -70.205 -158.605 -69.875 -158.275 ;
        RECT -70.205 -159.965 -69.875 -159.635 ;
        RECT -70.205 -161.325 -69.875 -160.995 ;
        RECT -70.205 -162.685 -69.875 -162.355 ;
        RECT -70.205 -164.045 -69.875 -163.715 ;
        RECT -70.205 -165.405 -69.875 -165.075 ;
        RECT -70.205 -166.765 -69.875 -166.435 ;
        RECT -70.205 -168.125 -69.875 -167.795 ;
        RECT -70.205 -169.485 -69.875 -169.155 ;
        RECT -70.205 -170.845 -69.875 -170.515 ;
        RECT -70.205 -172.205 -69.875 -171.875 ;
        RECT -70.205 -173.565 -69.875 -173.235 ;
        RECT -70.205 -174.925 -69.875 -174.595 ;
        RECT -70.205 -176.285 -69.875 -175.955 ;
        RECT -70.205 -177.645 -69.875 -177.315 ;
        RECT -70.205 -179.005 -69.875 -178.675 ;
        RECT -70.205 -180.365 -69.875 -180.035 ;
        RECT -70.205 -181.725 -69.875 -181.395 ;
        RECT -70.205 -183.085 -69.875 -182.755 ;
        RECT -70.205 -184.445 -69.875 -184.115 ;
        RECT -70.205 -185.805 -69.875 -185.475 ;
        RECT -70.205 -187.165 -69.875 -186.835 ;
        RECT -70.205 -188.525 -69.875 -188.195 ;
        RECT -70.205 -189.885 -69.875 -189.555 ;
        RECT -70.205 -191.245 -69.875 -190.915 ;
        RECT -70.205 -192.605 -69.875 -192.275 ;
        RECT -70.205 -193.965 -69.875 -193.635 ;
        RECT -70.205 -195.325 -69.875 -194.995 ;
        RECT -70.205 -196.685 -69.875 -196.355 ;
        RECT -70.205 -198.045 -69.875 -197.715 ;
        RECT -70.205 -199.405 -69.875 -199.075 ;
        RECT -70.205 -200.765 -69.875 -200.435 ;
        RECT -70.205 -202.125 -69.875 -201.795 ;
        RECT -70.205 -203.485 -69.875 -203.155 ;
        RECT -70.205 -204.845 -69.875 -204.515 ;
        RECT -70.205 -206.205 -69.875 -205.875 ;
        RECT -70.205 -207.565 -69.875 -207.235 ;
        RECT -70.205 -208.925 -69.875 -208.595 ;
        RECT -70.205 -210.285 -69.875 -209.955 ;
        RECT -70.205 -211.645 -69.875 -211.315 ;
        RECT -70.205 -213.005 -69.875 -212.675 ;
        RECT -70.205 -214.365 -69.875 -214.035 ;
        RECT -70.205 -215.725 -69.875 -215.395 ;
        RECT -70.205 -217.085 -69.875 -216.755 ;
        RECT -70.205 -218.445 -69.875 -218.115 ;
        RECT -70.205 -219.805 -69.875 -219.475 ;
        RECT -70.205 -221.165 -69.875 -220.835 ;
        RECT -70.205 -222.525 -69.875 -222.195 ;
        RECT -70.205 -223.885 -69.875 -223.555 ;
        RECT -70.205 -225.245 -69.875 -224.915 ;
        RECT -70.205 -227.965 -69.875 -227.635 ;
        RECT -70.205 -230.685 -69.875 -230.355 ;
        RECT -70.205 -232.045 -69.875 -231.715 ;
        RECT -70.205 -233.225 -69.875 -232.895 ;
        RECT -70.205 -234.765 -69.875 -234.435 ;
        RECT -70.205 -236.125 -69.875 -235.795 ;
        RECT -70.205 -237.485 -69.875 -237.155 ;
        RECT -70.205 -238.845 -69.875 -238.515 ;
        RECT -70.205 -241.09 -69.875 -239.96 ;
        RECT -70.2 -241.205 -69.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.845 -158.605 -68.515 -158.275 ;
        RECT -68.845 -159.965 -68.515 -159.635 ;
        RECT -68.845 -161.325 -68.515 -160.995 ;
        RECT -68.845 -162.685 -68.515 -162.355 ;
        RECT -68.845 -164.045 -68.515 -163.715 ;
        RECT -68.845 -165.405 -68.515 -165.075 ;
        RECT -68.845 -166.765 -68.515 -166.435 ;
        RECT -68.845 -168.125 -68.515 -167.795 ;
        RECT -68.845 -169.485 -68.515 -169.155 ;
        RECT -68.845 -170.845 -68.515 -170.515 ;
        RECT -68.845 -172.205 -68.515 -171.875 ;
        RECT -68.845 -173.565 -68.515 -173.235 ;
        RECT -68.845 -174.925 -68.515 -174.595 ;
        RECT -68.845 -176.285 -68.515 -175.955 ;
        RECT -68.845 -177.645 -68.515 -177.315 ;
        RECT -68.845 -179.005 -68.515 -178.675 ;
        RECT -68.845 -180.365 -68.515 -180.035 ;
        RECT -68.845 -181.725 -68.515 -181.395 ;
        RECT -68.845 -183.085 -68.515 -182.755 ;
        RECT -68.845 -184.445 -68.515 -184.115 ;
        RECT -68.845 -185.805 -68.515 -185.475 ;
        RECT -68.845 -187.165 -68.515 -186.835 ;
        RECT -68.845 -188.525 -68.515 -188.195 ;
        RECT -68.845 -189.885 -68.515 -189.555 ;
        RECT -68.845 -191.245 -68.515 -190.915 ;
        RECT -68.845 -192.605 -68.515 -192.275 ;
        RECT -68.845 -193.965 -68.515 -193.635 ;
        RECT -68.845 -195.325 -68.515 -194.995 ;
        RECT -68.845 -196.685 -68.515 -196.355 ;
        RECT -68.845 -198.045 -68.515 -197.715 ;
        RECT -68.845 -199.405 -68.515 -199.075 ;
        RECT -68.845 -200.765 -68.515 -200.435 ;
        RECT -68.845 -202.125 -68.515 -201.795 ;
        RECT -68.845 -203.485 -68.515 -203.155 ;
        RECT -68.845 -204.845 -68.515 -204.515 ;
        RECT -68.845 -206.205 -68.515 -205.875 ;
        RECT -68.845 -207.565 -68.515 -207.235 ;
        RECT -68.845 -208.925 -68.515 -208.595 ;
        RECT -68.845 -210.285 -68.515 -209.955 ;
        RECT -68.845 -211.645 -68.515 -211.315 ;
        RECT -68.845 -213.005 -68.515 -212.675 ;
        RECT -68.845 -214.365 -68.515 -214.035 ;
        RECT -68.845 -215.725 -68.515 -215.395 ;
        RECT -68.845 -217.085 -68.515 -216.755 ;
        RECT -68.845 -218.445 -68.515 -218.115 ;
        RECT -68.845 -219.805 -68.515 -219.475 ;
        RECT -68.845 -221.165 -68.515 -220.835 ;
        RECT -68.845 -222.525 -68.515 -222.195 ;
        RECT -68.845 -223.885 -68.515 -223.555 ;
        RECT -68.845 -225.245 -68.515 -224.915 ;
        RECT -68.845 -227.965 -68.515 -227.635 ;
        RECT -68.845 -230.685 -68.515 -230.355 ;
        RECT -68.845 -232.045 -68.515 -231.715 ;
        RECT -68.845 -233.225 -68.515 -232.895 ;
        RECT -68.845 -234.765 -68.515 -234.435 ;
        RECT -68.845 -236.125 -68.515 -235.795 ;
        RECT -68.845 -237.485 -68.515 -237.155 ;
        RECT -68.845 -238.845 -68.515 -238.515 ;
        RECT -68.845 -241.09 -68.515 -239.96 ;
        RECT -68.84 -241.205 -68.52 245.285 ;
        RECT -68.845 244.04 -68.515 245.17 ;
        RECT -68.845 242.595 -68.515 242.925 ;
        RECT -68.845 241.235 -68.515 241.565 ;
        RECT -68.845 239.875 -68.515 240.205 ;
        RECT -68.845 238.515 -68.515 238.845 ;
        RECT -68.845 237.155 -68.515 237.485 ;
        RECT -68.845 235.795 -68.515 236.125 ;
        RECT -68.845 234.435 -68.515 234.765 ;
        RECT -68.845 233.075 -68.515 233.405 ;
        RECT -68.845 231.715 -68.515 232.045 ;
        RECT -68.845 230.355 -68.515 230.685 ;
        RECT -68.845 228.995 -68.515 229.325 ;
        RECT -68.845 227.635 -68.515 227.965 ;
        RECT -68.845 226.275 -68.515 226.605 ;
        RECT -68.845 224.915 -68.515 225.245 ;
        RECT -68.845 223.555 -68.515 223.885 ;
        RECT -68.845 222.195 -68.515 222.525 ;
        RECT -68.845 220.835 -68.515 221.165 ;
        RECT -68.845 219.475 -68.515 219.805 ;
        RECT -68.845 218.115 -68.515 218.445 ;
        RECT -68.845 216.755 -68.515 217.085 ;
        RECT -68.845 215.395 -68.515 215.725 ;
        RECT -68.845 214.035 -68.515 214.365 ;
        RECT -68.845 212.675 -68.515 213.005 ;
        RECT -68.845 211.315 -68.515 211.645 ;
        RECT -68.845 209.955 -68.515 210.285 ;
        RECT -68.845 208.595 -68.515 208.925 ;
        RECT -68.845 207.235 -68.515 207.565 ;
        RECT -68.845 205.875 -68.515 206.205 ;
        RECT -68.845 204.515 -68.515 204.845 ;
        RECT -68.845 203.155 -68.515 203.485 ;
        RECT -68.845 201.795 -68.515 202.125 ;
        RECT -68.845 200.435 -68.515 200.765 ;
        RECT -68.845 199.075 -68.515 199.405 ;
        RECT -68.845 197.715 -68.515 198.045 ;
        RECT -68.845 196.355 -68.515 196.685 ;
        RECT -68.845 194.995 -68.515 195.325 ;
        RECT -68.845 193.635 -68.515 193.965 ;
        RECT -68.845 192.275 -68.515 192.605 ;
        RECT -68.845 190.915 -68.515 191.245 ;
        RECT -68.845 189.555 -68.515 189.885 ;
        RECT -68.845 188.195 -68.515 188.525 ;
        RECT -68.845 186.835 -68.515 187.165 ;
        RECT -68.845 185.475 -68.515 185.805 ;
        RECT -68.845 184.115 -68.515 184.445 ;
        RECT -68.845 182.755 -68.515 183.085 ;
        RECT -68.845 181.395 -68.515 181.725 ;
        RECT -68.845 180.035 -68.515 180.365 ;
        RECT -68.845 178.675 -68.515 179.005 ;
        RECT -68.845 177.315 -68.515 177.645 ;
        RECT -68.845 175.955 -68.515 176.285 ;
        RECT -68.845 174.595 -68.515 174.925 ;
        RECT -68.845 173.235 -68.515 173.565 ;
        RECT -68.845 171.875 -68.515 172.205 ;
        RECT -68.845 170.515 -68.515 170.845 ;
        RECT -68.845 169.155 -68.515 169.485 ;
        RECT -68.845 167.795 -68.515 168.125 ;
        RECT -68.845 166.435 -68.515 166.765 ;
        RECT -68.845 165.075 -68.515 165.405 ;
        RECT -68.845 163.715 -68.515 164.045 ;
        RECT -68.845 162.355 -68.515 162.685 ;
        RECT -68.845 160.995 -68.515 161.325 ;
        RECT -68.845 159.635 -68.515 159.965 ;
        RECT -68.845 158.275 -68.515 158.605 ;
        RECT -68.845 156.915 -68.515 157.245 ;
        RECT -68.845 155.555 -68.515 155.885 ;
        RECT -68.845 154.195 -68.515 154.525 ;
        RECT -68.845 152.835 -68.515 153.165 ;
        RECT -68.845 151.475 -68.515 151.805 ;
        RECT -68.845 150.115 -68.515 150.445 ;
        RECT -68.845 148.755 -68.515 149.085 ;
        RECT -68.845 147.395 -68.515 147.725 ;
        RECT -68.845 146.035 -68.515 146.365 ;
        RECT -68.845 144.675 -68.515 145.005 ;
        RECT -68.845 143.315 -68.515 143.645 ;
        RECT -68.845 141.955 -68.515 142.285 ;
        RECT -68.845 140.595 -68.515 140.925 ;
        RECT -68.845 139.235 -68.515 139.565 ;
        RECT -68.845 137.875 -68.515 138.205 ;
        RECT -68.845 136.515 -68.515 136.845 ;
        RECT -68.845 135.155 -68.515 135.485 ;
        RECT -68.845 133.795 -68.515 134.125 ;
        RECT -68.845 132.435 -68.515 132.765 ;
        RECT -68.845 131.075 -68.515 131.405 ;
        RECT -68.845 129.715 -68.515 130.045 ;
        RECT -68.845 128.355 -68.515 128.685 ;
        RECT -68.845 126.995 -68.515 127.325 ;
        RECT -68.845 125.635 -68.515 125.965 ;
        RECT -68.845 124.275 -68.515 124.605 ;
        RECT -68.845 122.915 -68.515 123.245 ;
        RECT -68.845 121.555 -68.515 121.885 ;
        RECT -68.845 120.195 -68.515 120.525 ;
        RECT -68.845 118.835 -68.515 119.165 ;
        RECT -68.845 117.475 -68.515 117.805 ;
        RECT -68.845 116.115 -68.515 116.445 ;
        RECT -68.845 114.755 -68.515 115.085 ;
        RECT -68.845 113.395 -68.515 113.725 ;
        RECT -68.845 112.035 -68.515 112.365 ;
        RECT -68.845 110.675 -68.515 111.005 ;
        RECT -68.845 109.315 -68.515 109.645 ;
        RECT -68.845 107.955 -68.515 108.285 ;
        RECT -68.845 106.595 -68.515 106.925 ;
        RECT -68.845 105.235 -68.515 105.565 ;
        RECT -68.845 103.875 -68.515 104.205 ;
        RECT -68.845 102.515 -68.515 102.845 ;
        RECT -68.845 101.155 -68.515 101.485 ;
        RECT -68.845 99.795 -68.515 100.125 ;
        RECT -68.845 98.435 -68.515 98.765 ;
        RECT -68.845 97.075 -68.515 97.405 ;
        RECT -68.845 95.715 -68.515 96.045 ;
        RECT -68.845 94.355 -68.515 94.685 ;
        RECT -68.845 92.995 -68.515 93.325 ;
        RECT -68.845 91.635 -68.515 91.965 ;
        RECT -68.845 90.275 -68.515 90.605 ;
        RECT -68.845 88.915 -68.515 89.245 ;
        RECT -68.845 87.555 -68.515 87.885 ;
        RECT -68.845 86.195 -68.515 86.525 ;
        RECT -68.845 84.835 -68.515 85.165 ;
        RECT -68.845 83.475 -68.515 83.805 ;
        RECT -68.845 82.115 -68.515 82.445 ;
        RECT -68.845 80.755 -68.515 81.085 ;
        RECT -68.845 79.395 -68.515 79.725 ;
        RECT -68.845 78.035 -68.515 78.365 ;
        RECT -68.845 76.675 -68.515 77.005 ;
        RECT -68.845 75.315 -68.515 75.645 ;
        RECT -68.845 73.955 -68.515 74.285 ;
        RECT -68.845 72.595 -68.515 72.925 ;
        RECT -68.845 71.235 -68.515 71.565 ;
        RECT -68.845 69.875 -68.515 70.205 ;
        RECT -68.845 68.515 -68.515 68.845 ;
        RECT -68.845 67.155 -68.515 67.485 ;
        RECT -68.845 65.795 -68.515 66.125 ;
        RECT -68.845 64.435 -68.515 64.765 ;
        RECT -68.845 63.075 -68.515 63.405 ;
        RECT -68.845 61.715 -68.515 62.045 ;
        RECT -68.845 60.355 -68.515 60.685 ;
        RECT -68.845 58.995 -68.515 59.325 ;
        RECT -68.845 57.635 -68.515 57.965 ;
        RECT -68.845 56.275 -68.515 56.605 ;
        RECT -68.845 54.915 -68.515 55.245 ;
        RECT -68.845 53.555 -68.515 53.885 ;
        RECT -68.845 52.195 -68.515 52.525 ;
        RECT -68.845 50.835 -68.515 51.165 ;
        RECT -68.845 49.475 -68.515 49.805 ;
        RECT -68.845 48.115 -68.515 48.445 ;
        RECT -68.845 46.755 -68.515 47.085 ;
        RECT -68.845 45.395 -68.515 45.725 ;
        RECT -68.845 44.035 -68.515 44.365 ;
        RECT -68.845 42.675 -68.515 43.005 ;
        RECT -68.845 41.315 -68.515 41.645 ;
        RECT -68.845 39.955 -68.515 40.285 ;
        RECT -68.845 38.595 -68.515 38.925 ;
        RECT -68.845 37.235 -68.515 37.565 ;
        RECT -68.845 35.875 -68.515 36.205 ;
        RECT -68.845 34.515 -68.515 34.845 ;
        RECT -68.845 33.155 -68.515 33.485 ;
        RECT -68.845 31.795 -68.515 32.125 ;
        RECT -68.845 30.435 -68.515 30.765 ;
        RECT -68.845 29.075 -68.515 29.405 ;
        RECT -68.845 27.715 -68.515 28.045 ;
        RECT -68.845 26.355 -68.515 26.685 ;
        RECT -68.845 24.995 -68.515 25.325 ;
        RECT -68.845 23.635 -68.515 23.965 ;
        RECT -68.845 22.275 -68.515 22.605 ;
        RECT -68.845 20.915 -68.515 21.245 ;
        RECT -68.845 19.555 -68.515 19.885 ;
        RECT -68.845 18.195 -68.515 18.525 ;
        RECT -68.845 16.835 -68.515 17.165 ;
        RECT -68.845 15.475 -68.515 15.805 ;
        RECT -68.845 14.115 -68.515 14.445 ;
        RECT -68.845 12.755 -68.515 13.085 ;
        RECT -68.845 11.395 -68.515 11.725 ;
        RECT -68.845 10.035 -68.515 10.365 ;
        RECT -68.845 8.675 -68.515 9.005 ;
        RECT -68.845 7.315 -68.515 7.645 ;
        RECT -68.845 5.955 -68.515 6.285 ;
        RECT -68.845 4.595 -68.515 4.925 ;
        RECT -68.845 3.235 -68.515 3.565 ;
        RECT -68.845 1.875 -68.515 2.205 ;
        RECT -68.845 0.515 -68.515 0.845 ;
        RECT -68.845 -0.845 -68.515 -0.515 ;
        RECT -68.845 -2.205 -68.515 -1.875 ;
        RECT -68.845 -3.565 -68.515 -3.235 ;
        RECT -68.845 -4.925 -68.515 -4.595 ;
        RECT -68.845 -6.285 -68.515 -5.955 ;
        RECT -68.845 -7.645 -68.515 -7.315 ;
        RECT -68.845 -9.005 -68.515 -8.675 ;
        RECT -68.845 -10.365 -68.515 -10.035 ;
        RECT -68.845 -11.725 -68.515 -11.395 ;
        RECT -68.845 -13.085 -68.515 -12.755 ;
        RECT -68.845 -14.445 -68.515 -14.115 ;
        RECT -68.845 -15.805 -68.515 -15.475 ;
        RECT -68.845 -17.165 -68.515 -16.835 ;
        RECT -68.845 -18.525 -68.515 -18.195 ;
        RECT -68.845 -19.885 -68.515 -19.555 ;
        RECT -68.845 -21.245 -68.515 -20.915 ;
        RECT -68.845 -22.605 -68.515 -22.275 ;
        RECT -68.845 -23.965 -68.515 -23.635 ;
        RECT -68.845 -25.325 -68.515 -24.995 ;
        RECT -68.845 -26.685 -68.515 -26.355 ;
        RECT -68.845 -28.045 -68.515 -27.715 ;
        RECT -68.845 -29.405 -68.515 -29.075 ;
        RECT -68.845 -30.765 -68.515 -30.435 ;
        RECT -68.845 -32.125 -68.515 -31.795 ;
        RECT -68.845 -33.485 -68.515 -33.155 ;
        RECT -68.845 -34.845 -68.515 -34.515 ;
        RECT -68.845 -36.205 -68.515 -35.875 ;
        RECT -68.845 -37.565 -68.515 -37.235 ;
        RECT -68.845 -38.925 -68.515 -38.595 ;
        RECT -68.845 -40.285 -68.515 -39.955 ;
        RECT -68.845 -41.645 -68.515 -41.315 ;
        RECT -68.845 -43.005 -68.515 -42.675 ;
        RECT -68.845 -44.365 -68.515 -44.035 ;
        RECT -68.845 -45.725 -68.515 -45.395 ;
        RECT -68.845 -47.085 -68.515 -46.755 ;
        RECT -68.845 -48.445 -68.515 -48.115 ;
        RECT -68.845 -49.805 -68.515 -49.475 ;
        RECT -68.845 -51.165 -68.515 -50.835 ;
        RECT -68.845 -52.525 -68.515 -52.195 ;
        RECT -68.845 -53.885 -68.515 -53.555 ;
        RECT -68.845 -55.245 -68.515 -54.915 ;
        RECT -68.845 -56.605 -68.515 -56.275 ;
        RECT -68.845 -57.965 -68.515 -57.635 ;
        RECT -68.845 -59.325 -68.515 -58.995 ;
        RECT -68.845 -60.685 -68.515 -60.355 ;
        RECT -68.845 -62.045 -68.515 -61.715 ;
        RECT -68.845 -63.405 -68.515 -63.075 ;
        RECT -68.845 -64.765 -68.515 -64.435 ;
        RECT -68.845 -66.125 -68.515 -65.795 ;
        RECT -68.845 -67.485 -68.515 -67.155 ;
        RECT -68.845 -68.845 -68.515 -68.515 ;
        RECT -68.845 -70.205 -68.515 -69.875 ;
        RECT -68.845 -71.565 -68.515 -71.235 ;
        RECT -68.845 -72.925 -68.515 -72.595 ;
        RECT -68.845 -74.285 -68.515 -73.955 ;
        RECT -68.845 -75.645 -68.515 -75.315 ;
        RECT -68.845 -77.005 -68.515 -76.675 ;
        RECT -68.845 -78.365 -68.515 -78.035 ;
        RECT -68.845 -79.725 -68.515 -79.395 ;
        RECT -68.845 -81.085 -68.515 -80.755 ;
        RECT -68.845 -82.445 -68.515 -82.115 ;
        RECT -68.845 -83.805 -68.515 -83.475 ;
        RECT -68.845 -85.165 -68.515 -84.835 ;
        RECT -68.845 -86.525 -68.515 -86.195 ;
        RECT -68.845 -87.885 -68.515 -87.555 ;
        RECT -68.845 -89.245 -68.515 -88.915 ;
        RECT -68.845 -90.605 -68.515 -90.275 ;
        RECT -68.845 -91.965 -68.515 -91.635 ;
        RECT -68.845 -93.325 -68.515 -92.995 ;
        RECT -68.845 -94.685 -68.515 -94.355 ;
        RECT -68.845 -96.045 -68.515 -95.715 ;
        RECT -68.845 -97.405 -68.515 -97.075 ;
        RECT -68.845 -98.765 -68.515 -98.435 ;
        RECT -68.845 -100.125 -68.515 -99.795 ;
        RECT -68.845 -101.485 -68.515 -101.155 ;
        RECT -68.845 -102.845 -68.515 -102.515 ;
        RECT -68.845 -104.205 -68.515 -103.875 ;
        RECT -68.845 -105.565 -68.515 -105.235 ;
        RECT -68.845 -106.925 -68.515 -106.595 ;
        RECT -68.845 -108.285 -68.515 -107.955 ;
        RECT -68.845 -109.645 -68.515 -109.315 ;
        RECT -68.845 -111.005 -68.515 -110.675 ;
        RECT -68.845 -112.365 -68.515 -112.035 ;
        RECT -68.845 -113.725 -68.515 -113.395 ;
        RECT -68.845 -115.085 -68.515 -114.755 ;
        RECT -68.845 -116.445 -68.515 -116.115 ;
        RECT -68.845 -117.805 -68.515 -117.475 ;
        RECT -68.845 -119.165 -68.515 -118.835 ;
        RECT -68.845 -120.525 -68.515 -120.195 ;
        RECT -68.845 -121.885 -68.515 -121.555 ;
        RECT -68.845 -123.245 -68.515 -122.915 ;
        RECT -68.845 -124.605 -68.515 -124.275 ;
        RECT -68.845 -125.965 -68.515 -125.635 ;
        RECT -68.845 -127.325 -68.515 -126.995 ;
        RECT -68.845 -128.685 -68.515 -128.355 ;
        RECT -68.845 -130.045 -68.515 -129.715 ;
        RECT -68.845 -132.765 -68.515 -132.435 ;
        RECT -68.845 -134.125 -68.515 -133.795 ;
        RECT -68.845 -135.485 -68.515 -135.155 ;
        RECT -68.845 -136.845 -68.515 -136.515 ;
        RECT -68.845 -138.205 -68.515 -137.875 ;
        RECT -68.845 -139.39 -68.515 -139.06 ;
        RECT -68.845 -140.925 -68.515 -140.595 ;
        RECT -68.845 -142.285 -68.515 -141.955 ;
        RECT -68.845 -145.005 -68.515 -144.675 ;
        RECT -68.845 -146.365 -68.515 -146.035 ;
        RECT -68.845 -148.03 -68.515 -147.7 ;
        RECT -68.845 -149.085 -68.515 -148.755 ;
        RECT -68.845 -153.165 -68.515 -152.835 ;
        RECT -68.845 -154.525 -68.515 -154.195 ;
        RECT -68.845 -155.885 -68.515 -155.555 ;
        RECT -68.845 -157.245 -68.515 -156.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -75.645 244.04 -75.315 245.17 ;
        RECT -75.645 242.595 -75.315 242.925 ;
        RECT -75.645 241.235 -75.315 241.565 ;
        RECT -75.645 239.875 -75.315 240.205 ;
        RECT -75.645 238.515 -75.315 238.845 ;
        RECT -75.645 237.155 -75.315 237.485 ;
        RECT -75.645 235.795 -75.315 236.125 ;
        RECT -75.645 234.435 -75.315 234.765 ;
        RECT -75.645 233.075 -75.315 233.405 ;
        RECT -75.645 231.715 -75.315 232.045 ;
        RECT -75.645 230.355 -75.315 230.685 ;
        RECT -75.645 228.995 -75.315 229.325 ;
        RECT -75.645 227.635 -75.315 227.965 ;
        RECT -75.645 226.275 -75.315 226.605 ;
        RECT -75.645 224.915 -75.315 225.245 ;
        RECT -75.645 223.555 -75.315 223.885 ;
        RECT -75.645 222.195 -75.315 222.525 ;
        RECT -75.645 220.835 -75.315 221.165 ;
        RECT -75.645 219.475 -75.315 219.805 ;
        RECT -75.645 218.115 -75.315 218.445 ;
        RECT -75.645 216.755 -75.315 217.085 ;
        RECT -75.645 215.395 -75.315 215.725 ;
        RECT -75.645 214.035 -75.315 214.365 ;
        RECT -75.645 212.675 -75.315 213.005 ;
        RECT -75.645 211.315 -75.315 211.645 ;
        RECT -75.645 209.955 -75.315 210.285 ;
        RECT -75.645 208.595 -75.315 208.925 ;
        RECT -75.645 207.235 -75.315 207.565 ;
        RECT -75.645 205.875 -75.315 206.205 ;
        RECT -75.645 204.515 -75.315 204.845 ;
        RECT -75.645 203.155 -75.315 203.485 ;
        RECT -75.645 201.795 -75.315 202.125 ;
        RECT -75.645 200.435 -75.315 200.765 ;
        RECT -75.645 199.075 -75.315 199.405 ;
        RECT -75.645 197.715 -75.315 198.045 ;
        RECT -75.645 196.355 -75.315 196.685 ;
        RECT -75.645 194.995 -75.315 195.325 ;
        RECT -75.645 193.635 -75.315 193.965 ;
        RECT -75.645 192.275 -75.315 192.605 ;
        RECT -75.645 190.915 -75.315 191.245 ;
        RECT -75.645 189.555 -75.315 189.885 ;
        RECT -75.645 188.195 -75.315 188.525 ;
        RECT -75.645 186.835 -75.315 187.165 ;
        RECT -75.645 185.475 -75.315 185.805 ;
        RECT -75.645 184.115 -75.315 184.445 ;
        RECT -75.645 182.755 -75.315 183.085 ;
        RECT -75.645 181.395 -75.315 181.725 ;
        RECT -75.645 180.035 -75.315 180.365 ;
        RECT -75.645 178.675 -75.315 179.005 ;
        RECT -75.645 177.315 -75.315 177.645 ;
        RECT -75.645 175.955 -75.315 176.285 ;
        RECT -75.645 174.595 -75.315 174.925 ;
        RECT -75.645 173.235 -75.315 173.565 ;
        RECT -75.645 171.875 -75.315 172.205 ;
        RECT -75.645 170.515 -75.315 170.845 ;
        RECT -75.645 169.155 -75.315 169.485 ;
        RECT -75.645 167.795 -75.315 168.125 ;
        RECT -75.645 166.435 -75.315 166.765 ;
        RECT -75.645 165.075 -75.315 165.405 ;
        RECT -75.645 163.715 -75.315 164.045 ;
        RECT -75.645 162.355 -75.315 162.685 ;
        RECT -75.645 160.995 -75.315 161.325 ;
        RECT -75.645 159.635 -75.315 159.965 ;
        RECT -75.645 158.275 -75.315 158.605 ;
        RECT -75.645 156.915 -75.315 157.245 ;
        RECT -75.645 155.555 -75.315 155.885 ;
        RECT -75.645 154.195 -75.315 154.525 ;
        RECT -75.645 152.835 -75.315 153.165 ;
        RECT -75.645 151.475 -75.315 151.805 ;
        RECT -75.645 150.115 -75.315 150.445 ;
        RECT -75.645 148.755 -75.315 149.085 ;
        RECT -75.645 147.395 -75.315 147.725 ;
        RECT -75.645 146.035 -75.315 146.365 ;
        RECT -75.645 144.675 -75.315 145.005 ;
        RECT -75.645 143.315 -75.315 143.645 ;
        RECT -75.645 141.955 -75.315 142.285 ;
        RECT -75.645 140.595 -75.315 140.925 ;
        RECT -75.645 139.235 -75.315 139.565 ;
        RECT -75.645 137.875 -75.315 138.205 ;
        RECT -75.645 136.515 -75.315 136.845 ;
        RECT -75.645 135.155 -75.315 135.485 ;
        RECT -75.645 133.795 -75.315 134.125 ;
        RECT -75.645 132.435 -75.315 132.765 ;
        RECT -75.645 131.075 -75.315 131.405 ;
        RECT -75.645 129.715 -75.315 130.045 ;
        RECT -75.645 128.355 -75.315 128.685 ;
        RECT -75.645 126.995 -75.315 127.325 ;
        RECT -75.645 125.635 -75.315 125.965 ;
        RECT -75.645 124.275 -75.315 124.605 ;
        RECT -75.645 122.915 -75.315 123.245 ;
        RECT -75.645 121.555 -75.315 121.885 ;
        RECT -75.645 120.195 -75.315 120.525 ;
        RECT -75.645 118.835 -75.315 119.165 ;
        RECT -75.645 117.475 -75.315 117.805 ;
        RECT -75.645 116.115 -75.315 116.445 ;
        RECT -75.645 114.755 -75.315 115.085 ;
        RECT -75.645 113.395 -75.315 113.725 ;
        RECT -75.645 112.035 -75.315 112.365 ;
        RECT -75.645 110.675 -75.315 111.005 ;
        RECT -75.645 109.315 -75.315 109.645 ;
        RECT -75.645 107.955 -75.315 108.285 ;
        RECT -75.645 106.595 -75.315 106.925 ;
        RECT -75.645 105.235 -75.315 105.565 ;
        RECT -75.645 103.875 -75.315 104.205 ;
        RECT -75.645 102.515 -75.315 102.845 ;
        RECT -75.645 101.155 -75.315 101.485 ;
        RECT -75.645 99.795 -75.315 100.125 ;
        RECT -75.645 98.435 -75.315 98.765 ;
        RECT -75.645 97.075 -75.315 97.405 ;
        RECT -75.645 95.715 -75.315 96.045 ;
        RECT -75.645 94.355 -75.315 94.685 ;
        RECT -75.645 92.995 -75.315 93.325 ;
        RECT -75.645 91.635 -75.315 91.965 ;
        RECT -75.645 90.275 -75.315 90.605 ;
        RECT -75.645 88.915 -75.315 89.245 ;
        RECT -75.645 87.555 -75.315 87.885 ;
        RECT -75.645 86.195 -75.315 86.525 ;
        RECT -75.645 84.835 -75.315 85.165 ;
        RECT -75.645 83.475 -75.315 83.805 ;
        RECT -75.645 82.115 -75.315 82.445 ;
        RECT -75.645 80.755 -75.315 81.085 ;
        RECT -75.645 79.395 -75.315 79.725 ;
        RECT -75.645 78.035 -75.315 78.365 ;
        RECT -75.645 76.675 -75.315 77.005 ;
        RECT -75.645 75.315 -75.315 75.645 ;
        RECT -75.645 73.955 -75.315 74.285 ;
        RECT -75.645 72.595 -75.315 72.925 ;
        RECT -75.645 71.235 -75.315 71.565 ;
        RECT -75.645 69.875 -75.315 70.205 ;
        RECT -75.645 68.515 -75.315 68.845 ;
        RECT -75.645 67.155 -75.315 67.485 ;
        RECT -75.645 65.795 -75.315 66.125 ;
        RECT -75.645 64.435 -75.315 64.765 ;
        RECT -75.645 63.075 -75.315 63.405 ;
        RECT -75.645 61.715 -75.315 62.045 ;
        RECT -75.645 60.355 -75.315 60.685 ;
        RECT -75.645 58.995 -75.315 59.325 ;
        RECT -75.645 57.635 -75.315 57.965 ;
        RECT -75.645 56.275 -75.315 56.605 ;
        RECT -75.645 54.915 -75.315 55.245 ;
        RECT -75.645 53.555 -75.315 53.885 ;
        RECT -75.645 52.195 -75.315 52.525 ;
        RECT -75.645 50.835 -75.315 51.165 ;
        RECT -75.645 49.475 -75.315 49.805 ;
        RECT -75.645 48.115 -75.315 48.445 ;
        RECT -75.645 46.755 -75.315 47.085 ;
        RECT -75.645 45.395 -75.315 45.725 ;
        RECT -75.645 44.035 -75.315 44.365 ;
        RECT -75.645 42.675 -75.315 43.005 ;
        RECT -75.645 41.315 -75.315 41.645 ;
        RECT -75.645 39.955 -75.315 40.285 ;
        RECT -75.645 38.595 -75.315 38.925 ;
        RECT -75.645 37.235 -75.315 37.565 ;
        RECT -75.645 35.875 -75.315 36.205 ;
        RECT -75.645 34.515 -75.315 34.845 ;
        RECT -75.645 33.155 -75.315 33.485 ;
        RECT -75.645 31.795 -75.315 32.125 ;
        RECT -75.645 30.435 -75.315 30.765 ;
        RECT -75.645 29.075 -75.315 29.405 ;
        RECT -75.645 27.715 -75.315 28.045 ;
        RECT -75.645 26.355 -75.315 26.685 ;
        RECT -75.645 24.995 -75.315 25.325 ;
        RECT -75.645 23.635 -75.315 23.965 ;
        RECT -75.645 22.275 -75.315 22.605 ;
        RECT -75.645 20.915 -75.315 21.245 ;
        RECT -75.645 19.555 -75.315 19.885 ;
        RECT -75.645 18.195 -75.315 18.525 ;
        RECT -75.645 16.835 -75.315 17.165 ;
        RECT -75.645 15.475 -75.315 15.805 ;
        RECT -75.645 14.115 -75.315 14.445 ;
        RECT -75.645 12.755 -75.315 13.085 ;
        RECT -75.645 11.395 -75.315 11.725 ;
        RECT -75.645 10.035 -75.315 10.365 ;
        RECT -75.645 8.675 -75.315 9.005 ;
        RECT -75.645 7.315 -75.315 7.645 ;
        RECT -75.645 5.955 -75.315 6.285 ;
        RECT -75.645 4.595 -75.315 4.925 ;
        RECT -75.645 3.235 -75.315 3.565 ;
        RECT -75.645 1.875 -75.315 2.205 ;
        RECT -75.645 0.515 -75.315 0.845 ;
        RECT -75.645 -0.845 -75.315 -0.515 ;
        RECT -75.645 -2.205 -75.315 -1.875 ;
        RECT -75.645 -3.565 -75.315 -3.235 ;
        RECT -75.645 -4.925 -75.315 -4.595 ;
        RECT -75.645 -6.285 -75.315 -5.955 ;
        RECT -75.645 -7.645 -75.315 -7.315 ;
        RECT -75.645 -9.005 -75.315 -8.675 ;
        RECT -75.645 -10.365 -75.315 -10.035 ;
        RECT -75.645 -11.725 -75.315 -11.395 ;
        RECT -75.645 -13.085 -75.315 -12.755 ;
        RECT -75.645 -14.445 -75.315 -14.115 ;
        RECT -75.645 -15.805 -75.315 -15.475 ;
        RECT -75.645 -17.165 -75.315 -16.835 ;
        RECT -75.645 -18.525 -75.315 -18.195 ;
        RECT -75.645 -19.885 -75.315 -19.555 ;
        RECT -75.645 -21.245 -75.315 -20.915 ;
        RECT -75.645 -22.605 -75.315 -22.275 ;
        RECT -75.645 -23.965 -75.315 -23.635 ;
        RECT -75.645 -25.325 -75.315 -24.995 ;
        RECT -75.645 -26.685 -75.315 -26.355 ;
        RECT -75.645 -28.045 -75.315 -27.715 ;
        RECT -75.645 -29.405 -75.315 -29.075 ;
        RECT -75.645 -30.765 -75.315 -30.435 ;
        RECT -75.645 -32.125 -75.315 -31.795 ;
        RECT -75.645 -33.485 -75.315 -33.155 ;
        RECT -75.645 -34.845 -75.315 -34.515 ;
        RECT -75.645 -36.205 -75.315 -35.875 ;
        RECT -75.645 -37.565 -75.315 -37.235 ;
        RECT -75.645 -38.925 -75.315 -38.595 ;
        RECT -75.645 -40.285 -75.315 -39.955 ;
        RECT -75.645 -41.645 -75.315 -41.315 ;
        RECT -75.645 -43.005 -75.315 -42.675 ;
        RECT -75.645 -44.365 -75.315 -44.035 ;
        RECT -75.645 -45.725 -75.315 -45.395 ;
        RECT -75.645 -47.085 -75.315 -46.755 ;
        RECT -75.645 -48.445 -75.315 -48.115 ;
        RECT -75.645 -49.805 -75.315 -49.475 ;
        RECT -75.645 -51.165 -75.315 -50.835 ;
        RECT -75.645 -52.525 -75.315 -52.195 ;
        RECT -75.645 -53.885 -75.315 -53.555 ;
        RECT -75.645 -55.245 -75.315 -54.915 ;
        RECT -75.645 -56.605 -75.315 -56.275 ;
        RECT -75.645 -57.965 -75.315 -57.635 ;
        RECT -75.645 -59.325 -75.315 -58.995 ;
        RECT -75.645 -60.685 -75.315 -60.355 ;
        RECT -75.645 -62.045 -75.315 -61.715 ;
        RECT -75.645 -63.405 -75.315 -63.075 ;
        RECT -75.645 -64.765 -75.315 -64.435 ;
        RECT -75.645 -66.125 -75.315 -65.795 ;
        RECT -75.645 -67.485 -75.315 -67.155 ;
        RECT -75.645 -68.845 -75.315 -68.515 ;
        RECT -75.645 -70.205 -75.315 -69.875 ;
        RECT -75.645 -71.565 -75.315 -71.235 ;
        RECT -75.645 -72.925 -75.315 -72.595 ;
        RECT -75.645 -74.285 -75.315 -73.955 ;
        RECT -75.645 -75.645 -75.315 -75.315 ;
        RECT -75.645 -77.005 -75.315 -76.675 ;
        RECT -75.645 -78.365 -75.315 -78.035 ;
        RECT -75.645 -79.725 -75.315 -79.395 ;
        RECT -75.645 -81.085 -75.315 -80.755 ;
        RECT -75.645 -82.445 -75.315 -82.115 ;
        RECT -75.645 -83.805 -75.315 -83.475 ;
        RECT -75.645 -85.165 -75.315 -84.835 ;
        RECT -75.645 -86.525 -75.315 -86.195 ;
        RECT -75.645 -87.885 -75.315 -87.555 ;
        RECT -75.645 -89.245 -75.315 -88.915 ;
        RECT -75.645 -90.605 -75.315 -90.275 ;
        RECT -75.645 -91.965 -75.315 -91.635 ;
        RECT -75.645 -93.325 -75.315 -92.995 ;
        RECT -75.645 -94.685 -75.315 -94.355 ;
        RECT -75.645 -96.045 -75.315 -95.715 ;
        RECT -75.645 -97.405 -75.315 -97.075 ;
        RECT -75.645 -98.765 -75.315 -98.435 ;
        RECT -75.645 -100.125 -75.315 -99.795 ;
        RECT -75.645 -101.485 -75.315 -101.155 ;
        RECT -75.645 -102.845 -75.315 -102.515 ;
        RECT -75.645 -104.205 -75.315 -103.875 ;
        RECT -75.645 -105.565 -75.315 -105.235 ;
        RECT -75.645 -106.925 -75.315 -106.595 ;
        RECT -75.645 -108.285 -75.315 -107.955 ;
        RECT -75.645 -109.645 -75.315 -109.315 ;
        RECT -75.645 -111.005 -75.315 -110.675 ;
        RECT -75.645 -112.365 -75.315 -112.035 ;
        RECT -75.645 -113.725 -75.315 -113.395 ;
        RECT -75.645 -115.085 -75.315 -114.755 ;
        RECT -75.645 -116.445 -75.315 -116.115 ;
        RECT -75.645 -117.805 -75.315 -117.475 ;
        RECT -75.645 -119.165 -75.315 -118.835 ;
        RECT -75.645 -120.525 -75.315 -120.195 ;
        RECT -75.645 -121.885 -75.315 -121.555 ;
        RECT -75.645 -123.245 -75.315 -122.915 ;
        RECT -75.645 -124.605 -75.315 -124.275 ;
        RECT -75.645 -125.965 -75.315 -125.635 ;
        RECT -75.645 -127.325 -75.315 -126.995 ;
        RECT -75.645 -128.685 -75.315 -128.355 ;
        RECT -75.645 -130.045 -75.315 -129.715 ;
        RECT -75.645 -131.405 -75.315 -131.075 ;
        RECT -75.645 -132.765 -75.315 -132.435 ;
        RECT -75.645 -134.125 -75.315 -133.795 ;
        RECT -75.645 -135.485 -75.315 -135.155 ;
        RECT -75.645 -136.845 -75.315 -136.515 ;
        RECT -75.645 -138.205 -75.315 -137.875 ;
        RECT -75.645 -139.565 -75.315 -139.235 ;
        RECT -75.645 -140.925 -75.315 -140.595 ;
        RECT -75.645 -142.285 -75.315 -141.955 ;
        RECT -75.645 -143.645 -75.315 -143.315 ;
        RECT -75.645 -145.005 -75.315 -144.675 ;
        RECT -75.645 -146.365 -75.315 -146.035 ;
        RECT -75.645 -147.725 -75.315 -147.395 ;
        RECT -75.645 -149.085 -75.315 -148.755 ;
        RECT -75.645 -150.445 -75.315 -150.115 ;
        RECT -75.645 -151.805 -75.315 -151.475 ;
        RECT -75.645 -153.165 -75.315 -152.835 ;
        RECT -75.645 -154.525 -75.315 -154.195 ;
        RECT -75.645 -155.885 -75.315 -155.555 ;
        RECT -75.645 -157.245 -75.315 -156.915 ;
        RECT -75.645 -158.605 -75.315 -158.275 ;
        RECT -75.645 -159.965 -75.315 -159.635 ;
        RECT -75.645 -161.325 -75.315 -160.995 ;
        RECT -75.645 -162.685 -75.315 -162.355 ;
        RECT -75.645 -164.045 -75.315 -163.715 ;
        RECT -75.645 -165.405 -75.315 -165.075 ;
        RECT -75.645 -166.765 -75.315 -166.435 ;
        RECT -75.645 -168.125 -75.315 -167.795 ;
        RECT -75.645 -169.485 -75.315 -169.155 ;
        RECT -75.645 -170.845 -75.315 -170.515 ;
        RECT -75.645 -172.205 -75.315 -171.875 ;
        RECT -75.645 -173.565 -75.315 -173.235 ;
        RECT -75.645 -174.925 -75.315 -174.595 ;
        RECT -75.645 -176.285 -75.315 -175.955 ;
        RECT -75.645 -177.645 -75.315 -177.315 ;
        RECT -75.645 -179.005 -75.315 -178.675 ;
        RECT -75.645 -180.365 -75.315 -180.035 ;
        RECT -75.645 -181.725 -75.315 -181.395 ;
        RECT -75.645 -183.085 -75.315 -182.755 ;
        RECT -75.645 -184.445 -75.315 -184.115 ;
        RECT -75.645 -185.805 -75.315 -185.475 ;
        RECT -75.645 -187.165 -75.315 -186.835 ;
        RECT -75.645 -188.525 -75.315 -188.195 ;
        RECT -75.645 -189.885 -75.315 -189.555 ;
        RECT -75.645 -191.245 -75.315 -190.915 ;
        RECT -75.645 -192.605 -75.315 -192.275 ;
        RECT -75.645 -193.965 -75.315 -193.635 ;
        RECT -75.645 -195.325 -75.315 -194.995 ;
        RECT -75.645 -196.685 -75.315 -196.355 ;
        RECT -75.645 -198.045 -75.315 -197.715 ;
        RECT -75.645 -199.405 -75.315 -199.075 ;
        RECT -75.645 -200.765 -75.315 -200.435 ;
        RECT -75.645 -202.125 -75.315 -201.795 ;
        RECT -75.645 -203.485 -75.315 -203.155 ;
        RECT -75.645 -204.845 -75.315 -204.515 ;
        RECT -75.645 -206.205 -75.315 -205.875 ;
        RECT -75.645 -207.565 -75.315 -207.235 ;
        RECT -75.645 -208.925 -75.315 -208.595 ;
        RECT -75.645 -210.285 -75.315 -209.955 ;
        RECT -75.645 -211.645 -75.315 -211.315 ;
        RECT -75.645 -213.005 -75.315 -212.675 ;
        RECT -75.645 -214.365 -75.315 -214.035 ;
        RECT -75.645 -215.725 -75.315 -215.395 ;
        RECT -75.645 -217.085 -75.315 -216.755 ;
        RECT -75.645 -218.445 -75.315 -218.115 ;
        RECT -75.645 -219.805 -75.315 -219.475 ;
        RECT -75.645 -221.165 -75.315 -220.835 ;
        RECT -75.645 -222.525 -75.315 -222.195 ;
        RECT -75.645 -223.885 -75.315 -223.555 ;
        RECT -75.645 -225.245 -75.315 -224.915 ;
        RECT -75.645 -227.965 -75.315 -227.635 ;
        RECT -75.645 -230.685 -75.315 -230.355 ;
        RECT -75.645 -232.045 -75.315 -231.715 ;
        RECT -75.645 -233.225 -75.315 -232.895 ;
        RECT -75.645 -234.765 -75.315 -234.435 ;
        RECT -75.645 -236.125 -75.315 -235.795 ;
        RECT -75.645 -237.485 -75.315 -237.155 ;
        RECT -75.645 -238.845 -75.315 -238.515 ;
        RECT -75.645 -241.09 -75.315 -239.96 ;
        RECT -75.64 -241.205 -75.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.285 244.04 -73.955 245.17 ;
        RECT -74.285 242.595 -73.955 242.925 ;
        RECT -74.285 241.235 -73.955 241.565 ;
        RECT -74.285 239.875 -73.955 240.205 ;
        RECT -74.285 238.515 -73.955 238.845 ;
        RECT -74.285 237.155 -73.955 237.485 ;
        RECT -74.285 235.795 -73.955 236.125 ;
        RECT -74.285 234.435 -73.955 234.765 ;
        RECT -74.285 233.075 -73.955 233.405 ;
        RECT -74.285 231.715 -73.955 232.045 ;
        RECT -74.285 230.355 -73.955 230.685 ;
        RECT -74.285 228.995 -73.955 229.325 ;
        RECT -74.285 227.635 -73.955 227.965 ;
        RECT -74.285 226.275 -73.955 226.605 ;
        RECT -74.285 224.915 -73.955 225.245 ;
        RECT -74.285 223.555 -73.955 223.885 ;
        RECT -74.285 222.195 -73.955 222.525 ;
        RECT -74.285 220.835 -73.955 221.165 ;
        RECT -74.285 219.475 -73.955 219.805 ;
        RECT -74.285 218.115 -73.955 218.445 ;
        RECT -74.285 216.755 -73.955 217.085 ;
        RECT -74.285 215.395 -73.955 215.725 ;
        RECT -74.285 214.035 -73.955 214.365 ;
        RECT -74.285 212.675 -73.955 213.005 ;
        RECT -74.285 211.315 -73.955 211.645 ;
        RECT -74.285 209.955 -73.955 210.285 ;
        RECT -74.285 208.595 -73.955 208.925 ;
        RECT -74.285 207.235 -73.955 207.565 ;
        RECT -74.285 205.875 -73.955 206.205 ;
        RECT -74.285 204.515 -73.955 204.845 ;
        RECT -74.285 203.155 -73.955 203.485 ;
        RECT -74.285 201.795 -73.955 202.125 ;
        RECT -74.285 200.435 -73.955 200.765 ;
        RECT -74.285 199.075 -73.955 199.405 ;
        RECT -74.285 197.715 -73.955 198.045 ;
        RECT -74.285 196.355 -73.955 196.685 ;
        RECT -74.285 194.995 -73.955 195.325 ;
        RECT -74.285 193.635 -73.955 193.965 ;
        RECT -74.285 192.275 -73.955 192.605 ;
        RECT -74.285 190.915 -73.955 191.245 ;
        RECT -74.285 189.555 -73.955 189.885 ;
        RECT -74.285 188.195 -73.955 188.525 ;
        RECT -74.285 186.835 -73.955 187.165 ;
        RECT -74.285 185.475 -73.955 185.805 ;
        RECT -74.285 184.115 -73.955 184.445 ;
        RECT -74.285 182.755 -73.955 183.085 ;
        RECT -74.285 181.395 -73.955 181.725 ;
        RECT -74.285 180.035 -73.955 180.365 ;
        RECT -74.285 178.675 -73.955 179.005 ;
        RECT -74.285 177.315 -73.955 177.645 ;
        RECT -74.285 175.955 -73.955 176.285 ;
        RECT -74.285 174.595 -73.955 174.925 ;
        RECT -74.285 173.235 -73.955 173.565 ;
        RECT -74.285 171.875 -73.955 172.205 ;
        RECT -74.285 170.515 -73.955 170.845 ;
        RECT -74.285 169.155 -73.955 169.485 ;
        RECT -74.285 167.795 -73.955 168.125 ;
        RECT -74.285 166.435 -73.955 166.765 ;
        RECT -74.285 165.075 -73.955 165.405 ;
        RECT -74.285 163.715 -73.955 164.045 ;
        RECT -74.285 162.355 -73.955 162.685 ;
        RECT -74.285 160.995 -73.955 161.325 ;
        RECT -74.285 159.635 -73.955 159.965 ;
        RECT -74.285 158.275 -73.955 158.605 ;
        RECT -74.285 156.915 -73.955 157.245 ;
        RECT -74.285 155.555 -73.955 155.885 ;
        RECT -74.285 154.195 -73.955 154.525 ;
        RECT -74.285 152.835 -73.955 153.165 ;
        RECT -74.285 151.475 -73.955 151.805 ;
        RECT -74.285 150.115 -73.955 150.445 ;
        RECT -74.285 148.755 -73.955 149.085 ;
        RECT -74.285 147.395 -73.955 147.725 ;
        RECT -74.285 146.035 -73.955 146.365 ;
        RECT -74.285 144.675 -73.955 145.005 ;
        RECT -74.285 143.315 -73.955 143.645 ;
        RECT -74.285 141.955 -73.955 142.285 ;
        RECT -74.285 140.595 -73.955 140.925 ;
        RECT -74.285 139.235 -73.955 139.565 ;
        RECT -74.285 137.875 -73.955 138.205 ;
        RECT -74.285 136.515 -73.955 136.845 ;
        RECT -74.285 135.155 -73.955 135.485 ;
        RECT -74.285 133.795 -73.955 134.125 ;
        RECT -74.285 132.435 -73.955 132.765 ;
        RECT -74.285 131.075 -73.955 131.405 ;
        RECT -74.285 129.715 -73.955 130.045 ;
        RECT -74.285 128.355 -73.955 128.685 ;
        RECT -74.285 126.995 -73.955 127.325 ;
        RECT -74.285 125.635 -73.955 125.965 ;
        RECT -74.285 124.275 -73.955 124.605 ;
        RECT -74.285 122.915 -73.955 123.245 ;
        RECT -74.285 121.555 -73.955 121.885 ;
        RECT -74.285 120.195 -73.955 120.525 ;
        RECT -74.285 118.835 -73.955 119.165 ;
        RECT -74.285 117.475 -73.955 117.805 ;
        RECT -74.285 116.115 -73.955 116.445 ;
        RECT -74.285 114.755 -73.955 115.085 ;
        RECT -74.285 113.395 -73.955 113.725 ;
        RECT -74.285 112.035 -73.955 112.365 ;
        RECT -74.285 110.675 -73.955 111.005 ;
        RECT -74.285 109.315 -73.955 109.645 ;
        RECT -74.285 107.955 -73.955 108.285 ;
        RECT -74.285 106.595 -73.955 106.925 ;
        RECT -74.285 105.235 -73.955 105.565 ;
        RECT -74.285 103.875 -73.955 104.205 ;
        RECT -74.285 102.515 -73.955 102.845 ;
        RECT -74.285 101.155 -73.955 101.485 ;
        RECT -74.285 99.795 -73.955 100.125 ;
        RECT -74.285 98.435 -73.955 98.765 ;
        RECT -74.285 97.075 -73.955 97.405 ;
        RECT -74.285 95.715 -73.955 96.045 ;
        RECT -74.285 94.355 -73.955 94.685 ;
        RECT -74.285 92.995 -73.955 93.325 ;
        RECT -74.285 91.635 -73.955 91.965 ;
        RECT -74.285 90.275 -73.955 90.605 ;
        RECT -74.285 88.915 -73.955 89.245 ;
        RECT -74.285 87.555 -73.955 87.885 ;
        RECT -74.285 86.195 -73.955 86.525 ;
        RECT -74.285 84.835 -73.955 85.165 ;
        RECT -74.285 83.475 -73.955 83.805 ;
        RECT -74.285 82.115 -73.955 82.445 ;
        RECT -74.285 80.755 -73.955 81.085 ;
        RECT -74.285 79.395 -73.955 79.725 ;
        RECT -74.285 78.035 -73.955 78.365 ;
        RECT -74.285 76.675 -73.955 77.005 ;
        RECT -74.285 75.315 -73.955 75.645 ;
        RECT -74.285 73.955 -73.955 74.285 ;
        RECT -74.285 72.595 -73.955 72.925 ;
        RECT -74.285 71.235 -73.955 71.565 ;
        RECT -74.285 69.875 -73.955 70.205 ;
        RECT -74.285 68.515 -73.955 68.845 ;
        RECT -74.285 67.155 -73.955 67.485 ;
        RECT -74.285 65.795 -73.955 66.125 ;
        RECT -74.285 64.435 -73.955 64.765 ;
        RECT -74.285 63.075 -73.955 63.405 ;
        RECT -74.285 61.715 -73.955 62.045 ;
        RECT -74.285 60.355 -73.955 60.685 ;
        RECT -74.285 58.995 -73.955 59.325 ;
        RECT -74.285 57.635 -73.955 57.965 ;
        RECT -74.285 56.275 -73.955 56.605 ;
        RECT -74.285 54.915 -73.955 55.245 ;
        RECT -74.285 53.555 -73.955 53.885 ;
        RECT -74.285 52.195 -73.955 52.525 ;
        RECT -74.285 50.835 -73.955 51.165 ;
        RECT -74.285 49.475 -73.955 49.805 ;
        RECT -74.285 48.115 -73.955 48.445 ;
        RECT -74.285 46.755 -73.955 47.085 ;
        RECT -74.285 45.395 -73.955 45.725 ;
        RECT -74.285 44.035 -73.955 44.365 ;
        RECT -74.285 42.675 -73.955 43.005 ;
        RECT -74.285 41.315 -73.955 41.645 ;
        RECT -74.285 39.955 -73.955 40.285 ;
        RECT -74.285 38.595 -73.955 38.925 ;
        RECT -74.285 37.235 -73.955 37.565 ;
        RECT -74.285 35.875 -73.955 36.205 ;
        RECT -74.285 34.515 -73.955 34.845 ;
        RECT -74.285 33.155 -73.955 33.485 ;
        RECT -74.285 31.795 -73.955 32.125 ;
        RECT -74.285 30.435 -73.955 30.765 ;
        RECT -74.285 29.075 -73.955 29.405 ;
        RECT -74.285 27.715 -73.955 28.045 ;
        RECT -74.285 26.355 -73.955 26.685 ;
        RECT -74.285 24.995 -73.955 25.325 ;
        RECT -74.285 23.635 -73.955 23.965 ;
        RECT -74.285 22.275 -73.955 22.605 ;
        RECT -74.285 20.915 -73.955 21.245 ;
        RECT -74.285 19.555 -73.955 19.885 ;
        RECT -74.285 18.195 -73.955 18.525 ;
        RECT -74.285 16.835 -73.955 17.165 ;
        RECT -74.285 15.475 -73.955 15.805 ;
        RECT -74.285 14.115 -73.955 14.445 ;
        RECT -74.285 12.755 -73.955 13.085 ;
        RECT -74.285 11.395 -73.955 11.725 ;
        RECT -74.285 10.035 -73.955 10.365 ;
        RECT -74.285 8.675 -73.955 9.005 ;
        RECT -74.285 7.315 -73.955 7.645 ;
        RECT -74.285 5.955 -73.955 6.285 ;
        RECT -74.285 4.595 -73.955 4.925 ;
        RECT -74.285 3.235 -73.955 3.565 ;
        RECT -74.285 1.875 -73.955 2.205 ;
        RECT -74.285 0.515 -73.955 0.845 ;
        RECT -74.285 -0.845 -73.955 -0.515 ;
        RECT -74.285 -2.205 -73.955 -1.875 ;
        RECT -74.285 -3.565 -73.955 -3.235 ;
        RECT -74.285 -4.925 -73.955 -4.595 ;
        RECT -74.285 -6.285 -73.955 -5.955 ;
        RECT -74.285 -7.645 -73.955 -7.315 ;
        RECT -74.285 -9.005 -73.955 -8.675 ;
        RECT -74.285 -10.365 -73.955 -10.035 ;
        RECT -74.285 -11.725 -73.955 -11.395 ;
        RECT -74.285 -13.085 -73.955 -12.755 ;
        RECT -74.285 -14.445 -73.955 -14.115 ;
        RECT -74.285 -15.805 -73.955 -15.475 ;
        RECT -74.285 -17.165 -73.955 -16.835 ;
        RECT -74.285 -18.525 -73.955 -18.195 ;
        RECT -74.285 -19.885 -73.955 -19.555 ;
        RECT -74.285 -21.245 -73.955 -20.915 ;
        RECT -74.285 -22.605 -73.955 -22.275 ;
        RECT -74.285 -23.965 -73.955 -23.635 ;
        RECT -74.285 -25.325 -73.955 -24.995 ;
        RECT -74.285 -26.685 -73.955 -26.355 ;
        RECT -74.285 -28.045 -73.955 -27.715 ;
        RECT -74.285 -29.405 -73.955 -29.075 ;
        RECT -74.285 -30.765 -73.955 -30.435 ;
        RECT -74.285 -32.125 -73.955 -31.795 ;
        RECT -74.285 -33.485 -73.955 -33.155 ;
        RECT -74.285 -34.845 -73.955 -34.515 ;
        RECT -74.285 -36.205 -73.955 -35.875 ;
        RECT -74.285 -37.565 -73.955 -37.235 ;
        RECT -74.285 -38.925 -73.955 -38.595 ;
        RECT -74.285 -40.285 -73.955 -39.955 ;
        RECT -74.285 -41.645 -73.955 -41.315 ;
        RECT -74.285 -43.005 -73.955 -42.675 ;
        RECT -74.285 -44.365 -73.955 -44.035 ;
        RECT -74.285 -45.725 -73.955 -45.395 ;
        RECT -74.285 -47.085 -73.955 -46.755 ;
        RECT -74.285 -48.445 -73.955 -48.115 ;
        RECT -74.285 -49.805 -73.955 -49.475 ;
        RECT -74.285 -51.165 -73.955 -50.835 ;
        RECT -74.285 -52.525 -73.955 -52.195 ;
        RECT -74.285 -53.885 -73.955 -53.555 ;
        RECT -74.285 -55.245 -73.955 -54.915 ;
        RECT -74.285 -56.605 -73.955 -56.275 ;
        RECT -74.285 -57.965 -73.955 -57.635 ;
        RECT -74.285 -59.325 -73.955 -58.995 ;
        RECT -74.285 -60.685 -73.955 -60.355 ;
        RECT -74.285 -62.045 -73.955 -61.715 ;
        RECT -74.285 -63.405 -73.955 -63.075 ;
        RECT -74.285 -64.765 -73.955 -64.435 ;
        RECT -74.285 -66.125 -73.955 -65.795 ;
        RECT -74.285 -67.485 -73.955 -67.155 ;
        RECT -74.285 -68.845 -73.955 -68.515 ;
        RECT -74.285 -70.205 -73.955 -69.875 ;
        RECT -74.285 -71.565 -73.955 -71.235 ;
        RECT -74.285 -72.925 -73.955 -72.595 ;
        RECT -74.285 -74.285 -73.955 -73.955 ;
        RECT -74.285 -75.645 -73.955 -75.315 ;
        RECT -74.285 -77.005 -73.955 -76.675 ;
        RECT -74.285 -78.365 -73.955 -78.035 ;
        RECT -74.285 -79.725 -73.955 -79.395 ;
        RECT -74.285 -81.085 -73.955 -80.755 ;
        RECT -74.285 -82.445 -73.955 -82.115 ;
        RECT -74.285 -83.805 -73.955 -83.475 ;
        RECT -74.285 -85.165 -73.955 -84.835 ;
        RECT -74.285 -86.525 -73.955 -86.195 ;
        RECT -74.285 -87.885 -73.955 -87.555 ;
        RECT -74.285 -89.245 -73.955 -88.915 ;
        RECT -74.285 -90.605 -73.955 -90.275 ;
        RECT -74.285 -91.965 -73.955 -91.635 ;
        RECT -74.285 -93.325 -73.955 -92.995 ;
        RECT -74.285 -94.685 -73.955 -94.355 ;
        RECT -74.285 -96.045 -73.955 -95.715 ;
        RECT -74.285 -97.405 -73.955 -97.075 ;
        RECT -74.285 -98.765 -73.955 -98.435 ;
        RECT -74.285 -100.125 -73.955 -99.795 ;
        RECT -74.285 -101.485 -73.955 -101.155 ;
        RECT -74.285 -102.845 -73.955 -102.515 ;
        RECT -74.285 -104.205 -73.955 -103.875 ;
        RECT -74.285 -105.565 -73.955 -105.235 ;
        RECT -74.285 -106.925 -73.955 -106.595 ;
        RECT -74.285 -108.285 -73.955 -107.955 ;
        RECT -74.285 -109.645 -73.955 -109.315 ;
        RECT -74.285 -111.005 -73.955 -110.675 ;
        RECT -74.285 -112.365 -73.955 -112.035 ;
        RECT -74.285 -113.725 -73.955 -113.395 ;
        RECT -74.285 -115.085 -73.955 -114.755 ;
        RECT -74.285 -116.445 -73.955 -116.115 ;
        RECT -74.285 -117.805 -73.955 -117.475 ;
        RECT -74.285 -119.165 -73.955 -118.835 ;
        RECT -74.285 -120.525 -73.955 -120.195 ;
        RECT -74.285 -121.885 -73.955 -121.555 ;
        RECT -74.285 -123.245 -73.955 -122.915 ;
        RECT -74.285 -124.605 -73.955 -124.275 ;
        RECT -74.285 -125.965 -73.955 -125.635 ;
        RECT -74.285 -127.325 -73.955 -126.995 ;
        RECT -74.285 -128.685 -73.955 -128.355 ;
        RECT -74.285 -130.045 -73.955 -129.715 ;
        RECT -74.285 -131.405 -73.955 -131.075 ;
        RECT -74.285 -132.765 -73.955 -132.435 ;
        RECT -74.285 -134.125 -73.955 -133.795 ;
        RECT -74.285 -135.485 -73.955 -135.155 ;
        RECT -74.285 -136.845 -73.955 -136.515 ;
        RECT -74.285 -138.205 -73.955 -137.875 ;
        RECT -74.285 -139.565 -73.955 -139.235 ;
        RECT -74.285 -140.925 -73.955 -140.595 ;
        RECT -74.285 -142.285 -73.955 -141.955 ;
        RECT -74.285 -143.645 -73.955 -143.315 ;
        RECT -74.285 -145.005 -73.955 -144.675 ;
        RECT -74.285 -146.365 -73.955 -146.035 ;
        RECT -74.285 -147.725 -73.955 -147.395 ;
        RECT -74.285 -149.085 -73.955 -148.755 ;
        RECT -74.285 -150.445 -73.955 -150.115 ;
        RECT -74.285 -151.805 -73.955 -151.475 ;
        RECT -74.285 -153.165 -73.955 -152.835 ;
        RECT -74.285 -154.525 -73.955 -154.195 ;
        RECT -74.285 -155.885 -73.955 -155.555 ;
        RECT -74.285 -157.245 -73.955 -156.915 ;
        RECT -74.285 -158.605 -73.955 -158.275 ;
        RECT -74.285 -159.965 -73.955 -159.635 ;
        RECT -74.285 -161.325 -73.955 -160.995 ;
        RECT -74.285 -162.685 -73.955 -162.355 ;
        RECT -74.285 -164.045 -73.955 -163.715 ;
        RECT -74.285 -165.405 -73.955 -165.075 ;
        RECT -74.285 -166.765 -73.955 -166.435 ;
        RECT -74.285 -168.125 -73.955 -167.795 ;
        RECT -74.285 -169.485 -73.955 -169.155 ;
        RECT -74.285 -170.845 -73.955 -170.515 ;
        RECT -74.285 -172.205 -73.955 -171.875 ;
        RECT -74.285 -173.565 -73.955 -173.235 ;
        RECT -74.285 -174.925 -73.955 -174.595 ;
        RECT -74.285 -176.285 -73.955 -175.955 ;
        RECT -74.285 -177.645 -73.955 -177.315 ;
        RECT -74.285 -179.005 -73.955 -178.675 ;
        RECT -74.285 -180.365 -73.955 -180.035 ;
        RECT -74.285 -181.725 -73.955 -181.395 ;
        RECT -74.285 -183.085 -73.955 -182.755 ;
        RECT -74.285 -184.445 -73.955 -184.115 ;
        RECT -74.285 -185.805 -73.955 -185.475 ;
        RECT -74.285 -187.165 -73.955 -186.835 ;
        RECT -74.285 -188.525 -73.955 -188.195 ;
        RECT -74.285 -189.885 -73.955 -189.555 ;
        RECT -74.285 -191.245 -73.955 -190.915 ;
        RECT -74.285 -192.605 -73.955 -192.275 ;
        RECT -74.285 -193.965 -73.955 -193.635 ;
        RECT -74.285 -195.325 -73.955 -194.995 ;
        RECT -74.285 -196.685 -73.955 -196.355 ;
        RECT -74.285 -198.045 -73.955 -197.715 ;
        RECT -74.285 -199.405 -73.955 -199.075 ;
        RECT -74.285 -200.765 -73.955 -200.435 ;
        RECT -74.285 -202.125 -73.955 -201.795 ;
        RECT -74.285 -203.485 -73.955 -203.155 ;
        RECT -74.285 -204.845 -73.955 -204.515 ;
        RECT -74.285 -206.205 -73.955 -205.875 ;
        RECT -74.285 -207.565 -73.955 -207.235 ;
        RECT -74.285 -208.925 -73.955 -208.595 ;
        RECT -74.285 -210.285 -73.955 -209.955 ;
        RECT -74.285 -211.645 -73.955 -211.315 ;
        RECT -74.285 -213.005 -73.955 -212.675 ;
        RECT -74.285 -214.365 -73.955 -214.035 ;
        RECT -74.285 -215.725 -73.955 -215.395 ;
        RECT -74.285 -217.085 -73.955 -216.755 ;
        RECT -74.285 -218.445 -73.955 -218.115 ;
        RECT -74.285 -219.805 -73.955 -219.475 ;
        RECT -74.285 -221.165 -73.955 -220.835 ;
        RECT -74.285 -222.525 -73.955 -222.195 ;
        RECT -74.285 -223.885 -73.955 -223.555 ;
        RECT -74.285 -225.245 -73.955 -224.915 ;
        RECT -74.285 -227.965 -73.955 -227.635 ;
        RECT -74.285 -230.685 -73.955 -230.355 ;
        RECT -74.285 -232.045 -73.955 -231.715 ;
        RECT -74.285 -233.225 -73.955 -232.895 ;
        RECT -74.285 -234.765 -73.955 -234.435 ;
        RECT -74.285 -236.125 -73.955 -235.795 ;
        RECT -74.285 -237.485 -73.955 -237.155 ;
        RECT -74.285 -238.845 -73.955 -238.515 ;
        RECT -74.285 -241.09 -73.955 -239.96 ;
        RECT -74.28 -241.205 -73.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.925 -81.085 -72.595 -80.755 ;
        RECT -72.925 -82.445 -72.595 -82.115 ;
        RECT -72.925 -83.805 -72.595 -83.475 ;
        RECT -72.925 -85.165 -72.595 -84.835 ;
        RECT -72.925 -86.525 -72.595 -86.195 ;
        RECT -72.925 -87.885 -72.595 -87.555 ;
        RECT -72.925 -89.245 -72.595 -88.915 ;
        RECT -72.925 -90.605 -72.595 -90.275 ;
        RECT -72.925 -91.965 -72.595 -91.635 ;
        RECT -72.925 -93.325 -72.595 -92.995 ;
        RECT -72.925 -94.685 -72.595 -94.355 ;
        RECT -72.925 -96.045 -72.595 -95.715 ;
        RECT -72.925 -97.405 -72.595 -97.075 ;
        RECT -72.925 -98.765 -72.595 -98.435 ;
        RECT -72.925 -100.125 -72.595 -99.795 ;
        RECT -72.925 -101.485 -72.595 -101.155 ;
        RECT -72.925 -102.845 -72.595 -102.515 ;
        RECT -72.925 -104.205 -72.595 -103.875 ;
        RECT -72.925 -105.565 -72.595 -105.235 ;
        RECT -72.925 -106.925 -72.595 -106.595 ;
        RECT -72.925 -108.285 -72.595 -107.955 ;
        RECT -72.925 -109.645 -72.595 -109.315 ;
        RECT -72.925 -111.005 -72.595 -110.675 ;
        RECT -72.925 -112.365 -72.595 -112.035 ;
        RECT -72.925 -113.725 -72.595 -113.395 ;
        RECT -72.925 -115.085 -72.595 -114.755 ;
        RECT -72.925 -116.445 -72.595 -116.115 ;
        RECT -72.925 -117.805 -72.595 -117.475 ;
        RECT -72.925 -119.165 -72.595 -118.835 ;
        RECT -72.925 -120.525 -72.595 -120.195 ;
        RECT -72.925 -121.885 -72.595 -121.555 ;
        RECT -72.925 -123.245 -72.595 -122.915 ;
        RECT -72.925 -124.605 -72.595 -124.275 ;
        RECT -72.925 -125.965 -72.595 -125.635 ;
        RECT -72.925 -127.325 -72.595 -126.995 ;
        RECT -72.925 -128.685 -72.595 -128.355 ;
        RECT -72.925 -130.045 -72.595 -129.715 ;
        RECT -72.925 -131.405 -72.595 -131.075 ;
        RECT -72.925 -132.765 -72.595 -132.435 ;
        RECT -72.925 -134.125 -72.595 -133.795 ;
        RECT -72.925 -135.485 -72.595 -135.155 ;
        RECT -72.925 -136.845 -72.595 -136.515 ;
        RECT -72.925 -138.205 -72.595 -137.875 ;
        RECT -72.925 -139.565 -72.595 -139.235 ;
        RECT -72.925 -140.925 -72.595 -140.595 ;
        RECT -72.925 -142.285 -72.595 -141.955 ;
        RECT -72.925 -143.645 -72.595 -143.315 ;
        RECT -72.925 -145.005 -72.595 -144.675 ;
        RECT -72.925 -146.365 -72.595 -146.035 ;
        RECT -72.925 -147.725 -72.595 -147.395 ;
        RECT -72.925 -149.085 -72.595 -148.755 ;
        RECT -72.92 -149.76 -72.6 245.285 ;
        RECT -72.925 244.04 -72.595 245.17 ;
        RECT -72.925 242.595 -72.595 242.925 ;
        RECT -72.925 241.235 -72.595 241.565 ;
        RECT -72.925 239.875 -72.595 240.205 ;
        RECT -72.925 238.515 -72.595 238.845 ;
        RECT -72.925 237.155 -72.595 237.485 ;
        RECT -72.925 235.795 -72.595 236.125 ;
        RECT -72.925 234.435 -72.595 234.765 ;
        RECT -72.925 233.075 -72.595 233.405 ;
        RECT -72.925 231.715 -72.595 232.045 ;
        RECT -72.925 230.355 -72.595 230.685 ;
        RECT -72.925 228.995 -72.595 229.325 ;
        RECT -72.925 227.635 -72.595 227.965 ;
        RECT -72.925 226.275 -72.595 226.605 ;
        RECT -72.925 224.915 -72.595 225.245 ;
        RECT -72.925 223.555 -72.595 223.885 ;
        RECT -72.925 222.195 -72.595 222.525 ;
        RECT -72.925 220.835 -72.595 221.165 ;
        RECT -72.925 219.475 -72.595 219.805 ;
        RECT -72.925 218.115 -72.595 218.445 ;
        RECT -72.925 216.755 -72.595 217.085 ;
        RECT -72.925 215.395 -72.595 215.725 ;
        RECT -72.925 214.035 -72.595 214.365 ;
        RECT -72.925 212.675 -72.595 213.005 ;
        RECT -72.925 211.315 -72.595 211.645 ;
        RECT -72.925 209.955 -72.595 210.285 ;
        RECT -72.925 208.595 -72.595 208.925 ;
        RECT -72.925 207.235 -72.595 207.565 ;
        RECT -72.925 205.875 -72.595 206.205 ;
        RECT -72.925 204.515 -72.595 204.845 ;
        RECT -72.925 203.155 -72.595 203.485 ;
        RECT -72.925 201.795 -72.595 202.125 ;
        RECT -72.925 200.435 -72.595 200.765 ;
        RECT -72.925 199.075 -72.595 199.405 ;
        RECT -72.925 197.715 -72.595 198.045 ;
        RECT -72.925 196.355 -72.595 196.685 ;
        RECT -72.925 194.995 -72.595 195.325 ;
        RECT -72.925 193.635 -72.595 193.965 ;
        RECT -72.925 192.275 -72.595 192.605 ;
        RECT -72.925 190.915 -72.595 191.245 ;
        RECT -72.925 189.555 -72.595 189.885 ;
        RECT -72.925 188.195 -72.595 188.525 ;
        RECT -72.925 186.835 -72.595 187.165 ;
        RECT -72.925 185.475 -72.595 185.805 ;
        RECT -72.925 184.115 -72.595 184.445 ;
        RECT -72.925 182.755 -72.595 183.085 ;
        RECT -72.925 181.395 -72.595 181.725 ;
        RECT -72.925 180.035 -72.595 180.365 ;
        RECT -72.925 178.675 -72.595 179.005 ;
        RECT -72.925 177.315 -72.595 177.645 ;
        RECT -72.925 175.955 -72.595 176.285 ;
        RECT -72.925 174.595 -72.595 174.925 ;
        RECT -72.925 173.235 -72.595 173.565 ;
        RECT -72.925 171.875 -72.595 172.205 ;
        RECT -72.925 170.515 -72.595 170.845 ;
        RECT -72.925 169.155 -72.595 169.485 ;
        RECT -72.925 167.795 -72.595 168.125 ;
        RECT -72.925 166.435 -72.595 166.765 ;
        RECT -72.925 165.075 -72.595 165.405 ;
        RECT -72.925 163.715 -72.595 164.045 ;
        RECT -72.925 162.355 -72.595 162.685 ;
        RECT -72.925 160.995 -72.595 161.325 ;
        RECT -72.925 159.635 -72.595 159.965 ;
        RECT -72.925 158.275 -72.595 158.605 ;
        RECT -72.925 156.915 -72.595 157.245 ;
        RECT -72.925 155.555 -72.595 155.885 ;
        RECT -72.925 154.195 -72.595 154.525 ;
        RECT -72.925 152.835 -72.595 153.165 ;
        RECT -72.925 151.475 -72.595 151.805 ;
        RECT -72.925 150.115 -72.595 150.445 ;
        RECT -72.925 148.755 -72.595 149.085 ;
        RECT -72.925 147.395 -72.595 147.725 ;
        RECT -72.925 146.035 -72.595 146.365 ;
        RECT -72.925 144.675 -72.595 145.005 ;
        RECT -72.925 143.315 -72.595 143.645 ;
        RECT -72.925 141.955 -72.595 142.285 ;
        RECT -72.925 140.595 -72.595 140.925 ;
        RECT -72.925 139.235 -72.595 139.565 ;
        RECT -72.925 137.875 -72.595 138.205 ;
        RECT -72.925 136.515 -72.595 136.845 ;
        RECT -72.925 135.155 -72.595 135.485 ;
        RECT -72.925 133.795 -72.595 134.125 ;
        RECT -72.925 132.435 -72.595 132.765 ;
        RECT -72.925 131.075 -72.595 131.405 ;
        RECT -72.925 129.715 -72.595 130.045 ;
        RECT -72.925 128.355 -72.595 128.685 ;
        RECT -72.925 126.995 -72.595 127.325 ;
        RECT -72.925 125.635 -72.595 125.965 ;
        RECT -72.925 124.275 -72.595 124.605 ;
        RECT -72.925 122.915 -72.595 123.245 ;
        RECT -72.925 121.555 -72.595 121.885 ;
        RECT -72.925 120.195 -72.595 120.525 ;
        RECT -72.925 118.835 -72.595 119.165 ;
        RECT -72.925 117.475 -72.595 117.805 ;
        RECT -72.925 116.115 -72.595 116.445 ;
        RECT -72.925 114.755 -72.595 115.085 ;
        RECT -72.925 113.395 -72.595 113.725 ;
        RECT -72.925 112.035 -72.595 112.365 ;
        RECT -72.925 110.675 -72.595 111.005 ;
        RECT -72.925 109.315 -72.595 109.645 ;
        RECT -72.925 107.955 -72.595 108.285 ;
        RECT -72.925 106.595 -72.595 106.925 ;
        RECT -72.925 105.235 -72.595 105.565 ;
        RECT -72.925 103.875 -72.595 104.205 ;
        RECT -72.925 102.515 -72.595 102.845 ;
        RECT -72.925 101.155 -72.595 101.485 ;
        RECT -72.925 99.795 -72.595 100.125 ;
        RECT -72.925 98.435 -72.595 98.765 ;
        RECT -72.925 97.075 -72.595 97.405 ;
        RECT -72.925 95.715 -72.595 96.045 ;
        RECT -72.925 94.355 -72.595 94.685 ;
        RECT -72.925 92.995 -72.595 93.325 ;
        RECT -72.925 91.635 -72.595 91.965 ;
        RECT -72.925 90.275 -72.595 90.605 ;
        RECT -72.925 88.915 -72.595 89.245 ;
        RECT -72.925 87.555 -72.595 87.885 ;
        RECT -72.925 86.195 -72.595 86.525 ;
        RECT -72.925 84.835 -72.595 85.165 ;
        RECT -72.925 83.475 -72.595 83.805 ;
        RECT -72.925 82.115 -72.595 82.445 ;
        RECT -72.925 80.755 -72.595 81.085 ;
        RECT -72.925 79.395 -72.595 79.725 ;
        RECT -72.925 78.035 -72.595 78.365 ;
        RECT -72.925 76.675 -72.595 77.005 ;
        RECT -72.925 75.315 -72.595 75.645 ;
        RECT -72.925 73.955 -72.595 74.285 ;
        RECT -72.925 72.595 -72.595 72.925 ;
        RECT -72.925 71.235 -72.595 71.565 ;
        RECT -72.925 69.875 -72.595 70.205 ;
        RECT -72.925 68.515 -72.595 68.845 ;
        RECT -72.925 67.155 -72.595 67.485 ;
        RECT -72.925 65.795 -72.595 66.125 ;
        RECT -72.925 64.435 -72.595 64.765 ;
        RECT -72.925 63.075 -72.595 63.405 ;
        RECT -72.925 61.715 -72.595 62.045 ;
        RECT -72.925 60.355 -72.595 60.685 ;
        RECT -72.925 58.995 -72.595 59.325 ;
        RECT -72.925 57.635 -72.595 57.965 ;
        RECT -72.925 56.275 -72.595 56.605 ;
        RECT -72.925 54.915 -72.595 55.245 ;
        RECT -72.925 53.555 -72.595 53.885 ;
        RECT -72.925 52.195 -72.595 52.525 ;
        RECT -72.925 50.835 -72.595 51.165 ;
        RECT -72.925 49.475 -72.595 49.805 ;
        RECT -72.925 48.115 -72.595 48.445 ;
        RECT -72.925 46.755 -72.595 47.085 ;
        RECT -72.925 45.395 -72.595 45.725 ;
        RECT -72.925 44.035 -72.595 44.365 ;
        RECT -72.925 42.675 -72.595 43.005 ;
        RECT -72.925 41.315 -72.595 41.645 ;
        RECT -72.925 39.955 -72.595 40.285 ;
        RECT -72.925 38.595 -72.595 38.925 ;
        RECT -72.925 37.235 -72.595 37.565 ;
        RECT -72.925 35.875 -72.595 36.205 ;
        RECT -72.925 34.515 -72.595 34.845 ;
        RECT -72.925 33.155 -72.595 33.485 ;
        RECT -72.925 31.795 -72.595 32.125 ;
        RECT -72.925 30.435 -72.595 30.765 ;
        RECT -72.925 29.075 -72.595 29.405 ;
        RECT -72.925 27.715 -72.595 28.045 ;
        RECT -72.925 26.355 -72.595 26.685 ;
        RECT -72.925 24.995 -72.595 25.325 ;
        RECT -72.925 23.635 -72.595 23.965 ;
        RECT -72.925 22.275 -72.595 22.605 ;
        RECT -72.925 20.915 -72.595 21.245 ;
        RECT -72.925 19.555 -72.595 19.885 ;
        RECT -72.925 18.195 -72.595 18.525 ;
        RECT -72.925 16.835 -72.595 17.165 ;
        RECT -72.925 15.475 -72.595 15.805 ;
        RECT -72.925 14.115 -72.595 14.445 ;
        RECT -72.925 12.755 -72.595 13.085 ;
        RECT -72.925 11.395 -72.595 11.725 ;
        RECT -72.925 10.035 -72.595 10.365 ;
        RECT -72.925 8.675 -72.595 9.005 ;
        RECT -72.925 7.315 -72.595 7.645 ;
        RECT -72.925 5.955 -72.595 6.285 ;
        RECT -72.925 4.595 -72.595 4.925 ;
        RECT -72.925 3.235 -72.595 3.565 ;
        RECT -72.925 1.875 -72.595 2.205 ;
        RECT -72.925 0.515 -72.595 0.845 ;
        RECT -72.925 -0.845 -72.595 -0.515 ;
        RECT -72.925 -2.205 -72.595 -1.875 ;
        RECT -72.925 -3.565 -72.595 -3.235 ;
        RECT -72.925 -4.925 -72.595 -4.595 ;
        RECT -72.925 -6.285 -72.595 -5.955 ;
        RECT -72.925 -7.645 -72.595 -7.315 ;
        RECT -72.925 -9.005 -72.595 -8.675 ;
        RECT -72.925 -10.365 -72.595 -10.035 ;
        RECT -72.925 -11.725 -72.595 -11.395 ;
        RECT -72.925 -13.085 -72.595 -12.755 ;
        RECT -72.925 -14.445 -72.595 -14.115 ;
        RECT -72.925 -15.805 -72.595 -15.475 ;
        RECT -72.925 -17.165 -72.595 -16.835 ;
        RECT -72.925 -18.525 -72.595 -18.195 ;
        RECT -72.925 -19.885 -72.595 -19.555 ;
        RECT -72.925 -21.245 -72.595 -20.915 ;
        RECT -72.925 -22.605 -72.595 -22.275 ;
        RECT -72.925 -23.965 -72.595 -23.635 ;
        RECT -72.925 -25.325 -72.595 -24.995 ;
        RECT -72.925 -26.685 -72.595 -26.355 ;
        RECT -72.925 -28.045 -72.595 -27.715 ;
        RECT -72.925 -29.405 -72.595 -29.075 ;
        RECT -72.925 -30.765 -72.595 -30.435 ;
        RECT -72.925 -32.125 -72.595 -31.795 ;
        RECT -72.925 -33.485 -72.595 -33.155 ;
        RECT -72.925 -34.845 -72.595 -34.515 ;
        RECT -72.925 -36.205 -72.595 -35.875 ;
        RECT -72.925 -37.565 -72.595 -37.235 ;
        RECT -72.925 -38.925 -72.595 -38.595 ;
        RECT -72.925 -40.285 -72.595 -39.955 ;
        RECT -72.925 -41.645 -72.595 -41.315 ;
        RECT -72.925 -43.005 -72.595 -42.675 ;
        RECT -72.925 -44.365 -72.595 -44.035 ;
        RECT -72.925 -45.725 -72.595 -45.395 ;
        RECT -72.925 -47.085 -72.595 -46.755 ;
        RECT -72.925 -48.445 -72.595 -48.115 ;
        RECT -72.925 -49.805 -72.595 -49.475 ;
        RECT -72.925 -51.165 -72.595 -50.835 ;
        RECT -72.925 -52.525 -72.595 -52.195 ;
        RECT -72.925 -53.885 -72.595 -53.555 ;
        RECT -72.925 -55.245 -72.595 -54.915 ;
        RECT -72.925 -56.605 -72.595 -56.275 ;
        RECT -72.925 -57.965 -72.595 -57.635 ;
        RECT -72.925 -59.325 -72.595 -58.995 ;
        RECT -72.925 -60.685 -72.595 -60.355 ;
        RECT -72.925 -62.045 -72.595 -61.715 ;
        RECT -72.925 -63.405 -72.595 -63.075 ;
        RECT -72.925 -64.765 -72.595 -64.435 ;
        RECT -72.925 -66.125 -72.595 -65.795 ;
        RECT -72.925 -67.485 -72.595 -67.155 ;
        RECT -72.925 -68.845 -72.595 -68.515 ;
        RECT -72.925 -70.205 -72.595 -69.875 ;
        RECT -72.925 -71.565 -72.595 -71.235 ;
        RECT -72.925 -72.925 -72.595 -72.595 ;
        RECT -72.925 -74.285 -72.595 -73.955 ;
        RECT -72.925 -75.645 -72.595 -75.315 ;
        RECT -72.925 -77.005 -72.595 -76.675 ;
        RECT -72.925 -78.365 -72.595 -78.035 ;
        RECT -72.925 -79.725 -72.595 -79.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.725 244.04 -79.395 245.17 ;
        RECT -79.725 242.595 -79.395 242.925 ;
        RECT -79.725 241.235 -79.395 241.565 ;
        RECT -79.725 239.875 -79.395 240.205 ;
        RECT -79.725 238.515 -79.395 238.845 ;
        RECT -79.725 237.155 -79.395 237.485 ;
        RECT -79.725 235.795 -79.395 236.125 ;
        RECT -79.725 234.435 -79.395 234.765 ;
        RECT -79.725 233.075 -79.395 233.405 ;
        RECT -79.725 231.715 -79.395 232.045 ;
        RECT -79.725 230.355 -79.395 230.685 ;
        RECT -79.725 228.995 -79.395 229.325 ;
        RECT -79.725 227.635 -79.395 227.965 ;
        RECT -79.725 226.275 -79.395 226.605 ;
        RECT -79.725 224.915 -79.395 225.245 ;
        RECT -79.725 223.555 -79.395 223.885 ;
        RECT -79.725 222.195 -79.395 222.525 ;
        RECT -79.725 220.835 -79.395 221.165 ;
        RECT -79.725 219.475 -79.395 219.805 ;
        RECT -79.725 218.115 -79.395 218.445 ;
        RECT -79.725 216.755 -79.395 217.085 ;
        RECT -79.725 215.395 -79.395 215.725 ;
        RECT -79.725 214.035 -79.395 214.365 ;
        RECT -79.725 212.675 -79.395 213.005 ;
        RECT -79.725 211.315 -79.395 211.645 ;
        RECT -79.725 209.955 -79.395 210.285 ;
        RECT -79.725 208.595 -79.395 208.925 ;
        RECT -79.725 207.235 -79.395 207.565 ;
        RECT -79.725 205.875 -79.395 206.205 ;
        RECT -79.725 204.515 -79.395 204.845 ;
        RECT -79.725 203.155 -79.395 203.485 ;
        RECT -79.725 201.795 -79.395 202.125 ;
        RECT -79.725 200.435 -79.395 200.765 ;
        RECT -79.725 199.075 -79.395 199.405 ;
        RECT -79.725 197.715 -79.395 198.045 ;
        RECT -79.725 196.355 -79.395 196.685 ;
        RECT -79.725 194.995 -79.395 195.325 ;
        RECT -79.725 193.635 -79.395 193.965 ;
        RECT -79.725 192.275 -79.395 192.605 ;
        RECT -79.725 190.915 -79.395 191.245 ;
        RECT -79.725 189.555 -79.395 189.885 ;
        RECT -79.725 188.195 -79.395 188.525 ;
        RECT -79.725 186.835 -79.395 187.165 ;
        RECT -79.725 185.475 -79.395 185.805 ;
        RECT -79.725 184.115 -79.395 184.445 ;
        RECT -79.725 182.755 -79.395 183.085 ;
        RECT -79.725 181.395 -79.395 181.725 ;
        RECT -79.725 180.035 -79.395 180.365 ;
        RECT -79.725 178.675 -79.395 179.005 ;
        RECT -79.725 177.315 -79.395 177.645 ;
        RECT -79.725 175.955 -79.395 176.285 ;
        RECT -79.725 174.595 -79.395 174.925 ;
        RECT -79.725 173.235 -79.395 173.565 ;
        RECT -79.725 171.875 -79.395 172.205 ;
        RECT -79.725 170.515 -79.395 170.845 ;
        RECT -79.725 169.155 -79.395 169.485 ;
        RECT -79.725 167.795 -79.395 168.125 ;
        RECT -79.725 166.435 -79.395 166.765 ;
        RECT -79.725 165.075 -79.395 165.405 ;
        RECT -79.725 163.715 -79.395 164.045 ;
        RECT -79.725 162.355 -79.395 162.685 ;
        RECT -79.725 160.995 -79.395 161.325 ;
        RECT -79.725 159.635 -79.395 159.965 ;
        RECT -79.725 158.275 -79.395 158.605 ;
        RECT -79.725 156.915 -79.395 157.245 ;
        RECT -79.725 155.555 -79.395 155.885 ;
        RECT -79.725 154.195 -79.395 154.525 ;
        RECT -79.725 152.835 -79.395 153.165 ;
        RECT -79.725 151.475 -79.395 151.805 ;
        RECT -79.725 150.115 -79.395 150.445 ;
        RECT -79.725 148.755 -79.395 149.085 ;
        RECT -79.725 147.395 -79.395 147.725 ;
        RECT -79.725 146.035 -79.395 146.365 ;
        RECT -79.725 144.675 -79.395 145.005 ;
        RECT -79.725 143.315 -79.395 143.645 ;
        RECT -79.725 141.955 -79.395 142.285 ;
        RECT -79.725 140.595 -79.395 140.925 ;
        RECT -79.725 139.235 -79.395 139.565 ;
        RECT -79.725 137.875 -79.395 138.205 ;
        RECT -79.725 136.515 -79.395 136.845 ;
        RECT -79.725 135.155 -79.395 135.485 ;
        RECT -79.725 133.795 -79.395 134.125 ;
        RECT -79.725 132.435 -79.395 132.765 ;
        RECT -79.725 131.075 -79.395 131.405 ;
        RECT -79.725 129.715 -79.395 130.045 ;
        RECT -79.725 128.355 -79.395 128.685 ;
        RECT -79.725 126.995 -79.395 127.325 ;
        RECT -79.725 125.635 -79.395 125.965 ;
        RECT -79.725 124.275 -79.395 124.605 ;
        RECT -79.725 122.915 -79.395 123.245 ;
        RECT -79.725 121.555 -79.395 121.885 ;
        RECT -79.725 120.195 -79.395 120.525 ;
        RECT -79.725 118.835 -79.395 119.165 ;
        RECT -79.725 117.475 -79.395 117.805 ;
        RECT -79.725 116.115 -79.395 116.445 ;
        RECT -79.725 114.755 -79.395 115.085 ;
        RECT -79.725 113.395 -79.395 113.725 ;
        RECT -79.725 112.035 -79.395 112.365 ;
        RECT -79.725 110.675 -79.395 111.005 ;
        RECT -79.725 109.315 -79.395 109.645 ;
        RECT -79.725 107.955 -79.395 108.285 ;
        RECT -79.725 106.595 -79.395 106.925 ;
        RECT -79.725 105.235 -79.395 105.565 ;
        RECT -79.725 103.875 -79.395 104.205 ;
        RECT -79.725 102.515 -79.395 102.845 ;
        RECT -79.725 101.155 -79.395 101.485 ;
        RECT -79.725 99.795 -79.395 100.125 ;
        RECT -79.725 98.435 -79.395 98.765 ;
        RECT -79.725 97.075 -79.395 97.405 ;
        RECT -79.725 95.715 -79.395 96.045 ;
        RECT -79.725 94.355 -79.395 94.685 ;
        RECT -79.725 92.995 -79.395 93.325 ;
        RECT -79.725 91.635 -79.395 91.965 ;
        RECT -79.725 90.275 -79.395 90.605 ;
        RECT -79.725 88.915 -79.395 89.245 ;
        RECT -79.725 87.555 -79.395 87.885 ;
        RECT -79.725 86.195 -79.395 86.525 ;
        RECT -79.725 84.835 -79.395 85.165 ;
        RECT -79.725 83.475 -79.395 83.805 ;
        RECT -79.725 82.115 -79.395 82.445 ;
        RECT -79.725 80.755 -79.395 81.085 ;
        RECT -79.725 79.395 -79.395 79.725 ;
        RECT -79.725 78.035 -79.395 78.365 ;
        RECT -79.725 76.675 -79.395 77.005 ;
        RECT -79.725 75.315 -79.395 75.645 ;
        RECT -79.725 73.955 -79.395 74.285 ;
        RECT -79.725 72.595 -79.395 72.925 ;
        RECT -79.725 71.235 -79.395 71.565 ;
        RECT -79.725 69.875 -79.395 70.205 ;
        RECT -79.725 68.515 -79.395 68.845 ;
        RECT -79.725 67.155 -79.395 67.485 ;
        RECT -79.725 65.795 -79.395 66.125 ;
        RECT -79.725 64.435 -79.395 64.765 ;
        RECT -79.725 63.075 -79.395 63.405 ;
        RECT -79.725 61.715 -79.395 62.045 ;
        RECT -79.725 60.355 -79.395 60.685 ;
        RECT -79.725 58.995 -79.395 59.325 ;
        RECT -79.725 57.635 -79.395 57.965 ;
        RECT -79.725 56.275 -79.395 56.605 ;
        RECT -79.725 54.915 -79.395 55.245 ;
        RECT -79.725 53.555 -79.395 53.885 ;
        RECT -79.725 52.195 -79.395 52.525 ;
        RECT -79.725 50.835 -79.395 51.165 ;
        RECT -79.725 49.475 -79.395 49.805 ;
        RECT -79.725 48.115 -79.395 48.445 ;
        RECT -79.725 46.755 -79.395 47.085 ;
        RECT -79.725 45.395 -79.395 45.725 ;
        RECT -79.725 44.035 -79.395 44.365 ;
        RECT -79.725 42.675 -79.395 43.005 ;
        RECT -79.725 41.315 -79.395 41.645 ;
        RECT -79.725 39.955 -79.395 40.285 ;
        RECT -79.725 38.595 -79.395 38.925 ;
        RECT -79.725 37.235 -79.395 37.565 ;
        RECT -79.725 35.875 -79.395 36.205 ;
        RECT -79.725 34.515 -79.395 34.845 ;
        RECT -79.725 33.155 -79.395 33.485 ;
        RECT -79.725 31.795 -79.395 32.125 ;
        RECT -79.725 30.435 -79.395 30.765 ;
        RECT -79.725 29.075 -79.395 29.405 ;
        RECT -79.725 27.715 -79.395 28.045 ;
        RECT -79.725 26.355 -79.395 26.685 ;
        RECT -79.725 24.995 -79.395 25.325 ;
        RECT -79.725 23.635 -79.395 23.965 ;
        RECT -79.725 22.275 -79.395 22.605 ;
        RECT -79.725 20.915 -79.395 21.245 ;
        RECT -79.725 19.555 -79.395 19.885 ;
        RECT -79.725 18.195 -79.395 18.525 ;
        RECT -79.725 16.835 -79.395 17.165 ;
        RECT -79.725 15.475 -79.395 15.805 ;
        RECT -79.725 14.115 -79.395 14.445 ;
        RECT -79.725 12.755 -79.395 13.085 ;
        RECT -79.725 11.395 -79.395 11.725 ;
        RECT -79.725 10.035 -79.395 10.365 ;
        RECT -79.725 8.675 -79.395 9.005 ;
        RECT -79.725 7.315 -79.395 7.645 ;
        RECT -79.725 5.955 -79.395 6.285 ;
        RECT -79.725 4.595 -79.395 4.925 ;
        RECT -79.725 3.235 -79.395 3.565 ;
        RECT -79.725 1.875 -79.395 2.205 ;
        RECT -79.725 0.515 -79.395 0.845 ;
        RECT -79.725 -0.845 -79.395 -0.515 ;
        RECT -79.725 -2.205 -79.395 -1.875 ;
        RECT -79.725 -3.565 -79.395 -3.235 ;
        RECT -79.725 -4.925 -79.395 -4.595 ;
        RECT -79.725 -6.285 -79.395 -5.955 ;
        RECT -79.725 -7.645 -79.395 -7.315 ;
        RECT -79.725 -9.005 -79.395 -8.675 ;
        RECT -79.725 -10.365 -79.395 -10.035 ;
        RECT -79.725 -11.725 -79.395 -11.395 ;
        RECT -79.725 -13.085 -79.395 -12.755 ;
        RECT -79.725 -14.445 -79.395 -14.115 ;
        RECT -79.725 -15.805 -79.395 -15.475 ;
        RECT -79.725 -17.165 -79.395 -16.835 ;
        RECT -79.725 -18.525 -79.395 -18.195 ;
        RECT -79.725 -19.885 -79.395 -19.555 ;
        RECT -79.725 -21.245 -79.395 -20.915 ;
        RECT -79.725 -22.605 -79.395 -22.275 ;
        RECT -79.725 -23.965 -79.395 -23.635 ;
        RECT -79.725 -25.325 -79.395 -24.995 ;
        RECT -79.725 -26.685 -79.395 -26.355 ;
        RECT -79.725 -28.045 -79.395 -27.715 ;
        RECT -79.725 -29.405 -79.395 -29.075 ;
        RECT -79.725 -30.765 -79.395 -30.435 ;
        RECT -79.725 -32.125 -79.395 -31.795 ;
        RECT -79.725 -33.485 -79.395 -33.155 ;
        RECT -79.725 -34.845 -79.395 -34.515 ;
        RECT -79.725 -36.205 -79.395 -35.875 ;
        RECT -79.725 -37.565 -79.395 -37.235 ;
        RECT -79.725 -38.925 -79.395 -38.595 ;
        RECT -79.725 -40.285 -79.395 -39.955 ;
        RECT -79.725 -41.645 -79.395 -41.315 ;
        RECT -79.725 -43.005 -79.395 -42.675 ;
        RECT -79.725 -44.365 -79.395 -44.035 ;
        RECT -79.725 -45.725 -79.395 -45.395 ;
        RECT -79.725 -47.085 -79.395 -46.755 ;
        RECT -79.725 -48.445 -79.395 -48.115 ;
        RECT -79.725 -49.805 -79.395 -49.475 ;
        RECT -79.725 -51.165 -79.395 -50.835 ;
        RECT -79.725 -52.525 -79.395 -52.195 ;
        RECT -79.725 -53.885 -79.395 -53.555 ;
        RECT -79.725 -55.245 -79.395 -54.915 ;
        RECT -79.725 -56.605 -79.395 -56.275 ;
        RECT -79.725 -57.965 -79.395 -57.635 ;
        RECT -79.725 -59.325 -79.395 -58.995 ;
        RECT -79.725 -60.685 -79.395 -60.355 ;
        RECT -79.725 -62.045 -79.395 -61.715 ;
        RECT -79.725 -63.405 -79.395 -63.075 ;
        RECT -79.725 -64.765 -79.395 -64.435 ;
        RECT -79.725 -66.125 -79.395 -65.795 ;
        RECT -79.725 -67.485 -79.395 -67.155 ;
        RECT -79.725 -68.845 -79.395 -68.515 ;
        RECT -79.725 -70.205 -79.395 -69.875 ;
        RECT -79.725 -71.565 -79.395 -71.235 ;
        RECT -79.725 -72.925 -79.395 -72.595 ;
        RECT -79.725 -74.285 -79.395 -73.955 ;
        RECT -79.725 -75.645 -79.395 -75.315 ;
        RECT -79.725 -77.005 -79.395 -76.675 ;
        RECT -79.725 -78.365 -79.395 -78.035 ;
        RECT -79.725 -79.725 -79.395 -79.395 ;
        RECT -79.725 -81.085 -79.395 -80.755 ;
        RECT -79.725 -82.445 -79.395 -82.115 ;
        RECT -79.725 -83.805 -79.395 -83.475 ;
        RECT -79.725 -85.165 -79.395 -84.835 ;
        RECT -79.725 -86.525 -79.395 -86.195 ;
        RECT -79.725 -87.885 -79.395 -87.555 ;
        RECT -79.725 -89.245 -79.395 -88.915 ;
        RECT -79.725 -90.605 -79.395 -90.275 ;
        RECT -79.725 -91.965 -79.395 -91.635 ;
        RECT -79.725 -93.325 -79.395 -92.995 ;
        RECT -79.725 -94.685 -79.395 -94.355 ;
        RECT -79.725 -96.045 -79.395 -95.715 ;
        RECT -79.725 -97.405 -79.395 -97.075 ;
        RECT -79.725 -98.765 -79.395 -98.435 ;
        RECT -79.725 -100.125 -79.395 -99.795 ;
        RECT -79.725 -101.485 -79.395 -101.155 ;
        RECT -79.725 -102.845 -79.395 -102.515 ;
        RECT -79.725 -104.205 -79.395 -103.875 ;
        RECT -79.725 -105.565 -79.395 -105.235 ;
        RECT -79.725 -106.925 -79.395 -106.595 ;
        RECT -79.725 -108.285 -79.395 -107.955 ;
        RECT -79.725 -109.645 -79.395 -109.315 ;
        RECT -79.725 -111.005 -79.395 -110.675 ;
        RECT -79.725 -112.365 -79.395 -112.035 ;
        RECT -79.725 -113.725 -79.395 -113.395 ;
        RECT -79.725 -115.085 -79.395 -114.755 ;
        RECT -79.725 -116.445 -79.395 -116.115 ;
        RECT -79.725 -117.805 -79.395 -117.475 ;
        RECT -79.725 -119.165 -79.395 -118.835 ;
        RECT -79.725 -120.525 -79.395 -120.195 ;
        RECT -79.725 -121.885 -79.395 -121.555 ;
        RECT -79.725 -123.245 -79.395 -122.915 ;
        RECT -79.725 -124.605 -79.395 -124.275 ;
        RECT -79.725 -125.965 -79.395 -125.635 ;
        RECT -79.725 -127.325 -79.395 -126.995 ;
        RECT -79.725 -128.685 -79.395 -128.355 ;
        RECT -79.725 -130.045 -79.395 -129.715 ;
        RECT -79.725 -131.405 -79.395 -131.075 ;
        RECT -79.725 -132.765 -79.395 -132.435 ;
        RECT -79.725 -134.125 -79.395 -133.795 ;
        RECT -79.725 -135.485 -79.395 -135.155 ;
        RECT -79.725 -136.845 -79.395 -136.515 ;
        RECT -79.725 -138.205 -79.395 -137.875 ;
        RECT -79.725 -139.565 -79.395 -139.235 ;
        RECT -79.725 -140.925 -79.395 -140.595 ;
        RECT -79.725 -142.285 -79.395 -141.955 ;
        RECT -79.725 -143.645 -79.395 -143.315 ;
        RECT -79.725 -145.005 -79.395 -144.675 ;
        RECT -79.725 -146.365 -79.395 -146.035 ;
        RECT -79.725 -147.725 -79.395 -147.395 ;
        RECT -79.725 -149.085 -79.395 -148.755 ;
        RECT -79.725 -150.445 -79.395 -150.115 ;
        RECT -79.725 -151.805 -79.395 -151.475 ;
        RECT -79.725 -153.165 -79.395 -152.835 ;
        RECT -79.725 -154.525 -79.395 -154.195 ;
        RECT -79.725 -155.885 -79.395 -155.555 ;
        RECT -79.725 -157.245 -79.395 -156.915 ;
        RECT -79.725 -158.605 -79.395 -158.275 ;
        RECT -79.725 -159.965 -79.395 -159.635 ;
        RECT -79.725 -161.325 -79.395 -160.995 ;
        RECT -79.725 -162.685 -79.395 -162.355 ;
        RECT -79.725 -164.045 -79.395 -163.715 ;
        RECT -79.725 -165.405 -79.395 -165.075 ;
        RECT -79.725 -166.765 -79.395 -166.435 ;
        RECT -79.725 -168.125 -79.395 -167.795 ;
        RECT -79.725 -169.485 -79.395 -169.155 ;
        RECT -79.725 -170.845 -79.395 -170.515 ;
        RECT -79.725 -172.205 -79.395 -171.875 ;
        RECT -79.725 -173.565 -79.395 -173.235 ;
        RECT -79.725 -174.925 -79.395 -174.595 ;
        RECT -79.725 -176.285 -79.395 -175.955 ;
        RECT -79.725 -177.645 -79.395 -177.315 ;
        RECT -79.725 -179.005 -79.395 -178.675 ;
        RECT -79.725 -180.365 -79.395 -180.035 ;
        RECT -79.725 -181.725 -79.395 -181.395 ;
        RECT -79.725 -183.085 -79.395 -182.755 ;
        RECT -79.725 -184.445 -79.395 -184.115 ;
        RECT -79.725 -185.805 -79.395 -185.475 ;
        RECT -79.725 -187.165 -79.395 -186.835 ;
        RECT -79.725 -188.525 -79.395 -188.195 ;
        RECT -79.725 -189.885 -79.395 -189.555 ;
        RECT -79.725 -191.245 -79.395 -190.915 ;
        RECT -79.725 -192.605 -79.395 -192.275 ;
        RECT -79.725 -193.965 -79.395 -193.635 ;
        RECT -79.725 -195.325 -79.395 -194.995 ;
        RECT -79.725 -196.685 -79.395 -196.355 ;
        RECT -79.725 -198.045 -79.395 -197.715 ;
        RECT -79.725 -199.405 -79.395 -199.075 ;
        RECT -79.725 -200.765 -79.395 -200.435 ;
        RECT -79.725 -202.125 -79.395 -201.795 ;
        RECT -79.725 -203.485 -79.395 -203.155 ;
        RECT -79.725 -204.845 -79.395 -204.515 ;
        RECT -79.725 -206.205 -79.395 -205.875 ;
        RECT -79.725 -207.565 -79.395 -207.235 ;
        RECT -79.725 -208.925 -79.395 -208.595 ;
        RECT -79.725 -210.285 -79.395 -209.955 ;
        RECT -79.725 -211.645 -79.395 -211.315 ;
        RECT -79.725 -213.005 -79.395 -212.675 ;
        RECT -79.725 -214.365 -79.395 -214.035 ;
        RECT -79.725 -215.725 -79.395 -215.395 ;
        RECT -79.725 -217.085 -79.395 -216.755 ;
        RECT -79.725 -218.445 -79.395 -218.115 ;
        RECT -79.725 -219.805 -79.395 -219.475 ;
        RECT -79.725 -221.165 -79.395 -220.835 ;
        RECT -79.725 -222.525 -79.395 -222.195 ;
        RECT -79.725 -223.885 -79.395 -223.555 ;
        RECT -79.725 -225.245 -79.395 -224.915 ;
        RECT -79.725 -226.605 -79.395 -226.275 ;
        RECT -79.725 -227.965 -79.395 -227.635 ;
        RECT -79.725 -229.325 -79.395 -228.995 ;
        RECT -79.725 -230.685 -79.395 -230.355 ;
        RECT -79.725 -232.045 -79.395 -231.715 ;
        RECT -79.725 -233.405 -79.395 -233.075 ;
        RECT -79.725 -234.765 -79.395 -234.435 ;
        RECT -79.725 -236.125 -79.395 -235.795 ;
        RECT -79.725 -237.485 -79.395 -237.155 ;
        RECT -79.725 -238.845 -79.395 -238.515 ;
        RECT -79.725 -241.09 -79.395 -239.96 ;
        RECT -79.72 -241.205 -79.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -78.365 244.04 -78.035 245.17 ;
        RECT -78.365 242.595 -78.035 242.925 ;
        RECT -78.365 241.235 -78.035 241.565 ;
        RECT -78.365 239.875 -78.035 240.205 ;
        RECT -78.365 238.515 -78.035 238.845 ;
        RECT -78.365 237.155 -78.035 237.485 ;
        RECT -78.365 235.795 -78.035 236.125 ;
        RECT -78.365 234.435 -78.035 234.765 ;
        RECT -78.365 233.075 -78.035 233.405 ;
        RECT -78.365 231.715 -78.035 232.045 ;
        RECT -78.365 230.355 -78.035 230.685 ;
        RECT -78.365 228.995 -78.035 229.325 ;
        RECT -78.365 227.635 -78.035 227.965 ;
        RECT -78.365 226.275 -78.035 226.605 ;
        RECT -78.365 224.915 -78.035 225.245 ;
        RECT -78.365 223.555 -78.035 223.885 ;
        RECT -78.365 222.195 -78.035 222.525 ;
        RECT -78.365 220.835 -78.035 221.165 ;
        RECT -78.365 219.475 -78.035 219.805 ;
        RECT -78.365 218.115 -78.035 218.445 ;
        RECT -78.365 216.755 -78.035 217.085 ;
        RECT -78.365 215.395 -78.035 215.725 ;
        RECT -78.365 214.035 -78.035 214.365 ;
        RECT -78.365 212.675 -78.035 213.005 ;
        RECT -78.365 211.315 -78.035 211.645 ;
        RECT -78.365 209.955 -78.035 210.285 ;
        RECT -78.365 208.595 -78.035 208.925 ;
        RECT -78.365 207.235 -78.035 207.565 ;
        RECT -78.365 205.875 -78.035 206.205 ;
        RECT -78.365 204.515 -78.035 204.845 ;
        RECT -78.365 203.155 -78.035 203.485 ;
        RECT -78.365 201.795 -78.035 202.125 ;
        RECT -78.365 200.435 -78.035 200.765 ;
        RECT -78.365 199.075 -78.035 199.405 ;
        RECT -78.365 197.715 -78.035 198.045 ;
        RECT -78.365 196.355 -78.035 196.685 ;
        RECT -78.365 194.995 -78.035 195.325 ;
        RECT -78.365 193.635 -78.035 193.965 ;
        RECT -78.365 192.275 -78.035 192.605 ;
        RECT -78.365 190.915 -78.035 191.245 ;
        RECT -78.365 189.555 -78.035 189.885 ;
        RECT -78.365 188.195 -78.035 188.525 ;
        RECT -78.365 186.835 -78.035 187.165 ;
        RECT -78.365 185.475 -78.035 185.805 ;
        RECT -78.365 184.115 -78.035 184.445 ;
        RECT -78.365 182.755 -78.035 183.085 ;
        RECT -78.365 181.395 -78.035 181.725 ;
        RECT -78.365 180.035 -78.035 180.365 ;
        RECT -78.365 178.675 -78.035 179.005 ;
        RECT -78.365 177.315 -78.035 177.645 ;
        RECT -78.365 175.955 -78.035 176.285 ;
        RECT -78.365 174.595 -78.035 174.925 ;
        RECT -78.365 173.235 -78.035 173.565 ;
        RECT -78.365 171.875 -78.035 172.205 ;
        RECT -78.365 170.515 -78.035 170.845 ;
        RECT -78.365 169.155 -78.035 169.485 ;
        RECT -78.365 167.795 -78.035 168.125 ;
        RECT -78.365 166.435 -78.035 166.765 ;
        RECT -78.365 165.075 -78.035 165.405 ;
        RECT -78.365 163.715 -78.035 164.045 ;
        RECT -78.365 162.355 -78.035 162.685 ;
        RECT -78.365 160.995 -78.035 161.325 ;
        RECT -78.365 159.635 -78.035 159.965 ;
        RECT -78.365 158.275 -78.035 158.605 ;
        RECT -78.365 156.915 -78.035 157.245 ;
        RECT -78.365 155.555 -78.035 155.885 ;
        RECT -78.365 154.195 -78.035 154.525 ;
        RECT -78.365 152.835 -78.035 153.165 ;
        RECT -78.365 151.475 -78.035 151.805 ;
        RECT -78.365 150.115 -78.035 150.445 ;
        RECT -78.365 148.755 -78.035 149.085 ;
        RECT -78.365 147.395 -78.035 147.725 ;
        RECT -78.365 146.035 -78.035 146.365 ;
        RECT -78.365 144.675 -78.035 145.005 ;
        RECT -78.365 143.315 -78.035 143.645 ;
        RECT -78.365 141.955 -78.035 142.285 ;
        RECT -78.365 140.595 -78.035 140.925 ;
        RECT -78.365 139.235 -78.035 139.565 ;
        RECT -78.365 137.875 -78.035 138.205 ;
        RECT -78.365 136.515 -78.035 136.845 ;
        RECT -78.365 135.155 -78.035 135.485 ;
        RECT -78.365 133.795 -78.035 134.125 ;
        RECT -78.365 132.435 -78.035 132.765 ;
        RECT -78.365 131.075 -78.035 131.405 ;
        RECT -78.365 129.715 -78.035 130.045 ;
        RECT -78.365 128.355 -78.035 128.685 ;
        RECT -78.365 126.995 -78.035 127.325 ;
        RECT -78.365 125.635 -78.035 125.965 ;
        RECT -78.365 124.275 -78.035 124.605 ;
        RECT -78.365 122.915 -78.035 123.245 ;
        RECT -78.365 121.555 -78.035 121.885 ;
        RECT -78.365 120.195 -78.035 120.525 ;
        RECT -78.365 118.835 -78.035 119.165 ;
        RECT -78.365 117.475 -78.035 117.805 ;
        RECT -78.365 116.115 -78.035 116.445 ;
        RECT -78.365 114.755 -78.035 115.085 ;
        RECT -78.365 113.395 -78.035 113.725 ;
        RECT -78.365 112.035 -78.035 112.365 ;
        RECT -78.365 110.675 -78.035 111.005 ;
        RECT -78.365 109.315 -78.035 109.645 ;
        RECT -78.365 107.955 -78.035 108.285 ;
        RECT -78.365 106.595 -78.035 106.925 ;
        RECT -78.365 105.235 -78.035 105.565 ;
        RECT -78.365 103.875 -78.035 104.205 ;
        RECT -78.365 102.515 -78.035 102.845 ;
        RECT -78.365 101.155 -78.035 101.485 ;
        RECT -78.365 99.795 -78.035 100.125 ;
        RECT -78.365 98.435 -78.035 98.765 ;
        RECT -78.365 97.075 -78.035 97.405 ;
        RECT -78.365 95.715 -78.035 96.045 ;
        RECT -78.365 94.355 -78.035 94.685 ;
        RECT -78.365 92.995 -78.035 93.325 ;
        RECT -78.365 91.635 -78.035 91.965 ;
        RECT -78.365 90.275 -78.035 90.605 ;
        RECT -78.365 88.915 -78.035 89.245 ;
        RECT -78.365 87.555 -78.035 87.885 ;
        RECT -78.365 86.195 -78.035 86.525 ;
        RECT -78.365 84.835 -78.035 85.165 ;
        RECT -78.365 83.475 -78.035 83.805 ;
        RECT -78.365 82.115 -78.035 82.445 ;
        RECT -78.365 80.755 -78.035 81.085 ;
        RECT -78.365 79.395 -78.035 79.725 ;
        RECT -78.365 78.035 -78.035 78.365 ;
        RECT -78.365 76.675 -78.035 77.005 ;
        RECT -78.365 75.315 -78.035 75.645 ;
        RECT -78.365 73.955 -78.035 74.285 ;
        RECT -78.365 72.595 -78.035 72.925 ;
        RECT -78.365 71.235 -78.035 71.565 ;
        RECT -78.365 69.875 -78.035 70.205 ;
        RECT -78.365 68.515 -78.035 68.845 ;
        RECT -78.365 67.155 -78.035 67.485 ;
        RECT -78.365 65.795 -78.035 66.125 ;
        RECT -78.365 64.435 -78.035 64.765 ;
        RECT -78.365 63.075 -78.035 63.405 ;
        RECT -78.365 61.715 -78.035 62.045 ;
        RECT -78.365 60.355 -78.035 60.685 ;
        RECT -78.365 58.995 -78.035 59.325 ;
        RECT -78.365 57.635 -78.035 57.965 ;
        RECT -78.365 56.275 -78.035 56.605 ;
        RECT -78.365 54.915 -78.035 55.245 ;
        RECT -78.365 53.555 -78.035 53.885 ;
        RECT -78.365 52.195 -78.035 52.525 ;
        RECT -78.365 50.835 -78.035 51.165 ;
        RECT -78.365 49.475 -78.035 49.805 ;
        RECT -78.365 48.115 -78.035 48.445 ;
        RECT -78.365 46.755 -78.035 47.085 ;
        RECT -78.365 45.395 -78.035 45.725 ;
        RECT -78.365 44.035 -78.035 44.365 ;
        RECT -78.365 42.675 -78.035 43.005 ;
        RECT -78.365 41.315 -78.035 41.645 ;
        RECT -78.365 39.955 -78.035 40.285 ;
        RECT -78.365 38.595 -78.035 38.925 ;
        RECT -78.365 37.235 -78.035 37.565 ;
        RECT -78.365 35.875 -78.035 36.205 ;
        RECT -78.365 34.515 -78.035 34.845 ;
        RECT -78.365 33.155 -78.035 33.485 ;
        RECT -78.365 31.795 -78.035 32.125 ;
        RECT -78.365 30.435 -78.035 30.765 ;
        RECT -78.365 29.075 -78.035 29.405 ;
        RECT -78.365 27.715 -78.035 28.045 ;
        RECT -78.365 26.355 -78.035 26.685 ;
        RECT -78.365 24.995 -78.035 25.325 ;
        RECT -78.365 23.635 -78.035 23.965 ;
        RECT -78.365 22.275 -78.035 22.605 ;
        RECT -78.365 20.915 -78.035 21.245 ;
        RECT -78.365 19.555 -78.035 19.885 ;
        RECT -78.365 18.195 -78.035 18.525 ;
        RECT -78.365 16.835 -78.035 17.165 ;
        RECT -78.365 15.475 -78.035 15.805 ;
        RECT -78.365 14.115 -78.035 14.445 ;
        RECT -78.365 12.755 -78.035 13.085 ;
        RECT -78.365 11.395 -78.035 11.725 ;
        RECT -78.365 10.035 -78.035 10.365 ;
        RECT -78.365 8.675 -78.035 9.005 ;
        RECT -78.365 7.315 -78.035 7.645 ;
        RECT -78.365 5.955 -78.035 6.285 ;
        RECT -78.365 4.595 -78.035 4.925 ;
        RECT -78.365 3.235 -78.035 3.565 ;
        RECT -78.365 1.875 -78.035 2.205 ;
        RECT -78.365 0.515 -78.035 0.845 ;
        RECT -78.365 -0.845 -78.035 -0.515 ;
        RECT -78.365 -2.205 -78.035 -1.875 ;
        RECT -78.365 -3.565 -78.035 -3.235 ;
        RECT -78.365 -4.925 -78.035 -4.595 ;
        RECT -78.365 -6.285 -78.035 -5.955 ;
        RECT -78.365 -7.645 -78.035 -7.315 ;
        RECT -78.365 -9.005 -78.035 -8.675 ;
        RECT -78.365 -10.365 -78.035 -10.035 ;
        RECT -78.365 -11.725 -78.035 -11.395 ;
        RECT -78.365 -13.085 -78.035 -12.755 ;
        RECT -78.365 -14.445 -78.035 -14.115 ;
        RECT -78.365 -15.805 -78.035 -15.475 ;
        RECT -78.365 -17.165 -78.035 -16.835 ;
        RECT -78.365 -18.525 -78.035 -18.195 ;
        RECT -78.365 -19.885 -78.035 -19.555 ;
        RECT -78.365 -21.245 -78.035 -20.915 ;
        RECT -78.365 -22.605 -78.035 -22.275 ;
        RECT -78.365 -23.965 -78.035 -23.635 ;
        RECT -78.365 -25.325 -78.035 -24.995 ;
        RECT -78.365 -26.685 -78.035 -26.355 ;
        RECT -78.365 -28.045 -78.035 -27.715 ;
        RECT -78.365 -29.405 -78.035 -29.075 ;
        RECT -78.365 -30.765 -78.035 -30.435 ;
        RECT -78.365 -32.125 -78.035 -31.795 ;
        RECT -78.365 -33.485 -78.035 -33.155 ;
        RECT -78.365 -34.845 -78.035 -34.515 ;
        RECT -78.365 -36.205 -78.035 -35.875 ;
        RECT -78.365 -37.565 -78.035 -37.235 ;
        RECT -78.365 -38.925 -78.035 -38.595 ;
        RECT -78.365 -40.285 -78.035 -39.955 ;
        RECT -78.365 -41.645 -78.035 -41.315 ;
        RECT -78.365 -43.005 -78.035 -42.675 ;
        RECT -78.365 -44.365 -78.035 -44.035 ;
        RECT -78.365 -45.725 -78.035 -45.395 ;
        RECT -78.365 -47.085 -78.035 -46.755 ;
        RECT -78.365 -48.445 -78.035 -48.115 ;
        RECT -78.365 -49.805 -78.035 -49.475 ;
        RECT -78.365 -51.165 -78.035 -50.835 ;
        RECT -78.365 -52.525 -78.035 -52.195 ;
        RECT -78.365 -53.885 -78.035 -53.555 ;
        RECT -78.365 -55.245 -78.035 -54.915 ;
        RECT -78.365 -56.605 -78.035 -56.275 ;
        RECT -78.365 -57.965 -78.035 -57.635 ;
        RECT -78.365 -59.325 -78.035 -58.995 ;
        RECT -78.365 -60.685 -78.035 -60.355 ;
        RECT -78.365 -62.045 -78.035 -61.715 ;
        RECT -78.365 -63.405 -78.035 -63.075 ;
        RECT -78.365 -64.765 -78.035 -64.435 ;
        RECT -78.365 -66.125 -78.035 -65.795 ;
        RECT -78.365 -67.485 -78.035 -67.155 ;
        RECT -78.365 -68.845 -78.035 -68.515 ;
        RECT -78.365 -70.205 -78.035 -69.875 ;
        RECT -78.365 -71.565 -78.035 -71.235 ;
        RECT -78.365 -72.925 -78.035 -72.595 ;
        RECT -78.365 -74.285 -78.035 -73.955 ;
        RECT -78.365 -75.645 -78.035 -75.315 ;
        RECT -78.365 -77.005 -78.035 -76.675 ;
        RECT -78.365 -78.365 -78.035 -78.035 ;
        RECT -78.365 -79.725 -78.035 -79.395 ;
        RECT -78.365 -81.085 -78.035 -80.755 ;
        RECT -78.365 -82.445 -78.035 -82.115 ;
        RECT -78.365 -83.805 -78.035 -83.475 ;
        RECT -78.365 -85.165 -78.035 -84.835 ;
        RECT -78.365 -86.525 -78.035 -86.195 ;
        RECT -78.365 -87.885 -78.035 -87.555 ;
        RECT -78.365 -89.245 -78.035 -88.915 ;
        RECT -78.365 -90.605 -78.035 -90.275 ;
        RECT -78.365 -91.965 -78.035 -91.635 ;
        RECT -78.365 -93.325 -78.035 -92.995 ;
        RECT -78.365 -94.685 -78.035 -94.355 ;
        RECT -78.365 -96.045 -78.035 -95.715 ;
        RECT -78.365 -97.405 -78.035 -97.075 ;
        RECT -78.365 -98.765 -78.035 -98.435 ;
        RECT -78.365 -100.125 -78.035 -99.795 ;
        RECT -78.365 -101.485 -78.035 -101.155 ;
        RECT -78.365 -102.845 -78.035 -102.515 ;
        RECT -78.365 -104.205 -78.035 -103.875 ;
        RECT -78.365 -105.565 -78.035 -105.235 ;
        RECT -78.365 -106.925 -78.035 -106.595 ;
        RECT -78.365 -108.285 -78.035 -107.955 ;
        RECT -78.365 -109.645 -78.035 -109.315 ;
        RECT -78.365 -111.005 -78.035 -110.675 ;
        RECT -78.365 -112.365 -78.035 -112.035 ;
        RECT -78.365 -113.725 -78.035 -113.395 ;
        RECT -78.365 -115.085 -78.035 -114.755 ;
        RECT -78.365 -116.445 -78.035 -116.115 ;
        RECT -78.365 -117.805 -78.035 -117.475 ;
        RECT -78.365 -119.165 -78.035 -118.835 ;
        RECT -78.365 -120.525 -78.035 -120.195 ;
        RECT -78.365 -121.885 -78.035 -121.555 ;
        RECT -78.365 -123.245 -78.035 -122.915 ;
        RECT -78.365 -124.605 -78.035 -124.275 ;
        RECT -78.365 -125.965 -78.035 -125.635 ;
        RECT -78.365 -127.325 -78.035 -126.995 ;
        RECT -78.365 -128.685 -78.035 -128.355 ;
        RECT -78.365 -130.045 -78.035 -129.715 ;
        RECT -78.365 -131.405 -78.035 -131.075 ;
        RECT -78.365 -132.765 -78.035 -132.435 ;
        RECT -78.365 -134.125 -78.035 -133.795 ;
        RECT -78.365 -135.485 -78.035 -135.155 ;
        RECT -78.365 -136.845 -78.035 -136.515 ;
        RECT -78.365 -138.205 -78.035 -137.875 ;
        RECT -78.365 -139.565 -78.035 -139.235 ;
        RECT -78.365 -140.925 -78.035 -140.595 ;
        RECT -78.365 -142.285 -78.035 -141.955 ;
        RECT -78.365 -143.645 -78.035 -143.315 ;
        RECT -78.365 -145.005 -78.035 -144.675 ;
        RECT -78.365 -146.365 -78.035 -146.035 ;
        RECT -78.365 -147.725 -78.035 -147.395 ;
        RECT -78.365 -149.085 -78.035 -148.755 ;
        RECT -78.365 -150.445 -78.035 -150.115 ;
        RECT -78.365 -151.805 -78.035 -151.475 ;
        RECT -78.365 -153.165 -78.035 -152.835 ;
        RECT -78.365 -154.525 -78.035 -154.195 ;
        RECT -78.365 -155.885 -78.035 -155.555 ;
        RECT -78.365 -157.245 -78.035 -156.915 ;
        RECT -78.365 -158.605 -78.035 -158.275 ;
        RECT -78.365 -159.965 -78.035 -159.635 ;
        RECT -78.365 -161.325 -78.035 -160.995 ;
        RECT -78.365 -162.685 -78.035 -162.355 ;
        RECT -78.365 -164.045 -78.035 -163.715 ;
        RECT -78.365 -165.405 -78.035 -165.075 ;
        RECT -78.365 -166.765 -78.035 -166.435 ;
        RECT -78.365 -168.125 -78.035 -167.795 ;
        RECT -78.365 -169.485 -78.035 -169.155 ;
        RECT -78.365 -170.845 -78.035 -170.515 ;
        RECT -78.365 -172.205 -78.035 -171.875 ;
        RECT -78.365 -173.565 -78.035 -173.235 ;
        RECT -78.365 -174.925 -78.035 -174.595 ;
        RECT -78.365 -176.285 -78.035 -175.955 ;
        RECT -78.365 -177.645 -78.035 -177.315 ;
        RECT -78.365 -179.005 -78.035 -178.675 ;
        RECT -78.365 -180.365 -78.035 -180.035 ;
        RECT -78.365 -181.725 -78.035 -181.395 ;
        RECT -78.365 -183.085 -78.035 -182.755 ;
        RECT -78.365 -184.445 -78.035 -184.115 ;
        RECT -78.365 -185.805 -78.035 -185.475 ;
        RECT -78.365 -187.165 -78.035 -186.835 ;
        RECT -78.365 -188.525 -78.035 -188.195 ;
        RECT -78.365 -189.885 -78.035 -189.555 ;
        RECT -78.365 -191.245 -78.035 -190.915 ;
        RECT -78.365 -192.605 -78.035 -192.275 ;
        RECT -78.365 -193.965 -78.035 -193.635 ;
        RECT -78.365 -195.325 -78.035 -194.995 ;
        RECT -78.365 -196.685 -78.035 -196.355 ;
        RECT -78.365 -198.045 -78.035 -197.715 ;
        RECT -78.365 -199.405 -78.035 -199.075 ;
        RECT -78.365 -200.765 -78.035 -200.435 ;
        RECT -78.365 -202.125 -78.035 -201.795 ;
        RECT -78.365 -203.485 -78.035 -203.155 ;
        RECT -78.365 -204.845 -78.035 -204.515 ;
        RECT -78.365 -206.205 -78.035 -205.875 ;
        RECT -78.365 -207.565 -78.035 -207.235 ;
        RECT -78.365 -208.925 -78.035 -208.595 ;
        RECT -78.365 -210.285 -78.035 -209.955 ;
        RECT -78.365 -211.645 -78.035 -211.315 ;
        RECT -78.365 -213.005 -78.035 -212.675 ;
        RECT -78.365 -214.365 -78.035 -214.035 ;
        RECT -78.365 -215.725 -78.035 -215.395 ;
        RECT -78.365 -217.085 -78.035 -216.755 ;
        RECT -78.365 -218.445 -78.035 -218.115 ;
        RECT -78.365 -219.805 -78.035 -219.475 ;
        RECT -78.365 -221.165 -78.035 -220.835 ;
        RECT -78.365 -222.525 -78.035 -222.195 ;
        RECT -78.365 -223.885 -78.035 -223.555 ;
        RECT -78.365 -225.245 -78.035 -224.915 ;
        RECT -78.365 -227.965 -78.035 -227.635 ;
        RECT -78.365 -229.325 -78.035 -228.995 ;
        RECT -78.365 -230.685 -78.035 -230.355 ;
        RECT -78.365 -232.045 -78.035 -231.715 ;
        RECT -78.365 -234.765 -78.035 -234.435 ;
        RECT -78.365 -236.125 -78.035 -235.795 ;
        RECT -78.365 -237.485 -78.035 -237.155 ;
        RECT -78.365 -238.845 -78.035 -238.515 ;
        RECT -78.365 -241.09 -78.035 -239.96 ;
        RECT -78.36 -241.205 -78.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -77.005 -77.005 -76.675 -76.675 ;
        RECT -77.005 -78.365 -76.675 -78.035 ;
        RECT -77.005 -79.725 -76.675 -79.395 ;
        RECT -77.005 -81.085 -76.675 -80.755 ;
        RECT -77.005 -82.445 -76.675 -82.115 ;
        RECT -77.005 -83.805 -76.675 -83.475 ;
        RECT -77.005 -85.165 -76.675 -84.835 ;
        RECT -77.005 -86.525 -76.675 -86.195 ;
        RECT -77.005 -87.885 -76.675 -87.555 ;
        RECT -77.005 -89.245 -76.675 -88.915 ;
        RECT -77.005 -90.605 -76.675 -90.275 ;
        RECT -77.005 -91.965 -76.675 -91.635 ;
        RECT -77.005 -93.325 -76.675 -92.995 ;
        RECT -77.005 -94.685 -76.675 -94.355 ;
        RECT -77.005 -96.045 -76.675 -95.715 ;
        RECT -77.005 -97.405 -76.675 -97.075 ;
        RECT -77.005 -98.765 -76.675 -98.435 ;
        RECT -77.005 -100.125 -76.675 -99.795 ;
        RECT -77.005 -101.485 -76.675 -101.155 ;
        RECT -77.005 -102.845 -76.675 -102.515 ;
        RECT -77.005 -104.205 -76.675 -103.875 ;
        RECT -77.005 -105.565 -76.675 -105.235 ;
        RECT -77.005 -106.925 -76.675 -106.595 ;
        RECT -77.005 -108.285 -76.675 -107.955 ;
        RECT -77.005 -109.645 -76.675 -109.315 ;
        RECT -77.005 -111.005 -76.675 -110.675 ;
        RECT -77.005 -112.365 -76.675 -112.035 ;
        RECT -77.005 -113.725 -76.675 -113.395 ;
        RECT -77.005 -115.085 -76.675 -114.755 ;
        RECT -77.005 -116.445 -76.675 -116.115 ;
        RECT -77.005 -117.805 -76.675 -117.475 ;
        RECT -77.005 -119.165 -76.675 -118.835 ;
        RECT -77.005 -120.525 -76.675 -120.195 ;
        RECT -77.005 -121.885 -76.675 -121.555 ;
        RECT -77.005 -123.245 -76.675 -122.915 ;
        RECT -77.005 -124.605 -76.675 -124.275 ;
        RECT -77.005 -125.965 -76.675 -125.635 ;
        RECT -77.005 -127.325 -76.675 -126.995 ;
        RECT -77.005 -128.685 -76.675 -128.355 ;
        RECT -77.005 -130.045 -76.675 -129.715 ;
        RECT -77.005 -131.405 -76.675 -131.075 ;
        RECT -77.005 -132.765 -76.675 -132.435 ;
        RECT -77.005 -134.125 -76.675 -133.795 ;
        RECT -77.005 -135.485 -76.675 -135.155 ;
        RECT -77.005 -136.845 -76.675 -136.515 ;
        RECT -77.005 -138.205 -76.675 -137.875 ;
        RECT -77.005 -139.565 -76.675 -139.235 ;
        RECT -77.005 -140.925 -76.675 -140.595 ;
        RECT -77.005 -142.285 -76.675 -141.955 ;
        RECT -77.005 -143.645 -76.675 -143.315 ;
        RECT -77.005 -145.005 -76.675 -144.675 ;
        RECT -77.005 -146.365 -76.675 -146.035 ;
        RECT -77.005 -147.725 -76.675 -147.395 ;
        RECT -77.005 -149.085 -76.675 -148.755 ;
        RECT -77.005 -150.445 -76.675 -150.115 ;
        RECT -77.005 -151.805 -76.675 -151.475 ;
        RECT -77.005 -153.165 -76.675 -152.835 ;
        RECT -77.005 -154.525 -76.675 -154.195 ;
        RECT -77.005 -155.885 -76.675 -155.555 ;
        RECT -77.005 -157.245 -76.675 -156.915 ;
        RECT -77.005 -158.605 -76.675 -158.275 ;
        RECT -77.005 -159.965 -76.675 -159.635 ;
        RECT -77.005 -161.325 -76.675 -160.995 ;
        RECT -77.005 -162.685 -76.675 -162.355 ;
        RECT -77.005 -164.045 -76.675 -163.715 ;
        RECT -77.005 -165.405 -76.675 -165.075 ;
        RECT -77.005 -166.765 -76.675 -166.435 ;
        RECT -77.005 -168.125 -76.675 -167.795 ;
        RECT -77.005 -169.485 -76.675 -169.155 ;
        RECT -77.005 -170.845 -76.675 -170.515 ;
        RECT -77.005 -172.205 -76.675 -171.875 ;
        RECT -77.005 -173.565 -76.675 -173.235 ;
        RECT -77.005 -174.925 -76.675 -174.595 ;
        RECT -77.005 -176.285 -76.675 -175.955 ;
        RECT -77.005 -177.645 -76.675 -177.315 ;
        RECT -77.005 -179.005 -76.675 -178.675 ;
        RECT -77.005 -180.365 -76.675 -180.035 ;
        RECT -77.005 -181.725 -76.675 -181.395 ;
        RECT -77.005 -183.085 -76.675 -182.755 ;
        RECT -77.005 -184.445 -76.675 -184.115 ;
        RECT -77.005 -185.805 -76.675 -185.475 ;
        RECT -77.005 -187.165 -76.675 -186.835 ;
        RECT -77.005 -188.525 -76.675 -188.195 ;
        RECT -77.005 -189.885 -76.675 -189.555 ;
        RECT -77.005 -191.245 -76.675 -190.915 ;
        RECT -77.005 -192.605 -76.675 -192.275 ;
        RECT -77.005 -193.965 -76.675 -193.635 ;
        RECT -77.005 -195.325 -76.675 -194.995 ;
        RECT -77.005 -196.685 -76.675 -196.355 ;
        RECT -77.005 -198.045 -76.675 -197.715 ;
        RECT -77.005 -199.405 -76.675 -199.075 ;
        RECT -77.005 -200.765 -76.675 -200.435 ;
        RECT -77.005 -202.125 -76.675 -201.795 ;
        RECT -77.005 -203.485 -76.675 -203.155 ;
        RECT -77.005 -204.845 -76.675 -204.515 ;
        RECT -77.005 -206.205 -76.675 -205.875 ;
        RECT -77.005 -207.565 -76.675 -207.235 ;
        RECT -77.005 -208.925 -76.675 -208.595 ;
        RECT -77.005 -210.285 -76.675 -209.955 ;
        RECT -77.005 -211.645 -76.675 -211.315 ;
        RECT -77.005 -213.005 -76.675 -212.675 ;
        RECT -77.005 -214.365 -76.675 -214.035 ;
        RECT -77.005 -215.725 -76.675 -215.395 ;
        RECT -77.005 -217.085 -76.675 -216.755 ;
        RECT -77.005 -218.445 -76.675 -218.115 ;
        RECT -77.005 -219.805 -76.675 -219.475 ;
        RECT -77.005 -221.165 -76.675 -220.835 ;
        RECT -77.005 -222.525 -76.675 -222.195 ;
        RECT -77.005 -223.885 -76.675 -223.555 ;
        RECT -77.005 -225.245 -76.675 -224.915 ;
        RECT -77.005 -227.965 -76.675 -227.635 ;
        RECT -77.005 -232.045 -76.675 -231.715 ;
        RECT -77.005 -233.225 -76.675 -232.895 ;
        RECT -77.005 -234.765 -76.675 -234.435 ;
        RECT -77.005 -236.125 -76.675 -235.795 ;
        RECT -77.005 -237.485 -76.675 -237.155 ;
        RECT -77.005 -238.845 -76.675 -238.515 ;
        RECT -77.005 -241.09 -76.675 -239.96 ;
        RECT -77 -241.205 -76.68 245.285 ;
        RECT -77.005 244.04 -76.675 245.17 ;
        RECT -77.005 242.595 -76.675 242.925 ;
        RECT -77.005 241.235 -76.675 241.565 ;
        RECT -77.005 239.875 -76.675 240.205 ;
        RECT -77.005 238.515 -76.675 238.845 ;
        RECT -77.005 237.155 -76.675 237.485 ;
        RECT -77.005 235.795 -76.675 236.125 ;
        RECT -77.005 234.435 -76.675 234.765 ;
        RECT -77.005 233.075 -76.675 233.405 ;
        RECT -77.005 231.715 -76.675 232.045 ;
        RECT -77.005 230.355 -76.675 230.685 ;
        RECT -77.005 228.995 -76.675 229.325 ;
        RECT -77.005 227.635 -76.675 227.965 ;
        RECT -77.005 226.275 -76.675 226.605 ;
        RECT -77.005 224.915 -76.675 225.245 ;
        RECT -77.005 223.555 -76.675 223.885 ;
        RECT -77.005 222.195 -76.675 222.525 ;
        RECT -77.005 220.835 -76.675 221.165 ;
        RECT -77.005 219.475 -76.675 219.805 ;
        RECT -77.005 218.115 -76.675 218.445 ;
        RECT -77.005 216.755 -76.675 217.085 ;
        RECT -77.005 215.395 -76.675 215.725 ;
        RECT -77.005 214.035 -76.675 214.365 ;
        RECT -77.005 212.675 -76.675 213.005 ;
        RECT -77.005 211.315 -76.675 211.645 ;
        RECT -77.005 209.955 -76.675 210.285 ;
        RECT -77.005 208.595 -76.675 208.925 ;
        RECT -77.005 207.235 -76.675 207.565 ;
        RECT -77.005 205.875 -76.675 206.205 ;
        RECT -77.005 204.515 -76.675 204.845 ;
        RECT -77.005 203.155 -76.675 203.485 ;
        RECT -77.005 201.795 -76.675 202.125 ;
        RECT -77.005 200.435 -76.675 200.765 ;
        RECT -77.005 199.075 -76.675 199.405 ;
        RECT -77.005 197.715 -76.675 198.045 ;
        RECT -77.005 196.355 -76.675 196.685 ;
        RECT -77.005 194.995 -76.675 195.325 ;
        RECT -77.005 193.635 -76.675 193.965 ;
        RECT -77.005 192.275 -76.675 192.605 ;
        RECT -77.005 190.915 -76.675 191.245 ;
        RECT -77.005 189.555 -76.675 189.885 ;
        RECT -77.005 188.195 -76.675 188.525 ;
        RECT -77.005 186.835 -76.675 187.165 ;
        RECT -77.005 185.475 -76.675 185.805 ;
        RECT -77.005 184.115 -76.675 184.445 ;
        RECT -77.005 182.755 -76.675 183.085 ;
        RECT -77.005 181.395 -76.675 181.725 ;
        RECT -77.005 180.035 -76.675 180.365 ;
        RECT -77.005 178.675 -76.675 179.005 ;
        RECT -77.005 177.315 -76.675 177.645 ;
        RECT -77.005 175.955 -76.675 176.285 ;
        RECT -77.005 174.595 -76.675 174.925 ;
        RECT -77.005 173.235 -76.675 173.565 ;
        RECT -77.005 171.875 -76.675 172.205 ;
        RECT -77.005 170.515 -76.675 170.845 ;
        RECT -77.005 169.155 -76.675 169.485 ;
        RECT -77.005 167.795 -76.675 168.125 ;
        RECT -77.005 166.435 -76.675 166.765 ;
        RECT -77.005 165.075 -76.675 165.405 ;
        RECT -77.005 163.715 -76.675 164.045 ;
        RECT -77.005 162.355 -76.675 162.685 ;
        RECT -77.005 160.995 -76.675 161.325 ;
        RECT -77.005 159.635 -76.675 159.965 ;
        RECT -77.005 158.275 -76.675 158.605 ;
        RECT -77.005 156.915 -76.675 157.245 ;
        RECT -77.005 155.555 -76.675 155.885 ;
        RECT -77.005 154.195 -76.675 154.525 ;
        RECT -77.005 152.835 -76.675 153.165 ;
        RECT -77.005 151.475 -76.675 151.805 ;
        RECT -77.005 150.115 -76.675 150.445 ;
        RECT -77.005 148.755 -76.675 149.085 ;
        RECT -77.005 147.395 -76.675 147.725 ;
        RECT -77.005 146.035 -76.675 146.365 ;
        RECT -77.005 144.675 -76.675 145.005 ;
        RECT -77.005 143.315 -76.675 143.645 ;
        RECT -77.005 141.955 -76.675 142.285 ;
        RECT -77.005 140.595 -76.675 140.925 ;
        RECT -77.005 139.235 -76.675 139.565 ;
        RECT -77.005 137.875 -76.675 138.205 ;
        RECT -77.005 136.515 -76.675 136.845 ;
        RECT -77.005 135.155 -76.675 135.485 ;
        RECT -77.005 133.795 -76.675 134.125 ;
        RECT -77.005 132.435 -76.675 132.765 ;
        RECT -77.005 131.075 -76.675 131.405 ;
        RECT -77.005 129.715 -76.675 130.045 ;
        RECT -77.005 128.355 -76.675 128.685 ;
        RECT -77.005 126.995 -76.675 127.325 ;
        RECT -77.005 125.635 -76.675 125.965 ;
        RECT -77.005 124.275 -76.675 124.605 ;
        RECT -77.005 122.915 -76.675 123.245 ;
        RECT -77.005 121.555 -76.675 121.885 ;
        RECT -77.005 120.195 -76.675 120.525 ;
        RECT -77.005 118.835 -76.675 119.165 ;
        RECT -77.005 117.475 -76.675 117.805 ;
        RECT -77.005 116.115 -76.675 116.445 ;
        RECT -77.005 114.755 -76.675 115.085 ;
        RECT -77.005 113.395 -76.675 113.725 ;
        RECT -77.005 112.035 -76.675 112.365 ;
        RECT -77.005 110.675 -76.675 111.005 ;
        RECT -77.005 109.315 -76.675 109.645 ;
        RECT -77.005 107.955 -76.675 108.285 ;
        RECT -77.005 106.595 -76.675 106.925 ;
        RECT -77.005 105.235 -76.675 105.565 ;
        RECT -77.005 103.875 -76.675 104.205 ;
        RECT -77.005 102.515 -76.675 102.845 ;
        RECT -77.005 101.155 -76.675 101.485 ;
        RECT -77.005 99.795 -76.675 100.125 ;
        RECT -77.005 98.435 -76.675 98.765 ;
        RECT -77.005 97.075 -76.675 97.405 ;
        RECT -77.005 95.715 -76.675 96.045 ;
        RECT -77.005 94.355 -76.675 94.685 ;
        RECT -77.005 92.995 -76.675 93.325 ;
        RECT -77.005 91.635 -76.675 91.965 ;
        RECT -77.005 90.275 -76.675 90.605 ;
        RECT -77.005 88.915 -76.675 89.245 ;
        RECT -77.005 87.555 -76.675 87.885 ;
        RECT -77.005 86.195 -76.675 86.525 ;
        RECT -77.005 84.835 -76.675 85.165 ;
        RECT -77.005 83.475 -76.675 83.805 ;
        RECT -77.005 82.115 -76.675 82.445 ;
        RECT -77.005 80.755 -76.675 81.085 ;
        RECT -77.005 79.395 -76.675 79.725 ;
        RECT -77.005 78.035 -76.675 78.365 ;
        RECT -77.005 76.675 -76.675 77.005 ;
        RECT -77.005 75.315 -76.675 75.645 ;
        RECT -77.005 73.955 -76.675 74.285 ;
        RECT -77.005 72.595 -76.675 72.925 ;
        RECT -77.005 71.235 -76.675 71.565 ;
        RECT -77.005 69.875 -76.675 70.205 ;
        RECT -77.005 68.515 -76.675 68.845 ;
        RECT -77.005 67.155 -76.675 67.485 ;
        RECT -77.005 65.795 -76.675 66.125 ;
        RECT -77.005 64.435 -76.675 64.765 ;
        RECT -77.005 63.075 -76.675 63.405 ;
        RECT -77.005 61.715 -76.675 62.045 ;
        RECT -77.005 60.355 -76.675 60.685 ;
        RECT -77.005 58.995 -76.675 59.325 ;
        RECT -77.005 57.635 -76.675 57.965 ;
        RECT -77.005 56.275 -76.675 56.605 ;
        RECT -77.005 54.915 -76.675 55.245 ;
        RECT -77.005 53.555 -76.675 53.885 ;
        RECT -77.005 52.195 -76.675 52.525 ;
        RECT -77.005 50.835 -76.675 51.165 ;
        RECT -77.005 49.475 -76.675 49.805 ;
        RECT -77.005 48.115 -76.675 48.445 ;
        RECT -77.005 46.755 -76.675 47.085 ;
        RECT -77.005 45.395 -76.675 45.725 ;
        RECT -77.005 44.035 -76.675 44.365 ;
        RECT -77.005 42.675 -76.675 43.005 ;
        RECT -77.005 41.315 -76.675 41.645 ;
        RECT -77.005 39.955 -76.675 40.285 ;
        RECT -77.005 38.595 -76.675 38.925 ;
        RECT -77.005 37.235 -76.675 37.565 ;
        RECT -77.005 35.875 -76.675 36.205 ;
        RECT -77.005 34.515 -76.675 34.845 ;
        RECT -77.005 33.155 -76.675 33.485 ;
        RECT -77.005 31.795 -76.675 32.125 ;
        RECT -77.005 30.435 -76.675 30.765 ;
        RECT -77.005 29.075 -76.675 29.405 ;
        RECT -77.005 27.715 -76.675 28.045 ;
        RECT -77.005 26.355 -76.675 26.685 ;
        RECT -77.005 24.995 -76.675 25.325 ;
        RECT -77.005 23.635 -76.675 23.965 ;
        RECT -77.005 22.275 -76.675 22.605 ;
        RECT -77.005 20.915 -76.675 21.245 ;
        RECT -77.005 19.555 -76.675 19.885 ;
        RECT -77.005 18.195 -76.675 18.525 ;
        RECT -77.005 16.835 -76.675 17.165 ;
        RECT -77.005 15.475 -76.675 15.805 ;
        RECT -77.005 14.115 -76.675 14.445 ;
        RECT -77.005 12.755 -76.675 13.085 ;
        RECT -77.005 11.395 -76.675 11.725 ;
        RECT -77.005 10.035 -76.675 10.365 ;
        RECT -77.005 8.675 -76.675 9.005 ;
        RECT -77.005 7.315 -76.675 7.645 ;
        RECT -77.005 5.955 -76.675 6.285 ;
        RECT -77.005 4.595 -76.675 4.925 ;
        RECT -77.005 3.235 -76.675 3.565 ;
        RECT -77.005 1.875 -76.675 2.205 ;
        RECT -77.005 0.515 -76.675 0.845 ;
        RECT -77.005 -0.845 -76.675 -0.515 ;
        RECT -77.005 -2.205 -76.675 -1.875 ;
        RECT -77.005 -3.565 -76.675 -3.235 ;
        RECT -77.005 -4.925 -76.675 -4.595 ;
        RECT -77.005 -6.285 -76.675 -5.955 ;
        RECT -77.005 -7.645 -76.675 -7.315 ;
        RECT -77.005 -9.005 -76.675 -8.675 ;
        RECT -77.005 -10.365 -76.675 -10.035 ;
        RECT -77.005 -11.725 -76.675 -11.395 ;
        RECT -77.005 -13.085 -76.675 -12.755 ;
        RECT -77.005 -14.445 -76.675 -14.115 ;
        RECT -77.005 -15.805 -76.675 -15.475 ;
        RECT -77.005 -17.165 -76.675 -16.835 ;
        RECT -77.005 -18.525 -76.675 -18.195 ;
        RECT -77.005 -19.885 -76.675 -19.555 ;
        RECT -77.005 -21.245 -76.675 -20.915 ;
        RECT -77.005 -22.605 -76.675 -22.275 ;
        RECT -77.005 -23.965 -76.675 -23.635 ;
        RECT -77.005 -25.325 -76.675 -24.995 ;
        RECT -77.005 -26.685 -76.675 -26.355 ;
        RECT -77.005 -28.045 -76.675 -27.715 ;
        RECT -77.005 -29.405 -76.675 -29.075 ;
        RECT -77.005 -30.765 -76.675 -30.435 ;
        RECT -77.005 -32.125 -76.675 -31.795 ;
        RECT -77.005 -33.485 -76.675 -33.155 ;
        RECT -77.005 -34.845 -76.675 -34.515 ;
        RECT -77.005 -36.205 -76.675 -35.875 ;
        RECT -77.005 -37.565 -76.675 -37.235 ;
        RECT -77.005 -38.925 -76.675 -38.595 ;
        RECT -77.005 -40.285 -76.675 -39.955 ;
        RECT -77.005 -41.645 -76.675 -41.315 ;
        RECT -77.005 -43.005 -76.675 -42.675 ;
        RECT -77.005 -44.365 -76.675 -44.035 ;
        RECT -77.005 -45.725 -76.675 -45.395 ;
        RECT -77.005 -47.085 -76.675 -46.755 ;
        RECT -77.005 -48.445 -76.675 -48.115 ;
        RECT -77.005 -49.805 -76.675 -49.475 ;
        RECT -77.005 -51.165 -76.675 -50.835 ;
        RECT -77.005 -52.525 -76.675 -52.195 ;
        RECT -77.005 -53.885 -76.675 -53.555 ;
        RECT -77.005 -55.245 -76.675 -54.915 ;
        RECT -77.005 -56.605 -76.675 -56.275 ;
        RECT -77.005 -57.965 -76.675 -57.635 ;
        RECT -77.005 -59.325 -76.675 -58.995 ;
        RECT -77.005 -60.685 -76.675 -60.355 ;
        RECT -77.005 -62.045 -76.675 -61.715 ;
        RECT -77.005 -63.405 -76.675 -63.075 ;
        RECT -77.005 -64.765 -76.675 -64.435 ;
        RECT -77.005 -66.125 -76.675 -65.795 ;
        RECT -77.005 -67.485 -76.675 -67.155 ;
        RECT -77.005 -68.845 -76.675 -68.515 ;
        RECT -77.005 -70.205 -76.675 -69.875 ;
        RECT -77.005 -71.565 -76.675 -71.235 ;
        RECT -77.005 -72.925 -76.675 -72.595 ;
        RECT -77.005 -74.285 -76.675 -73.955 ;
        RECT -77.005 -75.645 -76.675 -75.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -83.805 244.04 -83.475 245.17 ;
        RECT -83.805 242.595 -83.475 242.925 ;
        RECT -83.805 241.235 -83.475 241.565 ;
        RECT -83.805 239.875 -83.475 240.205 ;
        RECT -83.805 238.515 -83.475 238.845 ;
        RECT -83.805 237.155 -83.475 237.485 ;
        RECT -83.805 235.795 -83.475 236.125 ;
        RECT -83.805 234.435 -83.475 234.765 ;
        RECT -83.805 233.075 -83.475 233.405 ;
        RECT -83.805 231.715 -83.475 232.045 ;
        RECT -83.805 230.355 -83.475 230.685 ;
        RECT -83.805 228.995 -83.475 229.325 ;
        RECT -83.805 227.635 -83.475 227.965 ;
        RECT -83.805 226.275 -83.475 226.605 ;
        RECT -83.805 224.915 -83.475 225.245 ;
        RECT -83.805 223.555 -83.475 223.885 ;
        RECT -83.805 222.195 -83.475 222.525 ;
        RECT -83.805 220.835 -83.475 221.165 ;
        RECT -83.805 219.475 -83.475 219.805 ;
        RECT -83.805 218.115 -83.475 218.445 ;
        RECT -83.805 216.755 -83.475 217.085 ;
        RECT -83.805 215.395 -83.475 215.725 ;
        RECT -83.805 214.035 -83.475 214.365 ;
        RECT -83.805 212.675 -83.475 213.005 ;
        RECT -83.805 211.315 -83.475 211.645 ;
        RECT -83.805 209.955 -83.475 210.285 ;
        RECT -83.805 208.595 -83.475 208.925 ;
        RECT -83.805 207.235 -83.475 207.565 ;
        RECT -83.805 205.875 -83.475 206.205 ;
        RECT -83.805 204.515 -83.475 204.845 ;
        RECT -83.805 203.155 -83.475 203.485 ;
        RECT -83.805 201.795 -83.475 202.125 ;
        RECT -83.805 200.435 -83.475 200.765 ;
        RECT -83.805 199.075 -83.475 199.405 ;
        RECT -83.805 197.715 -83.475 198.045 ;
        RECT -83.805 196.355 -83.475 196.685 ;
        RECT -83.805 194.995 -83.475 195.325 ;
        RECT -83.805 193.635 -83.475 193.965 ;
        RECT -83.805 192.275 -83.475 192.605 ;
        RECT -83.805 190.915 -83.475 191.245 ;
        RECT -83.805 189.555 -83.475 189.885 ;
        RECT -83.805 188.195 -83.475 188.525 ;
        RECT -83.805 186.835 -83.475 187.165 ;
        RECT -83.805 185.475 -83.475 185.805 ;
        RECT -83.805 184.115 -83.475 184.445 ;
        RECT -83.805 182.755 -83.475 183.085 ;
        RECT -83.805 181.395 -83.475 181.725 ;
        RECT -83.805 180.035 -83.475 180.365 ;
        RECT -83.805 178.675 -83.475 179.005 ;
        RECT -83.805 177.315 -83.475 177.645 ;
        RECT -83.805 175.955 -83.475 176.285 ;
        RECT -83.805 174.595 -83.475 174.925 ;
        RECT -83.805 173.235 -83.475 173.565 ;
        RECT -83.805 171.875 -83.475 172.205 ;
        RECT -83.805 170.515 -83.475 170.845 ;
        RECT -83.805 169.155 -83.475 169.485 ;
        RECT -83.805 167.795 -83.475 168.125 ;
        RECT -83.805 166.435 -83.475 166.765 ;
        RECT -83.805 165.075 -83.475 165.405 ;
        RECT -83.805 163.715 -83.475 164.045 ;
        RECT -83.805 162.355 -83.475 162.685 ;
        RECT -83.805 160.995 -83.475 161.325 ;
        RECT -83.805 159.635 -83.475 159.965 ;
        RECT -83.805 158.275 -83.475 158.605 ;
        RECT -83.805 156.915 -83.475 157.245 ;
        RECT -83.805 155.555 -83.475 155.885 ;
        RECT -83.805 154.195 -83.475 154.525 ;
        RECT -83.805 152.835 -83.475 153.165 ;
        RECT -83.805 151.475 -83.475 151.805 ;
        RECT -83.805 150.115 -83.475 150.445 ;
        RECT -83.805 148.755 -83.475 149.085 ;
        RECT -83.805 147.395 -83.475 147.725 ;
        RECT -83.805 146.035 -83.475 146.365 ;
        RECT -83.805 144.675 -83.475 145.005 ;
        RECT -83.805 143.315 -83.475 143.645 ;
        RECT -83.805 141.955 -83.475 142.285 ;
        RECT -83.805 140.595 -83.475 140.925 ;
        RECT -83.805 139.235 -83.475 139.565 ;
        RECT -83.805 137.875 -83.475 138.205 ;
        RECT -83.805 136.515 -83.475 136.845 ;
        RECT -83.805 135.155 -83.475 135.485 ;
        RECT -83.805 133.795 -83.475 134.125 ;
        RECT -83.805 132.435 -83.475 132.765 ;
        RECT -83.805 131.075 -83.475 131.405 ;
        RECT -83.805 129.715 -83.475 130.045 ;
        RECT -83.805 128.355 -83.475 128.685 ;
        RECT -83.805 126.995 -83.475 127.325 ;
        RECT -83.805 125.635 -83.475 125.965 ;
        RECT -83.805 124.275 -83.475 124.605 ;
        RECT -83.805 122.915 -83.475 123.245 ;
        RECT -83.805 121.555 -83.475 121.885 ;
        RECT -83.805 120.195 -83.475 120.525 ;
        RECT -83.805 118.835 -83.475 119.165 ;
        RECT -83.805 117.475 -83.475 117.805 ;
        RECT -83.805 116.115 -83.475 116.445 ;
        RECT -83.805 114.755 -83.475 115.085 ;
        RECT -83.805 113.395 -83.475 113.725 ;
        RECT -83.805 112.035 -83.475 112.365 ;
        RECT -83.805 110.675 -83.475 111.005 ;
        RECT -83.805 109.315 -83.475 109.645 ;
        RECT -83.805 107.955 -83.475 108.285 ;
        RECT -83.805 106.595 -83.475 106.925 ;
        RECT -83.805 105.235 -83.475 105.565 ;
        RECT -83.805 103.875 -83.475 104.205 ;
        RECT -83.805 102.515 -83.475 102.845 ;
        RECT -83.805 101.155 -83.475 101.485 ;
        RECT -83.805 99.795 -83.475 100.125 ;
        RECT -83.805 98.435 -83.475 98.765 ;
        RECT -83.805 97.075 -83.475 97.405 ;
        RECT -83.805 95.715 -83.475 96.045 ;
        RECT -83.805 94.355 -83.475 94.685 ;
        RECT -83.805 92.995 -83.475 93.325 ;
        RECT -83.805 91.635 -83.475 91.965 ;
        RECT -83.805 90.275 -83.475 90.605 ;
        RECT -83.805 88.915 -83.475 89.245 ;
        RECT -83.805 87.555 -83.475 87.885 ;
        RECT -83.805 86.195 -83.475 86.525 ;
        RECT -83.805 84.835 -83.475 85.165 ;
        RECT -83.805 83.475 -83.475 83.805 ;
        RECT -83.805 82.115 -83.475 82.445 ;
        RECT -83.805 80.755 -83.475 81.085 ;
        RECT -83.805 79.395 -83.475 79.725 ;
        RECT -83.805 78.035 -83.475 78.365 ;
        RECT -83.805 76.675 -83.475 77.005 ;
        RECT -83.805 75.315 -83.475 75.645 ;
        RECT -83.805 73.955 -83.475 74.285 ;
        RECT -83.805 72.595 -83.475 72.925 ;
        RECT -83.805 71.235 -83.475 71.565 ;
        RECT -83.805 69.875 -83.475 70.205 ;
        RECT -83.805 68.515 -83.475 68.845 ;
        RECT -83.805 67.155 -83.475 67.485 ;
        RECT -83.805 65.795 -83.475 66.125 ;
        RECT -83.805 64.435 -83.475 64.765 ;
        RECT -83.805 63.075 -83.475 63.405 ;
        RECT -83.805 61.715 -83.475 62.045 ;
        RECT -83.805 60.355 -83.475 60.685 ;
        RECT -83.805 58.995 -83.475 59.325 ;
        RECT -83.805 57.635 -83.475 57.965 ;
        RECT -83.805 56.275 -83.475 56.605 ;
        RECT -83.805 54.915 -83.475 55.245 ;
        RECT -83.805 53.555 -83.475 53.885 ;
        RECT -83.805 52.195 -83.475 52.525 ;
        RECT -83.805 50.835 -83.475 51.165 ;
        RECT -83.805 49.475 -83.475 49.805 ;
        RECT -83.805 48.115 -83.475 48.445 ;
        RECT -83.805 46.755 -83.475 47.085 ;
        RECT -83.805 45.395 -83.475 45.725 ;
        RECT -83.805 44.035 -83.475 44.365 ;
        RECT -83.805 42.675 -83.475 43.005 ;
        RECT -83.805 41.315 -83.475 41.645 ;
        RECT -83.805 39.955 -83.475 40.285 ;
        RECT -83.805 38.595 -83.475 38.925 ;
        RECT -83.805 37.235 -83.475 37.565 ;
        RECT -83.805 35.875 -83.475 36.205 ;
        RECT -83.805 34.515 -83.475 34.845 ;
        RECT -83.805 33.155 -83.475 33.485 ;
        RECT -83.805 31.795 -83.475 32.125 ;
        RECT -83.805 30.435 -83.475 30.765 ;
        RECT -83.805 29.075 -83.475 29.405 ;
        RECT -83.805 27.715 -83.475 28.045 ;
        RECT -83.805 26.355 -83.475 26.685 ;
        RECT -83.805 24.995 -83.475 25.325 ;
        RECT -83.805 23.635 -83.475 23.965 ;
        RECT -83.805 22.275 -83.475 22.605 ;
        RECT -83.805 20.915 -83.475 21.245 ;
        RECT -83.805 19.555 -83.475 19.885 ;
        RECT -83.805 18.195 -83.475 18.525 ;
        RECT -83.805 16.835 -83.475 17.165 ;
        RECT -83.805 15.475 -83.475 15.805 ;
        RECT -83.805 14.115 -83.475 14.445 ;
        RECT -83.805 12.755 -83.475 13.085 ;
        RECT -83.805 11.395 -83.475 11.725 ;
        RECT -83.805 10.035 -83.475 10.365 ;
        RECT -83.805 8.675 -83.475 9.005 ;
        RECT -83.805 7.315 -83.475 7.645 ;
        RECT -83.805 5.955 -83.475 6.285 ;
        RECT -83.805 4.595 -83.475 4.925 ;
        RECT -83.805 3.235 -83.475 3.565 ;
        RECT -83.805 1.875 -83.475 2.205 ;
        RECT -83.805 0.515 -83.475 0.845 ;
        RECT -83.805 -0.845 -83.475 -0.515 ;
        RECT -83.805 -2.205 -83.475 -1.875 ;
        RECT -83.805 -3.565 -83.475 -3.235 ;
        RECT -83.805 -4.925 -83.475 -4.595 ;
        RECT -83.805 -6.285 -83.475 -5.955 ;
        RECT -83.805 -7.645 -83.475 -7.315 ;
        RECT -83.805 -9.005 -83.475 -8.675 ;
        RECT -83.805 -10.365 -83.475 -10.035 ;
        RECT -83.805 -11.725 -83.475 -11.395 ;
        RECT -83.805 -13.085 -83.475 -12.755 ;
        RECT -83.805 -14.445 -83.475 -14.115 ;
        RECT -83.805 -15.805 -83.475 -15.475 ;
        RECT -83.805 -17.165 -83.475 -16.835 ;
        RECT -83.805 -18.525 -83.475 -18.195 ;
        RECT -83.805 -19.885 -83.475 -19.555 ;
        RECT -83.805 -21.245 -83.475 -20.915 ;
        RECT -83.805 -22.605 -83.475 -22.275 ;
        RECT -83.805 -23.965 -83.475 -23.635 ;
        RECT -83.805 -25.325 -83.475 -24.995 ;
        RECT -83.805 -26.685 -83.475 -26.355 ;
        RECT -83.805 -28.045 -83.475 -27.715 ;
        RECT -83.805 -29.405 -83.475 -29.075 ;
        RECT -83.805 -30.765 -83.475 -30.435 ;
        RECT -83.805 -32.125 -83.475 -31.795 ;
        RECT -83.805 -33.485 -83.475 -33.155 ;
        RECT -83.805 -34.845 -83.475 -34.515 ;
        RECT -83.805 -36.205 -83.475 -35.875 ;
        RECT -83.805 -37.565 -83.475 -37.235 ;
        RECT -83.805 -38.925 -83.475 -38.595 ;
        RECT -83.805 -40.285 -83.475 -39.955 ;
        RECT -83.805 -41.645 -83.475 -41.315 ;
        RECT -83.805 -43.005 -83.475 -42.675 ;
        RECT -83.805 -44.365 -83.475 -44.035 ;
        RECT -83.805 -45.725 -83.475 -45.395 ;
        RECT -83.805 -47.085 -83.475 -46.755 ;
        RECT -83.805 -48.445 -83.475 -48.115 ;
        RECT -83.805 -49.805 -83.475 -49.475 ;
        RECT -83.805 -51.165 -83.475 -50.835 ;
        RECT -83.805 -52.525 -83.475 -52.195 ;
        RECT -83.805 -53.885 -83.475 -53.555 ;
        RECT -83.805 -55.245 -83.475 -54.915 ;
        RECT -83.805 -56.605 -83.475 -56.275 ;
        RECT -83.805 -57.965 -83.475 -57.635 ;
        RECT -83.805 -59.325 -83.475 -58.995 ;
        RECT -83.805 -60.685 -83.475 -60.355 ;
        RECT -83.805 -62.045 -83.475 -61.715 ;
        RECT -83.805 -63.405 -83.475 -63.075 ;
        RECT -83.805 -64.765 -83.475 -64.435 ;
        RECT -83.805 -66.125 -83.475 -65.795 ;
        RECT -83.805 -67.485 -83.475 -67.155 ;
        RECT -83.805 -68.845 -83.475 -68.515 ;
        RECT -83.805 -70.205 -83.475 -69.875 ;
        RECT -83.805 -71.565 -83.475 -71.235 ;
        RECT -83.805 -72.925 -83.475 -72.595 ;
        RECT -83.805 -74.285 -83.475 -73.955 ;
        RECT -83.805 -75.645 -83.475 -75.315 ;
        RECT -83.805 -77.005 -83.475 -76.675 ;
        RECT -83.805 -78.365 -83.475 -78.035 ;
        RECT -83.805 -79.725 -83.475 -79.395 ;
        RECT -83.805 -81.085 -83.475 -80.755 ;
        RECT -83.805 -82.445 -83.475 -82.115 ;
        RECT -83.805 -83.805 -83.475 -83.475 ;
        RECT -83.805 -85.165 -83.475 -84.835 ;
        RECT -83.805 -86.525 -83.475 -86.195 ;
        RECT -83.805 -87.885 -83.475 -87.555 ;
        RECT -83.805 -89.245 -83.475 -88.915 ;
        RECT -83.805 -90.605 -83.475 -90.275 ;
        RECT -83.805 -91.965 -83.475 -91.635 ;
        RECT -83.805 -93.325 -83.475 -92.995 ;
        RECT -83.805 -94.685 -83.475 -94.355 ;
        RECT -83.805 -96.045 -83.475 -95.715 ;
        RECT -83.805 -97.405 -83.475 -97.075 ;
        RECT -83.805 -98.765 -83.475 -98.435 ;
        RECT -83.805 -100.125 -83.475 -99.795 ;
        RECT -83.805 -101.485 -83.475 -101.155 ;
        RECT -83.805 -102.845 -83.475 -102.515 ;
        RECT -83.805 -104.205 -83.475 -103.875 ;
        RECT -83.805 -105.565 -83.475 -105.235 ;
        RECT -83.805 -106.925 -83.475 -106.595 ;
        RECT -83.805 -108.285 -83.475 -107.955 ;
        RECT -83.805 -109.645 -83.475 -109.315 ;
        RECT -83.805 -111.005 -83.475 -110.675 ;
        RECT -83.805 -112.365 -83.475 -112.035 ;
        RECT -83.805 -113.725 -83.475 -113.395 ;
        RECT -83.805 -115.085 -83.475 -114.755 ;
        RECT -83.805 -116.445 -83.475 -116.115 ;
        RECT -83.805 -117.805 -83.475 -117.475 ;
        RECT -83.805 -119.165 -83.475 -118.835 ;
        RECT -83.805 -120.525 -83.475 -120.195 ;
        RECT -83.805 -121.885 -83.475 -121.555 ;
        RECT -83.805 -123.245 -83.475 -122.915 ;
        RECT -83.805 -124.605 -83.475 -124.275 ;
        RECT -83.805 -125.965 -83.475 -125.635 ;
        RECT -83.805 -127.325 -83.475 -126.995 ;
        RECT -83.805 -128.685 -83.475 -128.355 ;
        RECT -83.805 -130.045 -83.475 -129.715 ;
        RECT -83.805 -131.405 -83.475 -131.075 ;
        RECT -83.805 -132.765 -83.475 -132.435 ;
        RECT -83.805 -134.125 -83.475 -133.795 ;
        RECT -83.805 -135.485 -83.475 -135.155 ;
        RECT -83.805 -136.845 -83.475 -136.515 ;
        RECT -83.805 -138.205 -83.475 -137.875 ;
        RECT -83.805 -139.565 -83.475 -139.235 ;
        RECT -83.805 -140.925 -83.475 -140.595 ;
        RECT -83.805 -142.285 -83.475 -141.955 ;
        RECT -83.805 -143.645 -83.475 -143.315 ;
        RECT -83.805 -145.005 -83.475 -144.675 ;
        RECT -83.805 -146.365 -83.475 -146.035 ;
        RECT -83.805 -147.725 -83.475 -147.395 ;
        RECT -83.805 -149.085 -83.475 -148.755 ;
        RECT -83.805 -150.445 -83.475 -150.115 ;
        RECT -83.805 -151.805 -83.475 -151.475 ;
        RECT -83.805 -153.165 -83.475 -152.835 ;
        RECT -83.805 -154.525 -83.475 -154.195 ;
        RECT -83.805 -155.885 -83.475 -155.555 ;
        RECT -83.805 -157.245 -83.475 -156.915 ;
        RECT -83.805 -158.605 -83.475 -158.275 ;
        RECT -83.805 -159.965 -83.475 -159.635 ;
        RECT -83.805 -161.325 -83.475 -160.995 ;
        RECT -83.805 -162.685 -83.475 -162.355 ;
        RECT -83.805 -164.045 -83.475 -163.715 ;
        RECT -83.805 -165.405 -83.475 -165.075 ;
        RECT -83.805 -166.765 -83.475 -166.435 ;
        RECT -83.805 -168.125 -83.475 -167.795 ;
        RECT -83.805 -169.485 -83.475 -169.155 ;
        RECT -83.805 -170.845 -83.475 -170.515 ;
        RECT -83.805 -172.205 -83.475 -171.875 ;
        RECT -83.805 -173.565 -83.475 -173.235 ;
        RECT -83.805 -174.925 -83.475 -174.595 ;
        RECT -83.805 -176.285 -83.475 -175.955 ;
        RECT -83.805 -177.645 -83.475 -177.315 ;
        RECT -83.805 -179.005 -83.475 -178.675 ;
        RECT -83.805 -180.365 -83.475 -180.035 ;
        RECT -83.805 -181.725 -83.475 -181.395 ;
        RECT -83.805 -183.085 -83.475 -182.755 ;
        RECT -83.805 -184.445 -83.475 -184.115 ;
        RECT -83.805 -185.805 -83.475 -185.475 ;
        RECT -83.805 -187.165 -83.475 -186.835 ;
        RECT -83.805 -188.525 -83.475 -188.195 ;
        RECT -83.805 -189.885 -83.475 -189.555 ;
        RECT -83.805 -191.245 -83.475 -190.915 ;
        RECT -83.805 -192.605 -83.475 -192.275 ;
        RECT -83.805 -193.965 -83.475 -193.635 ;
        RECT -83.805 -195.325 -83.475 -194.995 ;
        RECT -83.805 -196.685 -83.475 -196.355 ;
        RECT -83.805 -198.045 -83.475 -197.715 ;
        RECT -83.805 -199.405 -83.475 -199.075 ;
        RECT -83.805 -200.765 -83.475 -200.435 ;
        RECT -83.805 -202.125 -83.475 -201.795 ;
        RECT -83.805 -203.485 -83.475 -203.155 ;
        RECT -83.805 -204.845 -83.475 -204.515 ;
        RECT -83.805 -206.205 -83.475 -205.875 ;
        RECT -83.805 -207.565 -83.475 -207.235 ;
        RECT -83.805 -208.925 -83.475 -208.595 ;
        RECT -83.805 -210.285 -83.475 -209.955 ;
        RECT -83.805 -211.645 -83.475 -211.315 ;
        RECT -83.805 -213.005 -83.475 -212.675 ;
        RECT -83.805 -214.365 -83.475 -214.035 ;
        RECT -83.805 -215.725 -83.475 -215.395 ;
        RECT -83.805 -217.085 -83.475 -216.755 ;
        RECT -83.805 -218.445 -83.475 -218.115 ;
        RECT -83.805 -219.805 -83.475 -219.475 ;
        RECT -83.805 -221.165 -83.475 -220.835 ;
        RECT -83.805 -222.525 -83.475 -222.195 ;
        RECT -83.805 -223.885 -83.475 -223.555 ;
        RECT -83.805 -225.245 -83.475 -224.915 ;
        RECT -83.805 -226.605 -83.475 -226.275 ;
        RECT -83.805 -227.965 -83.475 -227.635 ;
        RECT -83.805 -229.325 -83.475 -228.995 ;
        RECT -83.805 -230.685 -83.475 -230.355 ;
        RECT -83.805 -232.045 -83.475 -231.715 ;
        RECT -83.805 -233.405 -83.475 -233.075 ;
        RECT -83.805 -234.765 -83.475 -234.435 ;
        RECT -83.805 -236.125 -83.475 -235.795 ;
        RECT -83.805 -237.485 -83.475 -237.155 ;
        RECT -83.805 -238.845 -83.475 -238.515 ;
        RECT -83.805 -241.09 -83.475 -239.96 ;
        RECT -83.8 -241.205 -83.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -82.445 244.04 -82.115 245.17 ;
        RECT -82.445 242.595 -82.115 242.925 ;
        RECT -82.445 241.235 -82.115 241.565 ;
        RECT -82.445 239.875 -82.115 240.205 ;
        RECT -82.445 238.515 -82.115 238.845 ;
        RECT -82.445 237.155 -82.115 237.485 ;
        RECT -82.445 235.795 -82.115 236.125 ;
        RECT -82.445 234.435 -82.115 234.765 ;
        RECT -82.445 233.075 -82.115 233.405 ;
        RECT -82.445 231.715 -82.115 232.045 ;
        RECT -82.445 230.355 -82.115 230.685 ;
        RECT -82.445 228.995 -82.115 229.325 ;
        RECT -82.445 227.635 -82.115 227.965 ;
        RECT -82.445 226.275 -82.115 226.605 ;
        RECT -82.445 224.915 -82.115 225.245 ;
        RECT -82.445 223.555 -82.115 223.885 ;
        RECT -82.445 222.195 -82.115 222.525 ;
        RECT -82.445 220.835 -82.115 221.165 ;
        RECT -82.445 219.475 -82.115 219.805 ;
        RECT -82.445 218.115 -82.115 218.445 ;
        RECT -82.445 216.755 -82.115 217.085 ;
        RECT -82.445 215.395 -82.115 215.725 ;
        RECT -82.445 214.035 -82.115 214.365 ;
        RECT -82.445 212.675 -82.115 213.005 ;
        RECT -82.445 211.315 -82.115 211.645 ;
        RECT -82.445 209.955 -82.115 210.285 ;
        RECT -82.445 208.595 -82.115 208.925 ;
        RECT -82.445 207.235 -82.115 207.565 ;
        RECT -82.445 205.875 -82.115 206.205 ;
        RECT -82.445 204.515 -82.115 204.845 ;
        RECT -82.445 203.155 -82.115 203.485 ;
        RECT -82.445 201.795 -82.115 202.125 ;
        RECT -82.445 200.435 -82.115 200.765 ;
        RECT -82.445 199.075 -82.115 199.405 ;
        RECT -82.445 197.715 -82.115 198.045 ;
        RECT -82.445 196.355 -82.115 196.685 ;
        RECT -82.445 194.995 -82.115 195.325 ;
        RECT -82.445 193.635 -82.115 193.965 ;
        RECT -82.445 192.275 -82.115 192.605 ;
        RECT -82.445 190.915 -82.115 191.245 ;
        RECT -82.445 189.555 -82.115 189.885 ;
        RECT -82.445 188.195 -82.115 188.525 ;
        RECT -82.445 186.835 -82.115 187.165 ;
        RECT -82.445 185.475 -82.115 185.805 ;
        RECT -82.445 184.115 -82.115 184.445 ;
        RECT -82.445 182.755 -82.115 183.085 ;
        RECT -82.445 181.395 -82.115 181.725 ;
        RECT -82.445 180.035 -82.115 180.365 ;
        RECT -82.445 178.675 -82.115 179.005 ;
        RECT -82.445 177.315 -82.115 177.645 ;
        RECT -82.445 175.955 -82.115 176.285 ;
        RECT -82.445 174.595 -82.115 174.925 ;
        RECT -82.445 173.235 -82.115 173.565 ;
        RECT -82.445 171.875 -82.115 172.205 ;
        RECT -82.445 170.515 -82.115 170.845 ;
        RECT -82.445 169.155 -82.115 169.485 ;
        RECT -82.445 167.795 -82.115 168.125 ;
        RECT -82.445 166.435 -82.115 166.765 ;
        RECT -82.445 165.075 -82.115 165.405 ;
        RECT -82.445 163.715 -82.115 164.045 ;
        RECT -82.445 162.355 -82.115 162.685 ;
        RECT -82.445 160.995 -82.115 161.325 ;
        RECT -82.445 159.635 -82.115 159.965 ;
        RECT -82.445 158.275 -82.115 158.605 ;
        RECT -82.445 156.915 -82.115 157.245 ;
        RECT -82.445 155.555 -82.115 155.885 ;
        RECT -82.445 154.195 -82.115 154.525 ;
        RECT -82.445 152.835 -82.115 153.165 ;
        RECT -82.445 151.475 -82.115 151.805 ;
        RECT -82.445 150.115 -82.115 150.445 ;
        RECT -82.445 148.755 -82.115 149.085 ;
        RECT -82.445 147.395 -82.115 147.725 ;
        RECT -82.445 146.035 -82.115 146.365 ;
        RECT -82.445 144.675 -82.115 145.005 ;
        RECT -82.445 143.315 -82.115 143.645 ;
        RECT -82.445 141.955 -82.115 142.285 ;
        RECT -82.445 140.595 -82.115 140.925 ;
        RECT -82.445 139.235 -82.115 139.565 ;
        RECT -82.445 137.875 -82.115 138.205 ;
        RECT -82.445 136.515 -82.115 136.845 ;
        RECT -82.445 135.155 -82.115 135.485 ;
        RECT -82.445 133.795 -82.115 134.125 ;
        RECT -82.445 132.435 -82.115 132.765 ;
        RECT -82.445 131.075 -82.115 131.405 ;
        RECT -82.445 129.715 -82.115 130.045 ;
        RECT -82.445 128.355 -82.115 128.685 ;
        RECT -82.445 126.995 -82.115 127.325 ;
        RECT -82.445 125.635 -82.115 125.965 ;
        RECT -82.445 124.275 -82.115 124.605 ;
        RECT -82.445 122.915 -82.115 123.245 ;
        RECT -82.445 121.555 -82.115 121.885 ;
        RECT -82.445 120.195 -82.115 120.525 ;
        RECT -82.445 118.835 -82.115 119.165 ;
        RECT -82.445 117.475 -82.115 117.805 ;
        RECT -82.445 116.115 -82.115 116.445 ;
        RECT -82.445 114.755 -82.115 115.085 ;
        RECT -82.445 113.395 -82.115 113.725 ;
        RECT -82.445 112.035 -82.115 112.365 ;
        RECT -82.445 110.675 -82.115 111.005 ;
        RECT -82.445 109.315 -82.115 109.645 ;
        RECT -82.445 107.955 -82.115 108.285 ;
        RECT -82.445 106.595 -82.115 106.925 ;
        RECT -82.445 105.235 -82.115 105.565 ;
        RECT -82.445 103.875 -82.115 104.205 ;
        RECT -82.445 102.515 -82.115 102.845 ;
        RECT -82.445 101.155 -82.115 101.485 ;
        RECT -82.445 99.795 -82.115 100.125 ;
        RECT -82.445 98.435 -82.115 98.765 ;
        RECT -82.445 97.075 -82.115 97.405 ;
        RECT -82.445 95.715 -82.115 96.045 ;
        RECT -82.445 94.355 -82.115 94.685 ;
        RECT -82.445 92.995 -82.115 93.325 ;
        RECT -82.445 91.635 -82.115 91.965 ;
        RECT -82.445 90.275 -82.115 90.605 ;
        RECT -82.445 88.915 -82.115 89.245 ;
        RECT -82.445 87.555 -82.115 87.885 ;
        RECT -82.445 86.195 -82.115 86.525 ;
        RECT -82.445 84.835 -82.115 85.165 ;
        RECT -82.445 83.475 -82.115 83.805 ;
        RECT -82.445 82.115 -82.115 82.445 ;
        RECT -82.445 80.755 -82.115 81.085 ;
        RECT -82.445 79.395 -82.115 79.725 ;
        RECT -82.445 78.035 -82.115 78.365 ;
        RECT -82.445 76.675 -82.115 77.005 ;
        RECT -82.445 75.315 -82.115 75.645 ;
        RECT -82.445 73.955 -82.115 74.285 ;
        RECT -82.445 72.595 -82.115 72.925 ;
        RECT -82.445 71.235 -82.115 71.565 ;
        RECT -82.445 69.875 -82.115 70.205 ;
        RECT -82.445 68.515 -82.115 68.845 ;
        RECT -82.445 67.155 -82.115 67.485 ;
        RECT -82.445 65.795 -82.115 66.125 ;
        RECT -82.445 64.435 -82.115 64.765 ;
        RECT -82.445 63.075 -82.115 63.405 ;
        RECT -82.445 61.715 -82.115 62.045 ;
        RECT -82.445 60.355 -82.115 60.685 ;
        RECT -82.445 58.995 -82.115 59.325 ;
        RECT -82.445 57.635 -82.115 57.965 ;
        RECT -82.445 56.275 -82.115 56.605 ;
        RECT -82.445 54.915 -82.115 55.245 ;
        RECT -82.445 53.555 -82.115 53.885 ;
        RECT -82.445 52.195 -82.115 52.525 ;
        RECT -82.445 50.835 -82.115 51.165 ;
        RECT -82.445 49.475 -82.115 49.805 ;
        RECT -82.445 48.115 -82.115 48.445 ;
        RECT -82.445 46.755 -82.115 47.085 ;
        RECT -82.445 45.395 -82.115 45.725 ;
        RECT -82.445 44.035 -82.115 44.365 ;
        RECT -82.445 42.675 -82.115 43.005 ;
        RECT -82.445 41.315 -82.115 41.645 ;
        RECT -82.445 39.955 -82.115 40.285 ;
        RECT -82.445 38.595 -82.115 38.925 ;
        RECT -82.445 37.235 -82.115 37.565 ;
        RECT -82.445 35.875 -82.115 36.205 ;
        RECT -82.445 34.515 -82.115 34.845 ;
        RECT -82.445 33.155 -82.115 33.485 ;
        RECT -82.445 31.795 -82.115 32.125 ;
        RECT -82.445 30.435 -82.115 30.765 ;
        RECT -82.445 29.075 -82.115 29.405 ;
        RECT -82.445 27.715 -82.115 28.045 ;
        RECT -82.445 26.355 -82.115 26.685 ;
        RECT -82.445 24.995 -82.115 25.325 ;
        RECT -82.445 23.635 -82.115 23.965 ;
        RECT -82.445 22.275 -82.115 22.605 ;
        RECT -82.445 20.915 -82.115 21.245 ;
        RECT -82.445 19.555 -82.115 19.885 ;
        RECT -82.445 18.195 -82.115 18.525 ;
        RECT -82.445 16.835 -82.115 17.165 ;
        RECT -82.445 15.475 -82.115 15.805 ;
        RECT -82.445 14.115 -82.115 14.445 ;
        RECT -82.445 12.755 -82.115 13.085 ;
        RECT -82.445 11.395 -82.115 11.725 ;
        RECT -82.445 10.035 -82.115 10.365 ;
        RECT -82.445 8.675 -82.115 9.005 ;
        RECT -82.445 7.315 -82.115 7.645 ;
        RECT -82.445 5.955 -82.115 6.285 ;
        RECT -82.445 4.595 -82.115 4.925 ;
        RECT -82.445 3.235 -82.115 3.565 ;
        RECT -82.445 1.875 -82.115 2.205 ;
        RECT -82.445 0.515 -82.115 0.845 ;
        RECT -82.445 -0.845 -82.115 -0.515 ;
        RECT -82.445 -2.205 -82.115 -1.875 ;
        RECT -82.445 -3.565 -82.115 -3.235 ;
        RECT -82.445 -4.925 -82.115 -4.595 ;
        RECT -82.445 -6.285 -82.115 -5.955 ;
        RECT -82.445 -7.645 -82.115 -7.315 ;
        RECT -82.445 -9.005 -82.115 -8.675 ;
        RECT -82.445 -10.365 -82.115 -10.035 ;
        RECT -82.445 -11.725 -82.115 -11.395 ;
        RECT -82.445 -13.085 -82.115 -12.755 ;
        RECT -82.445 -14.445 -82.115 -14.115 ;
        RECT -82.445 -15.805 -82.115 -15.475 ;
        RECT -82.445 -17.165 -82.115 -16.835 ;
        RECT -82.445 -18.525 -82.115 -18.195 ;
        RECT -82.445 -19.885 -82.115 -19.555 ;
        RECT -82.445 -21.245 -82.115 -20.915 ;
        RECT -82.445 -22.605 -82.115 -22.275 ;
        RECT -82.445 -23.965 -82.115 -23.635 ;
        RECT -82.445 -25.325 -82.115 -24.995 ;
        RECT -82.445 -26.685 -82.115 -26.355 ;
        RECT -82.445 -28.045 -82.115 -27.715 ;
        RECT -82.445 -29.405 -82.115 -29.075 ;
        RECT -82.445 -30.765 -82.115 -30.435 ;
        RECT -82.445 -32.125 -82.115 -31.795 ;
        RECT -82.445 -33.485 -82.115 -33.155 ;
        RECT -82.445 -34.845 -82.115 -34.515 ;
        RECT -82.445 -36.205 -82.115 -35.875 ;
        RECT -82.445 -37.565 -82.115 -37.235 ;
        RECT -82.445 -38.925 -82.115 -38.595 ;
        RECT -82.445 -40.285 -82.115 -39.955 ;
        RECT -82.445 -41.645 -82.115 -41.315 ;
        RECT -82.445 -43.005 -82.115 -42.675 ;
        RECT -82.445 -44.365 -82.115 -44.035 ;
        RECT -82.445 -45.725 -82.115 -45.395 ;
        RECT -82.445 -47.085 -82.115 -46.755 ;
        RECT -82.445 -48.445 -82.115 -48.115 ;
        RECT -82.445 -49.805 -82.115 -49.475 ;
        RECT -82.445 -51.165 -82.115 -50.835 ;
        RECT -82.445 -52.525 -82.115 -52.195 ;
        RECT -82.445 -53.885 -82.115 -53.555 ;
        RECT -82.445 -55.245 -82.115 -54.915 ;
        RECT -82.445 -56.605 -82.115 -56.275 ;
        RECT -82.445 -57.965 -82.115 -57.635 ;
        RECT -82.445 -59.325 -82.115 -58.995 ;
        RECT -82.445 -60.685 -82.115 -60.355 ;
        RECT -82.445 -62.045 -82.115 -61.715 ;
        RECT -82.445 -63.405 -82.115 -63.075 ;
        RECT -82.445 -64.765 -82.115 -64.435 ;
        RECT -82.445 -66.125 -82.115 -65.795 ;
        RECT -82.445 -67.485 -82.115 -67.155 ;
        RECT -82.445 -68.845 -82.115 -68.515 ;
        RECT -82.445 -70.205 -82.115 -69.875 ;
        RECT -82.445 -71.565 -82.115 -71.235 ;
        RECT -82.445 -72.925 -82.115 -72.595 ;
        RECT -82.445 -74.285 -82.115 -73.955 ;
        RECT -82.445 -75.645 -82.115 -75.315 ;
        RECT -82.445 -77.005 -82.115 -76.675 ;
        RECT -82.445 -78.365 -82.115 -78.035 ;
        RECT -82.445 -79.725 -82.115 -79.395 ;
        RECT -82.445 -81.085 -82.115 -80.755 ;
        RECT -82.445 -82.445 -82.115 -82.115 ;
        RECT -82.445 -83.805 -82.115 -83.475 ;
        RECT -82.445 -85.165 -82.115 -84.835 ;
        RECT -82.445 -86.525 -82.115 -86.195 ;
        RECT -82.445 -87.885 -82.115 -87.555 ;
        RECT -82.445 -89.245 -82.115 -88.915 ;
        RECT -82.445 -90.605 -82.115 -90.275 ;
        RECT -82.445 -91.965 -82.115 -91.635 ;
        RECT -82.445 -93.325 -82.115 -92.995 ;
        RECT -82.445 -94.685 -82.115 -94.355 ;
        RECT -82.445 -96.045 -82.115 -95.715 ;
        RECT -82.445 -97.405 -82.115 -97.075 ;
        RECT -82.445 -98.765 -82.115 -98.435 ;
        RECT -82.445 -100.125 -82.115 -99.795 ;
        RECT -82.445 -101.485 -82.115 -101.155 ;
        RECT -82.445 -102.845 -82.115 -102.515 ;
        RECT -82.445 -104.205 -82.115 -103.875 ;
        RECT -82.445 -105.565 -82.115 -105.235 ;
        RECT -82.445 -106.925 -82.115 -106.595 ;
        RECT -82.445 -108.285 -82.115 -107.955 ;
        RECT -82.445 -109.645 -82.115 -109.315 ;
        RECT -82.445 -111.005 -82.115 -110.675 ;
        RECT -82.445 -112.365 -82.115 -112.035 ;
        RECT -82.445 -113.725 -82.115 -113.395 ;
        RECT -82.445 -115.085 -82.115 -114.755 ;
        RECT -82.445 -116.445 -82.115 -116.115 ;
        RECT -82.445 -117.805 -82.115 -117.475 ;
        RECT -82.445 -119.165 -82.115 -118.835 ;
        RECT -82.445 -120.525 -82.115 -120.195 ;
        RECT -82.445 -121.885 -82.115 -121.555 ;
        RECT -82.445 -123.245 -82.115 -122.915 ;
        RECT -82.445 -124.605 -82.115 -124.275 ;
        RECT -82.445 -125.965 -82.115 -125.635 ;
        RECT -82.445 -127.325 -82.115 -126.995 ;
        RECT -82.445 -128.685 -82.115 -128.355 ;
        RECT -82.445 -130.045 -82.115 -129.715 ;
        RECT -82.445 -131.405 -82.115 -131.075 ;
        RECT -82.445 -132.765 -82.115 -132.435 ;
        RECT -82.445 -134.125 -82.115 -133.795 ;
        RECT -82.445 -135.485 -82.115 -135.155 ;
        RECT -82.445 -136.845 -82.115 -136.515 ;
        RECT -82.445 -138.205 -82.115 -137.875 ;
        RECT -82.445 -139.565 -82.115 -139.235 ;
        RECT -82.445 -140.925 -82.115 -140.595 ;
        RECT -82.445 -142.285 -82.115 -141.955 ;
        RECT -82.445 -143.645 -82.115 -143.315 ;
        RECT -82.445 -145.005 -82.115 -144.675 ;
        RECT -82.445 -146.365 -82.115 -146.035 ;
        RECT -82.445 -147.725 -82.115 -147.395 ;
        RECT -82.445 -149.085 -82.115 -148.755 ;
        RECT -82.445 -150.445 -82.115 -150.115 ;
        RECT -82.445 -151.805 -82.115 -151.475 ;
        RECT -82.445 -153.165 -82.115 -152.835 ;
        RECT -82.445 -154.525 -82.115 -154.195 ;
        RECT -82.445 -155.885 -82.115 -155.555 ;
        RECT -82.445 -157.245 -82.115 -156.915 ;
        RECT -82.445 -158.605 -82.115 -158.275 ;
        RECT -82.445 -159.965 -82.115 -159.635 ;
        RECT -82.445 -161.325 -82.115 -160.995 ;
        RECT -82.445 -162.685 -82.115 -162.355 ;
        RECT -82.445 -164.045 -82.115 -163.715 ;
        RECT -82.445 -165.405 -82.115 -165.075 ;
        RECT -82.445 -166.765 -82.115 -166.435 ;
        RECT -82.445 -168.125 -82.115 -167.795 ;
        RECT -82.445 -169.485 -82.115 -169.155 ;
        RECT -82.445 -170.845 -82.115 -170.515 ;
        RECT -82.445 -172.205 -82.115 -171.875 ;
        RECT -82.445 -173.565 -82.115 -173.235 ;
        RECT -82.445 -174.925 -82.115 -174.595 ;
        RECT -82.445 -176.285 -82.115 -175.955 ;
        RECT -82.445 -177.645 -82.115 -177.315 ;
        RECT -82.445 -179.005 -82.115 -178.675 ;
        RECT -82.445 -180.365 -82.115 -180.035 ;
        RECT -82.445 -181.725 -82.115 -181.395 ;
        RECT -82.445 -183.085 -82.115 -182.755 ;
        RECT -82.445 -184.445 -82.115 -184.115 ;
        RECT -82.445 -185.805 -82.115 -185.475 ;
        RECT -82.445 -187.165 -82.115 -186.835 ;
        RECT -82.445 -188.525 -82.115 -188.195 ;
        RECT -82.445 -189.885 -82.115 -189.555 ;
        RECT -82.445 -191.245 -82.115 -190.915 ;
        RECT -82.445 -192.605 -82.115 -192.275 ;
        RECT -82.445 -193.965 -82.115 -193.635 ;
        RECT -82.445 -195.325 -82.115 -194.995 ;
        RECT -82.445 -196.685 -82.115 -196.355 ;
        RECT -82.445 -198.045 -82.115 -197.715 ;
        RECT -82.445 -199.405 -82.115 -199.075 ;
        RECT -82.445 -200.765 -82.115 -200.435 ;
        RECT -82.445 -202.125 -82.115 -201.795 ;
        RECT -82.445 -203.485 -82.115 -203.155 ;
        RECT -82.445 -204.845 -82.115 -204.515 ;
        RECT -82.445 -206.205 -82.115 -205.875 ;
        RECT -82.445 -207.565 -82.115 -207.235 ;
        RECT -82.445 -208.925 -82.115 -208.595 ;
        RECT -82.445 -210.285 -82.115 -209.955 ;
        RECT -82.445 -211.645 -82.115 -211.315 ;
        RECT -82.445 -213.005 -82.115 -212.675 ;
        RECT -82.445 -214.365 -82.115 -214.035 ;
        RECT -82.445 -215.725 -82.115 -215.395 ;
        RECT -82.445 -217.085 -82.115 -216.755 ;
        RECT -82.445 -218.445 -82.115 -218.115 ;
        RECT -82.445 -219.805 -82.115 -219.475 ;
        RECT -82.445 -221.165 -82.115 -220.835 ;
        RECT -82.445 -222.525 -82.115 -222.195 ;
        RECT -82.445 -223.885 -82.115 -223.555 ;
        RECT -82.445 -225.245 -82.115 -224.915 ;
        RECT -82.445 -226.605 -82.115 -226.275 ;
        RECT -82.445 -227.965 -82.115 -227.635 ;
        RECT -82.445 -229.325 -82.115 -228.995 ;
        RECT -82.445 -230.685 -82.115 -230.355 ;
        RECT -82.445 -232.045 -82.115 -231.715 ;
        RECT -82.445 -233.405 -82.115 -233.075 ;
        RECT -82.445 -234.765 -82.115 -234.435 ;
        RECT -82.445 -236.125 -82.115 -235.795 ;
        RECT -82.445 -237.485 -82.115 -237.155 ;
        RECT -82.445 -238.845 -82.115 -238.515 ;
        RECT -82.445 -241.09 -82.115 -239.96 ;
        RECT -82.44 -241.205 -82.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -81.085 16.835 -80.755 17.165 ;
        RECT -81.085 15.475 -80.755 15.805 ;
        RECT -81.085 14.115 -80.755 14.445 ;
        RECT -81.085 12.755 -80.755 13.085 ;
        RECT -81.085 11.395 -80.755 11.725 ;
        RECT -81.085 10.035 -80.755 10.365 ;
        RECT -81.085 8.675 -80.755 9.005 ;
        RECT -81.085 7.315 -80.755 7.645 ;
        RECT -81.085 5.955 -80.755 6.285 ;
        RECT -81.085 4.595 -80.755 4.925 ;
        RECT -81.085 3.235 -80.755 3.565 ;
        RECT -81.085 1.875 -80.755 2.205 ;
        RECT -81.085 0.515 -80.755 0.845 ;
        RECT -81.085 -0.845 -80.755 -0.515 ;
        RECT -81.085 -2.205 -80.755 -1.875 ;
        RECT -81.085 -3.565 -80.755 -3.235 ;
        RECT -81.085 -4.925 -80.755 -4.595 ;
        RECT -81.085 -6.285 -80.755 -5.955 ;
        RECT -81.085 -7.645 -80.755 -7.315 ;
        RECT -81.085 -9.005 -80.755 -8.675 ;
        RECT -81.085 -10.365 -80.755 -10.035 ;
        RECT -81.085 -11.725 -80.755 -11.395 ;
        RECT -81.085 -13.085 -80.755 -12.755 ;
        RECT -81.085 -14.445 -80.755 -14.115 ;
        RECT -81.085 -15.805 -80.755 -15.475 ;
        RECT -81.085 -17.165 -80.755 -16.835 ;
        RECT -81.085 -18.525 -80.755 -18.195 ;
        RECT -81.085 -19.885 -80.755 -19.555 ;
        RECT -81.085 -21.245 -80.755 -20.915 ;
        RECT -81.085 -22.605 -80.755 -22.275 ;
        RECT -81.085 -23.965 -80.755 -23.635 ;
        RECT -81.085 -25.325 -80.755 -24.995 ;
        RECT -81.085 -26.685 -80.755 -26.355 ;
        RECT -81.085 -28.045 -80.755 -27.715 ;
        RECT -81.085 -29.405 -80.755 -29.075 ;
        RECT -81.085 -30.765 -80.755 -30.435 ;
        RECT -81.085 -32.125 -80.755 -31.795 ;
        RECT -81.085 -33.485 -80.755 -33.155 ;
        RECT -81.085 -34.845 -80.755 -34.515 ;
        RECT -81.085 -36.205 -80.755 -35.875 ;
        RECT -81.085 -37.565 -80.755 -37.235 ;
        RECT -81.085 -38.925 -80.755 -38.595 ;
        RECT -81.085 -40.285 -80.755 -39.955 ;
        RECT -81.085 -41.645 -80.755 -41.315 ;
        RECT -81.085 -43.005 -80.755 -42.675 ;
        RECT -81.085 -44.365 -80.755 -44.035 ;
        RECT -81.085 -45.725 -80.755 -45.395 ;
        RECT -81.085 -47.085 -80.755 -46.755 ;
        RECT -81.085 -48.445 -80.755 -48.115 ;
        RECT -81.085 -49.805 -80.755 -49.475 ;
        RECT -81.085 -51.165 -80.755 -50.835 ;
        RECT -81.085 -52.525 -80.755 -52.195 ;
        RECT -81.085 -53.885 -80.755 -53.555 ;
        RECT -81.085 -55.245 -80.755 -54.915 ;
        RECT -81.085 -56.605 -80.755 -56.275 ;
        RECT -81.085 -57.965 -80.755 -57.635 ;
        RECT -81.085 -59.325 -80.755 -58.995 ;
        RECT -81.085 -60.685 -80.755 -60.355 ;
        RECT -81.085 -62.045 -80.755 -61.715 ;
        RECT -81.085 -63.405 -80.755 -63.075 ;
        RECT -81.085 -64.765 -80.755 -64.435 ;
        RECT -81.085 -66.125 -80.755 -65.795 ;
        RECT -81.085 -67.485 -80.755 -67.155 ;
        RECT -81.085 -68.845 -80.755 -68.515 ;
        RECT -81.085 -70.205 -80.755 -69.875 ;
        RECT -81.085 -71.565 -80.755 -71.235 ;
        RECT -81.085 -72.925 -80.755 -72.595 ;
        RECT -81.085 -74.285 -80.755 -73.955 ;
        RECT -81.085 -75.645 -80.755 -75.315 ;
        RECT -81.085 -77.005 -80.755 -76.675 ;
        RECT -81.085 -78.365 -80.755 -78.035 ;
        RECT -81.085 -79.725 -80.755 -79.395 ;
        RECT -81.085 -81.085 -80.755 -80.755 ;
        RECT -81.085 -82.445 -80.755 -82.115 ;
        RECT -81.085 -83.805 -80.755 -83.475 ;
        RECT -81.085 -85.165 -80.755 -84.835 ;
        RECT -81.085 -86.525 -80.755 -86.195 ;
        RECT -81.085 -87.885 -80.755 -87.555 ;
        RECT -81.085 -89.245 -80.755 -88.915 ;
        RECT -81.085 -90.605 -80.755 -90.275 ;
        RECT -81.085 -91.965 -80.755 -91.635 ;
        RECT -81.085 -93.325 -80.755 -92.995 ;
        RECT -81.085 -94.685 -80.755 -94.355 ;
        RECT -81.085 -96.045 -80.755 -95.715 ;
        RECT -81.085 -97.405 -80.755 -97.075 ;
        RECT -81.085 -98.765 -80.755 -98.435 ;
        RECT -81.085 -100.125 -80.755 -99.795 ;
        RECT -81.085 -101.485 -80.755 -101.155 ;
        RECT -81.085 -102.845 -80.755 -102.515 ;
        RECT -81.085 -104.205 -80.755 -103.875 ;
        RECT -81.085 -105.565 -80.755 -105.235 ;
        RECT -81.085 -106.925 -80.755 -106.595 ;
        RECT -81.085 -108.285 -80.755 -107.955 ;
        RECT -81.085 -109.645 -80.755 -109.315 ;
        RECT -81.085 -111.005 -80.755 -110.675 ;
        RECT -81.085 -112.365 -80.755 -112.035 ;
        RECT -81.085 -113.725 -80.755 -113.395 ;
        RECT -81.085 -115.085 -80.755 -114.755 ;
        RECT -81.085 -116.445 -80.755 -116.115 ;
        RECT -81.085 -117.805 -80.755 -117.475 ;
        RECT -81.085 -119.165 -80.755 -118.835 ;
        RECT -81.085 -120.525 -80.755 -120.195 ;
        RECT -81.085 -121.885 -80.755 -121.555 ;
        RECT -81.085 -123.245 -80.755 -122.915 ;
        RECT -81.085 -124.605 -80.755 -124.275 ;
        RECT -81.085 -125.965 -80.755 -125.635 ;
        RECT -81.085 -127.325 -80.755 -126.995 ;
        RECT -81.085 -128.685 -80.755 -128.355 ;
        RECT -81.085 -130.045 -80.755 -129.715 ;
        RECT -81.085 -131.405 -80.755 -131.075 ;
        RECT -81.085 -132.765 -80.755 -132.435 ;
        RECT -81.085 -134.125 -80.755 -133.795 ;
        RECT -81.085 -135.485 -80.755 -135.155 ;
        RECT -81.085 -136.845 -80.755 -136.515 ;
        RECT -81.085 -138.205 -80.755 -137.875 ;
        RECT -81.085 -139.565 -80.755 -139.235 ;
        RECT -81.085 -140.925 -80.755 -140.595 ;
        RECT -81.085 -142.285 -80.755 -141.955 ;
        RECT -81.085 -143.645 -80.755 -143.315 ;
        RECT -81.085 -145.005 -80.755 -144.675 ;
        RECT -81.085 -146.365 -80.755 -146.035 ;
        RECT -81.085 -147.725 -80.755 -147.395 ;
        RECT -81.085 -149.085 -80.755 -148.755 ;
        RECT -81.085 -150.445 -80.755 -150.115 ;
        RECT -81.085 -151.805 -80.755 -151.475 ;
        RECT -81.085 -153.165 -80.755 -152.835 ;
        RECT -81.085 -154.525 -80.755 -154.195 ;
        RECT -81.085 -155.885 -80.755 -155.555 ;
        RECT -81.085 -157.245 -80.755 -156.915 ;
        RECT -81.085 -158.605 -80.755 -158.275 ;
        RECT -81.085 -159.965 -80.755 -159.635 ;
        RECT -81.085 -161.325 -80.755 -160.995 ;
        RECT -81.085 -162.685 -80.755 -162.355 ;
        RECT -81.085 -164.045 -80.755 -163.715 ;
        RECT -81.085 -165.405 -80.755 -165.075 ;
        RECT -81.085 -166.765 -80.755 -166.435 ;
        RECT -81.085 -168.125 -80.755 -167.795 ;
        RECT -81.085 -169.485 -80.755 -169.155 ;
        RECT -81.085 -170.845 -80.755 -170.515 ;
        RECT -81.085 -172.205 -80.755 -171.875 ;
        RECT -81.085 -173.565 -80.755 -173.235 ;
        RECT -81.085 -174.925 -80.755 -174.595 ;
        RECT -81.085 -176.285 -80.755 -175.955 ;
        RECT -81.085 -177.645 -80.755 -177.315 ;
        RECT -81.085 -179.005 -80.755 -178.675 ;
        RECT -81.085 -180.365 -80.755 -180.035 ;
        RECT -81.085 -181.725 -80.755 -181.395 ;
        RECT -81.085 -183.085 -80.755 -182.755 ;
        RECT -81.085 -184.445 -80.755 -184.115 ;
        RECT -81.085 -185.805 -80.755 -185.475 ;
        RECT -81.085 -187.165 -80.755 -186.835 ;
        RECT -81.085 -188.525 -80.755 -188.195 ;
        RECT -81.085 -189.885 -80.755 -189.555 ;
        RECT -81.085 -191.245 -80.755 -190.915 ;
        RECT -81.085 -192.605 -80.755 -192.275 ;
        RECT -81.085 -193.965 -80.755 -193.635 ;
        RECT -81.085 -195.325 -80.755 -194.995 ;
        RECT -81.085 -196.685 -80.755 -196.355 ;
        RECT -81.085 -198.045 -80.755 -197.715 ;
        RECT -81.085 -199.405 -80.755 -199.075 ;
        RECT -81.085 -200.765 -80.755 -200.435 ;
        RECT -81.085 -202.125 -80.755 -201.795 ;
        RECT -81.085 -203.485 -80.755 -203.155 ;
        RECT -81.085 -204.845 -80.755 -204.515 ;
        RECT -81.085 -206.205 -80.755 -205.875 ;
        RECT -81.085 -207.565 -80.755 -207.235 ;
        RECT -81.085 -208.925 -80.755 -208.595 ;
        RECT -81.085 -210.285 -80.755 -209.955 ;
        RECT -81.085 -211.645 -80.755 -211.315 ;
        RECT -81.085 -213.005 -80.755 -212.675 ;
        RECT -81.085 -214.365 -80.755 -214.035 ;
        RECT -81.085 -215.725 -80.755 -215.395 ;
        RECT -81.085 -217.085 -80.755 -216.755 ;
        RECT -81.085 -218.445 -80.755 -218.115 ;
        RECT -81.085 -219.805 -80.755 -219.475 ;
        RECT -81.085 -221.165 -80.755 -220.835 ;
        RECT -81.085 -222.525 -80.755 -222.195 ;
        RECT -81.085 -223.885 -80.755 -223.555 ;
        RECT -81.085 -225.245 -80.755 -224.915 ;
        RECT -81.085 -226.605 -80.755 -226.275 ;
        RECT -81.085 -227.965 -80.755 -227.635 ;
        RECT -81.085 -229.325 -80.755 -228.995 ;
        RECT -81.085 -230.685 -80.755 -230.355 ;
        RECT -81.085 -232.045 -80.755 -231.715 ;
        RECT -81.085 -233.405 -80.755 -233.075 ;
        RECT -81.085 -234.765 -80.755 -234.435 ;
        RECT -81.085 -236.125 -80.755 -235.795 ;
        RECT -81.085 -237.485 -80.755 -237.155 ;
        RECT -81.085 -238.845 -80.755 -238.515 ;
        RECT -81.085 -241.09 -80.755 -239.96 ;
        RECT -81.08 -241.205 -80.76 245.285 ;
        RECT -81.085 244.04 -80.755 245.17 ;
        RECT -81.085 242.595 -80.755 242.925 ;
        RECT -81.085 241.235 -80.755 241.565 ;
        RECT -81.085 239.875 -80.755 240.205 ;
        RECT -81.085 238.515 -80.755 238.845 ;
        RECT -81.085 237.155 -80.755 237.485 ;
        RECT -81.085 235.795 -80.755 236.125 ;
        RECT -81.085 234.435 -80.755 234.765 ;
        RECT -81.085 233.075 -80.755 233.405 ;
        RECT -81.085 231.715 -80.755 232.045 ;
        RECT -81.085 230.355 -80.755 230.685 ;
        RECT -81.085 228.995 -80.755 229.325 ;
        RECT -81.085 227.635 -80.755 227.965 ;
        RECT -81.085 226.275 -80.755 226.605 ;
        RECT -81.085 224.915 -80.755 225.245 ;
        RECT -81.085 223.555 -80.755 223.885 ;
        RECT -81.085 222.195 -80.755 222.525 ;
        RECT -81.085 220.835 -80.755 221.165 ;
        RECT -81.085 219.475 -80.755 219.805 ;
        RECT -81.085 218.115 -80.755 218.445 ;
        RECT -81.085 216.755 -80.755 217.085 ;
        RECT -81.085 215.395 -80.755 215.725 ;
        RECT -81.085 214.035 -80.755 214.365 ;
        RECT -81.085 212.675 -80.755 213.005 ;
        RECT -81.085 211.315 -80.755 211.645 ;
        RECT -81.085 209.955 -80.755 210.285 ;
        RECT -81.085 208.595 -80.755 208.925 ;
        RECT -81.085 207.235 -80.755 207.565 ;
        RECT -81.085 205.875 -80.755 206.205 ;
        RECT -81.085 204.515 -80.755 204.845 ;
        RECT -81.085 203.155 -80.755 203.485 ;
        RECT -81.085 201.795 -80.755 202.125 ;
        RECT -81.085 200.435 -80.755 200.765 ;
        RECT -81.085 199.075 -80.755 199.405 ;
        RECT -81.085 197.715 -80.755 198.045 ;
        RECT -81.085 196.355 -80.755 196.685 ;
        RECT -81.085 194.995 -80.755 195.325 ;
        RECT -81.085 193.635 -80.755 193.965 ;
        RECT -81.085 192.275 -80.755 192.605 ;
        RECT -81.085 190.915 -80.755 191.245 ;
        RECT -81.085 189.555 -80.755 189.885 ;
        RECT -81.085 188.195 -80.755 188.525 ;
        RECT -81.085 186.835 -80.755 187.165 ;
        RECT -81.085 185.475 -80.755 185.805 ;
        RECT -81.085 184.115 -80.755 184.445 ;
        RECT -81.085 182.755 -80.755 183.085 ;
        RECT -81.085 181.395 -80.755 181.725 ;
        RECT -81.085 180.035 -80.755 180.365 ;
        RECT -81.085 178.675 -80.755 179.005 ;
        RECT -81.085 177.315 -80.755 177.645 ;
        RECT -81.085 175.955 -80.755 176.285 ;
        RECT -81.085 174.595 -80.755 174.925 ;
        RECT -81.085 173.235 -80.755 173.565 ;
        RECT -81.085 171.875 -80.755 172.205 ;
        RECT -81.085 170.515 -80.755 170.845 ;
        RECT -81.085 169.155 -80.755 169.485 ;
        RECT -81.085 167.795 -80.755 168.125 ;
        RECT -81.085 166.435 -80.755 166.765 ;
        RECT -81.085 165.075 -80.755 165.405 ;
        RECT -81.085 163.715 -80.755 164.045 ;
        RECT -81.085 162.355 -80.755 162.685 ;
        RECT -81.085 160.995 -80.755 161.325 ;
        RECT -81.085 159.635 -80.755 159.965 ;
        RECT -81.085 158.275 -80.755 158.605 ;
        RECT -81.085 156.915 -80.755 157.245 ;
        RECT -81.085 155.555 -80.755 155.885 ;
        RECT -81.085 154.195 -80.755 154.525 ;
        RECT -81.085 152.835 -80.755 153.165 ;
        RECT -81.085 151.475 -80.755 151.805 ;
        RECT -81.085 150.115 -80.755 150.445 ;
        RECT -81.085 148.755 -80.755 149.085 ;
        RECT -81.085 147.395 -80.755 147.725 ;
        RECT -81.085 146.035 -80.755 146.365 ;
        RECT -81.085 144.675 -80.755 145.005 ;
        RECT -81.085 143.315 -80.755 143.645 ;
        RECT -81.085 141.955 -80.755 142.285 ;
        RECT -81.085 140.595 -80.755 140.925 ;
        RECT -81.085 139.235 -80.755 139.565 ;
        RECT -81.085 137.875 -80.755 138.205 ;
        RECT -81.085 136.515 -80.755 136.845 ;
        RECT -81.085 135.155 -80.755 135.485 ;
        RECT -81.085 133.795 -80.755 134.125 ;
        RECT -81.085 132.435 -80.755 132.765 ;
        RECT -81.085 131.075 -80.755 131.405 ;
        RECT -81.085 129.715 -80.755 130.045 ;
        RECT -81.085 128.355 -80.755 128.685 ;
        RECT -81.085 126.995 -80.755 127.325 ;
        RECT -81.085 125.635 -80.755 125.965 ;
        RECT -81.085 124.275 -80.755 124.605 ;
        RECT -81.085 122.915 -80.755 123.245 ;
        RECT -81.085 121.555 -80.755 121.885 ;
        RECT -81.085 120.195 -80.755 120.525 ;
        RECT -81.085 118.835 -80.755 119.165 ;
        RECT -81.085 117.475 -80.755 117.805 ;
        RECT -81.085 116.115 -80.755 116.445 ;
        RECT -81.085 114.755 -80.755 115.085 ;
        RECT -81.085 113.395 -80.755 113.725 ;
        RECT -81.085 112.035 -80.755 112.365 ;
        RECT -81.085 110.675 -80.755 111.005 ;
        RECT -81.085 109.315 -80.755 109.645 ;
        RECT -81.085 107.955 -80.755 108.285 ;
        RECT -81.085 106.595 -80.755 106.925 ;
        RECT -81.085 105.235 -80.755 105.565 ;
        RECT -81.085 103.875 -80.755 104.205 ;
        RECT -81.085 102.515 -80.755 102.845 ;
        RECT -81.085 101.155 -80.755 101.485 ;
        RECT -81.085 99.795 -80.755 100.125 ;
        RECT -81.085 98.435 -80.755 98.765 ;
        RECT -81.085 97.075 -80.755 97.405 ;
        RECT -81.085 95.715 -80.755 96.045 ;
        RECT -81.085 94.355 -80.755 94.685 ;
        RECT -81.085 92.995 -80.755 93.325 ;
        RECT -81.085 91.635 -80.755 91.965 ;
        RECT -81.085 90.275 -80.755 90.605 ;
        RECT -81.085 88.915 -80.755 89.245 ;
        RECT -81.085 87.555 -80.755 87.885 ;
        RECT -81.085 86.195 -80.755 86.525 ;
        RECT -81.085 84.835 -80.755 85.165 ;
        RECT -81.085 83.475 -80.755 83.805 ;
        RECT -81.085 82.115 -80.755 82.445 ;
        RECT -81.085 80.755 -80.755 81.085 ;
        RECT -81.085 79.395 -80.755 79.725 ;
        RECT -81.085 78.035 -80.755 78.365 ;
        RECT -81.085 76.675 -80.755 77.005 ;
        RECT -81.085 75.315 -80.755 75.645 ;
        RECT -81.085 73.955 -80.755 74.285 ;
        RECT -81.085 72.595 -80.755 72.925 ;
        RECT -81.085 71.235 -80.755 71.565 ;
        RECT -81.085 69.875 -80.755 70.205 ;
        RECT -81.085 68.515 -80.755 68.845 ;
        RECT -81.085 67.155 -80.755 67.485 ;
        RECT -81.085 65.795 -80.755 66.125 ;
        RECT -81.085 64.435 -80.755 64.765 ;
        RECT -81.085 63.075 -80.755 63.405 ;
        RECT -81.085 61.715 -80.755 62.045 ;
        RECT -81.085 60.355 -80.755 60.685 ;
        RECT -81.085 58.995 -80.755 59.325 ;
        RECT -81.085 57.635 -80.755 57.965 ;
        RECT -81.085 56.275 -80.755 56.605 ;
        RECT -81.085 54.915 -80.755 55.245 ;
        RECT -81.085 53.555 -80.755 53.885 ;
        RECT -81.085 52.195 -80.755 52.525 ;
        RECT -81.085 50.835 -80.755 51.165 ;
        RECT -81.085 49.475 -80.755 49.805 ;
        RECT -81.085 48.115 -80.755 48.445 ;
        RECT -81.085 46.755 -80.755 47.085 ;
        RECT -81.085 45.395 -80.755 45.725 ;
        RECT -81.085 44.035 -80.755 44.365 ;
        RECT -81.085 42.675 -80.755 43.005 ;
        RECT -81.085 41.315 -80.755 41.645 ;
        RECT -81.085 39.955 -80.755 40.285 ;
        RECT -81.085 38.595 -80.755 38.925 ;
        RECT -81.085 37.235 -80.755 37.565 ;
        RECT -81.085 35.875 -80.755 36.205 ;
        RECT -81.085 34.515 -80.755 34.845 ;
        RECT -81.085 33.155 -80.755 33.485 ;
        RECT -81.085 31.795 -80.755 32.125 ;
        RECT -81.085 30.435 -80.755 30.765 ;
        RECT -81.085 29.075 -80.755 29.405 ;
        RECT -81.085 27.715 -80.755 28.045 ;
        RECT -81.085 26.355 -80.755 26.685 ;
        RECT -81.085 24.995 -80.755 25.325 ;
        RECT -81.085 23.635 -80.755 23.965 ;
        RECT -81.085 22.275 -80.755 22.605 ;
        RECT -81.085 20.915 -80.755 21.245 ;
        RECT -81.085 19.555 -80.755 19.885 ;
        RECT -81.085 18.195 -80.755 18.525 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -21.92 -244.085 -21.6 -243.765 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.04 -244.085 -27.72 -243.765 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -34.16 -244.085 -33.84 -243.765 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -40.28 -244.085 -39.96 -243.765 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -46.4 -244.085 -46.08 -243.765 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -52.52 -244.085 -52.2 -243.765 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -58.64 -244.085 -58.32 -243.765 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -65.44 -244.085 -65.12 -243.765 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -71.56 -244.085 -71.24 -243.765 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -77.68 -244.085 -77.36 -243.765 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -9.68 -244.085 -9.36 -243.765 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.6 -244.085 6 -243.685 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 114.6 -244.085 115 -243.685 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 125.5 -244.085 125.9 -243.685 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.4 -244.085 136.8 -243.685 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 147.3 -244.085 147.7 -243.685 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.2 -244.085 158.6 -243.685 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 169.1 -244.085 169.5 -243.685 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 180 -244.085 180.4 -243.685 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 190.9 -244.085 191.3 -243.685 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.8 -244.085 202.2 -243.685 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.7 -244.085 213.1 -243.685 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.5 -244.085 16.9 -243.685 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 223.6 -244.085 224 -243.685 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 234.5 -244.085 234.9 -243.685 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 245.4 -244.085 245.8 -243.685 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.3 -244.085 256.7 -243.685 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 267.2 -244.085 267.6 -243.685 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 278.1 -244.085 278.5 -243.685 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 289 -244.085 289.4 -243.685 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 299.9 -244.085 300.3 -243.685 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 310.8 -244.085 311.2 -243.685 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 321.7 -244.085 322.1 -243.685 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 27.4 -244.085 27.8 -243.685 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 332.6 -244.085 333 -243.685 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 343.5 -244.085 343.9 -243.685 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 38.3 -244.085 38.7 -243.685 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 49.2 -244.085 49.6 -243.685 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.1 -244.085 60.5 -243.685 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71 -244.085 71.4 -243.685 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 81.9 -244.085 82.3 -243.685 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 92.8 -244.085 93.2 -243.685 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.7 -244.085 104.1 -243.685 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4 -244.085 4.4 -243.685 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113 -244.085 113.4 -243.685 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 123.9 -244.085 124.3 -243.685 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.8 -244.085 135.2 -243.685 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 145.7 -244.085 146.1 -243.685 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.6 -244.085 157 -243.685 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 167.5 -244.085 167.9 -243.685 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.4 -244.085 178.8 -243.685 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 189.3 -244.085 189.7 -243.685 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.2 -244.085 200.6 -243.685 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.1 -244.085 211.5 -243.685 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 14.9 -244.085 15.3 -243.685 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222 -244.085 222.4 -243.685 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.9 -244.085 233.3 -243.685 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 243.8 -244.085 244.2 -243.685 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.7 -244.085 255.1 -243.685 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 265.6 -244.085 266 -243.685 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.5 -244.085 276.9 -243.685 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 287.4 -244.085 287.8 -243.685 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 298.3 -244.085 298.7 -243.685 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 309.2 -244.085 309.6 -243.685 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 320.1 -244.085 320.5 -243.685 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.8 -244.085 26.2 -243.685 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 331 -244.085 331.4 -243.685 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 341.9 -244.085 342.3 -243.685 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.7 -244.085 37.1 -243.685 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 47.6 -244.085 48 -243.685 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.5 -244.085 58.9 -243.685 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 69.4 -244.085 69.8 -243.685 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.3 -244.085 80.7 -243.685 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 -244.085 91.6 -243.685 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.1 -244.085 102.5 -243.685 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -15.8 -244.085 -15.48 -243.765 ;
    END
  END we
  PIN wmask
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.4 -244.085 6.8 -243.685 ;
    END
  END wmask
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -89.065 -244.085 369.225 248.165 ;
    LAYER met2 SPACING 0.14 ;
      RECT -89.065 -244.085 369.225 248.165 ;
    LAYER met3 SPACING 0.3 ;
      RECT -1.525 -25.325 -1.195 -24.995 ;
      RECT -1.52 -134.805 -1.2 -24.995 ;
      RECT -1.525 -134.805 -1.195 -134.475 ;
      RECT -2.205 -23.965 -1.875 -23.635 ;
      RECT -2.2 -136.165 -1.88 -23.635 ;
      RECT -2.205 -136.165 -1.875 -135.835 ;
      RECT -2.885 -22.605 -2.555 -22.275 ;
      RECT -2.88 -137.525 -2.56 -22.275 ;
      RECT -2.885 -137.525 -2.555 -137.195 ;
      RECT -3.565 -21.245 -3.235 -20.915 ;
      RECT -3.56 -138.885 -3.24 -20.915 ;
      RECT -3.565 -138.885 -3.235 -138.555 ;
      RECT -9.685 -224.565 -9.355 -224.235 ;
      RECT -9.68 -243.275 -9.36 -224.235 ;
      RECT -9.685 -229.325 -9.355 -228.995 ;
      RECT -11.045 -225.245 -10.715 -224.915 ;
      RECT -11.04 -230.005 -10.72 -224.915 ;
      RECT -11.045 -230.005 -10.715 -229.675 ;
      RECT -12.405 -11.045 -12.075 -10.715 ;
      RECT -12.4 -161.325 -12.08 -10.715 ;
      RECT -12.405 -161.325 -12.075 -160.995 ;
      RECT -13.085 -117.805 -12.755 -117.475 ;
      RECT -13.08 -216.405 -12.76 -117.475 ;
      RECT -13.085 -216.405 -12.755 -216.075 ;
      RECT -15.8 -243.275 -15.48 -230.11 ;
      RECT -15.805 -230.56 -15.475 -230.23 ;
      RECT -16.485 -224.565 -16.155 -224.235 ;
      RECT -16.48 -231.365 -16.16 -224.235 ;
      RECT -16.485 -231.365 -16.155 -231.035 ;
      RECT -16.485 -71.565 -16.155 -71.235 ;
      RECT -16.48 -161.325 -16.16 -71.235 ;
      RECT -16.485 -161.325 -16.155 -160.995 ;
      RECT -17.165 -225.245 -16.835 -224.915 ;
      RECT -17.16 -230.005 -16.84 -224.915 ;
      RECT -17.165 -230.005 -16.835 -229.675 ;
      RECT -18.525 -148.73 -18.195 -148.4 ;
      RECT -18.52 -228.645 -18.2 -148.4 ;
      RECT -18.525 -228.645 -18.195 -228.315 ;
      RECT -18.525 -20.69 -18.195 -20.36 ;
      RECT -18.52 -128.005 -18.2 -20.36 ;
      RECT -18.525 -128.005 -18.195 -127.675 ;
      RECT -19.205 -149.21 -18.875 -148.88 ;
      RECT -19.2 -227.965 -18.88 -148.88 ;
      RECT -19.205 -227.965 -18.875 -227.635 ;
      RECT -19.205 -21.17 -18.875 -20.84 ;
      RECT -19.2 -127.325 -18.88 -20.84 ;
      RECT -19.205 -127.325 -18.875 -126.995 ;
      RECT -19.885 -149.69 -19.555 -149.36 ;
      RECT -19.88 -227.285 -19.56 -149.36 ;
      RECT -19.885 -227.285 -19.555 -226.955 ;
      RECT -19.885 -21.65 -19.555 -21.32 ;
      RECT -19.88 -126.645 -19.56 -21.32 ;
      RECT -19.885 -126.645 -19.555 -126.315 ;
      RECT -20.565 -150.17 -20.235 -149.84 ;
      RECT -20.56 -231.365 -20.24 -149.84 ;
      RECT -20.565 -231.365 -20.235 -231.035 ;
      RECT -20.565 -22.13 -20.235 -21.8 ;
      RECT -20.56 -125.965 -20.24 -21.8 ;
      RECT -20.565 -125.965 -20.235 -125.635 ;
      RECT -21.245 -150.65 -20.915 -150.32 ;
      RECT -21.24 -225.245 -20.92 -150.32 ;
      RECT -21.245 -225.245 -20.915 -224.915 ;
      RECT -21.245 -22.61 -20.915 -22.28 ;
      RECT -21.24 -125.285 -20.92 -22.28 ;
      RECT -21.245 -125.285 -20.915 -124.955 ;
      RECT -21.92 -243.275 -21.6 -230.11 ;
      RECT -21.925 -230.56 -21.595 -230.23 ;
      RECT -21.925 -151.13 -21.595 -150.8 ;
      RECT -21.92 -224.565 -21.6 -150.8 ;
      RECT -21.925 -224.565 -21.595 -224.235 ;
      RECT -21.925 -23.09 -21.595 -22.76 ;
      RECT -21.92 -123.245 -21.6 -22.76 ;
      RECT -21.925 -123.245 -21.595 -122.915 ;
      RECT -23.285 -227.285 -22.955 -226.955 ;
      RECT -23.28 -230.005 -22.96 -226.955 ;
      RECT -23.285 -230.005 -22.955 -229.675 ;
      RECT -28.04 -243.275 -27.72 -230.11 ;
      RECT -28.045 -230.56 -27.715 -230.23 ;
      RECT -28.725 -58.93 -28.395 -58.6 ;
      RECT -28.72 -121.885 -28.4 -58.6 ;
      RECT -28.725 -121.885 -28.395 -121.555 ;
      RECT -29.405 -228.645 -29.075 -228.315 ;
      RECT -29.4 -230.005 -29.08 -228.315 ;
      RECT -29.405 -230.005 -29.075 -229.675 ;
      RECT -29.405 -59.41 -29.075 -59.08 ;
      RECT -29.4 -122.565 -29.08 -59.08 ;
      RECT -29.405 -122.565 -29.075 -122.235 ;
      RECT -30.085 -227.965 -29.755 -227.635 ;
      RECT -30.08 -231.365 -29.76 -227.635 ;
      RECT -30.085 -231.365 -29.755 -231.035 ;
      RECT -30.085 -59.89 -29.755 -59.56 ;
      RECT -30.08 -121.205 -29.76 -59.56 ;
      RECT -30.085 -121.205 -29.755 -120.875 ;
      RECT -30.765 -60.37 -30.435 -60.04 ;
      RECT -30.76 -120.525 -30.44 -60.04 ;
      RECT -30.765 -120.525 -30.435 -120.195 ;
      RECT -34.16 -243.275 -33.84 -230.11 ;
      RECT -34.165 -230.56 -33.835 -230.23 ;
      RECT -35.525 -152.485 -35.195 -152.155 ;
      RECT -35.52 -230.005 -35.2 -152.155 ;
      RECT -35.525 -230.005 -35.195 -229.675 ;
      RECT -36.885 -2.205 -36.555 -1.875 ;
      RECT -36.88 -2.885 -36.56 -1.875 ;
      RECT -36.885 -2.885 -36.555 -2.555 ;
      RECT -38.925 -153.165 -38.595 -152.835 ;
      RECT -38.92 -231.365 -38.6 -152.835 ;
      RECT -38.925 -231.365 -38.595 -231.035 ;
      RECT -40.28 -243.275 -39.96 -230.11 ;
      RECT -40.285 -230.56 -39.955 -230.23 ;
      RECT -41.645 -152.485 -41.315 -152.155 ;
      RECT -41.64 -230.005 -41.32 -152.155 ;
      RECT -41.645 -230.005 -41.315 -229.675 ;
      RECT -42.325 -2.205 -41.995 -1.875 ;
      RECT -42.32 -6.965 -42 -1.875 ;
      RECT -42.325 -6.965 -41.995 -6.635 ;
      RECT -43.005 -58.93 -42.675 -58.6 ;
      RECT -43 -124.605 -42.68 -58.6 ;
      RECT -43.005 -124.605 -42.675 -124.275 ;
      RECT -43.685 -153.165 -43.355 -152.835 ;
      RECT -43.68 -231.365 -43.36 -152.835 ;
      RECT -43.685 -231.365 -43.355 -231.035 ;
      RECT -43.685 -59.41 -43.355 -59.08 ;
      RECT -43.68 -123.925 -43.36 -59.08 ;
      RECT -43.685 -123.925 -43.355 -123.595 ;
      RECT -44.365 -59.89 -44.035 -59.56 ;
      RECT -44.36 -122.565 -44.04 -59.56 ;
      RECT -44.365 -122.565 -44.035 -122.235 ;
      RECT -45.045 -60.37 -44.715 -60.04 ;
      RECT -45.04 -121.885 -44.72 -60.04 ;
      RECT -45.045 -121.885 -44.715 -121.555 ;
      RECT -46.4 -243.275 -46.08 -230.11 ;
      RECT -46.405 -230.56 -46.075 -230.23 ;
      RECT -46.405 -2.205 -46.075 -1.875 ;
      RECT -46.4 -27.365 -46.08 -1.875 ;
      RECT -46.405 -27.365 -46.075 -27.035 ;
      RECT -47.085 -2.205 -46.755 -1.875 ;
      RECT -47.08 -28.045 -46.76 -1.875 ;
      RECT -47.085 -28.045 -46.755 -27.715 ;
      RECT -47.765 -152.485 -47.435 -152.155 ;
      RECT -47.76 -230.005 -47.44 -152.155 ;
      RECT -47.765 -230.005 -47.435 -229.675 ;
      RECT -48.445 -150.445 -48.115 -150.115 ;
      RECT -48.44 -231.365 -48.12 -150.115 ;
      RECT -48.445 -231.365 -48.115 -231.035 ;
      RECT -50.08 116.48 -48.8 117.12 ;
      RECT -49.12 -158.605 -48.8 117.12 ;
      RECT -49.125 -158.605 -48.795 -158.275 ;
      RECT -52.52 -243.275 -52.2 -230.11 ;
      RECT -52.525 -230.56 -52.195 -230.23 ;
      RECT -53.205 -150.445 -52.875 -150.115 ;
      RECT -53.2 -231.365 -52.88 -150.115 ;
      RECT -53.205 -231.365 -52.875 -231.035 ;
      RECT -54.565 -152.485 -54.235 -152.155 ;
      RECT -54.56 -230.005 -54.24 -152.155 ;
      RECT -54.565 -230.005 -54.235 -229.675 ;
      RECT -55.925 86.875 -55.595 87.205 ;
      RECT -55.92 -11.045 -55.6 87.205 ;
      RECT -55.925 -11.045 -55.595 -10.715 ;
      RECT -56.605 86.195 -56.275 86.525 ;
      RECT -56.6 -161.325 -56.28 86.525 ;
      RECT -56.605 -161.325 -56.275 -160.995 ;
      RECT -57.965 -150.445 -57.635 -150.115 ;
      RECT -57.96 -231.365 -57.64 -150.115 ;
      RECT -57.965 -231.365 -57.635 -231.035 ;
      RECT -58.64 -243.275 -58.32 -230.11 ;
      RECT -58.645 -230.56 -58.315 -230.23 ;
      RECT -60.685 -152.485 -60.355 -152.155 ;
      RECT -60.68 -230.005 -60.36 -152.155 ;
      RECT -60.685 -230.005 -60.355 -229.675 ;
      RECT -63.405 -152.485 -63.075 -152.155 ;
      RECT -63.4 -231.365 -63.08 -152.155 ;
      RECT -63.405 -231.365 -63.075 -231.035 ;
      RECT -65.44 -243.275 -65.12 -230.11 ;
      RECT -65.445 -230.56 -65.115 -230.23 ;
      RECT -66.805 -150.445 -66.475 -150.115 ;
      RECT -66.8 -230.005 -66.48 -150.115 ;
      RECT -66.805 -230.005 -66.475 -229.675 ;
      RECT -68.165 -152.485 -67.835 -152.155 ;
      RECT -68.16 -231.365 -67.84 -152.155 ;
      RECT -68.165 -231.365 -67.835 -231.035 ;
      RECT -71.56 -243.275 -71.24 -230.11 ;
      RECT -71.565 -230.56 -71.235 -230.23 ;
      RECT -71.565 -151.805 -71.235 -151.475 ;
      RECT -71.56 -160.645 -71.24 -151.475 ;
      RECT -71.565 -160.645 -71.235 -160.315 ;
      RECT -72.925 -150.445 -72.595 -150.115 ;
      RECT -72.92 -230.005 -72.6 -150.115 ;
      RECT -72.925 -230.005 -72.595 -229.675 ;
      RECT -77.68 -243.275 -77.36 -230.11 ;
      RECT -77.685 -230.56 -77.355 -230.23 ;
      RECT 345.1 -111.675 345.5 -24.12 ;
      RECT 344.3 -110.815 344.7 -24.12 ;
      RECT 343.5 -243.195 343.9 -110.905 ;
      RECT 342.7 -94.96 343.1 -80.365 ;
      RECT 342.7 -76.54 343.1 -17.24 ;
      RECT 341.9 -243.195 342.3 -105.065 ;
      RECT 341.9 -95.46 342.3 -80.82 ;
      RECT 341.9 -76.97 342.3 -12.97 ;
      RECT 334.2 -111.675 334.6 -24.12 ;
      RECT 333.4 -110.815 333.8 -24.12 ;
      RECT 332.6 -243.195 333 -110.905 ;
      RECT 331.8 -94.96 332.2 -80.365 ;
      RECT 331.8 -76.54 332.2 -17.24 ;
      RECT 331 -243.195 331.4 -105.065 ;
      RECT 331 -95.46 331.4 -80.82 ;
      RECT 331 -76.97 331.4 -12.97 ;
      RECT 323.3 -111.675 323.7 -24.12 ;
      RECT 322.5 -110.815 322.9 -24.12 ;
      RECT 321.7 -243.195 322.1 -110.905 ;
      RECT 320.9 -94.96 321.3 -80.365 ;
      RECT 320.9 -76.54 321.3 -17.24 ;
      RECT 320.1 -243.195 320.5 -105.065 ;
      RECT 320.1 -95.46 320.5 -80.82 ;
      RECT 320.1 -76.97 320.5 -12.97 ;
      RECT 312.4 -111.675 312.8 -24.12 ;
      RECT 311.6 -110.815 312 -24.12 ;
      RECT 310.8 -243.195 311.2 -110.905 ;
      RECT 310 -94.96 310.4 -80.365 ;
      RECT 310 -76.54 310.4 -17.24 ;
      RECT 309.2 -243.195 309.6 -105.065 ;
      RECT 309.2 -95.46 309.6 -80.82 ;
      RECT 309.2 -76.97 309.6 -12.97 ;
      RECT 301.5 -111.675 301.9 -24.12 ;
      RECT 300.7 -110.815 301.1 -24.12 ;
      RECT 299.9 -243.195 300.3 -110.905 ;
      RECT 299.1 -94.96 299.5 -80.365 ;
      RECT 299.1 -76.54 299.5 -17.24 ;
      RECT 298.3 -243.195 298.7 -105.065 ;
      RECT 298.3 -95.46 298.7 -80.82 ;
      RECT 298.3 -76.97 298.7 -12.97 ;
      RECT 290.6 -111.675 291 -24.12 ;
      RECT 289.8 -110.815 290.2 -24.12 ;
      RECT 289 -243.195 289.4 -110.905 ;
      RECT 288.2 -94.96 288.6 -80.365 ;
      RECT 288.2 -76.54 288.6 -17.24 ;
      RECT 287.4 -243.195 287.8 -105.065 ;
      RECT 287.4 -95.46 287.8 -80.82 ;
      RECT 287.4 -76.97 287.8 -12.97 ;
      RECT 279.7 -111.675 280.1 -24.12 ;
      RECT 278.9 -110.815 279.3 -24.12 ;
      RECT 278.1 -243.195 278.5 -110.905 ;
      RECT 277.3 -94.96 277.7 -80.365 ;
      RECT 277.3 -76.54 277.7 -17.24 ;
      RECT 276.5 -243.195 276.9 -105.065 ;
      RECT 276.5 -95.46 276.9 -80.82 ;
      RECT 276.5 -76.97 276.9 -12.97 ;
      RECT 268.8 -111.675 269.2 -24.12 ;
      RECT 268 -110.815 268.4 -24.12 ;
      RECT 267.2 -243.195 267.6 -110.905 ;
      RECT 266.4 -94.96 266.8 -80.365 ;
      RECT 266.4 -76.54 266.8 -17.24 ;
      RECT 265.6 -243.195 266 -105.065 ;
      RECT 265.6 -95.46 266 -80.82 ;
      RECT 265.6 -76.97 266 -12.97 ;
      RECT 257.9 -111.675 258.3 -24.12 ;
      RECT 257.1 -110.815 257.5 -24.12 ;
      RECT 256.3 -243.195 256.7 -110.905 ;
      RECT 255.5 -94.96 255.9 -80.365 ;
      RECT 255.5 -76.54 255.9 -17.24 ;
      RECT 254.7 -243.195 255.1 -105.065 ;
      RECT 254.7 -95.46 255.1 -80.82 ;
      RECT 254.7 -76.97 255.1 -12.97 ;
      RECT 247 -111.675 247.4 -24.12 ;
      RECT 246.2 -110.815 246.6 -24.12 ;
      RECT 245.4 -243.195 245.8 -110.905 ;
      RECT 244.6 -94.96 245 -80.365 ;
      RECT 244.6 -76.54 245 -17.24 ;
      RECT 243.8 -243.195 244.2 -105.065 ;
      RECT 243.8 -95.46 244.2 -80.82 ;
      RECT 243.8 -76.97 244.2 -12.97 ;
      RECT 236.1 -111.675 236.5 -24.12 ;
      RECT 235.3 -110.815 235.7 -24.12 ;
      RECT 234.5 -243.195 234.9 -110.905 ;
      RECT 233.7 -94.96 234.1 -80.365 ;
      RECT 233.7 -76.54 234.1 -17.24 ;
      RECT 232.9 -243.195 233.3 -105.065 ;
      RECT 232.9 -95.46 233.3 -80.82 ;
      RECT 232.9 -76.97 233.3 -12.97 ;
      RECT 225.2 -111.675 225.6 -24.12 ;
      RECT 224.4 -110.815 224.8 -24.12 ;
      RECT 223.6 -243.195 224 -110.905 ;
      RECT 222.8 -94.96 223.2 -80.365 ;
      RECT 222.8 -76.54 223.2 -17.24 ;
      RECT 222 -243.195 222.4 -105.065 ;
      RECT 222 -95.46 222.4 -80.82 ;
      RECT 222 -76.97 222.4 -12.97 ;
      RECT 214.3 -111.675 214.7 -24.12 ;
      RECT 213.5 -110.815 213.9 -24.12 ;
      RECT 212.7 -243.195 213.1 -110.905 ;
      RECT 211.9 -94.96 212.3 -80.365 ;
      RECT 211.9 -76.54 212.3 -17.24 ;
      RECT 211.1 -243.195 211.5 -105.065 ;
      RECT 211.1 -95.46 211.5 -80.82 ;
      RECT 211.1 -76.97 211.5 -12.97 ;
      RECT 203.4 -111.675 203.8 -24.12 ;
      RECT 202.6 -110.815 203 -24.12 ;
      RECT 201.8 -243.195 202.2 -110.905 ;
      RECT 201 -94.96 201.4 -80.365 ;
      RECT 201 -76.54 201.4 -17.24 ;
      RECT 200.2 -243.195 200.6 -105.065 ;
      RECT 200.2 -95.46 200.6 -80.82 ;
      RECT 200.2 -76.97 200.6 -12.97 ;
      RECT 192.5 -111.675 192.9 -24.12 ;
      RECT 191.7 -110.815 192.1 -24.12 ;
      RECT 190.9 -243.195 191.3 -110.905 ;
      RECT 190.1 -94.96 190.5 -80.365 ;
      RECT 190.1 -76.54 190.5 -17.24 ;
      RECT 189.3 -243.195 189.7 -105.065 ;
      RECT 189.3 -95.46 189.7 -80.82 ;
      RECT 189.3 -76.97 189.7 -12.97 ;
      RECT 181.6 -111.675 182 -24.12 ;
      RECT 180.8 -110.815 181.2 -24.12 ;
      RECT 180 -243.195 180.4 -110.905 ;
      RECT 179.2 -94.96 179.6 -80.365 ;
      RECT 179.2 -76.54 179.6 -17.24 ;
      RECT 178.4 -243.195 178.8 -105.065 ;
      RECT 178.4 -95.46 178.8 -80.82 ;
      RECT 178.4 -76.97 178.8 -12.97 ;
      RECT 170.7 -111.675 171.1 -24.12 ;
      RECT 169.9 -110.815 170.3 -24.12 ;
      RECT 169.1 -243.195 169.5 -110.905 ;
      RECT 168.3 -94.96 168.7 -80.365 ;
      RECT 168.3 -76.54 168.7 -17.24 ;
      RECT 167.5 -243.195 167.9 -105.065 ;
      RECT 167.5 -95.46 167.9 -80.82 ;
      RECT 167.5 -76.97 167.9 -12.97 ;
      RECT 159.8 -111.675 160.2 -24.12 ;
      RECT 159 -110.815 159.4 -24.12 ;
      RECT 158.2 -243.195 158.6 -110.905 ;
      RECT 157.4 -94.96 157.8 -80.365 ;
      RECT 157.4 -76.54 157.8 -17.24 ;
      RECT 156.6 -243.195 157 -105.065 ;
      RECT 156.6 -95.46 157 -80.82 ;
      RECT 156.6 -76.97 157 -12.97 ;
      RECT 148.9 -111.675 149.3 -24.12 ;
      RECT 148.1 -110.815 148.5 -24.12 ;
      RECT 147.3 -243.195 147.7 -110.905 ;
      RECT 146.5 -94.96 146.9 -80.365 ;
      RECT 146.5 -76.54 146.9 -17.24 ;
      RECT 145.7 -243.195 146.1 -105.065 ;
      RECT 145.7 -95.46 146.1 -80.82 ;
      RECT 145.7 -76.97 146.1 -12.97 ;
      RECT 138 -111.675 138.4 -24.12 ;
      RECT 137.2 -110.815 137.6 -24.12 ;
      RECT 136.4 -243.195 136.8 -110.905 ;
      RECT 135.6 -94.96 136 -80.365 ;
      RECT 135.6 -76.54 136 -17.24 ;
      RECT 134.8 -243.195 135.2 -105.065 ;
      RECT 134.8 -95.46 135.2 -80.82 ;
      RECT 134.8 -76.97 135.2 -12.97 ;
      RECT 127.1 -111.675 127.5 -24.12 ;
      RECT 126.3 -110.815 126.7 -24.12 ;
      RECT 125.5 -243.195 125.9 -110.905 ;
      RECT 124.7 -94.96 125.1 -80.365 ;
      RECT 124.7 -76.54 125.1 -17.24 ;
      RECT 123.9 -243.195 124.3 -105.065 ;
      RECT 123.9 -95.46 124.3 -80.82 ;
      RECT 123.9 -76.97 124.3 -12.97 ;
      RECT 116.2 -111.675 116.6 -24.12 ;
      RECT 115.4 -110.815 115.8 -24.12 ;
      RECT 114.6 -243.195 115 -110.905 ;
      RECT 113.8 -94.96 114.2 -80.365 ;
      RECT 113.8 -76.54 114.2 -17.24 ;
      RECT 113 -243.195 113.4 -105.065 ;
      RECT 113 -95.46 113.4 -80.82 ;
      RECT 113 -76.97 113.4 -12.97 ;
      RECT 105.3 -111.675 105.7 -24.12 ;
      RECT 104.5 -110.815 104.9 -24.12 ;
      RECT 103.7 -243.195 104.1 -110.905 ;
      RECT 102.9 -94.96 103.3 -80.365 ;
      RECT 102.9 -76.54 103.3 -17.24 ;
      RECT 102.1 -243.195 102.5 -105.065 ;
      RECT 102.1 -95.46 102.5 -80.82 ;
      RECT 102.1 -76.97 102.5 -12.97 ;
      RECT 94.4 -111.675 94.8 -24.12 ;
      RECT 93.6 -110.815 94 -24.12 ;
      RECT 92.8 -243.195 93.2 -110.905 ;
      RECT 92 -94.96 92.4 -80.365 ;
      RECT 92 -76.54 92.4 -17.24 ;
      RECT 91.2 -243.195 91.6 -105.065 ;
      RECT 91.2 -95.46 91.6 -80.82 ;
      RECT 91.2 -76.97 91.6 -12.97 ;
      RECT 83.5 -111.675 83.9 -24.12 ;
      RECT 82.7 -110.815 83.1 -24.12 ;
      RECT 81.9 -243.195 82.3 -110.905 ;
      RECT 81.1 -94.96 81.5 -80.365 ;
      RECT 81.1 -76.54 81.5 -17.24 ;
      RECT 80.3 -243.195 80.7 -105.065 ;
      RECT 80.3 -95.46 80.7 -80.82 ;
      RECT 80.3 -76.97 80.7 -12.97 ;
      RECT 72.6 -111.675 73 -24.12 ;
      RECT 71.8 -110.815 72.2 -24.12 ;
      RECT 71 -243.195 71.4 -110.905 ;
      RECT 70.2 -94.96 70.6 -80.365 ;
      RECT 70.2 -76.54 70.6 -17.24 ;
      RECT 69.4 -243.195 69.8 -105.065 ;
      RECT 69.4 -95.46 69.8 -80.82 ;
      RECT 69.4 -76.97 69.8 -12.97 ;
      RECT 61.7 -111.675 62.1 -24.12 ;
      RECT 60.9 -110.815 61.3 -24.12 ;
      RECT 60.1 -243.195 60.5 -110.905 ;
      RECT 59.3 -94.96 59.7 -80.365 ;
      RECT 59.3 -76.54 59.7 -17.24 ;
      RECT 58.5 -243.195 58.9 -105.065 ;
      RECT 58.5 -95.46 58.9 -80.82 ;
      RECT 58.5 -76.97 58.9 -12.97 ;
      RECT 50.8 -111.675 51.2 -24.12 ;
      RECT 50 -110.815 50.4 -24.12 ;
      RECT 49.2 -243.195 49.6 -110.905 ;
      RECT 48.4 -94.96 48.8 -80.365 ;
      RECT 48.4 -76.54 48.8 -17.24 ;
      RECT 47.6 -243.195 48 -105.065 ;
      RECT 47.6 -95.46 48 -80.82 ;
      RECT 47.6 -76.97 48 -12.97 ;
      RECT 39.9 -111.675 40.3 -24.12 ;
      RECT 39.1 -110.815 39.5 -24.12 ;
      RECT 38.3 -243.195 38.7 -110.905 ;
      RECT 37.5 -94.96 37.9 -80.365 ;
      RECT 37.5 -76.54 37.9 -17.24 ;
      RECT 36.7 -243.195 37.1 -105.065 ;
      RECT 36.7 -95.46 37.1 -80.82 ;
      RECT 36.7 -76.97 37.1 -12.97 ;
      RECT 29 -111.675 29.4 -24.12 ;
      RECT 28.2 -110.815 28.6 -24.12 ;
      RECT 27.4 -243.195 27.8 -110.905 ;
      RECT 26.6 -94.96 27 -80.365 ;
      RECT 26.6 -76.54 27 -17.24 ;
      RECT 25.8 -243.195 26.2 -105.065 ;
      RECT 25.8 -95.46 26.2 -80.82 ;
      RECT 25.8 -76.97 26.2 -12.97 ;
      RECT 18.1 -111.675 18.5 -24.12 ;
      RECT 17.3 -110.815 17.7 -24.12 ;
      RECT 16.5 -243.195 16.9 -110.905 ;
      RECT 15.7 -94.96 16.1 -80.365 ;
      RECT 15.7 -76.54 16.1 -17.24 ;
      RECT 14.9 -243.195 15.3 -105.065 ;
      RECT 14.9 -95.46 15.3 -80.82 ;
      RECT 14.9 -76.97 15.3 -12.97 ;
      RECT 8 -118.52 8.4 -24.12 ;
      RECT 7.2 -111.675 7.6 -24.12 ;
      RECT 6.4 -243.195 6.8 -118.61 ;
      RECT 6.4 -110.815 6.8 -24.12 ;
      RECT 5.6 -243.195 6 -110.905 ;
      RECT 4.8 -94.96 5.2 -80.365 ;
      RECT 4.8 -76.54 5.2 -17.24 ;
      RECT 4 -243.195 4.4 -105.065 ;
      RECT 4 -95.46 4.4 -80.82 ;
      RECT 4 -76.97 4.4 -12.97 ;
  END
END sram22_1024x32m8w32

END LIBRARY
