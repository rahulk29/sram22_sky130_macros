* Substrate SPICE library
* This is a generated file. Be careful when editing manually: this file may be overwritten.


.SUBCKT sky130_fd_sc_hs__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 a_1800_291# a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X1 VGND CLK a_728_331# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Q a_2363_352# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR CLK a_728_331# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 a_1499_149# a_728_331# a_1586_149# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X5 a_536_81# a_331_392# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X6 a_156_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X7 a_298_294# a_818_418# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X8 a_70_74# a_728_331# a_298_294# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X9 a_331_392# a_728_331# a_1586_149# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 a_70_74# D a_156_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X11 a_818_418# a_728_331# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_818_418# a_728_331# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_1586_149# a_818_418# a_1755_389# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X14 Q_N a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 a_298_294# a_818_418# a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X16 VGND RESET_B a_536_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X17 a_1755_389# a_1800_291# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X18 a_1586_149# a_818_418# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Q a_2363_352# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 VGND a_1586_149# Q_N VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VGND a_1586_149# a_2363_352# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X22 VPWR a_298_294# a_331_392# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X23 a_298_294# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X24 a_1499_149# a_1800_291# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X25 VPWR a_331_392# a_683_485# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X26 VPWR D a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X27 VPWR RESET_B a_1800_291# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X28 a_1974_74# a_1586_149# a_1800_291# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X29 a_70_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X30 Q_N a_1586_149# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 VPWR a_1586_149# a_2363_352# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X32 VGND a_2363_352# Q VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X33 VPWR a_1586_149# Q_N VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND RESET_B a_1974_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X35 a_683_485# a_728_331# a_298_294# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X36 VGND a_298_294# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VPWR a_2363_352# Q VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__dfrbp_2

.SUBCKT sky130_fd_sc_hs__dfrbp_2_wrapper CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 CLK D RESET_B VGND VNB VPB VPWR Q Q_N sky130_fd_sc_hs__dfrbp_2

.ENDS sky130_fd_sc_hs__dfrbp_2_wrapper

.SUBCKT dff_array_8 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_8

.SUBCKT sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_2

.SUBCKT sky130_fd_sc_hs__inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_2

.ENDS sky130_fd_sc_hs__inv_2_wrapper

.SUBCKT sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_4

.SUBCKT sky130_fd_sc_hs__inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_4

.ENDS sky130_fd_sc_hs__inv_4_wrapper

.SUBCKT inv_chain_9 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_9

.SUBCKT sky130_fd_sc_hs__and2_4 A B VGND VNB VPB VPWR X

  X0 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X2 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X5 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X8 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X14 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X15 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_4

.SUBCKT sky130_fd_sc_hs__and2_4_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_4

.ENDS sky130_fd_sc_hs__and2_4_wrapper

.SUBCKT edge_detector din dout vdd vss

  Xdelay_chain din delayed vdd vss inv_chain_9
  Xand din delayed vss vss vdd vdd dout sky130_fd_sc_hs__and2_4_wrapper

.ENDS edge_detector

.SUBCKT sram_sp_horiz_wlstrap_p2 VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_horiz_wlstrap_p2

.SUBCKT sram_sp_horiz_wlstrap_p2_wrapper VSS VNB

  X0 VSS VNB sram_sp_horiz_wlstrap_p2

.ENDS sram_sp_horiz_wlstrap_p2_wrapper

.SUBCKT mos_w2640_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.640


.ENDS mos_w2640_l150_m1_nf1_id1

.SUBCKT mos_w1050_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.050


.ENDS mos_w1050_l150_m1_nf1_id0

.SUBCKT folded_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w2640_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1050_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2640_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1050_l150_m1_nf1_id0

.ENDS folded_inv_3

.SUBCKT sram_sp_colend BR VDD VSS BL VNB VPB

  X0 BR VNB BR VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_colend

.SUBCKT mos_w2540_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.540


.ENDS mos_w2540_l150_m1_nf1_id1

.SUBCKT mos_w1020_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.020


.ENDS mos_w1020_l150_m1_nf1_id0

.SUBCKT folded_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w2540_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1020_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2540_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1020_l150_m1_nf1_id0

.ENDS folded_inv_4

.SUBCKT sramgen_sp_sense_amp clk inn inp outn outp VDD VSS

  XSWOP outp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWON outn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMP midp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMN midn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XPFBP outp outn VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XPFBN outn outp VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XTAIL tail clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=4 w=1.680

  XNFBP outp outn midp VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XNFBN outn outp midn VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINP midn inp tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINN midp inn tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680


.ENDS sramgen_sp_sense_amp

.SUBCKT mos_w2000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.000


.ENDS mos_w2000_l150_m1_nf1_id0

.SUBCKT mos_w2500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.500


.ENDS mos_w2500_l150_m1_nf1_id1

.SUBCKT nand2 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2

.SUBCKT mos_w5000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=5.000


.ENDS mos_w5000_l150_m1_nf1_id1

.SUBCKT folded_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w2000_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w2000_l150_m1_nf1_id0

.ENDS folded_inv_1

.SUBCKT and2 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_1

.ENDS and2

.SUBCKT sky130_fd_sc_hs__and2_2 A B VGND VNB VPB VPWR X

  X0 a_31_74# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 X a_31_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 X a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_118_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 a_31_74# A a_118_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VPWR A a_31_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X6 VPWR a_31_74# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND a_31_74# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_2

.SUBCKT mos_w800_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.800


.ENDS mos_w800_l150_m1_nf1_id0

.SUBCKT mos_w3100_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=3.100


.ENDS mos_w3100_l150_m1_nf1_id0

.SUBCKT mos_w4500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=4.500


.ENDS mos_w4500_l150_m1_nf1_id1

.SUBCKT column_mos vdd vss bl

  Xgate_nmos vss bl vss vss mos_w800_l150_m1_nf1_id0
  Xdrain_nmos bl vss vss vss mos_w3100_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w4500_l150_m1_nf1_id1

.ENDS column_mos

.SUBCKT mos_w1250_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.250


.ENDS mos_w1250_l150_m1_nf1_id1

.SUBCKT mos_w500_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id0

.SUBCKT folded_inv vdd vss a y

  XMP0 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w500_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w500_l150_m1_nf1_id0

.ENDS folded_inv

.SUBCKT mos_w700_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id1

.SUBCKT mos_w700_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id0

.SUBCKT multi_finger_inv vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv

.SUBCKT multi_finger_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_1

.SUBCKT multi_finger_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_2

.SUBCKT multi_finger_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_3

.SUBCKT multi_finger_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_4

.SUBCKT decoder_stage_1 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv
  Xgate_2_0_0 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_2_0_1 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_2_0_2 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_3_0_0 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_1 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_2 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_3 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_4 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_5 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_6 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_7 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_8 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_9 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_4_0_0 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_1 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_2 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_3 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_4 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_5 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_6 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_7 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_8 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_9 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_10 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_11 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_12 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_13 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_14 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_15 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_16 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_17 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_18 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_19 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_20 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_21 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_5_0_0 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_1 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_2 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_3 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_4 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_5 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_6 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_7 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_8 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_9 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_10 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_11 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_12 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_13 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_14 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_15 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_16 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_17 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_18 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_19 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_20 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_21 vdd vss y_b y multi_finger_inv_4

.ENDS decoder_stage_1

.SUBCKT multi_finger_inv_8 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_8

.SUBCKT sramgen_svt_inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_2

.SUBCKT sramgen_svt_inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_2

.ENDS sramgen_svt_inv_2_wrapper

.SUBCKT sramgen_svt_inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_4

.SUBCKT sramgen_svt_inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_4

.ENDS sramgen_svt_inv_4_wrapper

.SUBCKT svt_inv_chain_30 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sramgen_svt_inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sramgen_svt_inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sramgen_svt_inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sramgen_svt_inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sramgen_svt_inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sramgen_svt_inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sramgen_svt_inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sramgen_svt_inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sramgen_svt_inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sramgen_svt_inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sramgen_svt_inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sramgen_svt_inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sramgen_svt_inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sramgen_svt_inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sramgen_svt_inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sramgen_svt_inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sramgen_svt_inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd x[17] sramgen_svt_inv_2_wrapper
  Xinv18 x[17] vss vss vdd vdd x[18] sramgen_svt_inv_2_wrapper
  Xinv19 x[18] vss vss vdd vdd x[19] sramgen_svt_inv_2_wrapper
  Xinv20 x[19] vss vss vdd vdd x[20] sramgen_svt_inv_2_wrapper
  Xinv21 x[20] vss vss vdd vdd x[21] sramgen_svt_inv_2_wrapper
  Xinv22 x[21] vss vss vdd vdd x[22] sramgen_svt_inv_2_wrapper
  Xinv23 x[22] vss vss vdd vdd x[23] sramgen_svt_inv_2_wrapper
  Xinv24 x[23] vss vss vdd vdd x[24] sramgen_svt_inv_2_wrapper
  Xinv25 x[24] vss vss vdd vdd x[25] sramgen_svt_inv_2_wrapper
  Xinv26 x[25] vss vss vdd vdd x[26] sramgen_svt_inv_2_wrapper
  Xinv27 x[26] vss vss vdd vdd x[27] sramgen_svt_inv_2_wrapper
  Xinv28 x[27] vss vss vdd vdd x[28] sramgen_svt_inv_2_wrapper
  Xinv29 x[28] vss vss vdd vdd dout sramgen_svt_inv_4_wrapper

.ENDS svt_inv_chain_30

.SUBCKT mos_w9900_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=9.900


.ENDS mos_w9900_l150_m1_nf1_id1

.SUBCKT mos_w5950_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=5.950


.ENDS mos_w5950_l150_m1_nf1_id1

.SUBCKT precharge_1 vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w9900_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w9900_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w5950_l150_m1_nf1_id1

.ENDS precharge_1

.SUBCKT multi_finger_inv_13 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_13

.SUBCKT sky130_fd_sc_hs__nand2_8 A B VGND VNB VPB VPWR Y

  X0 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nand2_8

.SUBCKT sram_sp_rowtapend_replica VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_rowtapend_replica

.SUBCKT sram_sp_rowtapend_replica_wrapper VSS VNB

  X0 VSS VNB sram_sp_rowtapend_replica

.ENDS sram_sp_rowtapend_replica_wrapper

.SUBCKT nand2_1 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2_1

.SUBCKT decoder_stage_8 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] predecode_0_0 predecode_0_1 predecode_0_2 predecode_0_3 predecode_1_0 predecode_1_1 predecode_1_2 predecode_1_3

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_1
  Xgate_0_0_1 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_1
  Xgate_0_1_1 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_2 predecode_1_0 y_b[2] nand2_1
  Xgate_0_2_1 vdd vss predecode_0_2 predecode_1_0 y_b[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_3 predecode_1_0 y_b[3] nand2_1
  Xgate_0_3_1 vdd vss predecode_0_3 predecode_1_0 y_b[3] nand2_1
  Xgate_0_4_0 vdd vss predecode_0_0 predecode_1_1 y_b[4] nand2_1
  Xgate_0_4_1 vdd vss predecode_0_0 predecode_1_1 y_b[4] nand2_1
  Xgate_0_5_0 vdd vss predecode_0_1 predecode_1_1 y_b[5] nand2_1
  Xgate_0_5_1 vdd vss predecode_0_1 predecode_1_1 y_b[5] nand2_1
  Xgate_0_6_0 vdd vss predecode_0_2 predecode_1_1 y_b[6] nand2_1
  Xgate_0_6_1 vdd vss predecode_0_2 predecode_1_1 y_b[6] nand2_1
  Xgate_0_7_0 vdd vss predecode_0_3 predecode_1_1 y_b[7] nand2_1
  Xgate_0_7_1 vdd vss predecode_0_3 predecode_1_1 y_b[7] nand2_1
  Xgate_0_8_0 vdd vss predecode_0_0 predecode_1_2 y_b[8] nand2_1
  Xgate_0_8_1 vdd vss predecode_0_0 predecode_1_2 y_b[8] nand2_1
  Xgate_0_9_0 vdd vss predecode_0_1 predecode_1_2 y_b[9] nand2_1
  Xgate_0_9_1 vdd vss predecode_0_1 predecode_1_2 y_b[9] nand2_1
  Xgate_0_10_0 vdd vss predecode_0_2 predecode_1_2 y_b[10] nand2_1
  Xgate_0_10_1 vdd vss predecode_0_2 predecode_1_2 y_b[10] nand2_1
  Xgate_0_11_0 vdd vss predecode_0_3 predecode_1_2 y_b[11] nand2_1
  Xgate_0_11_1 vdd vss predecode_0_3 predecode_1_2 y_b[11] nand2_1
  Xgate_0_12_0 vdd vss predecode_0_0 predecode_1_3 y_b[12] nand2_1
  Xgate_0_12_1 vdd vss predecode_0_0 predecode_1_3 y_b[12] nand2_1
  Xgate_0_13_0 vdd vss predecode_0_1 predecode_1_3 y_b[13] nand2_1
  Xgate_0_13_1 vdd vss predecode_0_1 predecode_1_3 y_b[13] nand2_1
  Xgate_0_14_0 vdd vss predecode_0_2 predecode_1_3 y_b[14] nand2_1
  Xgate_0_14_1 vdd vss predecode_0_2 predecode_1_3 y_b[14] nand2_1
  Xgate_0_15_0 vdd vss predecode_0_3 predecode_1_3 y_b[15] nand2_1
  Xgate_0_15_1 vdd vss predecode_0_3 predecode_1_3 y_b[15] nand2_1
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_4
  Xgate_1_0_1 vdd vss y_b[0] y[0] folded_inv_4
  Xgate_1_0_2 vdd vss y_b[0] y[0] folded_inv_4
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_4
  Xgate_1_1_1 vdd vss y_b[1] y[1] folded_inv_4
  Xgate_1_1_2 vdd vss y_b[1] y[1] folded_inv_4
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_4
  Xgate_1_2_1 vdd vss y_b[2] y[2] folded_inv_4
  Xgate_1_2_2 vdd vss y_b[2] y[2] folded_inv_4
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_4
  Xgate_1_3_1 vdd vss y_b[3] y[3] folded_inv_4
  Xgate_1_3_2 vdd vss y_b[3] y[3] folded_inv_4
  Xgate_1_4_0 vdd vss y_b[4] y[4] folded_inv_4
  Xgate_1_4_1 vdd vss y_b[4] y[4] folded_inv_4
  Xgate_1_4_2 vdd vss y_b[4] y[4] folded_inv_4
  Xgate_1_5_0 vdd vss y_b[5] y[5] folded_inv_4
  Xgate_1_5_1 vdd vss y_b[5] y[5] folded_inv_4
  Xgate_1_5_2 vdd vss y_b[5] y[5] folded_inv_4
  Xgate_1_6_0 vdd vss y_b[6] y[6] folded_inv_4
  Xgate_1_6_1 vdd vss y_b[6] y[6] folded_inv_4
  Xgate_1_6_2 vdd vss y_b[6] y[6] folded_inv_4
  Xgate_1_7_0 vdd vss y_b[7] y[7] folded_inv_4
  Xgate_1_7_1 vdd vss y_b[7] y[7] folded_inv_4
  Xgate_1_7_2 vdd vss y_b[7] y[7] folded_inv_4
  Xgate_1_8_0 vdd vss y_b[8] y[8] folded_inv_4
  Xgate_1_8_1 vdd vss y_b[8] y[8] folded_inv_4
  Xgate_1_8_2 vdd vss y_b[8] y[8] folded_inv_4
  Xgate_1_9_0 vdd vss y_b[9] y[9] folded_inv_4
  Xgate_1_9_1 vdd vss y_b[9] y[9] folded_inv_4
  Xgate_1_9_2 vdd vss y_b[9] y[9] folded_inv_4
  Xgate_1_10_0 vdd vss y_b[10] y[10] folded_inv_4
  Xgate_1_10_1 vdd vss y_b[10] y[10] folded_inv_4
  Xgate_1_10_2 vdd vss y_b[10] y[10] folded_inv_4
  Xgate_1_11_0 vdd vss y_b[11] y[11] folded_inv_4
  Xgate_1_11_1 vdd vss y_b[11] y[11] folded_inv_4
  Xgate_1_11_2 vdd vss y_b[11] y[11] folded_inv_4
  Xgate_1_12_0 vdd vss y_b[12] y[12] folded_inv_4
  Xgate_1_12_1 vdd vss y_b[12] y[12] folded_inv_4
  Xgate_1_12_2 vdd vss y_b[12] y[12] folded_inv_4
  Xgate_1_13_0 vdd vss y_b[13] y[13] folded_inv_4
  Xgate_1_13_1 vdd vss y_b[13] y[13] folded_inv_4
  Xgate_1_13_2 vdd vss y_b[13] y[13] folded_inv_4
  Xgate_1_14_0 vdd vss y_b[14] y[14] folded_inv_4
  Xgate_1_14_1 vdd vss y_b[14] y[14] folded_inv_4
  Xgate_1_14_2 vdd vss y_b[14] y[14] folded_inv_4
  Xgate_1_15_0 vdd vss y_b[15] y[15] folded_inv_4
  Xgate_1_15_1 vdd vss y_b[15] y[15] folded_inv_4
  Xgate_1_15_2 vdd vss y_b[15] y[15] folded_inv_4

.ENDS decoder_stage_8

.SUBCKT inv_chain_3 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_3

.SUBCKT mos_w2530_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.530


.ENDS mos_w2530_l150_m1_nf1_id1

.SUBCKT mos_w1000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id0

.SUBCKT folded_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w2530_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1000_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2530_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1000_l150_m1_nf1_id0

.ENDS folded_inv_2

.SUBCKT decoder_stage_7 vdd vss y y_b predecode_0_0 predecode_1_0

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 x_0 nand2_1
  Xgate_1_0_0 vdd vss x_0 x_1 folded_inv_2
  Xgate_2_0_0 vdd vss x_1 y_b folded_inv_3
  Xgate_2_0_1 vdd vss x_1 y_b folded_inv_3
  Xgate_3_0_0 vdd vss y_b y folded_inv_3
  Xgate_3_0_1 vdd vss y_b y folded_inv_3

.ENDS decoder_stage_7

.SUBCKT sky130_fd_sc_hs__nand2_8_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_8

.ENDS sky130_fd_sc_hs__nand2_8_wrapper

.SUBCKT sr_latch sb rb q qb vdd vss

  Xnand_set q0b sb vss vss vdd vdd q0 sky130_fd_sc_hs__nand2_8_wrapper
  Xnand_reset q0 rb vss vss vdd vdd q0b sky130_fd_sc_hs__nand2_8_wrapper
  Xqb_inv q0 vss vss vdd vdd qb sky130_fd_sc_hs__inv_2_wrapper
  Xq_inv q0b vss vss vdd vdd q sky130_fd_sc_hs__inv_2_wrapper

.ENDS sr_latch

.SUBCKT column_mos_1 vdd vss bl

  Xdrain_nmos bl vss vss vss mos_w3100_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w4500_l150_m1_nf1_id1

.ENDS column_mos_1

.SUBCKT multi_finger_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_6

.SUBCKT decoder_stage_3 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_6
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_6

.ENDS decoder_stage_3

.SUBCKT mos_w9850_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=9.850


.ENDS mos_w9850_l150_m1_nf1_id0

.SUBCKT mos_w9850_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=9.850


.ENDS mos_w9850_l150_m1_nf1_id1

.SUBCKT tristate_inv din en en_b din_b vdd vss

  Xmn_en din_b en nint vss mos_w9850_l150_m1_nf1_id0
  Xmn_pd nint din vss vss mos_w9850_l150_m1_nf1_id0
  Xmp_en din_b en_b pint vdd mos_w9850_l150_m1_nf1_id1
  Xmp_pu pint din vdd vdd mos_w9850_l150_m1_nf1_id1

.ENDS tristate_inv

.SUBCKT write_driver en en_b data data_b bl br vdd vss

  Xbldriver data_b en en_b bl vdd vss tristate_inv
  Xbrdriver data en en_b br vdd vss tristate_inv

.ENDS write_driver

.SUBCKT mos_w3000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=3.000


.ENDS mos_w3000_l150_m1_nf1_id0

.SUBCKT replica_column_mos vdd vss bl

  Xunit0 vdd vss bl column_mos
  Xunit1 vdd vss bl column_mos_1
  Xunit2 vdd vss bl column_mos_1
  Xunit3 vdd vss bl column_mos_1
  Xunit4 vdd vss bl column_mos_1

.ENDS replica_column_mos

.SUBCKT mos_w13900_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=13.900


.ENDS mos_w13900_l150_m1_nf1_id1

.SUBCKT mos_w9250_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=9.250


.ENDS mos_w9250_l150_m1_nf1_id0

.SUBCKT tgate_mux sel_b sel bl br bl_out br_out vdd vss

  XMPBL bl_out sel_b bl vdd mos_w13900_l150_m1_nf1_id1
  XMPBR br_out sel_b br vdd mos_w13900_l150_m1_nf1_id1
  XMNBL bl_out sel bl vss mos_w9250_l150_m1_nf1_id0
  XMNBR br_out sel br vss mos_w9250_l150_m1_nf1_id0

.ENDS tgate_mux

.SUBCKT sramgen_sp_sense_amp_wrapper clk inn inp outn outp VDD VSS

  X0 clk inn inp outn outp VDD VSS sramgen_sp_sense_amp

.ENDS sramgen_sp_sense_amp_wrapper

.SUBCKT mos_w1000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id1

.SUBCKT mos_w600_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.600


.ENDS mos_w600_l150_m1_nf1_id0

.SUBCKT folded_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w600_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w600_l150_m1_nf1_id0

.ENDS folded_inv_6

.SUBCKT diff_latch vdd vss din1 din2 dout1 dout2

  Xinbuf_1 vdd vss din1 rst folded_inv_6
  Xinbuf_2 vdd vss din2 set folded_inv_6
  Xoutbuf_1 vdd vss q dout2 folded_inv_6
  Xoutbuf_2 vdd vss qb dout1 folded_inv_6
  Xinvq_1 vdd vss q qb folded_inv_6
  Xinvq_2 vdd vss qb q folded_inv_6
  XMN10 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN11 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN20 qb set vss vss mos_w1000_l150_m1_nf1_id0
  XMN21 qb set vss vss mos_w1000_l150_m1_nf1_id0

.ENDS diff_latch

.SUBCKT column clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we we_b din dout sense_en

  Xprecharge_0 vdd bl[0] br[0] pc_b precharge_1
  Xmux_0 sel_b[0] sel[0] bl[0] br[0] bl_out br_out vdd vss tgate_mux
  Xprecharge_1 vdd bl[1] br[1] pc_b precharge_1
  Xmux_1 sel_b[1] sel[1] bl[1] br[1] bl_out br_out vdd vss tgate_mux
  Xprecharge_2 vdd bl[2] br[2] pc_b precharge_1
  Xmux_2 sel_b[2] sel[2] bl[2] br[2] bl_out br_out vdd vss tgate_mux
  Xprecharge_3 vdd bl[3] br[3] pc_b precharge_1
  Xmux_3 sel_b[3] sel[3] bl[3] br[3] bl_out br_out vdd vss tgate_mux
  Xprecharge_4 vdd bl[4] br[4] pc_b precharge_1
  Xmux_4 sel_b[4] sel[4] bl[4] br[4] bl_out br_out vdd vss tgate_mux
  Xprecharge_5 vdd bl[5] br[5] pc_b precharge_1
  Xmux_5 sel_b[5] sel[5] bl[5] br[5] bl_out br_out vdd vss tgate_mux
  Xprecharge_6 vdd bl[6] br[6] pc_b precharge_1
  Xmux_6 sel_b[6] sel[6] bl[6] br[6] bl_out br_out vdd vss tgate_mux
  Xprecharge_7 vdd bl[7] br[7] pc_b precharge_1
  Xmux_7 sel_b[7] sel[7] bl[7] br[7] bl_out br_out vdd vss tgate_mux
  Xwrite_driver we we_b q q_b bl_out br_out vdd vss write_driver
  Xsense_amp sense_en br_out bl_out sa_outn sa_outp vdd vss sramgen_sp_sense_amp_wrapper
  Xlatch vdd vss sa_outp sa_outn dout diff_latch_outn diff_latch
  Xdff clk din rstb vss vss vdd vdd q q_b sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS column

.SUBCKT col_peripherals clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7]

  Xwmask_dffs vdd vss clk rstb wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask_in[0] wmask_in[1] wmask_in[2] wmask_in[3] wmask_in[4] wmask_in[5] wmask_in[6] wmask_in[7] wmask_in_b[0] wmask_in_b[1] wmask_in_b[2] wmask_in_b[3] wmask_in_b[4] wmask_in_b[5] wmask_in_b[6] wmask_in_b[7] dff_array_8
  Xwmask_and_0 vdd vss we_i[0] we_ib[0] we wmask_in[0] decoder_stage_7
  Xwmask_and_1 vdd vss we_i[1] we_ib[1] we wmask_in[1] decoder_stage_7
  Xwmask_and_2 vdd vss we_i[2] we_ib[2] we wmask_in[2] decoder_stage_7
  Xwmask_and_3 vdd vss we_i[3] we_ib[3] we wmask_in[3] decoder_stage_7
  Xwmask_and_4 vdd vss we_i[4] we_ib[4] we wmask_in[4] decoder_stage_7
  Xwmask_and_5 vdd vss we_i[5] we_ib[5] we wmask_in[5] decoder_stage_7
  Xwmask_and_6 vdd vss we_i[6] we_ib[6] we wmask_in[6] decoder_stage_7
  Xwmask_and_7 vdd vss we_i[7] we_ib[7] we wmask_in[7] decoder_stage_7
  Xcol_group_0 clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[0] we_ib[0] din[0] dout[0] sense_en column
  Xcol_group_1 clk rstb vdd vss bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[1] we_ib[1] din[1] dout[1] sense_en column
  Xcol_group_2 clk rstb vdd vss bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[2] we_ib[2] din[2] dout[2] sense_en column
  Xcol_group_3 clk rstb vdd vss bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[3] we_ib[3] din[3] dout[3] sense_en column
  Xcol_group_4 clk rstb vdd vss bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[4] we_ib[4] din[4] dout[4] sense_en column
  Xcol_group_5 clk rstb vdd vss bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[5] we_ib[5] din[5] dout[5] sense_en column
  Xcol_group_6 clk rstb vdd vss bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[6] we_ib[6] din[6] dout[6] sense_en column
  Xcol_group_7 clk rstb vdd vss bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] pc_b sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel_b[0] sel_b[1] sel_b[2] sel_b[3] sel_b[4] sel_b[5] sel_b[6] sel_b[7] we_i[7] we_ib[7] din[7] dout[7] sense_en column

.ENDS col_peripherals

.SUBCKT multi_finger_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_5

.SUBCKT decoder_stage_2 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_5
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_5

.ENDS decoder_stage_2

.SUBCKT nand3 vdd vss a b c y

  Xn1 x1 a vss vss mos_w3000_l150_m1_nf1_id0
  Xn2 x2 b x1 vss mos_w3000_l150_m1_nf1_id0
  Xn3 y c x2 vss mos_w3000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp3 y c vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand3

.SUBCKT multi_finger_inv_10 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_10

.SUBCKT multi_finger_inv_11 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_11

.SUBCKT multi_finger_inv_12 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_12

.SUBCKT multi_finger_inv_14 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_14

.SUBCKT decoder_stage_6 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_0 x_0[0] nand3
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_0 x_0[1] nand3
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_0 x_0[2] nand3
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_0 x_0[3] nand3
  Xgate_0_4_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_1 x_0[4] nand3
  Xgate_0_5_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_1 x_0[5] nand3
  Xgate_0_6_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_1 x_0[6] nand3
  Xgate_0_7_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_1 x_0[7] nand3
  Xgate_1_0_0 vdd vss x_0[0] x_1[0] multi_finger_inv_10
  Xgate_1_1_0 vdd vss x_0[1] x_1[1] multi_finger_inv_10
  Xgate_1_2_0 vdd vss x_0[2] x_1[2] multi_finger_inv_10
  Xgate_1_3_0 vdd vss x_0[3] x_1[3] multi_finger_inv_10
  Xgate_1_4_0 vdd vss x_0[4] x_1[4] multi_finger_inv_10
  Xgate_1_5_0 vdd vss x_0[5] x_1[5] multi_finger_inv_10
  Xgate_1_6_0 vdd vss x_0[6] x_1[6] multi_finger_inv_10
  Xgate_1_7_0 vdd vss x_0[7] x_1[7] multi_finger_inv_10
  Xgate_2_0_0 vdd vss x_1[0] x_2[0] multi_finger_inv_11
  Xgate_2_0_1 vdd vss x_1[0] x_2[0] multi_finger_inv_11
  Xgate_2_1_0 vdd vss x_1[1] x_2[1] multi_finger_inv_11
  Xgate_2_1_1 vdd vss x_1[1] x_2[1] multi_finger_inv_11
  Xgate_2_2_0 vdd vss x_1[2] x_2[2] multi_finger_inv_11
  Xgate_2_2_1 vdd vss x_1[2] x_2[2] multi_finger_inv_11
  Xgate_2_3_0 vdd vss x_1[3] x_2[3] multi_finger_inv_11
  Xgate_2_3_1 vdd vss x_1[3] x_2[3] multi_finger_inv_11
  Xgate_2_4_0 vdd vss x_1[4] x_2[4] multi_finger_inv_11
  Xgate_2_4_1 vdd vss x_1[4] x_2[4] multi_finger_inv_11
  Xgate_2_5_0 vdd vss x_1[5] x_2[5] multi_finger_inv_11
  Xgate_2_5_1 vdd vss x_1[5] x_2[5] multi_finger_inv_11
  Xgate_2_6_0 vdd vss x_1[6] x_2[6] multi_finger_inv_11
  Xgate_2_6_1 vdd vss x_1[6] x_2[6] multi_finger_inv_11
  Xgate_2_7_0 vdd vss x_1[7] x_2[7] multi_finger_inv_11
  Xgate_2_7_1 vdd vss x_1[7] x_2[7] multi_finger_inv_11
  Xgate_3_0_0 vdd vss x_2[0] x_3[0] multi_finger_inv_12
  Xgate_3_0_1 vdd vss x_2[0] x_3[0] multi_finger_inv_12
  Xgate_3_0_2 vdd vss x_2[0] x_3[0] multi_finger_inv_12
  Xgate_3_0_3 vdd vss x_2[0] x_3[0] multi_finger_inv_12
  Xgate_3_1_0 vdd vss x_2[1] x_3[1] multi_finger_inv_12
  Xgate_3_1_1 vdd vss x_2[1] x_3[1] multi_finger_inv_12
  Xgate_3_1_2 vdd vss x_2[1] x_3[1] multi_finger_inv_12
  Xgate_3_1_3 vdd vss x_2[1] x_3[1] multi_finger_inv_12
  Xgate_3_2_0 vdd vss x_2[2] x_3[2] multi_finger_inv_12
  Xgate_3_2_1 vdd vss x_2[2] x_3[2] multi_finger_inv_12
  Xgate_3_2_2 vdd vss x_2[2] x_3[2] multi_finger_inv_12
  Xgate_3_2_3 vdd vss x_2[2] x_3[2] multi_finger_inv_12
  Xgate_3_3_0 vdd vss x_2[3] x_3[3] multi_finger_inv_12
  Xgate_3_3_1 vdd vss x_2[3] x_3[3] multi_finger_inv_12
  Xgate_3_3_2 vdd vss x_2[3] x_3[3] multi_finger_inv_12
  Xgate_3_3_3 vdd vss x_2[3] x_3[3] multi_finger_inv_12
  Xgate_3_4_0 vdd vss x_2[4] x_3[4] multi_finger_inv_12
  Xgate_3_4_1 vdd vss x_2[4] x_3[4] multi_finger_inv_12
  Xgate_3_4_2 vdd vss x_2[4] x_3[4] multi_finger_inv_12
  Xgate_3_4_3 vdd vss x_2[4] x_3[4] multi_finger_inv_12
  Xgate_3_5_0 vdd vss x_2[5] x_3[5] multi_finger_inv_12
  Xgate_3_5_1 vdd vss x_2[5] x_3[5] multi_finger_inv_12
  Xgate_3_5_2 vdd vss x_2[5] x_3[5] multi_finger_inv_12
  Xgate_3_5_3 vdd vss x_2[5] x_3[5] multi_finger_inv_12
  Xgate_3_6_0 vdd vss x_2[6] x_3[6] multi_finger_inv_12
  Xgate_3_6_1 vdd vss x_2[6] x_3[6] multi_finger_inv_12
  Xgate_3_6_2 vdd vss x_2[6] x_3[6] multi_finger_inv_12
  Xgate_3_6_3 vdd vss x_2[6] x_3[6] multi_finger_inv_12
  Xgate_3_7_0 vdd vss x_2[7] x_3[7] multi_finger_inv_12
  Xgate_3_7_1 vdd vss x_2[7] x_3[7] multi_finger_inv_12
  Xgate_3_7_2 vdd vss x_2[7] x_3[7] multi_finger_inv_12
  Xgate_3_7_3 vdd vss x_2[7] x_3[7] multi_finger_inv_12
  Xgate_4_0_0 vdd vss x_3[0] y_b[0] multi_finger_inv_13
  Xgate_4_0_1 vdd vss x_3[0] y_b[0] multi_finger_inv_13
  Xgate_4_0_2 vdd vss x_3[0] y_b[0] multi_finger_inv_13
  Xgate_4_0_3 vdd vss x_3[0] y_b[0] multi_finger_inv_13
  Xgate_4_1_0 vdd vss x_3[1] y_b[1] multi_finger_inv_13
  Xgate_4_1_1 vdd vss x_3[1] y_b[1] multi_finger_inv_13
  Xgate_4_1_2 vdd vss x_3[1] y_b[1] multi_finger_inv_13
  Xgate_4_1_3 vdd vss x_3[1] y_b[1] multi_finger_inv_13
  Xgate_4_2_0 vdd vss x_3[2] y_b[2] multi_finger_inv_13
  Xgate_4_2_1 vdd vss x_3[2] y_b[2] multi_finger_inv_13
  Xgate_4_2_2 vdd vss x_3[2] y_b[2] multi_finger_inv_13
  Xgate_4_2_3 vdd vss x_3[2] y_b[2] multi_finger_inv_13
  Xgate_4_3_0 vdd vss x_3[3] y_b[3] multi_finger_inv_13
  Xgate_4_3_1 vdd vss x_3[3] y_b[3] multi_finger_inv_13
  Xgate_4_3_2 vdd vss x_3[3] y_b[3] multi_finger_inv_13
  Xgate_4_3_3 vdd vss x_3[3] y_b[3] multi_finger_inv_13
  Xgate_4_4_0 vdd vss x_3[4] y_b[4] multi_finger_inv_13
  Xgate_4_4_1 vdd vss x_3[4] y_b[4] multi_finger_inv_13
  Xgate_4_4_2 vdd vss x_3[4] y_b[4] multi_finger_inv_13
  Xgate_4_4_3 vdd vss x_3[4] y_b[4] multi_finger_inv_13
  Xgate_4_5_0 vdd vss x_3[5] y_b[5] multi_finger_inv_13
  Xgate_4_5_1 vdd vss x_3[5] y_b[5] multi_finger_inv_13
  Xgate_4_5_2 vdd vss x_3[5] y_b[5] multi_finger_inv_13
  Xgate_4_5_3 vdd vss x_3[5] y_b[5] multi_finger_inv_13
  Xgate_4_6_0 vdd vss x_3[6] y_b[6] multi_finger_inv_13
  Xgate_4_6_1 vdd vss x_3[6] y_b[6] multi_finger_inv_13
  Xgate_4_6_2 vdd vss x_3[6] y_b[6] multi_finger_inv_13
  Xgate_4_6_3 vdd vss x_3[6] y_b[6] multi_finger_inv_13
  Xgate_4_7_0 vdd vss x_3[7] y_b[7] multi_finger_inv_13
  Xgate_4_7_1 vdd vss x_3[7] y_b[7] multi_finger_inv_13
  Xgate_4_7_2 vdd vss x_3[7] y_b[7] multi_finger_inv_13
  Xgate_4_7_3 vdd vss x_3[7] y_b[7] multi_finger_inv_13
  Xgate_5_0_0 vdd vss y_b[0] y[0] multi_finger_inv_14
  Xgate_5_0_1 vdd vss y_b[0] y[0] multi_finger_inv_14
  Xgate_5_0_2 vdd vss y_b[0] y[0] multi_finger_inv_14
  Xgate_5_0_3 vdd vss y_b[0] y[0] multi_finger_inv_14
  Xgate_5_1_0 vdd vss y_b[1] y[1] multi_finger_inv_14
  Xgate_5_1_1 vdd vss y_b[1] y[1] multi_finger_inv_14
  Xgate_5_1_2 vdd vss y_b[1] y[1] multi_finger_inv_14
  Xgate_5_1_3 vdd vss y_b[1] y[1] multi_finger_inv_14
  Xgate_5_2_0 vdd vss y_b[2] y[2] multi_finger_inv_14
  Xgate_5_2_1 vdd vss y_b[2] y[2] multi_finger_inv_14
  Xgate_5_2_2 vdd vss y_b[2] y[2] multi_finger_inv_14
  Xgate_5_2_3 vdd vss y_b[2] y[2] multi_finger_inv_14
  Xgate_5_3_0 vdd vss y_b[3] y[3] multi_finger_inv_14
  Xgate_5_3_1 vdd vss y_b[3] y[3] multi_finger_inv_14
  Xgate_5_3_2 vdd vss y_b[3] y[3] multi_finger_inv_14
  Xgate_5_3_3 vdd vss y_b[3] y[3] multi_finger_inv_14
  Xgate_5_4_0 vdd vss y_b[4] y[4] multi_finger_inv_14
  Xgate_5_4_1 vdd vss y_b[4] y[4] multi_finger_inv_14
  Xgate_5_4_2 vdd vss y_b[4] y[4] multi_finger_inv_14
  Xgate_5_4_3 vdd vss y_b[4] y[4] multi_finger_inv_14
  Xgate_5_5_0 vdd vss y_b[5] y[5] multi_finger_inv_14
  Xgate_5_5_1 vdd vss y_b[5] y[5] multi_finger_inv_14
  Xgate_5_5_2 vdd vss y_b[5] y[5] multi_finger_inv_14
  Xgate_5_5_3 vdd vss y_b[5] y[5] multi_finger_inv_14
  Xgate_5_6_0 vdd vss y_b[6] y[6] multi_finger_inv_14
  Xgate_5_6_1 vdd vss y_b[6] y[6] multi_finger_inv_14
  Xgate_5_6_2 vdd vss y_b[6] y[6] multi_finger_inv_14
  Xgate_5_6_3 vdd vss y_b[6] y[6] multi_finger_inv_14
  Xgate_5_7_0 vdd vss y_b[7] y[7] multi_finger_inv_14
  Xgate_5_7_1 vdd vss y_b[7] y[7] multi_finger_inv_14
  Xgate_5_7_2 vdd vss y_b[7] y[7] multi_finger_inv_14
  Xgate_5_7_3 vdd vss y_b[7] y[7] multi_finger_inv_14

.ENDS decoder_stage_6

.SUBCKT sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X18 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__inv_16

.SUBCKT sky130_fd_sc_hs__inv_16_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_16

.ENDS sky130_fd_sc_hs__inv_16_wrapper

.SUBCKT inv_chain_12 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_12

.SUBCKT sky130_fd_sc_hs__and2_2_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_2

.ENDS sky130_fd_sc_hs__and2_2_wrapper

.SUBCKT sky130_fd_sc_hs__buf_16 A VGND VNB VPB VPWR X

  X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X9 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X19 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X24 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X27 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X32 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X33 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X35 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X36 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X38 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X39 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X40 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X41 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X42 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X43 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__buf_16

.SUBCKT sky130_fd_sc_hs__buf_16_wrapper A VGND VNB VPB VPWR X

  X0 A VGND VNB VPB VPWR X sky130_fd_sc_hs__buf_16

.ENDS sky130_fd_sc_hs__buf_16_wrapper

.SUBCKT inv_chain_15 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sky130_fd_sc_hs__inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_15

.SUBCKT sky130_fd_sc_hs__mux2_4 A0 A1 S VGND VNB VPB VPWR X

  X0 a_27_368# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 a_722_391# A0 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X2 a_722_391# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X3 VGND a_27_368# a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_193_241# A1 a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X5 a_709_119# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 a_709_119# A1 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X7 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VPWR a_27_368# a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_193_241# A0 a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X12 a_937_119# A0 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_936_391# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X14 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VPWR S a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X17 a_936_391# A1 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X18 a_193_241# A0 a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X19 a_193_241# A1 a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X20 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X21 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X22 a_27_368# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X23 a_937_119# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X24 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND S a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640


.ENDS sky130_fd_sc_hs__mux2_4

.SUBCKT sky130_fd_sc_hs__mux2_4_wrapper A0 A1 S VGND VNB VPB VPWR X

  X0 A0 A1 S VGND VNB VPB VPWR X sky130_fd_sc_hs__mux2_4

.ENDS sky130_fd_sc_hs__mux2_4_wrapper

.SUBCKT inv_chain_14 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_14

.SUBCKT sky130_fd_sc_hs__nor2_4 A B VGND VNB VPB VPWR Y

  X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nor2_4

.SUBCKT sky130_fd_sc_hs__nor2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nor2_4

.ENDS sky130_fd_sc_hs__nor2_4_wrapper

.SUBCKT sky130_fd_sc_hs__nand2_4 A B VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__nand2_4

.SUBCKT sky130_fd_sc_hs__nand2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_4

.ENDS sky130_fd_sc_hs__nand2_4_wrapper

.SUBCKT inv_chain_2 din dout vdd vss

  Xinv0 din vss vss vdd vdd x sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_2

.SUBCKT control_logic_replica_v2 clk ce we rstb rbl saen pc_b rwl wlen wrdrven vdd vss

  Xreset_inv rstb vss vss vdd vdd reset sky130_fd_sc_hs__inv_16_wrapper
  Xclk_delay clk clkd vdd vss inv_chain_12
  Xclk_gate clkd ce vss vss vdd vdd clk_buf sky130_fd_sc_hs__and2_2_wrapper
  Xclk_pulse clk_buf clkp0 vdd vss edge_detector
  Xclk_pulse_buf clkp0 vss vss vdd vdd clkp sky130_fd_sc_hs__buf_16_wrapper
  Xclk_pulse_inv clkp vss vss vdd vdd clkp_b sky130_fd_sc_hs__inv_16_wrapper
  Xclkp_delay clkp_b clkpd vdd vss inv_chain_3
  Xclkpd_inv clkpd vss vss vdd vdd clkpd_b sky130_fd_sc_hs__inv_2_wrapper
  Xclkpd_delay clkpd_b clkpdd vdd vss inv_chain_15
  Xmux_wlen_rst rbl_b clkpdd we vss vss vdd vdd decrepstart sky130_fd_sc_hs__mux2_4_wrapper
  Xdecoder_replica decrepstart decrepend vdd vss svt_inv_chain_30
  Xdecoder_replica_delay decrepend wlen_rst_decoderd vdd vss inv_chain_14
  Xinv_we we vss vss vdd vdd we_b sky130_fd_sc_hs__inv_2_wrapper
  Xinv_rbl rbl vss vss vdd vdd rbl_b sky130_fd_sc_hs__inv_2_wrapper
  Xwlen_grst decrepstart reset vss vss vdd vdd wlen_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xpc_set wlen_rst_decoderd reset vss vss vdd vdd pc_set_b sky130_fd_sc_hs__nor2_4_wrapper
  Xwrdrven_grst decrepend reset vss vss vdd vdd wrdrven_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xclkp_grst clkp reset vss vss vdd vdd clkp_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xnand_sense_en we_b decrepend vss vss vdd vdd saen_set_b sky130_fd_sc_hs__nand2_4_wrapper
  Xnand_wlendb_web rbl_b we_b vss vss vdd vdd wlend sky130_fd_sc_hs__nand2_4_wrapper
  Xand_wlen wlen_q wlend vss vss vdd vdd wlen sky130_fd_sc_hs__and2_4_wrapper
  Xrwl_buf wlen_q vss vss vdd vdd rwl sky130_fd_sc_hs__buf_16_wrapper
  Xwl_ctl clkpd_b wlen_grst_b wlen_q wlen_b vdd vss sr_latch
  Xsaen_ctl saen_set_b clkp_grst_b saen saen_b vdd vss sr_latch
  Xpc_ctl pc_set_b clkp_b pc pc_b0 vdd vss sr_latch
  Xpc_b_buf pc_b0 vss vss vdd vdd pc_b sky130_fd_sc_hs__buf_16_wrapper
  Xwrdrven_set clkpd we vss vss vdd vdd wrdrven_set_b0 sky130_fd_sc_hs__nand2_4_wrapper
  Xwrdrven_set_delay wrdrven_set_b0 wrdrven_set_b vdd vss inv_chain_2
  Xwrdrven_ctl wrdrven_set_b wrdrven_grst_b wrdrven wrdrven_b vdd vss sr_latch

.ENDS control_logic_replica_v2

.SUBCKT mos_w3800_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.800


.ENDS mos_w3800_l150_m1_nf1_id1

.SUBCKT mos_w1530_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.530


.ENDS mos_w1530_l150_m1_nf1_id0

.SUBCKT folded_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w3800_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1530_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w3800_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1530_l150_m1_nf1_id0

.ENDS folded_inv_7

.SUBCKT decoder_stage_9 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 y_b[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 y_b[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 y_b[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 y_b[3] nand2_1
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_7
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_7
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_7
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_7

.ENDS decoder_stage_9

.SUBCKT decoder_3 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  X0 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_stage_9

.ENDS decoder_3

.SUBCKT decoder_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1

  X0 vdd vss child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_noconn_0[0] child_noconn_0[1] child_noconn_0[2] child_noconn_0[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_3
  X0_1 vdd vss child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_noconn_1[0] child_noconn_1[1] child_noconn_1[2] child_noconn_1[3] predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 decoder_3
  X0_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] decoder_stage_8

.ENDS decoder_2

.SUBCKT mos_w2800_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.800


.ENDS mos_w2800_l150_m1_nf1_id1

.SUBCKT mos_w1130_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.130


.ENDS mos_w1130_l150_m1_nf1_id0

.SUBCKT folded_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w2800_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1130_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2800_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1130_l150_m1_nf1_id0

.ENDS folded_inv_5

.SUBCKT and2_1 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_5

.ENDS and2_1

.SUBCKT multi_finger_inv_9 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_9

.SUBCKT decoder_stage_5 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y[128] y[129] y[130] y[131] y[132] y[133] y[134] y[135] y[136] y[137] y[138] y[139] y[140] y[141] y[142] y[143] y[144] y[145] y[146] y[147] y[148] y[149] y[150] y[151] y[152] y[153] y[154] y[155] y[156] y[157] y[158] y[159] y[160] y[161] y[162] y[163] y[164] y[165] y[166] y[167] y[168] y[169] y[170] y[171] y[172] y[173] y[174] y[175] y[176] y[177] y[178] y[179] y[180] y[181] y[182] y[183] y[184] y[185] y[186] y[187] y[188] y[189] y[190] y[191] y[192] y[193] y[194] y[195] y[196] y[197] y[198] y[199] y[200] y[201] y[202] y[203] y[204] y[205] y[206] y[207] y[208] y[209] y[210] y[211] y[212] y[213] y[214] y[215] y[216] y[217] y[218] y[219] y[220] y[221] y[222] y[223] y[224] y[225] y[226] y[227] y[228] y[229] y[230] y[231] y[232] y[233] y[234] y[235] y[236] y[237] y[238] y[239] y[240] y[241] y[242] y[243] y[244] y[245] y[246] y[247] y[248] y[249] y[250] y[251] y[252] y[253] y[254] y[255] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] y_b[128] y_b[129] y_b[130] y_b[131] y_b[132] y_b[133] y_b[134] y_b[135] y_b[136] y_b[137] y_b[138] y_b[139] y_b[140] y_b[141] y_b[142] y_b[143] y_b[144] y_b[145] y_b[146] y_b[147] y_b[148] y_b[149] y_b[150] y_b[151] y_b[152] y_b[153] y_b[154] y_b[155] y_b[156] y_b[157] y_b[158] y_b[159] y_b[160] y_b[161] y_b[162] y_b[163] y_b[164] y_b[165] y_b[166] y_b[167] y_b[168] y_b[169] y_b[170] y_b[171] y_b[172] y_b[173] y_b[174] y_b[175] y_b[176] y_b[177] y_b[178] y_b[179] y_b[180] y_b[181] y_b[182] y_b[183] y_b[184] y_b[185] y_b[186] y_b[187] y_b[188] y_b[189] y_b[190] y_b[191] y_b[192] y_b[193] y_b[194] y_b[195] y_b[196] y_b[197] y_b[198] y_b[199] y_b[200] y_b[201] y_b[202] y_b[203] y_b[204] y_b[205] y_b[206] y_b[207] y_b[208] y_b[209] y_b[210] y_b[211] y_b[212] y_b[213] y_b[214] y_b[215] y_b[216] y_b[217] y_b[218] y_b[219] y_b[220] y_b[221] y_b[222] y_b[223] y_b[224] y_b[225] y_b[226] y_b[227] y_b[228] y_b[229] y_b[230] y_b[231] y_b[232] y_b[233] y_b[234] y_b[235] y_b[236] y_b[237] y_b[238] y_b[239] y_b[240] y_b[241] y_b[242] y_b[243] y_b[244] y_b[245] y_b[246] y_b[247] y_b[248] y_b[249] y_b[250] y_b[251] y_b[252] y_b[253] y_b[254] y_b[255] predecode_0_0 predecode_0_1 predecode_0_2 predecode_0_3 predecode_0_4 predecode_0_5 predecode_0_6 predecode_0_7 predecode_0_8 predecode_0_9 predecode_0_10 predecode_0_11 predecode_0_12 predecode_0_13 predecode_0_14 predecode_0_15 predecode_1_0 predecode_1_1 predecode_1_2 predecode_1_3 predecode_1_4 predecode_1_5 predecode_1_6 predecode_1_7 predecode_1_8 predecode_1_9 predecode_1_10 predecode_1_11 predecode_1_12 predecode_1_13 predecode_1_14 predecode_1_15

  Xgate_0_0_0 vdd predecode_0_0 predecode_1_0 x_0[0] y_b_noconn_0_0_0 vss and2_1
  Xgate_0_1_0 vdd predecode_0_1 predecode_1_0 x_0[1] y_b_noconn_0_1_0 vss and2_1
  Xgate_0_2_0 vdd predecode_0_2 predecode_1_0 x_0[2] y_b_noconn_0_2_0 vss and2_1
  Xgate_0_3_0 vdd predecode_0_3 predecode_1_0 x_0[3] y_b_noconn_0_3_0 vss and2_1
  Xgate_0_4_0 vdd predecode_0_4 predecode_1_0 x_0[4] y_b_noconn_0_4_0 vss and2_1
  Xgate_0_5_0 vdd predecode_0_5 predecode_1_0 x_0[5] y_b_noconn_0_5_0 vss and2_1
  Xgate_0_6_0 vdd predecode_0_6 predecode_1_0 x_0[6] y_b_noconn_0_6_0 vss and2_1
  Xgate_0_7_0 vdd predecode_0_7 predecode_1_0 x_0[7] y_b_noconn_0_7_0 vss and2_1
  Xgate_0_8_0 vdd predecode_0_8 predecode_1_0 x_0[8] y_b_noconn_0_8_0 vss and2_1
  Xgate_0_9_0 vdd predecode_0_9 predecode_1_0 x_0[9] y_b_noconn_0_9_0 vss and2_1
  Xgate_0_10_0 vdd predecode_0_10 predecode_1_0 x_0[10] y_b_noconn_0_10_0 vss and2_1
  Xgate_0_11_0 vdd predecode_0_11 predecode_1_0 x_0[11] y_b_noconn_0_11_0 vss and2_1
  Xgate_0_12_0 vdd predecode_0_12 predecode_1_0 x_0[12] y_b_noconn_0_12_0 vss and2_1
  Xgate_0_13_0 vdd predecode_0_13 predecode_1_0 x_0[13] y_b_noconn_0_13_0 vss and2_1
  Xgate_0_14_0 vdd predecode_0_14 predecode_1_0 x_0[14] y_b_noconn_0_14_0 vss and2_1
  Xgate_0_15_0 vdd predecode_0_15 predecode_1_0 x_0[15] y_b_noconn_0_15_0 vss and2_1
  Xgate_0_16_0 vdd predecode_0_0 predecode_1_1 x_0[16] y_b_noconn_0_16_0 vss and2_1
  Xgate_0_17_0 vdd predecode_0_1 predecode_1_1 x_0[17] y_b_noconn_0_17_0 vss and2_1
  Xgate_0_18_0 vdd predecode_0_2 predecode_1_1 x_0[18] y_b_noconn_0_18_0 vss and2_1
  Xgate_0_19_0 vdd predecode_0_3 predecode_1_1 x_0[19] y_b_noconn_0_19_0 vss and2_1
  Xgate_0_20_0 vdd predecode_0_4 predecode_1_1 x_0[20] y_b_noconn_0_20_0 vss and2_1
  Xgate_0_21_0 vdd predecode_0_5 predecode_1_1 x_0[21] y_b_noconn_0_21_0 vss and2_1
  Xgate_0_22_0 vdd predecode_0_6 predecode_1_1 x_0[22] y_b_noconn_0_22_0 vss and2_1
  Xgate_0_23_0 vdd predecode_0_7 predecode_1_1 x_0[23] y_b_noconn_0_23_0 vss and2_1
  Xgate_0_24_0 vdd predecode_0_8 predecode_1_1 x_0[24] y_b_noconn_0_24_0 vss and2_1
  Xgate_0_25_0 vdd predecode_0_9 predecode_1_1 x_0[25] y_b_noconn_0_25_0 vss and2_1
  Xgate_0_26_0 vdd predecode_0_10 predecode_1_1 x_0[26] y_b_noconn_0_26_0 vss and2_1
  Xgate_0_27_0 vdd predecode_0_11 predecode_1_1 x_0[27] y_b_noconn_0_27_0 vss and2_1
  Xgate_0_28_0 vdd predecode_0_12 predecode_1_1 x_0[28] y_b_noconn_0_28_0 vss and2_1
  Xgate_0_29_0 vdd predecode_0_13 predecode_1_1 x_0[29] y_b_noconn_0_29_0 vss and2_1
  Xgate_0_30_0 vdd predecode_0_14 predecode_1_1 x_0[30] y_b_noconn_0_30_0 vss and2_1
  Xgate_0_31_0 vdd predecode_0_15 predecode_1_1 x_0[31] y_b_noconn_0_31_0 vss and2_1
  Xgate_0_32_0 vdd predecode_0_0 predecode_1_2 x_0[32] y_b_noconn_0_32_0 vss and2_1
  Xgate_0_33_0 vdd predecode_0_1 predecode_1_2 x_0[33] y_b_noconn_0_33_0 vss and2_1
  Xgate_0_34_0 vdd predecode_0_2 predecode_1_2 x_0[34] y_b_noconn_0_34_0 vss and2_1
  Xgate_0_35_0 vdd predecode_0_3 predecode_1_2 x_0[35] y_b_noconn_0_35_0 vss and2_1
  Xgate_0_36_0 vdd predecode_0_4 predecode_1_2 x_0[36] y_b_noconn_0_36_0 vss and2_1
  Xgate_0_37_0 vdd predecode_0_5 predecode_1_2 x_0[37] y_b_noconn_0_37_0 vss and2_1
  Xgate_0_38_0 vdd predecode_0_6 predecode_1_2 x_0[38] y_b_noconn_0_38_0 vss and2_1
  Xgate_0_39_0 vdd predecode_0_7 predecode_1_2 x_0[39] y_b_noconn_0_39_0 vss and2_1
  Xgate_0_40_0 vdd predecode_0_8 predecode_1_2 x_0[40] y_b_noconn_0_40_0 vss and2_1
  Xgate_0_41_0 vdd predecode_0_9 predecode_1_2 x_0[41] y_b_noconn_0_41_0 vss and2_1
  Xgate_0_42_0 vdd predecode_0_10 predecode_1_2 x_0[42] y_b_noconn_0_42_0 vss and2_1
  Xgate_0_43_0 vdd predecode_0_11 predecode_1_2 x_0[43] y_b_noconn_0_43_0 vss and2_1
  Xgate_0_44_0 vdd predecode_0_12 predecode_1_2 x_0[44] y_b_noconn_0_44_0 vss and2_1
  Xgate_0_45_0 vdd predecode_0_13 predecode_1_2 x_0[45] y_b_noconn_0_45_0 vss and2_1
  Xgate_0_46_0 vdd predecode_0_14 predecode_1_2 x_0[46] y_b_noconn_0_46_0 vss and2_1
  Xgate_0_47_0 vdd predecode_0_15 predecode_1_2 x_0[47] y_b_noconn_0_47_0 vss and2_1
  Xgate_0_48_0 vdd predecode_0_0 predecode_1_3 x_0[48] y_b_noconn_0_48_0 vss and2_1
  Xgate_0_49_0 vdd predecode_0_1 predecode_1_3 x_0[49] y_b_noconn_0_49_0 vss and2_1
  Xgate_0_50_0 vdd predecode_0_2 predecode_1_3 x_0[50] y_b_noconn_0_50_0 vss and2_1
  Xgate_0_51_0 vdd predecode_0_3 predecode_1_3 x_0[51] y_b_noconn_0_51_0 vss and2_1
  Xgate_0_52_0 vdd predecode_0_4 predecode_1_3 x_0[52] y_b_noconn_0_52_0 vss and2_1
  Xgate_0_53_0 vdd predecode_0_5 predecode_1_3 x_0[53] y_b_noconn_0_53_0 vss and2_1
  Xgate_0_54_0 vdd predecode_0_6 predecode_1_3 x_0[54] y_b_noconn_0_54_0 vss and2_1
  Xgate_0_55_0 vdd predecode_0_7 predecode_1_3 x_0[55] y_b_noconn_0_55_0 vss and2_1
  Xgate_0_56_0 vdd predecode_0_8 predecode_1_3 x_0[56] y_b_noconn_0_56_0 vss and2_1
  Xgate_0_57_0 vdd predecode_0_9 predecode_1_3 x_0[57] y_b_noconn_0_57_0 vss and2_1
  Xgate_0_58_0 vdd predecode_0_10 predecode_1_3 x_0[58] y_b_noconn_0_58_0 vss and2_1
  Xgate_0_59_0 vdd predecode_0_11 predecode_1_3 x_0[59] y_b_noconn_0_59_0 vss and2_1
  Xgate_0_60_0 vdd predecode_0_12 predecode_1_3 x_0[60] y_b_noconn_0_60_0 vss and2_1
  Xgate_0_61_0 vdd predecode_0_13 predecode_1_3 x_0[61] y_b_noconn_0_61_0 vss and2_1
  Xgate_0_62_0 vdd predecode_0_14 predecode_1_3 x_0[62] y_b_noconn_0_62_0 vss and2_1
  Xgate_0_63_0 vdd predecode_0_15 predecode_1_3 x_0[63] y_b_noconn_0_63_0 vss and2_1
  Xgate_0_64_0 vdd predecode_0_0 predecode_1_4 x_0[64] y_b_noconn_0_64_0 vss and2_1
  Xgate_0_65_0 vdd predecode_0_1 predecode_1_4 x_0[65] y_b_noconn_0_65_0 vss and2_1
  Xgate_0_66_0 vdd predecode_0_2 predecode_1_4 x_0[66] y_b_noconn_0_66_0 vss and2_1
  Xgate_0_67_0 vdd predecode_0_3 predecode_1_4 x_0[67] y_b_noconn_0_67_0 vss and2_1
  Xgate_0_68_0 vdd predecode_0_4 predecode_1_4 x_0[68] y_b_noconn_0_68_0 vss and2_1
  Xgate_0_69_0 vdd predecode_0_5 predecode_1_4 x_0[69] y_b_noconn_0_69_0 vss and2_1
  Xgate_0_70_0 vdd predecode_0_6 predecode_1_4 x_0[70] y_b_noconn_0_70_0 vss and2_1
  Xgate_0_71_0 vdd predecode_0_7 predecode_1_4 x_0[71] y_b_noconn_0_71_0 vss and2_1
  Xgate_0_72_0 vdd predecode_0_8 predecode_1_4 x_0[72] y_b_noconn_0_72_0 vss and2_1
  Xgate_0_73_0 vdd predecode_0_9 predecode_1_4 x_0[73] y_b_noconn_0_73_0 vss and2_1
  Xgate_0_74_0 vdd predecode_0_10 predecode_1_4 x_0[74] y_b_noconn_0_74_0 vss and2_1
  Xgate_0_75_0 vdd predecode_0_11 predecode_1_4 x_0[75] y_b_noconn_0_75_0 vss and2_1
  Xgate_0_76_0 vdd predecode_0_12 predecode_1_4 x_0[76] y_b_noconn_0_76_0 vss and2_1
  Xgate_0_77_0 vdd predecode_0_13 predecode_1_4 x_0[77] y_b_noconn_0_77_0 vss and2_1
  Xgate_0_78_0 vdd predecode_0_14 predecode_1_4 x_0[78] y_b_noconn_0_78_0 vss and2_1
  Xgate_0_79_0 vdd predecode_0_15 predecode_1_4 x_0[79] y_b_noconn_0_79_0 vss and2_1
  Xgate_0_80_0 vdd predecode_0_0 predecode_1_5 x_0[80] y_b_noconn_0_80_0 vss and2_1
  Xgate_0_81_0 vdd predecode_0_1 predecode_1_5 x_0[81] y_b_noconn_0_81_0 vss and2_1
  Xgate_0_82_0 vdd predecode_0_2 predecode_1_5 x_0[82] y_b_noconn_0_82_0 vss and2_1
  Xgate_0_83_0 vdd predecode_0_3 predecode_1_5 x_0[83] y_b_noconn_0_83_0 vss and2_1
  Xgate_0_84_0 vdd predecode_0_4 predecode_1_5 x_0[84] y_b_noconn_0_84_0 vss and2_1
  Xgate_0_85_0 vdd predecode_0_5 predecode_1_5 x_0[85] y_b_noconn_0_85_0 vss and2_1
  Xgate_0_86_0 vdd predecode_0_6 predecode_1_5 x_0[86] y_b_noconn_0_86_0 vss and2_1
  Xgate_0_87_0 vdd predecode_0_7 predecode_1_5 x_0[87] y_b_noconn_0_87_0 vss and2_1
  Xgate_0_88_0 vdd predecode_0_8 predecode_1_5 x_0[88] y_b_noconn_0_88_0 vss and2_1
  Xgate_0_89_0 vdd predecode_0_9 predecode_1_5 x_0[89] y_b_noconn_0_89_0 vss and2_1
  Xgate_0_90_0 vdd predecode_0_10 predecode_1_5 x_0[90] y_b_noconn_0_90_0 vss and2_1
  Xgate_0_91_0 vdd predecode_0_11 predecode_1_5 x_0[91] y_b_noconn_0_91_0 vss and2_1
  Xgate_0_92_0 vdd predecode_0_12 predecode_1_5 x_0[92] y_b_noconn_0_92_0 vss and2_1
  Xgate_0_93_0 vdd predecode_0_13 predecode_1_5 x_0[93] y_b_noconn_0_93_0 vss and2_1
  Xgate_0_94_0 vdd predecode_0_14 predecode_1_5 x_0[94] y_b_noconn_0_94_0 vss and2_1
  Xgate_0_95_0 vdd predecode_0_15 predecode_1_5 x_0[95] y_b_noconn_0_95_0 vss and2_1
  Xgate_0_96_0 vdd predecode_0_0 predecode_1_6 x_0[96] y_b_noconn_0_96_0 vss and2_1
  Xgate_0_97_0 vdd predecode_0_1 predecode_1_6 x_0[97] y_b_noconn_0_97_0 vss and2_1
  Xgate_0_98_0 vdd predecode_0_2 predecode_1_6 x_0[98] y_b_noconn_0_98_0 vss and2_1
  Xgate_0_99_0 vdd predecode_0_3 predecode_1_6 x_0[99] y_b_noconn_0_99_0 vss and2_1
  Xgate_0_100_0 vdd predecode_0_4 predecode_1_6 x_0[100] y_b_noconn_0_100_0 vss and2_1
  Xgate_0_101_0 vdd predecode_0_5 predecode_1_6 x_0[101] y_b_noconn_0_101_0 vss and2_1
  Xgate_0_102_0 vdd predecode_0_6 predecode_1_6 x_0[102] y_b_noconn_0_102_0 vss and2_1
  Xgate_0_103_0 vdd predecode_0_7 predecode_1_6 x_0[103] y_b_noconn_0_103_0 vss and2_1
  Xgate_0_104_0 vdd predecode_0_8 predecode_1_6 x_0[104] y_b_noconn_0_104_0 vss and2_1
  Xgate_0_105_0 vdd predecode_0_9 predecode_1_6 x_0[105] y_b_noconn_0_105_0 vss and2_1
  Xgate_0_106_0 vdd predecode_0_10 predecode_1_6 x_0[106] y_b_noconn_0_106_0 vss and2_1
  Xgate_0_107_0 vdd predecode_0_11 predecode_1_6 x_0[107] y_b_noconn_0_107_0 vss and2_1
  Xgate_0_108_0 vdd predecode_0_12 predecode_1_6 x_0[108] y_b_noconn_0_108_0 vss and2_1
  Xgate_0_109_0 vdd predecode_0_13 predecode_1_6 x_0[109] y_b_noconn_0_109_0 vss and2_1
  Xgate_0_110_0 vdd predecode_0_14 predecode_1_6 x_0[110] y_b_noconn_0_110_0 vss and2_1
  Xgate_0_111_0 vdd predecode_0_15 predecode_1_6 x_0[111] y_b_noconn_0_111_0 vss and2_1
  Xgate_0_112_0 vdd predecode_0_0 predecode_1_7 x_0[112] y_b_noconn_0_112_0 vss and2_1
  Xgate_0_113_0 vdd predecode_0_1 predecode_1_7 x_0[113] y_b_noconn_0_113_0 vss and2_1
  Xgate_0_114_0 vdd predecode_0_2 predecode_1_7 x_0[114] y_b_noconn_0_114_0 vss and2_1
  Xgate_0_115_0 vdd predecode_0_3 predecode_1_7 x_0[115] y_b_noconn_0_115_0 vss and2_1
  Xgate_0_116_0 vdd predecode_0_4 predecode_1_7 x_0[116] y_b_noconn_0_116_0 vss and2_1
  Xgate_0_117_0 vdd predecode_0_5 predecode_1_7 x_0[117] y_b_noconn_0_117_0 vss and2_1
  Xgate_0_118_0 vdd predecode_0_6 predecode_1_7 x_0[118] y_b_noconn_0_118_0 vss and2_1
  Xgate_0_119_0 vdd predecode_0_7 predecode_1_7 x_0[119] y_b_noconn_0_119_0 vss and2_1
  Xgate_0_120_0 vdd predecode_0_8 predecode_1_7 x_0[120] y_b_noconn_0_120_0 vss and2_1
  Xgate_0_121_0 vdd predecode_0_9 predecode_1_7 x_0[121] y_b_noconn_0_121_0 vss and2_1
  Xgate_0_122_0 vdd predecode_0_10 predecode_1_7 x_0[122] y_b_noconn_0_122_0 vss and2_1
  Xgate_0_123_0 vdd predecode_0_11 predecode_1_7 x_0[123] y_b_noconn_0_123_0 vss and2_1
  Xgate_0_124_0 vdd predecode_0_12 predecode_1_7 x_0[124] y_b_noconn_0_124_0 vss and2_1
  Xgate_0_125_0 vdd predecode_0_13 predecode_1_7 x_0[125] y_b_noconn_0_125_0 vss and2_1
  Xgate_0_126_0 vdd predecode_0_14 predecode_1_7 x_0[126] y_b_noconn_0_126_0 vss and2_1
  Xgate_0_127_0 vdd predecode_0_15 predecode_1_7 x_0[127] y_b_noconn_0_127_0 vss and2_1
  Xgate_0_128_0 vdd predecode_0_0 predecode_1_8 x_0[128] y_b_noconn_0_128_0 vss and2_1
  Xgate_0_129_0 vdd predecode_0_1 predecode_1_8 x_0[129] y_b_noconn_0_129_0 vss and2_1
  Xgate_0_130_0 vdd predecode_0_2 predecode_1_8 x_0[130] y_b_noconn_0_130_0 vss and2_1
  Xgate_0_131_0 vdd predecode_0_3 predecode_1_8 x_0[131] y_b_noconn_0_131_0 vss and2_1
  Xgate_0_132_0 vdd predecode_0_4 predecode_1_8 x_0[132] y_b_noconn_0_132_0 vss and2_1
  Xgate_0_133_0 vdd predecode_0_5 predecode_1_8 x_0[133] y_b_noconn_0_133_0 vss and2_1
  Xgate_0_134_0 vdd predecode_0_6 predecode_1_8 x_0[134] y_b_noconn_0_134_0 vss and2_1
  Xgate_0_135_0 vdd predecode_0_7 predecode_1_8 x_0[135] y_b_noconn_0_135_0 vss and2_1
  Xgate_0_136_0 vdd predecode_0_8 predecode_1_8 x_0[136] y_b_noconn_0_136_0 vss and2_1
  Xgate_0_137_0 vdd predecode_0_9 predecode_1_8 x_0[137] y_b_noconn_0_137_0 vss and2_1
  Xgate_0_138_0 vdd predecode_0_10 predecode_1_8 x_0[138] y_b_noconn_0_138_0 vss and2_1
  Xgate_0_139_0 vdd predecode_0_11 predecode_1_8 x_0[139] y_b_noconn_0_139_0 vss and2_1
  Xgate_0_140_0 vdd predecode_0_12 predecode_1_8 x_0[140] y_b_noconn_0_140_0 vss and2_1
  Xgate_0_141_0 vdd predecode_0_13 predecode_1_8 x_0[141] y_b_noconn_0_141_0 vss and2_1
  Xgate_0_142_0 vdd predecode_0_14 predecode_1_8 x_0[142] y_b_noconn_0_142_0 vss and2_1
  Xgate_0_143_0 vdd predecode_0_15 predecode_1_8 x_0[143] y_b_noconn_0_143_0 vss and2_1
  Xgate_0_144_0 vdd predecode_0_0 predecode_1_9 x_0[144] y_b_noconn_0_144_0 vss and2_1
  Xgate_0_145_0 vdd predecode_0_1 predecode_1_9 x_0[145] y_b_noconn_0_145_0 vss and2_1
  Xgate_0_146_0 vdd predecode_0_2 predecode_1_9 x_0[146] y_b_noconn_0_146_0 vss and2_1
  Xgate_0_147_0 vdd predecode_0_3 predecode_1_9 x_0[147] y_b_noconn_0_147_0 vss and2_1
  Xgate_0_148_0 vdd predecode_0_4 predecode_1_9 x_0[148] y_b_noconn_0_148_0 vss and2_1
  Xgate_0_149_0 vdd predecode_0_5 predecode_1_9 x_0[149] y_b_noconn_0_149_0 vss and2_1
  Xgate_0_150_0 vdd predecode_0_6 predecode_1_9 x_0[150] y_b_noconn_0_150_0 vss and2_1
  Xgate_0_151_0 vdd predecode_0_7 predecode_1_9 x_0[151] y_b_noconn_0_151_0 vss and2_1
  Xgate_0_152_0 vdd predecode_0_8 predecode_1_9 x_0[152] y_b_noconn_0_152_0 vss and2_1
  Xgate_0_153_0 vdd predecode_0_9 predecode_1_9 x_0[153] y_b_noconn_0_153_0 vss and2_1
  Xgate_0_154_0 vdd predecode_0_10 predecode_1_9 x_0[154] y_b_noconn_0_154_0 vss and2_1
  Xgate_0_155_0 vdd predecode_0_11 predecode_1_9 x_0[155] y_b_noconn_0_155_0 vss and2_1
  Xgate_0_156_0 vdd predecode_0_12 predecode_1_9 x_0[156] y_b_noconn_0_156_0 vss and2_1
  Xgate_0_157_0 vdd predecode_0_13 predecode_1_9 x_0[157] y_b_noconn_0_157_0 vss and2_1
  Xgate_0_158_0 vdd predecode_0_14 predecode_1_9 x_0[158] y_b_noconn_0_158_0 vss and2_1
  Xgate_0_159_0 vdd predecode_0_15 predecode_1_9 x_0[159] y_b_noconn_0_159_0 vss and2_1
  Xgate_0_160_0 vdd predecode_0_0 predecode_1_10 x_0[160] y_b_noconn_0_160_0 vss and2_1
  Xgate_0_161_0 vdd predecode_0_1 predecode_1_10 x_0[161] y_b_noconn_0_161_0 vss and2_1
  Xgate_0_162_0 vdd predecode_0_2 predecode_1_10 x_0[162] y_b_noconn_0_162_0 vss and2_1
  Xgate_0_163_0 vdd predecode_0_3 predecode_1_10 x_0[163] y_b_noconn_0_163_0 vss and2_1
  Xgate_0_164_0 vdd predecode_0_4 predecode_1_10 x_0[164] y_b_noconn_0_164_0 vss and2_1
  Xgate_0_165_0 vdd predecode_0_5 predecode_1_10 x_0[165] y_b_noconn_0_165_0 vss and2_1
  Xgate_0_166_0 vdd predecode_0_6 predecode_1_10 x_0[166] y_b_noconn_0_166_0 vss and2_1
  Xgate_0_167_0 vdd predecode_0_7 predecode_1_10 x_0[167] y_b_noconn_0_167_0 vss and2_1
  Xgate_0_168_0 vdd predecode_0_8 predecode_1_10 x_0[168] y_b_noconn_0_168_0 vss and2_1
  Xgate_0_169_0 vdd predecode_0_9 predecode_1_10 x_0[169] y_b_noconn_0_169_0 vss and2_1
  Xgate_0_170_0 vdd predecode_0_10 predecode_1_10 x_0[170] y_b_noconn_0_170_0 vss and2_1
  Xgate_0_171_0 vdd predecode_0_11 predecode_1_10 x_0[171] y_b_noconn_0_171_0 vss and2_1
  Xgate_0_172_0 vdd predecode_0_12 predecode_1_10 x_0[172] y_b_noconn_0_172_0 vss and2_1
  Xgate_0_173_0 vdd predecode_0_13 predecode_1_10 x_0[173] y_b_noconn_0_173_0 vss and2_1
  Xgate_0_174_0 vdd predecode_0_14 predecode_1_10 x_0[174] y_b_noconn_0_174_0 vss and2_1
  Xgate_0_175_0 vdd predecode_0_15 predecode_1_10 x_0[175] y_b_noconn_0_175_0 vss and2_1
  Xgate_0_176_0 vdd predecode_0_0 predecode_1_11 x_0[176] y_b_noconn_0_176_0 vss and2_1
  Xgate_0_177_0 vdd predecode_0_1 predecode_1_11 x_0[177] y_b_noconn_0_177_0 vss and2_1
  Xgate_0_178_0 vdd predecode_0_2 predecode_1_11 x_0[178] y_b_noconn_0_178_0 vss and2_1
  Xgate_0_179_0 vdd predecode_0_3 predecode_1_11 x_0[179] y_b_noconn_0_179_0 vss and2_1
  Xgate_0_180_0 vdd predecode_0_4 predecode_1_11 x_0[180] y_b_noconn_0_180_0 vss and2_1
  Xgate_0_181_0 vdd predecode_0_5 predecode_1_11 x_0[181] y_b_noconn_0_181_0 vss and2_1
  Xgate_0_182_0 vdd predecode_0_6 predecode_1_11 x_0[182] y_b_noconn_0_182_0 vss and2_1
  Xgate_0_183_0 vdd predecode_0_7 predecode_1_11 x_0[183] y_b_noconn_0_183_0 vss and2_1
  Xgate_0_184_0 vdd predecode_0_8 predecode_1_11 x_0[184] y_b_noconn_0_184_0 vss and2_1
  Xgate_0_185_0 vdd predecode_0_9 predecode_1_11 x_0[185] y_b_noconn_0_185_0 vss and2_1
  Xgate_0_186_0 vdd predecode_0_10 predecode_1_11 x_0[186] y_b_noconn_0_186_0 vss and2_1
  Xgate_0_187_0 vdd predecode_0_11 predecode_1_11 x_0[187] y_b_noconn_0_187_0 vss and2_1
  Xgate_0_188_0 vdd predecode_0_12 predecode_1_11 x_0[188] y_b_noconn_0_188_0 vss and2_1
  Xgate_0_189_0 vdd predecode_0_13 predecode_1_11 x_0[189] y_b_noconn_0_189_0 vss and2_1
  Xgate_0_190_0 vdd predecode_0_14 predecode_1_11 x_0[190] y_b_noconn_0_190_0 vss and2_1
  Xgate_0_191_0 vdd predecode_0_15 predecode_1_11 x_0[191] y_b_noconn_0_191_0 vss and2_1
  Xgate_0_192_0 vdd predecode_0_0 predecode_1_12 x_0[192] y_b_noconn_0_192_0 vss and2_1
  Xgate_0_193_0 vdd predecode_0_1 predecode_1_12 x_0[193] y_b_noconn_0_193_0 vss and2_1
  Xgate_0_194_0 vdd predecode_0_2 predecode_1_12 x_0[194] y_b_noconn_0_194_0 vss and2_1
  Xgate_0_195_0 vdd predecode_0_3 predecode_1_12 x_0[195] y_b_noconn_0_195_0 vss and2_1
  Xgate_0_196_0 vdd predecode_0_4 predecode_1_12 x_0[196] y_b_noconn_0_196_0 vss and2_1
  Xgate_0_197_0 vdd predecode_0_5 predecode_1_12 x_0[197] y_b_noconn_0_197_0 vss and2_1
  Xgate_0_198_0 vdd predecode_0_6 predecode_1_12 x_0[198] y_b_noconn_0_198_0 vss and2_1
  Xgate_0_199_0 vdd predecode_0_7 predecode_1_12 x_0[199] y_b_noconn_0_199_0 vss and2_1
  Xgate_0_200_0 vdd predecode_0_8 predecode_1_12 x_0[200] y_b_noconn_0_200_0 vss and2_1
  Xgate_0_201_0 vdd predecode_0_9 predecode_1_12 x_0[201] y_b_noconn_0_201_0 vss and2_1
  Xgate_0_202_0 vdd predecode_0_10 predecode_1_12 x_0[202] y_b_noconn_0_202_0 vss and2_1
  Xgate_0_203_0 vdd predecode_0_11 predecode_1_12 x_0[203] y_b_noconn_0_203_0 vss and2_1
  Xgate_0_204_0 vdd predecode_0_12 predecode_1_12 x_0[204] y_b_noconn_0_204_0 vss and2_1
  Xgate_0_205_0 vdd predecode_0_13 predecode_1_12 x_0[205] y_b_noconn_0_205_0 vss and2_1
  Xgate_0_206_0 vdd predecode_0_14 predecode_1_12 x_0[206] y_b_noconn_0_206_0 vss and2_1
  Xgate_0_207_0 vdd predecode_0_15 predecode_1_12 x_0[207] y_b_noconn_0_207_0 vss and2_1
  Xgate_0_208_0 vdd predecode_0_0 predecode_1_13 x_0[208] y_b_noconn_0_208_0 vss and2_1
  Xgate_0_209_0 vdd predecode_0_1 predecode_1_13 x_0[209] y_b_noconn_0_209_0 vss and2_1
  Xgate_0_210_0 vdd predecode_0_2 predecode_1_13 x_0[210] y_b_noconn_0_210_0 vss and2_1
  Xgate_0_211_0 vdd predecode_0_3 predecode_1_13 x_0[211] y_b_noconn_0_211_0 vss and2_1
  Xgate_0_212_0 vdd predecode_0_4 predecode_1_13 x_0[212] y_b_noconn_0_212_0 vss and2_1
  Xgate_0_213_0 vdd predecode_0_5 predecode_1_13 x_0[213] y_b_noconn_0_213_0 vss and2_1
  Xgate_0_214_0 vdd predecode_0_6 predecode_1_13 x_0[214] y_b_noconn_0_214_0 vss and2_1
  Xgate_0_215_0 vdd predecode_0_7 predecode_1_13 x_0[215] y_b_noconn_0_215_0 vss and2_1
  Xgate_0_216_0 vdd predecode_0_8 predecode_1_13 x_0[216] y_b_noconn_0_216_0 vss and2_1
  Xgate_0_217_0 vdd predecode_0_9 predecode_1_13 x_0[217] y_b_noconn_0_217_0 vss and2_1
  Xgate_0_218_0 vdd predecode_0_10 predecode_1_13 x_0[218] y_b_noconn_0_218_0 vss and2_1
  Xgate_0_219_0 vdd predecode_0_11 predecode_1_13 x_0[219] y_b_noconn_0_219_0 vss and2_1
  Xgate_0_220_0 vdd predecode_0_12 predecode_1_13 x_0[220] y_b_noconn_0_220_0 vss and2_1
  Xgate_0_221_0 vdd predecode_0_13 predecode_1_13 x_0[221] y_b_noconn_0_221_0 vss and2_1
  Xgate_0_222_0 vdd predecode_0_14 predecode_1_13 x_0[222] y_b_noconn_0_222_0 vss and2_1
  Xgate_0_223_0 vdd predecode_0_15 predecode_1_13 x_0[223] y_b_noconn_0_223_0 vss and2_1
  Xgate_0_224_0 vdd predecode_0_0 predecode_1_14 x_0[224] y_b_noconn_0_224_0 vss and2_1
  Xgate_0_225_0 vdd predecode_0_1 predecode_1_14 x_0[225] y_b_noconn_0_225_0 vss and2_1
  Xgate_0_226_0 vdd predecode_0_2 predecode_1_14 x_0[226] y_b_noconn_0_226_0 vss and2_1
  Xgate_0_227_0 vdd predecode_0_3 predecode_1_14 x_0[227] y_b_noconn_0_227_0 vss and2_1
  Xgate_0_228_0 vdd predecode_0_4 predecode_1_14 x_0[228] y_b_noconn_0_228_0 vss and2_1
  Xgate_0_229_0 vdd predecode_0_5 predecode_1_14 x_0[229] y_b_noconn_0_229_0 vss and2_1
  Xgate_0_230_0 vdd predecode_0_6 predecode_1_14 x_0[230] y_b_noconn_0_230_0 vss and2_1
  Xgate_0_231_0 vdd predecode_0_7 predecode_1_14 x_0[231] y_b_noconn_0_231_0 vss and2_1
  Xgate_0_232_0 vdd predecode_0_8 predecode_1_14 x_0[232] y_b_noconn_0_232_0 vss and2_1
  Xgate_0_233_0 vdd predecode_0_9 predecode_1_14 x_0[233] y_b_noconn_0_233_0 vss and2_1
  Xgate_0_234_0 vdd predecode_0_10 predecode_1_14 x_0[234] y_b_noconn_0_234_0 vss and2_1
  Xgate_0_235_0 vdd predecode_0_11 predecode_1_14 x_0[235] y_b_noconn_0_235_0 vss and2_1
  Xgate_0_236_0 vdd predecode_0_12 predecode_1_14 x_0[236] y_b_noconn_0_236_0 vss and2_1
  Xgate_0_237_0 vdd predecode_0_13 predecode_1_14 x_0[237] y_b_noconn_0_237_0 vss and2_1
  Xgate_0_238_0 vdd predecode_0_14 predecode_1_14 x_0[238] y_b_noconn_0_238_0 vss and2_1
  Xgate_0_239_0 vdd predecode_0_15 predecode_1_14 x_0[239] y_b_noconn_0_239_0 vss and2_1
  Xgate_0_240_0 vdd predecode_0_0 predecode_1_15 x_0[240] y_b_noconn_0_240_0 vss and2_1
  Xgate_0_241_0 vdd predecode_0_1 predecode_1_15 x_0[241] y_b_noconn_0_241_0 vss and2_1
  Xgate_0_242_0 vdd predecode_0_2 predecode_1_15 x_0[242] y_b_noconn_0_242_0 vss and2_1
  Xgate_0_243_0 vdd predecode_0_3 predecode_1_15 x_0[243] y_b_noconn_0_243_0 vss and2_1
  Xgate_0_244_0 vdd predecode_0_4 predecode_1_15 x_0[244] y_b_noconn_0_244_0 vss and2_1
  Xgate_0_245_0 vdd predecode_0_5 predecode_1_15 x_0[245] y_b_noconn_0_245_0 vss and2_1
  Xgate_0_246_0 vdd predecode_0_6 predecode_1_15 x_0[246] y_b_noconn_0_246_0 vss and2_1
  Xgate_0_247_0 vdd predecode_0_7 predecode_1_15 x_0[247] y_b_noconn_0_247_0 vss and2_1
  Xgate_0_248_0 vdd predecode_0_8 predecode_1_15 x_0[248] y_b_noconn_0_248_0 vss and2_1
  Xgate_0_249_0 vdd predecode_0_9 predecode_1_15 x_0[249] y_b_noconn_0_249_0 vss and2_1
  Xgate_0_250_0 vdd predecode_0_10 predecode_1_15 x_0[250] y_b_noconn_0_250_0 vss and2_1
  Xgate_0_251_0 vdd predecode_0_11 predecode_1_15 x_0[251] y_b_noconn_0_251_0 vss and2_1
  Xgate_0_252_0 vdd predecode_0_12 predecode_1_15 x_0[252] y_b_noconn_0_252_0 vss and2_1
  Xgate_0_253_0 vdd predecode_0_13 predecode_1_15 x_0[253] y_b_noconn_0_253_0 vss and2_1
  Xgate_0_254_0 vdd predecode_0_14 predecode_1_15 x_0[254] y_b_noconn_0_254_0 vss and2_1
  Xgate_0_255_0 vdd predecode_0_15 predecode_1_15 x_0[255] y_b_noconn_0_255_0 vss and2_1
  Xgate_1_0_0 vdd vss x_0[0] y_b[0] multi_finger_inv_8
  Xgate_1_1_0 vdd vss x_0[1] y_b[1] multi_finger_inv_8
  Xgate_1_2_0 vdd vss x_0[2] y_b[2] multi_finger_inv_8
  Xgate_1_3_0 vdd vss x_0[3] y_b[3] multi_finger_inv_8
  Xgate_1_4_0 vdd vss x_0[4] y_b[4] multi_finger_inv_8
  Xgate_1_5_0 vdd vss x_0[5] y_b[5] multi_finger_inv_8
  Xgate_1_6_0 vdd vss x_0[6] y_b[6] multi_finger_inv_8
  Xgate_1_7_0 vdd vss x_0[7] y_b[7] multi_finger_inv_8
  Xgate_1_8_0 vdd vss x_0[8] y_b[8] multi_finger_inv_8
  Xgate_1_9_0 vdd vss x_0[9] y_b[9] multi_finger_inv_8
  Xgate_1_10_0 vdd vss x_0[10] y_b[10] multi_finger_inv_8
  Xgate_1_11_0 vdd vss x_0[11] y_b[11] multi_finger_inv_8
  Xgate_1_12_0 vdd vss x_0[12] y_b[12] multi_finger_inv_8
  Xgate_1_13_0 vdd vss x_0[13] y_b[13] multi_finger_inv_8
  Xgate_1_14_0 vdd vss x_0[14] y_b[14] multi_finger_inv_8
  Xgate_1_15_0 vdd vss x_0[15] y_b[15] multi_finger_inv_8
  Xgate_1_16_0 vdd vss x_0[16] y_b[16] multi_finger_inv_8
  Xgate_1_17_0 vdd vss x_0[17] y_b[17] multi_finger_inv_8
  Xgate_1_18_0 vdd vss x_0[18] y_b[18] multi_finger_inv_8
  Xgate_1_19_0 vdd vss x_0[19] y_b[19] multi_finger_inv_8
  Xgate_1_20_0 vdd vss x_0[20] y_b[20] multi_finger_inv_8
  Xgate_1_21_0 vdd vss x_0[21] y_b[21] multi_finger_inv_8
  Xgate_1_22_0 vdd vss x_0[22] y_b[22] multi_finger_inv_8
  Xgate_1_23_0 vdd vss x_0[23] y_b[23] multi_finger_inv_8
  Xgate_1_24_0 vdd vss x_0[24] y_b[24] multi_finger_inv_8
  Xgate_1_25_0 vdd vss x_0[25] y_b[25] multi_finger_inv_8
  Xgate_1_26_0 vdd vss x_0[26] y_b[26] multi_finger_inv_8
  Xgate_1_27_0 vdd vss x_0[27] y_b[27] multi_finger_inv_8
  Xgate_1_28_0 vdd vss x_0[28] y_b[28] multi_finger_inv_8
  Xgate_1_29_0 vdd vss x_0[29] y_b[29] multi_finger_inv_8
  Xgate_1_30_0 vdd vss x_0[30] y_b[30] multi_finger_inv_8
  Xgate_1_31_0 vdd vss x_0[31] y_b[31] multi_finger_inv_8
  Xgate_1_32_0 vdd vss x_0[32] y_b[32] multi_finger_inv_8
  Xgate_1_33_0 vdd vss x_0[33] y_b[33] multi_finger_inv_8
  Xgate_1_34_0 vdd vss x_0[34] y_b[34] multi_finger_inv_8
  Xgate_1_35_0 vdd vss x_0[35] y_b[35] multi_finger_inv_8
  Xgate_1_36_0 vdd vss x_0[36] y_b[36] multi_finger_inv_8
  Xgate_1_37_0 vdd vss x_0[37] y_b[37] multi_finger_inv_8
  Xgate_1_38_0 vdd vss x_0[38] y_b[38] multi_finger_inv_8
  Xgate_1_39_0 vdd vss x_0[39] y_b[39] multi_finger_inv_8
  Xgate_1_40_0 vdd vss x_0[40] y_b[40] multi_finger_inv_8
  Xgate_1_41_0 vdd vss x_0[41] y_b[41] multi_finger_inv_8
  Xgate_1_42_0 vdd vss x_0[42] y_b[42] multi_finger_inv_8
  Xgate_1_43_0 vdd vss x_0[43] y_b[43] multi_finger_inv_8
  Xgate_1_44_0 vdd vss x_0[44] y_b[44] multi_finger_inv_8
  Xgate_1_45_0 vdd vss x_0[45] y_b[45] multi_finger_inv_8
  Xgate_1_46_0 vdd vss x_0[46] y_b[46] multi_finger_inv_8
  Xgate_1_47_0 vdd vss x_0[47] y_b[47] multi_finger_inv_8
  Xgate_1_48_0 vdd vss x_0[48] y_b[48] multi_finger_inv_8
  Xgate_1_49_0 vdd vss x_0[49] y_b[49] multi_finger_inv_8
  Xgate_1_50_0 vdd vss x_0[50] y_b[50] multi_finger_inv_8
  Xgate_1_51_0 vdd vss x_0[51] y_b[51] multi_finger_inv_8
  Xgate_1_52_0 vdd vss x_0[52] y_b[52] multi_finger_inv_8
  Xgate_1_53_0 vdd vss x_0[53] y_b[53] multi_finger_inv_8
  Xgate_1_54_0 vdd vss x_0[54] y_b[54] multi_finger_inv_8
  Xgate_1_55_0 vdd vss x_0[55] y_b[55] multi_finger_inv_8
  Xgate_1_56_0 vdd vss x_0[56] y_b[56] multi_finger_inv_8
  Xgate_1_57_0 vdd vss x_0[57] y_b[57] multi_finger_inv_8
  Xgate_1_58_0 vdd vss x_0[58] y_b[58] multi_finger_inv_8
  Xgate_1_59_0 vdd vss x_0[59] y_b[59] multi_finger_inv_8
  Xgate_1_60_0 vdd vss x_0[60] y_b[60] multi_finger_inv_8
  Xgate_1_61_0 vdd vss x_0[61] y_b[61] multi_finger_inv_8
  Xgate_1_62_0 vdd vss x_0[62] y_b[62] multi_finger_inv_8
  Xgate_1_63_0 vdd vss x_0[63] y_b[63] multi_finger_inv_8
  Xgate_1_64_0 vdd vss x_0[64] y_b[64] multi_finger_inv_8
  Xgate_1_65_0 vdd vss x_0[65] y_b[65] multi_finger_inv_8
  Xgate_1_66_0 vdd vss x_0[66] y_b[66] multi_finger_inv_8
  Xgate_1_67_0 vdd vss x_0[67] y_b[67] multi_finger_inv_8
  Xgate_1_68_0 vdd vss x_0[68] y_b[68] multi_finger_inv_8
  Xgate_1_69_0 vdd vss x_0[69] y_b[69] multi_finger_inv_8
  Xgate_1_70_0 vdd vss x_0[70] y_b[70] multi_finger_inv_8
  Xgate_1_71_0 vdd vss x_0[71] y_b[71] multi_finger_inv_8
  Xgate_1_72_0 vdd vss x_0[72] y_b[72] multi_finger_inv_8
  Xgate_1_73_0 vdd vss x_0[73] y_b[73] multi_finger_inv_8
  Xgate_1_74_0 vdd vss x_0[74] y_b[74] multi_finger_inv_8
  Xgate_1_75_0 vdd vss x_0[75] y_b[75] multi_finger_inv_8
  Xgate_1_76_0 vdd vss x_0[76] y_b[76] multi_finger_inv_8
  Xgate_1_77_0 vdd vss x_0[77] y_b[77] multi_finger_inv_8
  Xgate_1_78_0 vdd vss x_0[78] y_b[78] multi_finger_inv_8
  Xgate_1_79_0 vdd vss x_0[79] y_b[79] multi_finger_inv_8
  Xgate_1_80_0 vdd vss x_0[80] y_b[80] multi_finger_inv_8
  Xgate_1_81_0 vdd vss x_0[81] y_b[81] multi_finger_inv_8
  Xgate_1_82_0 vdd vss x_0[82] y_b[82] multi_finger_inv_8
  Xgate_1_83_0 vdd vss x_0[83] y_b[83] multi_finger_inv_8
  Xgate_1_84_0 vdd vss x_0[84] y_b[84] multi_finger_inv_8
  Xgate_1_85_0 vdd vss x_0[85] y_b[85] multi_finger_inv_8
  Xgate_1_86_0 vdd vss x_0[86] y_b[86] multi_finger_inv_8
  Xgate_1_87_0 vdd vss x_0[87] y_b[87] multi_finger_inv_8
  Xgate_1_88_0 vdd vss x_0[88] y_b[88] multi_finger_inv_8
  Xgate_1_89_0 vdd vss x_0[89] y_b[89] multi_finger_inv_8
  Xgate_1_90_0 vdd vss x_0[90] y_b[90] multi_finger_inv_8
  Xgate_1_91_0 vdd vss x_0[91] y_b[91] multi_finger_inv_8
  Xgate_1_92_0 vdd vss x_0[92] y_b[92] multi_finger_inv_8
  Xgate_1_93_0 vdd vss x_0[93] y_b[93] multi_finger_inv_8
  Xgate_1_94_0 vdd vss x_0[94] y_b[94] multi_finger_inv_8
  Xgate_1_95_0 vdd vss x_0[95] y_b[95] multi_finger_inv_8
  Xgate_1_96_0 vdd vss x_0[96] y_b[96] multi_finger_inv_8
  Xgate_1_97_0 vdd vss x_0[97] y_b[97] multi_finger_inv_8
  Xgate_1_98_0 vdd vss x_0[98] y_b[98] multi_finger_inv_8
  Xgate_1_99_0 vdd vss x_0[99] y_b[99] multi_finger_inv_8
  Xgate_1_100_0 vdd vss x_0[100] y_b[100] multi_finger_inv_8
  Xgate_1_101_0 vdd vss x_0[101] y_b[101] multi_finger_inv_8
  Xgate_1_102_0 vdd vss x_0[102] y_b[102] multi_finger_inv_8
  Xgate_1_103_0 vdd vss x_0[103] y_b[103] multi_finger_inv_8
  Xgate_1_104_0 vdd vss x_0[104] y_b[104] multi_finger_inv_8
  Xgate_1_105_0 vdd vss x_0[105] y_b[105] multi_finger_inv_8
  Xgate_1_106_0 vdd vss x_0[106] y_b[106] multi_finger_inv_8
  Xgate_1_107_0 vdd vss x_0[107] y_b[107] multi_finger_inv_8
  Xgate_1_108_0 vdd vss x_0[108] y_b[108] multi_finger_inv_8
  Xgate_1_109_0 vdd vss x_0[109] y_b[109] multi_finger_inv_8
  Xgate_1_110_0 vdd vss x_0[110] y_b[110] multi_finger_inv_8
  Xgate_1_111_0 vdd vss x_0[111] y_b[111] multi_finger_inv_8
  Xgate_1_112_0 vdd vss x_0[112] y_b[112] multi_finger_inv_8
  Xgate_1_113_0 vdd vss x_0[113] y_b[113] multi_finger_inv_8
  Xgate_1_114_0 vdd vss x_0[114] y_b[114] multi_finger_inv_8
  Xgate_1_115_0 vdd vss x_0[115] y_b[115] multi_finger_inv_8
  Xgate_1_116_0 vdd vss x_0[116] y_b[116] multi_finger_inv_8
  Xgate_1_117_0 vdd vss x_0[117] y_b[117] multi_finger_inv_8
  Xgate_1_118_0 vdd vss x_0[118] y_b[118] multi_finger_inv_8
  Xgate_1_119_0 vdd vss x_0[119] y_b[119] multi_finger_inv_8
  Xgate_1_120_0 vdd vss x_0[120] y_b[120] multi_finger_inv_8
  Xgate_1_121_0 vdd vss x_0[121] y_b[121] multi_finger_inv_8
  Xgate_1_122_0 vdd vss x_0[122] y_b[122] multi_finger_inv_8
  Xgate_1_123_0 vdd vss x_0[123] y_b[123] multi_finger_inv_8
  Xgate_1_124_0 vdd vss x_0[124] y_b[124] multi_finger_inv_8
  Xgate_1_125_0 vdd vss x_0[125] y_b[125] multi_finger_inv_8
  Xgate_1_126_0 vdd vss x_0[126] y_b[126] multi_finger_inv_8
  Xgate_1_127_0 vdd vss x_0[127] y_b[127] multi_finger_inv_8
  Xgate_1_128_0 vdd vss x_0[128] y_b[128] multi_finger_inv_8
  Xgate_1_129_0 vdd vss x_0[129] y_b[129] multi_finger_inv_8
  Xgate_1_130_0 vdd vss x_0[130] y_b[130] multi_finger_inv_8
  Xgate_1_131_0 vdd vss x_0[131] y_b[131] multi_finger_inv_8
  Xgate_1_132_0 vdd vss x_0[132] y_b[132] multi_finger_inv_8
  Xgate_1_133_0 vdd vss x_0[133] y_b[133] multi_finger_inv_8
  Xgate_1_134_0 vdd vss x_0[134] y_b[134] multi_finger_inv_8
  Xgate_1_135_0 vdd vss x_0[135] y_b[135] multi_finger_inv_8
  Xgate_1_136_0 vdd vss x_0[136] y_b[136] multi_finger_inv_8
  Xgate_1_137_0 vdd vss x_0[137] y_b[137] multi_finger_inv_8
  Xgate_1_138_0 vdd vss x_0[138] y_b[138] multi_finger_inv_8
  Xgate_1_139_0 vdd vss x_0[139] y_b[139] multi_finger_inv_8
  Xgate_1_140_0 vdd vss x_0[140] y_b[140] multi_finger_inv_8
  Xgate_1_141_0 vdd vss x_0[141] y_b[141] multi_finger_inv_8
  Xgate_1_142_0 vdd vss x_0[142] y_b[142] multi_finger_inv_8
  Xgate_1_143_0 vdd vss x_0[143] y_b[143] multi_finger_inv_8
  Xgate_1_144_0 vdd vss x_0[144] y_b[144] multi_finger_inv_8
  Xgate_1_145_0 vdd vss x_0[145] y_b[145] multi_finger_inv_8
  Xgate_1_146_0 vdd vss x_0[146] y_b[146] multi_finger_inv_8
  Xgate_1_147_0 vdd vss x_0[147] y_b[147] multi_finger_inv_8
  Xgate_1_148_0 vdd vss x_0[148] y_b[148] multi_finger_inv_8
  Xgate_1_149_0 vdd vss x_0[149] y_b[149] multi_finger_inv_8
  Xgate_1_150_0 vdd vss x_0[150] y_b[150] multi_finger_inv_8
  Xgate_1_151_0 vdd vss x_0[151] y_b[151] multi_finger_inv_8
  Xgate_1_152_0 vdd vss x_0[152] y_b[152] multi_finger_inv_8
  Xgate_1_153_0 vdd vss x_0[153] y_b[153] multi_finger_inv_8
  Xgate_1_154_0 vdd vss x_0[154] y_b[154] multi_finger_inv_8
  Xgate_1_155_0 vdd vss x_0[155] y_b[155] multi_finger_inv_8
  Xgate_1_156_0 vdd vss x_0[156] y_b[156] multi_finger_inv_8
  Xgate_1_157_0 vdd vss x_0[157] y_b[157] multi_finger_inv_8
  Xgate_1_158_0 vdd vss x_0[158] y_b[158] multi_finger_inv_8
  Xgate_1_159_0 vdd vss x_0[159] y_b[159] multi_finger_inv_8
  Xgate_1_160_0 vdd vss x_0[160] y_b[160] multi_finger_inv_8
  Xgate_1_161_0 vdd vss x_0[161] y_b[161] multi_finger_inv_8
  Xgate_1_162_0 vdd vss x_0[162] y_b[162] multi_finger_inv_8
  Xgate_1_163_0 vdd vss x_0[163] y_b[163] multi_finger_inv_8
  Xgate_1_164_0 vdd vss x_0[164] y_b[164] multi_finger_inv_8
  Xgate_1_165_0 vdd vss x_0[165] y_b[165] multi_finger_inv_8
  Xgate_1_166_0 vdd vss x_0[166] y_b[166] multi_finger_inv_8
  Xgate_1_167_0 vdd vss x_0[167] y_b[167] multi_finger_inv_8
  Xgate_1_168_0 vdd vss x_0[168] y_b[168] multi_finger_inv_8
  Xgate_1_169_0 vdd vss x_0[169] y_b[169] multi_finger_inv_8
  Xgate_1_170_0 vdd vss x_0[170] y_b[170] multi_finger_inv_8
  Xgate_1_171_0 vdd vss x_0[171] y_b[171] multi_finger_inv_8
  Xgate_1_172_0 vdd vss x_0[172] y_b[172] multi_finger_inv_8
  Xgate_1_173_0 vdd vss x_0[173] y_b[173] multi_finger_inv_8
  Xgate_1_174_0 vdd vss x_0[174] y_b[174] multi_finger_inv_8
  Xgate_1_175_0 vdd vss x_0[175] y_b[175] multi_finger_inv_8
  Xgate_1_176_0 vdd vss x_0[176] y_b[176] multi_finger_inv_8
  Xgate_1_177_0 vdd vss x_0[177] y_b[177] multi_finger_inv_8
  Xgate_1_178_0 vdd vss x_0[178] y_b[178] multi_finger_inv_8
  Xgate_1_179_0 vdd vss x_0[179] y_b[179] multi_finger_inv_8
  Xgate_1_180_0 vdd vss x_0[180] y_b[180] multi_finger_inv_8
  Xgate_1_181_0 vdd vss x_0[181] y_b[181] multi_finger_inv_8
  Xgate_1_182_0 vdd vss x_0[182] y_b[182] multi_finger_inv_8
  Xgate_1_183_0 vdd vss x_0[183] y_b[183] multi_finger_inv_8
  Xgate_1_184_0 vdd vss x_0[184] y_b[184] multi_finger_inv_8
  Xgate_1_185_0 vdd vss x_0[185] y_b[185] multi_finger_inv_8
  Xgate_1_186_0 vdd vss x_0[186] y_b[186] multi_finger_inv_8
  Xgate_1_187_0 vdd vss x_0[187] y_b[187] multi_finger_inv_8
  Xgate_1_188_0 vdd vss x_0[188] y_b[188] multi_finger_inv_8
  Xgate_1_189_0 vdd vss x_0[189] y_b[189] multi_finger_inv_8
  Xgate_1_190_0 vdd vss x_0[190] y_b[190] multi_finger_inv_8
  Xgate_1_191_0 vdd vss x_0[191] y_b[191] multi_finger_inv_8
  Xgate_1_192_0 vdd vss x_0[192] y_b[192] multi_finger_inv_8
  Xgate_1_193_0 vdd vss x_0[193] y_b[193] multi_finger_inv_8
  Xgate_1_194_0 vdd vss x_0[194] y_b[194] multi_finger_inv_8
  Xgate_1_195_0 vdd vss x_0[195] y_b[195] multi_finger_inv_8
  Xgate_1_196_0 vdd vss x_0[196] y_b[196] multi_finger_inv_8
  Xgate_1_197_0 vdd vss x_0[197] y_b[197] multi_finger_inv_8
  Xgate_1_198_0 vdd vss x_0[198] y_b[198] multi_finger_inv_8
  Xgate_1_199_0 vdd vss x_0[199] y_b[199] multi_finger_inv_8
  Xgate_1_200_0 vdd vss x_0[200] y_b[200] multi_finger_inv_8
  Xgate_1_201_0 vdd vss x_0[201] y_b[201] multi_finger_inv_8
  Xgate_1_202_0 vdd vss x_0[202] y_b[202] multi_finger_inv_8
  Xgate_1_203_0 vdd vss x_0[203] y_b[203] multi_finger_inv_8
  Xgate_1_204_0 vdd vss x_0[204] y_b[204] multi_finger_inv_8
  Xgate_1_205_0 vdd vss x_0[205] y_b[205] multi_finger_inv_8
  Xgate_1_206_0 vdd vss x_0[206] y_b[206] multi_finger_inv_8
  Xgate_1_207_0 vdd vss x_0[207] y_b[207] multi_finger_inv_8
  Xgate_1_208_0 vdd vss x_0[208] y_b[208] multi_finger_inv_8
  Xgate_1_209_0 vdd vss x_0[209] y_b[209] multi_finger_inv_8
  Xgate_1_210_0 vdd vss x_0[210] y_b[210] multi_finger_inv_8
  Xgate_1_211_0 vdd vss x_0[211] y_b[211] multi_finger_inv_8
  Xgate_1_212_0 vdd vss x_0[212] y_b[212] multi_finger_inv_8
  Xgate_1_213_0 vdd vss x_0[213] y_b[213] multi_finger_inv_8
  Xgate_1_214_0 vdd vss x_0[214] y_b[214] multi_finger_inv_8
  Xgate_1_215_0 vdd vss x_0[215] y_b[215] multi_finger_inv_8
  Xgate_1_216_0 vdd vss x_0[216] y_b[216] multi_finger_inv_8
  Xgate_1_217_0 vdd vss x_0[217] y_b[217] multi_finger_inv_8
  Xgate_1_218_0 vdd vss x_0[218] y_b[218] multi_finger_inv_8
  Xgate_1_219_0 vdd vss x_0[219] y_b[219] multi_finger_inv_8
  Xgate_1_220_0 vdd vss x_0[220] y_b[220] multi_finger_inv_8
  Xgate_1_221_0 vdd vss x_0[221] y_b[221] multi_finger_inv_8
  Xgate_1_222_0 vdd vss x_0[222] y_b[222] multi_finger_inv_8
  Xgate_1_223_0 vdd vss x_0[223] y_b[223] multi_finger_inv_8
  Xgate_1_224_0 vdd vss x_0[224] y_b[224] multi_finger_inv_8
  Xgate_1_225_0 vdd vss x_0[225] y_b[225] multi_finger_inv_8
  Xgate_1_226_0 vdd vss x_0[226] y_b[226] multi_finger_inv_8
  Xgate_1_227_0 vdd vss x_0[227] y_b[227] multi_finger_inv_8
  Xgate_1_228_0 vdd vss x_0[228] y_b[228] multi_finger_inv_8
  Xgate_1_229_0 vdd vss x_0[229] y_b[229] multi_finger_inv_8
  Xgate_1_230_0 vdd vss x_0[230] y_b[230] multi_finger_inv_8
  Xgate_1_231_0 vdd vss x_0[231] y_b[231] multi_finger_inv_8
  Xgate_1_232_0 vdd vss x_0[232] y_b[232] multi_finger_inv_8
  Xgate_1_233_0 vdd vss x_0[233] y_b[233] multi_finger_inv_8
  Xgate_1_234_0 vdd vss x_0[234] y_b[234] multi_finger_inv_8
  Xgate_1_235_0 vdd vss x_0[235] y_b[235] multi_finger_inv_8
  Xgate_1_236_0 vdd vss x_0[236] y_b[236] multi_finger_inv_8
  Xgate_1_237_0 vdd vss x_0[237] y_b[237] multi_finger_inv_8
  Xgate_1_238_0 vdd vss x_0[238] y_b[238] multi_finger_inv_8
  Xgate_1_239_0 vdd vss x_0[239] y_b[239] multi_finger_inv_8
  Xgate_1_240_0 vdd vss x_0[240] y_b[240] multi_finger_inv_8
  Xgate_1_241_0 vdd vss x_0[241] y_b[241] multi_finger_inv_8
  Xgate_1_242_0 vdd vss x_0[242] y_b[242] multi_finger_inv_8
  Xgate_1_243_0 vdd vss x_0[243] y_b[243] multi_finger_inv_8
  Xgate_1_244_0 vdd vss x_0[244] y_b[244] multi_finger_inv_8
  Xgate_1_245_0 vdd vss x_0[245] y_b[245] multi_finger_inv_8
  Xgate_1_246_0 vdd vss x_0[246] y_b[246] multi_finger_inv_8
  Xgate_1_247_0 vdd vss x_0[247] y_b[247] multi_finger_inv_8
  Xgate_1_248_0 vdd vss x_0[248] y_b[248] multi_finger_inv_8
  Xgate_1_249_0 vdd vss x_0[249] y_b[249] multi_finger_inv_8
  Xgate_1_250_0 vdd vss x_0[250] y_b[250] multi_finger_inv_8
  Xgate_1_251_0 vdd vss x_0[251] y_b[251] multi_finger_inv_8
  Xgate_1_252_0 vdd vss x_0[252] y_b[252] multi_finger_inv_8
  Xgate_1_253_0 vdd vss x_0[253] y_b[253] multi_finger_inv_8
  Xgate_1_254_0 vdd vss x_0[254] y_b[254] multi_finger_inv_8
  Xgate_1_255_0 vdd vss x_0[255] y_b[255] multi_finger_inv_8
  Xgate_2_0_0 vdd vss y_b[0] y[0] multi_finger_inv_9
  Xgate_2_1_0 vdd vss y_b[1] y[1] multi_finger_inv_9
  Xgate_2_2_0 vdd vss y_b[2] y[2] multi_finger_inv_9
  Xgate_2_3_0 vdd vss y_b[3] y[3] multi_finger_inv_9
  Xgate_2_4_0 vdd vss y_b[4] y[4] multi_finger_inv_9
  Xgate_2_5_0 vdd vss y_b[5] y[5] multi_finger_inv_9
  Xgate_2_6_0 vdd vss y_b[6] y[6] multi_finger_inv_9
  Xgate_2_7_0 vdd vss y_b[7] y[7] multi_finger_inv_9
  Xgate_2_8_0 vdd vss y_b[8] y[8] multi_finger_inv_9
  Xgate_2_9_0 vdd vss y_b[9] y[9] multi_finger_inv_9
  Xgate_2_10_0 vdd vss y_b[10] y[10] multi_finger_inv_9
  Xgate_2_11_0 vdd vss y_b[11] y[11] multi_finger_inv_9
  Xgate_2_12_0 vdd vss y_b[12] y[12] multi_finger_inv_9
  Xgate_2_13_0 vdd vss y_b[13] y[13] multi_finger_inv_9
  Xgate_2_14_0 vdd vss y_b[14] y[14] multi_finger_inv_9
  Xgate_2_15_0 vdd vss y_b[15] y[15] multi_finger_inv_9
  Xgate_2_16_0 vdd vss y_b[16] y[16] multi_finger_inv_9
  Xgate_2_17_0 vdd vss y_b[17] y[17] multi_finger_inv_9
  Xgate_2_18_0 vdd vss y_b[18] y[18] multi_finger_inv_9
  Xgate_2_19_0 vdd vss y_b[19] y[19] multi_finger_inv_9
  Xgate_2_20_0 vdd vss y_b[20] y[20] multi_finger_inv_9
  Xgate_2_21_0 vdd vss y_b[21] y[21] multi_finger_inv_9
  Xgate_2_22_0 vdd vss y_b[22] y[22] multi_finger_inv_9
  Xgate_2_23_0 vdd vss y_b[23] y[23] multi_finger_inv_9
  Xgate_2_24_0 vdd vss y_b[24] y[24] multi_finger_inv_9
  Xgate_2_25_0 vdd vss y_b[25] y[25] multi_finger_inv_9
  Xgate_2_26_0 vdd vss y_b[26] y[26] multi_finger_inv_9
  Xgate_2_27_0 vdd vss y_b[27] y[27] multi_finger_inv_9
  Xgate_2_28_0 vdd vss y_b[28] y[28] multi_finger_inv_9
  Xgate_2_29_0 vdd vss y_b[29] y[29] multi_finger_inv_9
  Xgate_2_30_0 vdd vss y_b[30] y[30] multi_finger_inv_9
  Xgate_2_31_0 vdd vss y_b[31] y[31] multi_finger_inv_9
  Xgate_2_32_0 vdd vss y_b[32] y[32] multi_finger_inv_9
  Xgate_2_33_0 vdd vss y_b[33] y[33] multi_finger_inv_9
  Xgate_2_34_0 vdd vss y_b[34] y[34] multi_finger_inv_9
  Xgate_2_35_0 vdd vss y_b[35] y[35] multi_finger_inv_9
  Xgate_2_36_0 vdd vss y_b[36] y[36] multi_finger_inv_9
  Xgate_2_37_0 vdd vss y_b[37] y[37] multi_finger_inv_9
  Xgate_2_38_0 vdd vss y_b[38] y[38] multi_finger_inv_9
  Xgate_2_39_0 vdd vss y_b[39] y[39] multi_finger_inv_9
  Xgate_2_40_0 vdd vss y_b[40] y[40] multi_finger_inv_9
  Xgate_2_41_0 vdd vss y_b[41] y[41] multi_finger_inv_9
  Xgate_2_42_0 vdd vss y_b[42] y[42] multi_finger_inv_9
  Xgate_2_43_0 vdd vss y_b[43] y[43] multi_finger_inv_9
  Xgate_2_44_0 vdd vss y_b[44] y[44] multi_finger_inv_9
  Xgate_2_45_0 vdd vss y_b[45] y[45] multi_finger_inv_9
  Xgate_2_46_0 vdd vss y_b[46] y[46] multi_finger_inv_9
  Xgate_2_47_0 vdd vss y_b[47] y[47] multi_finger_inv_9
  Xgate_2_48_0 vdd vss y_b[48] y[48] multi_finger_inv_9
  Xgate_2_49_0 vdd vss y_b[49] y[49] multi_finger_inv_9
  Xgate_2_50_0 vdd vss y_b[50] y[50] multi_finger_inv_9
  Xgate_2_51_0 vdd vss y_b[51] y[51] multi_finger_inv_9
  Xgate_2_52_0 vdd vss y_b[52] y[52] multi_finger_inv_9
  Xgate_2_53_0 vdd vss y_b[53] y[53] multi_finger_inv_9
  Xgate_2_54_0 vdd vss y_b[54] y[54] multi_finger_inv_9
  Xgate_2_55_0 vdd vss y_b[55] y[55] multi_finger_inv_9
  Xgate_2_56_0 vdd vss y_b[56] y[56] multi_finger_inv_9
  Xgate_2_57_0 vdd vss y_b[57] y[57] multi_finger_inv_9
  Xgate_2_58_0 vdd vss y_b[58] y[58] multi_finger_inv_9
  Xgate_2_59_0 vdd vss y_b[59] y[59] multi_finger_inv_9
  Xgate_2_60_0 vdd vss y_b[60] y[60] multi_finger_inv_9
  Xgate_2_61_0 vdd vss y_b[61] y[61] multi_finger_inv_9
  Xgate_2_62_0 vdd vss y_b[62] y[62] multi_finger_inv_9
  Xgate_2_63_0 vdd vss y_b[63] y[63] multi_finger_inv_9
  Xgate_2_64_0 vdd vss y_b[64] y[64] multi_finger_inv_9
  Xgate_2_65_0 vdd vss y_b[65] y[65] multi_finger_inv_9
  Xgate_2_66_0 vdd vss y_b[66] y[66] multi_finger_inv_9
  Xgate_2_67_0 vdd vss y_b[67] y[67] multi_finger_inv_9
  Xgate_2_68_0 vdd vss y_b[68] y[68] multi_finger_inv_9
  Xgate_2_69_0 vdd vss y_b[69] y[69] multi_finger_inv_9
  Xgate_2_70_0 vdd vss y_b[70] y[70] multi_finger_inv_9
  Xgate_2_71_0 vdd vss y_b[71] y[71] multi_finger_inv_9
  Xgate_2_72_0 vdd vss y_b[72] y[72] multi_finger_inv_9
  Xgate_2_73_0 vdd vss y_b[73] y[73] multi_finger_inv_9
  Xgate_2_74_0 vdd vss y_b[74] y[74] multi_finger_inv_9
  Xgate_2_75_0 vdd vss y_b[75] y[75] multi_finger_inv_9
  Xgate_2_76_0 vdd vss y_b[76] y[76] multi_finger_inv_9
  Xgate_2_77_0 vdd vss y_b[77] y[77] multi_finger_inv_9
  Xgate_2_78_0 vdd vss y_b[78] y[78] multi_finger_inv_9
  Xgate_2_79_0 vdd vss y_b[79] y[79] multi_finger_inv_9
  Xgate_2_80_0 vdd vss y_b[80] y[80] multi_finger_inv_9
  Xgate_2_81_0 vdd vss y_b[81] y[81] multi_finger_inv_9
  Xgate_2_82_0 vdd vss y_b[82] y[82] multi_finger_inv_9
  Xgate_2_83_0 vdd vss y_b[83] y[83] multi_finger_inv_9
  Xgate_2_84_0 vdd vss y_b[84] y[84] multi_finger_inv_9
  Xgate_2_85_0 vdd vss y_b[85] y[85] multi_finger_inv_9
  Xgate_2_86_0 vdd vss y_b[86] y[86] multi_finger_inv_9
  Xgate_2_87_0 vdd vss y_b[87] y[87] multi_finger_inv_9
  Xgate_2_88_0 vdd vss y_b[88] y[88] multi_finger_inv_9
  Xgate_2_89_0 vdd vss y_b[89] y[89] multi_finger_inv_9
  Xgate_2_90_0 vdd vss y_b[90] y[90] multi_finger_inv_9
  Xgate_2_91_0 vdd vss y_b[91] y[91] multi_finger_inv_9
  Xgate_2_92_0 vdd vss y_b[92] y[92] multi_finger_inv_9
  Xgate_2_93_0 vdd vss y_b[93] y[93] multi_finger_inv_9
  Xgate_2_94_0 vdd vss y_b[94] y[94] multi_finger_inv_9
  Xgate_2_95_0 vdd vss y_b[95] y[95] multi_finger_inv_9
  Xgate_2_96_0 vdd vss y_b[96] y[96] multi_finger_inv_9
  Xgate_2_97_0 vdd vss y_b[97] y[97] multi_finger_inv_9
  Xgate_2_98_0 vdd vss y_b[98] y[98] multi_finger_inv_9
  Xgate_2_99_0 vdd vss y_b[99] y[99] multi_finger_inv_9
  Xgate_2_100_0 vdd vss y_b[100] y[100] multi_finger_inv_9
  Xgate_2_101_0 vdd vss y_b[101] y[101] multi_finger_inv_9
  Xgate_2_102_0 vdd vss y_b[102] y[102] multi_finger_inv_9
  Xgate_2_103_0 vdd vss y_b[103] y[103] multi_finger_inv_9
  Xgate_2_104_0 vdd vss y_b[104] y[104] multi_finger_inv_9
  Xgate_2_105_0 vdd vss y_b[105] y[105] multi_finger_inv_9
  Xgate_2_106_0 vdd vss y_b[106] y[106] multi_finger_inv_9
  Xgate_2_107_0 vdd vss y_b[107] y[107] multi_finger_inv_9
  Xgate_2_108_0 vdd vss y_b[108] y[108] multi_finger_inv_9
  Xgate_2_109_0 vdd vss y_b[109] y[109] multi_finger_inv_9
  Xgate_2_110_0 vdd vss y_b[110] y[110] multi_finger_inv_9
  Xgate_2_111_0 vdd vss y_b[111] y[111] multi_finger_inv_9
  Xgate_2_112_0 vdd vss y_b[112] y[112] multi_finger_inv_9
  Xgate_2_113_0 vdd vss y_b[113] y[113] multi_finger_inv_9
  Xgate_2_114_0 vdd vss y_b[114] y[114] multi_finger_inv_9
  Xgate_2_115_0 vdd vss y_b[115] y[115] multi_finger_inv_9
  Xgate_2_116_0 vdd vss y_b[116] y[116] multi_finger_inv_9
  Xgate_2_117_0 vdd vss y_b[117] y[117] multi_finger_inv_9
  Xgate_2_118_0 vdd vss y_b[118] y[118] multi_finger_inv_9
  Xgate_2_119_0 vdd vss y_b[119] y[119] multi_finger_inv_9
  Xgate_2_120_0 vdd vss y_b[120] y[120] multi_finger_inv_9
  Xgate_2_121_0 vdd vss y_b[121] y[121] multi_finger_inv_9
  Xgate_2_122_0 vdd vss y_b[122] y[122] multi_finger_inv_9
  Xgate_2_123_0 vdd vss y_b[123] y[123] multi_finger_inv_9
  Xgate_2_124_0 vdd vss y_b[124] y[124] multi_finger_inv_9
  Xgate_2_125_0 vdd vss y_b[125] y[125] multi_finger_inv_9
  Xgate_2_126_0 vdd vss y_b[126] y[126] multi_finger_inv_9
  Xgate_2_127_0 vdd vss y_b[127] y[127] multi_finger_inv_9
  Xgate_2_128_0 vdd vss y_b[128] y[128] multi_finger_inv_9
  Xgate_2_129_0 vdd vss y_b[129] y[129] multi_finger_inv_9
  Xgate_2_130_0 vdd vss y_b[130] y[130] multi_finger_inv_9
  Xgate_2_131_0 vdd vss y_b[131] y[131] multi_finger_inv_9
  Xgate_2_132_0 vdd vss y_b[132] y[132] multi_finger_inv_9
  Xgate_2_133_0 vdd vss y_b[133] y[133] multi_finger_inv_9
  Xgate_2_134_0 vdd vss y_b[134] y[134] multi_finger_inv_9
  Xgate_2_135_0 vdd vss y_b[135] y[135] multi_finger_inv_9
  Xgate_2_136_0 vdd vss y_b[136] y[136] multi_finger_inv_9
  Xgate_2_137_0 vdd vss y_b[137] y[137] multi_finger_inv_9
  Xgate_2_138_0 vdd vss y_b[138] y[138] multi_finger_inv_9
  Xgate_2_139_0 vdd vss y_b[139] y[139] multi_finger_inv_9
  Xgate_2_140_0 vdd vss y_b[140] y[140] multi_finger_inv_9
  Xgate_2_141_0 vdd vss y_b[141] y[141] multi_finger_inv_9
  Xgate_2_142_0 vdd vss y_b[142] y[142] multi_finger_inv_9
  Xgate_2_143_0 vdd vss y_b[143] y[143] multi_finger_inv_9
  Xgate_2_144_0 vdd vss y_b[144] y[144] multi_finger_inv_9
  Xgate_2_145_0 vdd vss y_b[145] y[145] multi_finger_inv_9
  Xgate_2_146_0 vdd vss y_b[146] y[146] multi_finger_inv_9
  Xgate_2_147_0 vdd vss y_b[147] y[147] multi_finger_inv_9
  Xgate_2_148_0 vdd vss y_b[148] y[148] multi_finger_inv_9
  Xgate_2_149_0 vdd vss y_b[149] y[149] multi_finger_inv_9
  Xgate_2_150_0 vdd vss y_b[150] y[150] multi_finger_inv_9
  Xgate_2_151_0 vdd vss y_b[151] y[151] multi_finger_inv_9
  Xgate_2_152_0 vdd vss y_b[152] y[152] multi_finger_inv_9
  Xgate_2_153_0 vdd vss y_b[153] y[153] multi_finger_inv_9
  Xgate_2_154_0 vdd vss y_b[154] y[154] multi_finger_inv_9
  Xgate_2_155_0 vdd vss y_b[155] y[155] multi_finger_inv_9
  Xgate_2_156_0 vdd vss y_b[156] y[156] multi_finger_inv_9
  Xgate_2_157_0 vdd vss y_b[157] y[157] multi_finger_inv_9
  Xgate_2_158_0 vdd vss y_b[158] y[158] multi_finger_inv_9
  Xgate_2_159_0 vdd vss y_b[159] y[159] multi_finger_inv_9
  Xgate_2_160_0 vdd vss y_b[160] y[160] multi_finger_inv_9
  Xgate_2_161_0 vdd vss y_b[161] y[161] multi_finger_inv_9
  Xgate_2_162_0 vdd vss y_b[162] y[162] multi_finger_inv_9
  Xgate_2_163_0 vdd vss y_b[163] y[163] multi_finger_inv_9
  Xgate_2_164_0 vdd vss y_b[164] y[164] multi_finger_inv_9
  Xgate_2_165_0 vdd vss y_b[165] y[165] multi_finger_inv_9
  Xgate_2_166_0 vdd vss y_b[166] y[166] multi_finger_inv_9
  Xgate_2_167_0 vdd vss y_b[167] y[167] multi_finger_inv_9
  Xgate_2_168_0 vdd vss y_b[168] y[168] multi_finger_inv_9
  Xgate_2_169_0 vdd vss y_b[169] y[169] multi_finger_inv_9
  Xgate_2_170_0 vdd vss y_b[170] y[170] multi_finger_inv_9
  Xgate_2_171_0 vdd vss y_b[171] y[171] multi_finger_inv_9
  Xgate_2_172_0 vdd vss y_b[172] y[172] multi_finger_inv_9
  Xgate_2_173_0 vdd vss y_b[173] y[173] multi_finger_inv_9
  Xgate_2_174_0 vdd vss y_b[174] y[174] multi_finger_inv_9
  Xgate_2_175_0 vdd vss y_b[175] y[175] multi_finger_inv_9
  Xgate_2_176_0 vdd vss y_b[176] y[176] multi_finger_inv_9
  Xgate_2_177_0 vdd vss y_b[177] y[177] multi_finger_inv_9
  Xgate_2_178_0 vdd vss y_b[178] y[178] multi_finger_inv_9
  Xgate_2_179_0 vdd vss y_b[179] y[179] multi_finger_inv_9
  Xgate_2_180_0 vdd vss y_b[180] y[180] multi_finger_inv_9
  Xgate_2_181_0 vdd vss y_b[181] y[181] multi_finger_inv_9
  Xgate_2_182_0 vdd vss y_b[182] y[182] multi_finger_inv_9
  Xgate_2_183_0 vdd vss y_b[183] y[183] multi_finger_inv_9
  Xgate_2_184_0 vdd vss y_b[184] y[184] multi_finger_inv_9
  Xgate_2_185_0 vdd vss y_b[185] y[185] multi_finger_inv_9
  Xgate_2_186_0 vdd vss y_b[186] y[186] multi_finger_inv_9
  Xgate_2_187_0 vdd vss y_b[187] y[187] multi_finger_inv_9
  Xgate_2_188_0 vdd vss y_b[188] y[188] multi_finger_inv_9
  Xgate_2_189_0 vdd vss y_b[189] y[189] multi_finger_inv_9
  Xgate_2_190_0 vdd vss y_b[190] y[190] multi_finger_inv_9
  Xgate_2_191_0 vdd vss y_b[191] y[191] multi_finger_inv_9
  Xgate_2_192_0 vdd vss y_b[192] y[192] multi_finger_inv_9
  Xgate_2_193_0 vdd vss y_b[193] y[193] multi_finger_inv_9
  Xgate_2_194_0 vdd vss y_b[194] y[194] multi_finger_inv_9
  Xgate_2_195_0 vdd vss y_b[195] y[195] multi_finger_inv_9
  Xgate_2_196_0 vdd vss y_b[196] y[196] multi_finger_inv_9
  Xgate_2_197_0 vdd vss y_b[197] y[197] multi_finger_inv_9
  Xgate_2_198_0 vdd vss y_b[198] y[198] multi_finger_inv_9
  Xgate_2_199_0 vdd vss y_b[199] y[199] multi_finger_inv_9
  Xgate_2_200_0 vdd vss y_b[200] y[200] multi_finger_inv_9
  Xgate_2_201_0 vdd vss y_b[201] y[201] multi_finger_inv_9
  Xgate_2_202_0 vdd vss y_b[202] y[202] multi_finger_inv_9
  Xgate_2_203_0 vdd vss y_b[203] y[203] multi_finger_inv_9
  Xgate_2_204_0 vdd vss y_b[204] y[204] multi_finger_inv_9
  Xgate_2_205_0 vdd vss y_b[205] y[205] multi_finger_inv_9
  Xgate_2_206_0 vdd vss y_b[206] y[206] multi_finger_inv_9
  Xgate_2_207_0 vdd vss y_b[207] y[207] multi_finger_inv_9
  Xgate_2_208_0 vdd vss y_b[208] y[208] multi_finger_inv_9
  Xgate_2_209_0 vdd vss y_b[209] y[209] multi_finger_inv_9
  Xgate_2_210_0 vdd vss y_b[210] y[210] multi_finger_inv_9
  Xgate_2_211_0 vdd vss y_b[211] y[211] multi_finger_inv_9
  Xgate_2_212_0 vdd vss y_b[212] y[212] multi_finger_inv_9
  Xgate_2_213_0 vdd vss y_b[213] y[213] multi_finger_inv_9
  Xgate_2_214_0 vdd vss y_b[214] y[214] multi_finger_inv_9
  Xgate_2_215_0 vdd vss y_b[215] y[215] multi_finger_inv_9
  Xgate_2_216_0 vdd vss y_b[216] y[216] multi_finger_inv_9
  Xgate_2_217_0 vdd vss y_b[217] y[217] multi_finger_inv_9
  Xgate_2_218_0 vdd vss y_b[218] y[218] multi_finger_inv_9
  Xgate_2_219_0 vdd vss y_b[219] y[219] multi_finger_inv_9
  Xgate_2_220_0 vdd vss y_b[220] y[220] multi_finger_inv_9
  Xgate_2_221_0 vdd vss y_b[221] y[221] multi_finger_inv_9
  Xgate_2_222_0 vdd vss y_b[222] y[222] multi_finger_inv_9
  Xgate_2_223_0 vdd vss y_b[223] y[223] multi_finger_inv_9
  Xgate_2_224_0 vdd vss y_b[224] y[224] multi_finger_inv_9
  Xgate_2_225_0 vdd vss y_b[225] y[225] multi_finger_inv_9
  Xgate_2_226_0 vdd vss y_b[226] y[226] multi_finger_inv_9
  Xgate_2_227_0 vdd vss y_b[227] y[227] multi_finger_inv_9
  Xgate_2_228_0 vdd vss y_b[228] y[228] multi_finger_inv_9
  Xgate_2_229_0 vdd vss y_b[229] y[229] multi_finger_inv_9
  Xgate_2_230_0 vdd vss y_b[230] y[230] multi_finger_inv_9
  Xgate_2_231_0 vdd vss y_b[231] y[231] multi_finger_inv_9
  Xgate_2_232_0 vdd vss y_b[232] y[232] multi_finger_inv_9
  Xgate_2_233_0 vdd vss y_b[233] y[233] multi_finger_inv_9
  Xgate_2_234_0 vdd vss y_b[234] y[234] multi_finger_inv_9
  Xgate_2_235_0 vdd vss y_b[235] y[235] multi_finger_inv_9
  Xgate_2_236_0 vdd vss y_b[236] y[236] multi_finger_inv_9
  Xgate_2_237_0 vdd vss y_b[237] y[237] multi_finger_inv_9
  Xgate_2_238_0 vdd vss y_b[238] y[238] multi_finger_inv_9
  Xgate_2_239_0 vdd vss y_b[239] y[239] multi_finger_inv_9
  Xgate_2_240_0 vdd vss y_b[240] y[240] multi_finger_inv_9
  Xgate_2_241_0 vdd vss y_b[241] y[241] multi_finger_inv_9
  Xgate_2_242_0 vdd vss y_b[242] y[242] multi_finger_inv_9
  Xgate_2_243_0 vdd vss y_b[243] y[243] multi_finger_inv_9
  Xgate_2_244_0 vdd vss y_b[244] y[244] multi_finger_inv_9
  Xgate_2_245_0 vdd vss y_b[245] y[245] multi_finger_inv_9
  Xgate_2_246_0 vdd vss y_b[246] y[246] multi_finger_inv_9
  Xgate_2_247_0 vdd vss y_b[247] y[247] multi_finger_inv_9
  Xgate_2_248_0 vdd vss y_b[248] y[248] multi_finger_inv_9
  Xgate_2_249_0 vdd vss y_b[249] y[249] multi_finger_inv_9
  Xgate_2_250_0 vdd vss y_b[250] y[250] multi_finger_inv_9
  Xgate_2_251_0 vdd vss y_b[251] y[251] multi_finger_inv_9
  Xgate_2_252_0 vdd vss y_b[252] y[252] multi_finger_inv_9
  Xgate_2_253_0 vdd vss y_b[253] y[253] multi_finger_inv_9
  Xgate_2_254_0 vdd vss y_b[254] y[254] multi_finger_inv_9
  Xgate_2_255_0 vdd vss y_b[255] y[255] multi_finger_inv_9

.ENDS decoder_stage_5

.SUBCKT decoder vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y[128] y[129] y[130] y[131] y[132] y[133] y[134] y[135] y[136] y[137] y[138] y[139] y[140] y[141] y[142] y[143] y[144] y[145] y[146] y[147] y[148] y[149] y[150] y[151] y[152] y[153] y[154] y[155] y[156] y[157] y[158] y[159] y[160] y[161] y[162] y[163] y[164] y[165] y[166] y[167] y[168] y[169] y[170] y[171] y[172] y[173] y[174] y[175] y[176] y[177] y[178] y[179] y[180] y[181] y[182] y[183] y[184] y[185] y[186] y[187] y[188] y[189] y[190] y[191] y[192] y[193] y[194] y[195] y[196] y[197] y[198] y[199] y[200] y[201] y[202] y[203] y[204] y[205] y[206] y[207] y[208] y[209] y[210] y[211] y[212] y[213] y[214] y[215] y[216] y[217] y[218] y[219] y[220] y[221] y[222] y[223] y[224] y[225] y[226] y[227] y[228] y[229] y[230] y[231] y[232] y[233] y[234] y[235] y[236] y[237] y[238] y[239] y[240] y[241] y[242] y[243] y[244] y[245] y[246] y[247] y[248] y[249] y[250] y[251] y[252] y[253] y[254] y[255] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] y_b[128] y_b[129] y_b[130] y_b[131] y_b[132] y_b[133] y_b[134] y_b[135] y_b[136] y_b[137] y_b[138] y_b[139] y_b[140] y_b[141] y_b[142] y_b[143] y_b[144] y_b[145] y_b[146] y_b[147] y_b[148] y_b[149] y_b[150] y_b[151] y_b[152] y_b[153] y_b[154] y_b[155] y_b[156] y_b[157] y_b[158] y_b[159] y_b[160] y_b[161] y_b[162] y_b[163] y_b[164] y_b[165] y_b[166] y_b[167] y_b[168] y_b[169] y_b[170] y_b[171] y_b[172] y_b[173] y_b[174] y_b[175] y_b[176] y_b[177] y_b[178] y_b[179] y_b[180] y_b[181] y_b[182] y_b[183] y_b[184] y_b[185] y_b[186] y_b[187] y_b[188] y_b[189] y_b[190] y_b[191] y_b[192] y_b[193] y_b[194] y_b[195] y_b[196] y_b[197] y_b[198] y_b[199] y_b[200] y_b[201] y_b[202] y_b[203] y_b[204] y_b[205] y_b[206] y_b[207] y_b[208] y_b[209] y_b[210] y_b[211] y_b[212] y_b[213] y_b[214] y_b[215] y_b[216] y_b[217] y_b[218] y_b[219] y_b[220] y_b[221] y_b[222] y_b[223] y_b[224] y_b[225] y_b[226] y_b[227] y_b[228] y_b[229] y_b[230] y_b[231] y_b[232] y_b[233] y_b[234] y_b[235] y_b[236] y_b[237] y_b[238] y_b[239] y_b[240] y_b[241] y_b[242] y_b[243] y_b[244] y_b[245] y_b[246] y_b[247] y_b[248] y_b[249] y_b[250] y_b[251] y_b[252] y_b[253] y_b[254] y_b[255] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 predecode_4_0 predecode_4_1 predecode_5_0 predecode_5_1 predecode_6_0 predecode_6_1 predecode_7_0 predecode_7_1

  X0 vdd vss child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_0[4] child_conn_0[5] child_conn_0[6] child_conn_0[7] child_conn_0[8] child_conn_0[9] child_conn_0[10] child_conn_0[11] child_conn_0[12] child_conn_0[13] child_conn_0[14] child_conn_0[15] child_noconn_0[0] child_noconn_0[1] child_noconn_0[2] child_noconn_0[3] child_noconn_0[4] child_noconn_0[5] child_noconn_0[6] child_noconn_0[7] child_noconn_0[8] child_noconn_0[9] child_noconn_0[10] child_noconn_0[11] child_noconn_0[12] child_noconn_0[13] child_noconn_0[14] child_noconn_0[15] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 decoder_2
  X0_1 vdd vss child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_conn_1[4] child_conn_1[5] child_conn_1[6] child_conn_1[7] child_conn_1[8] child_conn_1[9] child_conn_1[10] child_conn_1[11] child_conn_1[12] child_conn_1[13] child_conn_1[14] child_conn_1[15] child_noconn_1[0] child_noconn_1[1] child_noconn_1[2] child_noconn_1[3] child_noconn_1[4] child_noconn_1[5] child_noconn_1[6] child_noconn_1[7] child_noconn_1[8] child_noconn_1[9] child_noconn_1[10] child_noconn_1[11] child_noconn_1[12] child_noconn_1[13] child_noconn_1[14] child_noconn_1[15] predecode_4_0 predecode_4_1 predecode_5_0 predecode_5_1 predecode_6_0 predecode_6_1 predecode_7_0 predecode_7_1 decoder_2
  X0_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y[64] y[65] y[66] y[67] y[68] y[69] y[70] y[71] y[72] y[73] y[74] y[75] y[76] y[77] y[78] y[79] y[80] y[81] y[82] y[83] y[84] y[85] y[86] y[87] y[88] y[89] y[90] y[91] y[92] y[93] y[94] y[95] y[96] y[97] y[98] y[99] y[100] y[101] y[102] y[103] y[104] y[105] y[106] y[107] y[108] y[109] y[110] y[111] y[112] y[113] y[114] y[115] y[116] y[117] y[118] y[119] y[120] y[121] y[122] y[123] y[124] y[125] y[126] y[127] y[128] y[129] y[130] y[131] y[132] y[133] y[134] y[135] y[136] y[137] y[138] y[139] y[140] y[141] y[142] y[143] y[144] y[145] y[146] y[147] y[148] y[149] y[150] y[151] y[152] y[153] y[154] y[155] y[156] y[157] y[158] y[159] y[160] y[161] y[162] y[163] y[164] y[165] y[166] y[167] y[168] y[169] y[170] y[171] y[172] y[173] y[174] y[175] y[176] y[177] y[178] y[179] y[180] y[181] y[182] y[183] y[184] y[185] y[186] y[187] y[188] y[189] y[190] y[191] y[192] y[193] y[194] y[195] y[196] y[197] y[198] y[199] y[200] y[201] y[202] y[203] y[204] y[205] y[206] y[207] y[208] y[209] y[210] y[211] y[212] y[213] y[214] y[215] y[216] y[217] y[218] y[219] y[220] y[221] y[222] y[223] y[224] y[225] y[226] y[227] y[228] y[229] y[230] y[231] y[232] y[233] y[234] y[235] y[236] y[237] y[238] y[239] y[240] y[241] y[242] y[243] y[244] y[245] y[246] y[247] y[248] y[249] y[250] y[251] y[252] y[253] y[254] y[255] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] y_b[64] y_b[65] y_b[66] y_b[67] y_b[68] y_b[69] y_b[70] y_b[71] y_b[72] y_b[73] y_b[74] y_b[75] y_b[76] y_b[77] y_b[78] y_b[79] y_b[80] y_b[81] y_b[82] y_b[83] y_b[84] y_b[85] y_b[86] y_b[87] y_b[88] y_b[89] y_b[90] y_b[91] y_b[92] y_b[93] y_b[94] y_b[95] y_b[96] y_b[97] y_b[98] y_b[99] y_b[100] y_b[101] y_b[102] y_b[103] y_b[104] y_b[105] y_b[106] y_b[107] y_b[108] y_b[109] y_b[110] y_b[111] y_b[112] y_b[113] y_b[114] y_b[115] y_b[116] y_b[117] y_b[118] y_b[119] y_b[120] y_b[121] y_b[122] y_b[123] y_b[124] y_b[125] y_b[126] y_b[127] y_b[128] y_b[129] y_b[130] y_b[131] y_b[132] y_b[133] y_b[134] y_b[135] y_b[136] y_b[137] y_b[138] y_b[139] y_b[140] y_b[141] y_b[142] y_b[143] y_b[144] y_b[145] y_b[146] y_b[147] y_b[148] y_b[149] y_b[150] y_b[151] y_b[152] y_b[153] y_b[154] y_b[155] y_b[156] y_b[157] y_b[158] y_b[159] y_b[160] y_b[161] y_b[162] y_b[163] y_b[164] y_b[165] y_b[166] y_b[167] y_b[168] y_b[169] y_b[170] y_b[171] y_b[172] y_b[173] y_b[174] y_b[175] y_b[176] y_b[177] y_b[178] y_b[179] y_b[180] y_b[181] y_b[182] y_b[183] y_b[184] y_b[185] y_b[186] y_b[187] y_b[188] y_b[189] y_b[190] y_b[191] y_b[192] y_b[193] y_b[194] y_b[195] y_b[196] y_b[197] y_b[198] y_b[199] y_b[200] y_b[201] y_b[202] y_b[203] y_b[204] y_b[205] y_b[206] y_b[207] y_b[208] y_b[209] y_b[210] y_b[211] y_b[212] y_b[213] y_b[214] y_b[215] y_b[216] y_b[217] y_b[218] y_b[219] y_b[220] y_b[221] y_b[222] y_b[223] y_b[224] y_b[225] y_b[226] y_b[227] y_b[228] y_b[229] y_b[230] y_b[231] y_b[232] y_b[233] y_b[234] y_b[235] y_b[236] y_b[237] y_b[238] y_b[239] y_b[240] y_b[241] y_b[242] y_b[243] y_b[244] y_b[245] y_b[246] y_b[247] y_b[248] y_b[249] y_b[250] y_b[251] y_b[252] y_b[253] y_b[254] y_b[255] child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_0[4] child_conn_0[5] child_conn_0[6] child_conn_0[7] child_conn_0[8] child_conn_0[9] child_conn_0[10] child_conn_0[11] child_conn_0[12] child_conn_0[13] child_conn_0[14] child_conn_0[15] child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_conn_1[4] child_conn_1[5] child_conn_1[6] child_conn_1[7] child_conn_1[8] child_conn_1[9] child_conn_1[10] child_conn_1[11] child_conn_1[12] child_conn_1[13] child_conn_1[14] child_conn_1[15] decoder_stage_5

.ENDS decoder

.SUBCKT sram_sp_cell BL BR VDD VSS WL VNB VPB

  X0 QB WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q QB VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 QB WL QB VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q QB VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q QB VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q QB VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell

.SUBCKT decoder_1 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  X0 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 decoder_stage_6

.ENDS decoder_1

.SUBCKT sram_sp_cell_wrapper BL BR VDD VSS WL VNB VPB

  X0 BL BR VDD VSS WL VNB VPB sram_sp_cell

.ENDS sram_sp_cell_wrapper

.SUBCKT sram_sp_colend_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_colend

.ENDS sram_sp_colend_wrapper

.SUBCKT sram_sp_hstrap BR VDD VSS BL VNB VPB

  X0 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140

  X1 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_hstrap

.SUBCKT sram_sp_hstrap_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_hstrap

.ENDS sram_sp_hstrap_wrapper

.SUBCKT sp_cell_array vdd vss dummy_bl dummy_br bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255]

  Xcell_0_0 bl[0] br[0] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_1 bl[1] br[1] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_2 bl[2] br[2] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_3 bl[3] br[3] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_4 bl[4] br[4] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_5 bl[5] br[5] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_6 bl[6] br[6] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_7 bl[7] br[7] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_8 bl[8] br[8] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_9 bl[9] br[9] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_10 bl[10] br[10] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_11 bl[11] br[11] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_12 bl[12] br[12] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_13 bl[13] br[13] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_14 bl[14] br[14] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_15 bl[15] br[15] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_16 bl[16] br[16] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_17 bl[17] br[17] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_18 bl[18] br[18] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_19 bl[19] br[19] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_20 bl[20] br[20] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_21 bl[21] br[21] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_22 bl[22] br[22] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_23 bl[23] br[23] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_24 bl[24] br[24] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_25 bl[25] br[25] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_26 bl[26] br[26] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_27 bl[27] br[27] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_28 bl[28] br[28] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_29 bl[29] br[29] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_30 bl[30] br[30] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_31 bl[31] br[31] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_32 bl[32] br[32] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_33 bl[33] br[33] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_34 bl[34] br[34] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_35 bl[35] br[35] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_36 bl[36] br[36] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_37 bl[37] br[37] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_38 bl[38] br[38] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_39 bl[39] br[39] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_40 bl[40] br[40] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_41 bl[41] br[41] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_42 bl[42] br[42] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_43 bl[43] br[43] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_44 bl[44] br[44] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_45 bl[45] br[45] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_46 bl[46] br[46] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_47 bl[47] br[47] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_48 bl[48] br[48] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_49 bl[49] br[49] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_50 bl[50] br[50] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_51 bl[51] br[51] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_52 bl[52] br[52] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_53 bl[53] br[53] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_54 bl[54] br[54] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_55 bl[55] br[55] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_56 bl[56] br[56] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_57 bl[57] br[57] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_58 bl[58] br[58] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_59 bl[59] br[59] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_60 bl[60] br[60] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_61 bl[61] br[61] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_62 bl[62] br[62] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_63 bl[63] br[63] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_1_0 bl[0] br[0] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_1 bl[1] br[1] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_2 bl[2] br[2] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_3 bl[3] br[3] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_4 bl[4] br[4] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_5 bl[5] br[5] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_6 bl[6] br[6] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_7 bl[7] br[7] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_8 bl[8] br[8] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_9 bl[9] br[9] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_10 bl[10] br[10] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_11 bl[11] br[11] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_12 bl[12] br[12] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_13 bl[13] br[13] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_14 bl[14] br[14] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_15 bl[15] br[15] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_16 bl[16] br[16] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_17 bl[17] br[17] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_18 bl[18] br[18] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_19 bl[19] br[19] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_20 bl[20] br[20] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_21 bl[21] br[21] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_22 bl[22] br[22] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_23 bl[23] br[23] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_24 bl[24] br[24] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_25 bl[25] br[25] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_26 bl[26] br[26] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_27 bl[27] br[27] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_28 bl[28] br[28] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_29 bl[29] br[29] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_30 bl[30] br[30] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_31 bl[31] br[31] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_32 bl[32] br[32] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_33 bl[33] br[33] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_34 bl[34] br[34] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_35 bl[35] br[35] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_36 bl[36] br[36] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_37 bl[37] br[37] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_38 bl[38] br[38] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_39 bl[39] br[39] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_40 bl[40] br[40] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_41 bl[41] br[41] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_42 bl[42] br[42] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_43 bl[43] br[43] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_44 bl[44] br[44] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_45 bl[45] br[45] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_46 bl[46] br[46] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_47 bl[47] br[47] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_48 bl[48] br[48] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_49 bl[49] br[49] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_50 bl[50] br[50] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_51 bl[51] br[51] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_52 bl[52] br[52] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_53 bl[53] br[53] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_54 bl[54] br[54] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_55 bl[55] br[55] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_56 bl[56] br[56] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_57 bl[57] br[57] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_58 bl[58] br[58] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_59 bl[59] br[59] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_60 bl[60] br[60] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_61 bl[61] br[61] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_62 bl[62] br[62] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_63 bl[63] br[63] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_2_0 bl[0] br[0] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_1 bl[1] br[1] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_2 bl[2] br[2] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_3 bl[3] br[3] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_4 bl[4] br[4] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_5 bl[5] br[5] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_6 bl[6] br[6] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_7 bl[7] br[7] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_8 bl[8] br[8] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_9 bl[9] br[9] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_10 bl[10] br[10] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_11 bl[11] br[11] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_12 bl[12] br[12] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_13 bl[13] br[13] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_14 bl[14] br[14] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_15 bl[15] br[15] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_16 bl[16] br[16] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_17 bl[17] br[17] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_18 bl[18] br[18] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_19 bl[19] br[19] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_20 bl[20] br[20] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_21 bl[21] br[21] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_22 bl[22] br[22] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_23 bl[23] br[23] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_24 bl[24] br[24] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_25 bl[25] br[25] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_26 bl[26] br[26] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_27 bl[27] br[27] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_28 bl[28] br[28] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_29 bl[29] br[29] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_30 bl[30] br[30] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_31 bl[31] br[31] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_32 bl[32] br[32] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_33 bl[33] br[33] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_34 bl[34] br[34] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_35 bl[35] br[35] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_36 bl[36] br[36] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_37 bl[37] br[37] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_38 bl[38] br[38] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_39 bl[39] br[39] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_40 bl[40] br[40] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_41 bl[41] br[41] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_42 bl[42] br[42] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_43 bl[43] br[43] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_44 bl[44] br[44] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_45 bl[45] br[45] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_46 bl[46] br[46] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_47 bl[47] br[47] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_48 bl[48] br[48] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_49 bl[49] br[49] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_50 bl[50] br[50] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_51 bl[51] br[51] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_52 bl[52] br[52] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_53 bl[53] br[53] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_54 bl[54] br[54] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_55 bl[55] br[55] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_56 bl[56] br[56] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_57 bl[57] br[57] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_58 bl[58] br[58] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_59 bl[59] br[59] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_60 bl[60] br[60] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_61 bl[61] br[61] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_62 bl[62] br[62] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_63 bl[63] br[63] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_3_0 bl[0] br[0] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_1 bl[1] br[1] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_2 bl[2] br[2] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_3 bl[3] br[3] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_4 bl[4] br[4] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_5 bl[5] br[5] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_6 bl[6] br[6] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_7 bl[7] br[7] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_8 bl[8] br[8] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_9 bl[9] br[9] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_10 bl[10] br[10] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_11 bl[11] br[11] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_12 bl[12] br[12] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_13 bl[13] br[13] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_14 bl[14] br[14] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_15 bl[15] br[15] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_16 bl[16] br[16] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_17 bl[17] br[17] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_18 bl[18] br[18] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_19 bl[19] br[19] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_20 bl[20] br[20] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_21 bl[21] br[21] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_22 bl[22] br[22] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_23 bl[23] br[23] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_24 bl[24] br[24] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_25 bl[25] br[25] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_26 bl[26] br[26] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_27 bl[27] br[27] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_28 bl[28] br[28] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_29 bl[29] br[29] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_30 bl[30] br[30] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_31 bl[31] br[31] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_32 bl[32] br[32] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_33 bl[33] br[33] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_34 bl[34] br[34] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_35 bl[35] br[35] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_36 bl[36] br[36] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_37 bl[37] br[37] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_38 bl[38] br[38] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_39 bl[39] br[39] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_40 bl[40] br[40] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_41 bl[41] br[41] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_42 bl[42] br[42] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_43 bl[43] br[43] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_44 bl[44] br[44] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_45 bl[45] br[45] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_46 bl[46] br[46] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_47 bl[47] br[47] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_48 bl[48] br[48] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_49 bl[49] br[49] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_50 bl[50] br[50] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_51 bl[51] br[51] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_52 bl[52] br[52] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_53 bl[53] br[53] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_54 bl[54] br[54] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_55 bl[55] br[55] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_56 bl[56] br[56] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_57 bl[57] br[57] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_58 bl[58] br[58] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_59 bl[59] br[59] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_60 bl[60] br[60] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_61 bl[61] br[61] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_62 bl[62] br[62] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_63 bl[63] br[63] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_4_0 bl[0] br[0] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_1 bl[1] br[1] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_2 bl[2] br[2] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_3 bl[3] br[3] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_4 bl[4] br[4] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_5 bl[5] br[5] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_6 bl[6] br[6] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_7 bl[7] br[7] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_8 bl[8] br[8] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_9 bl[9] br[9] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_10 bl[10] br[10] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_11 bl[11] br[11] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_12 bl[12] br[12] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_13 bl[13] br[13] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_14 bl[14] br[14] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_15 bl[15] br[15] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_16 bl[16] br[16] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_17 bl[17] br[17] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_18 bl[18] br[18] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_19 bl[19] br[19] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_20 bl[20] br[20] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_21 bl[21] br[21] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_22 bl[22] br[22] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_23 bl[23] br[23] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_24 bl[24] br[24] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_25 bl[25] br[25] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_26 bl[26] br[26] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_27 bl[27] br[27] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_28 bl[28] br[28] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_29 bl[29] br[29] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_30 bl[30] br[30] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_31 bl[31] br[31] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_32 bl[32] br[32] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_33 bl[33] br[33] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_34 bl[34] br[34] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_35 bl[35] br[35] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_36 bl[36] br[36] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_37 bl[37] br[37] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_38 bl[38] br[38] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_39 bl[39] br[39] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_40 bl[40] br[40] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_41 bl[41] br[41] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_42 bl[42] br[42] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_43 bl[43] br[43] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_44 bl[44] br[44] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_45 bl[45] br[45] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_46 bl[46] br[46] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_47 bl[47] br[47] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_48 bl[48] br[48] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_49 bl[49] br[49] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_50 bl[50] br[50] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_51 bl[51] br[51] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_52 bl[52] br[52] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_53 bl[53] br[53] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_54 bl[54] br[54] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_55 bl[55] br[55] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_56 bl[56] br[56] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_57 bl[57] br[57] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_58 bl[58] br[58] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_59 bl[59] br[59] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_60 bl[60] br[60] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_61 bl[61] br[61] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_62 bl[62] br[62] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_63 bl[63] br[63] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_5_0 bl[0] br[0] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_1 bl[1] br[1] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_2 bl[2] br[2] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_3 bl[3] br[3] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_4 bl[4] br[4] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_5 bl[5] br[5] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_6 bl[6] br[6] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_7 bl[7] br[7] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_8 bl[8] br[8] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_9 bl[9] br[9] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_10 bl[10] br[10] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_11 bl[11] br[11] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_12 bl[12] br[12] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_13 bl[13] br[13] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_14 bl[14] br[14] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_15 bl[15] br[15] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_16 bl[16] br[16] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_17 bl[17] br[17] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_18 bl[18] br[18] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_19 bl[19] br[19] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_20 bl[20] br[20] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_21 bl[21] br[21] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_22 bl[22] br[22] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_23 bl[23] br[23] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_24 bl[24] br[24] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_25 bl[25] br[25] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_26 bl[26] br[26] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_27 bl[27] br[27] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_28 bl[28] br[28] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_29 bl[29] br[29] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_30 bl[30] br[30] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_31 bl[31] br[31] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_32 bl[32] br[32] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_33 bl[33] br[33] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_34 bl[34] br[34] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_35 bl[35] br[35] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_36 bl[36] br[36] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_37 bl[37] br[37] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_38 bl[38] br[38] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_39 bl[39] br[39] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_40 bl[40] br[40] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_41 bl[41] br[41] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_42 bl[42] br[42] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_43 bl[43] br[43] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_44 bl[44] br[44] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_45 bl[45] br[45] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_46 bl[46] br[46] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_47 bl[47] br[47] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_48 bl[48] br[48] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_49 bl[49] br[49] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_50 bl[50] br[50] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_51 bl[51] br[51] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_52 bl[52] br[52] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_53 bl[53] br[53] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_54 bl[54] br[54] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_55 bl[55] br[55] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_56 bl[56] br[56] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_57 bl[57] br[57] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_58 bl[58] br[58] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_59 bl[59] br[59] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_60 bl[60] br[60] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_61 bl[61] br[61] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_62 bl[62] br[62] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_63 bl[63] br[63] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_6_0 bl[0] br[0] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_1 bl[1] br[1] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_2 bl[2] br[2] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_3 bl[3] br[3] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_4 bl[4] br[4] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_5 bl[5] br[5] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_6 bl[6] br[6] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_7 bl[7] br[7] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_8 bl[8] br[8] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_9 bl[9] br[9] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_10 bl[10] br[10] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_11 bl[11] br[11] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_12 bl[12] br[12] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_13 bl[13] br[13] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_14 bl[14] br[14] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_15 bl[15] br[15] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_16 bl[16] br[16] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_17 bl[17] br[17] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_18 bl[18] br[18] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_19 bl[19] br[19] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_20 bl[20] br[20] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_21 bl[21] br[21] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_22 bl[22] br[22] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_23 bl[23] br[23] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_24 bl[24] br[24] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_25 bl[25] br[25] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_26 bl[26] br[26] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_27 bl[27] br[27] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_28 bl[28] br[28] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_29 bl[29] br[29] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_30 bl[30] br[30] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_31 bl[31] br[31] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_32 bl[32] br[32] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_33 bl[33] br[33] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_34 bl[34] br[34] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_35 bl[35] br[35] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_36 bl[36] br[36] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_37 bl[37] br[37] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_38 bl[38] br[38] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_39 bl[39] br[39] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_40 bl[40] br[40] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_41 bl[41] br[41] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_42 bl[42] br[42] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_43 bl[43] br[43] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_44 bl[44] br[44] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_45 bl[45] br[45] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_46 bl[46] br[46] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_47 bl[47] br[47] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_48 bl[48] br[48] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_49 bl[49] br[49] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_50 bl[50] br[50] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_51 bl[51] br[51] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_52 bl[52] br[52] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_53 bl[53] br[53] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_54 bl[54] br[54] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_55 bl[55] br[55] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_56 bl[56] br[56] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_57 bl[57] br[57] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_58 bl[58] br[58] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_59 bl[59] br[59] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_60 bl[60] br[60] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_61 bl[61] br[61] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_62 bl[62] br[62] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_63 bl[63] br[63] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_7_0 bl[0] br[0] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_1 bl[1] br[1] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_2 bl[2] br[2] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_3 bl[3] br[3] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_4 bl[4] br[4] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_5 bl[5] br[5] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_6 bl[6] br[6] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_7 bl[7] br[7] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_8 bl[8] br[8] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_9 bl[9] br[9] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_10 bl[10] br[10] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_11 bl[11] br[11] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_12 bl[12] br[12] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_13 bl[13] br[13] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_14 bl[14] br[14] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_15 bl[15] br[15] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_16 bl[16] br[16] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_17 bl[17] br[17] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_18 bl[18] br[18] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_19 bl[19] br[19] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_20 bl[20] br[20] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_21 bl[21] br[21] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_22 bl[22] br[22] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_23 bl[23] br[23] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_24 bl[24] br[24] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_25 bl[25] br[25] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_26 bl[26] br[26] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_27 bl[27] br[27] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_28 bl[28] br[28] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_29 bl[29] br[29] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_30 bl[30] br[30] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_31 bl[31] br[31] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_32 bl[32] br[32] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_33 bl[33] br[33] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_34 bl[34] br[34] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_35 bl[35] br[35] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_36 bl[36] br[36] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_37 bl[37] br[37] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_38 bl[38] br[38] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_39 bl[39] br[39] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_40 bl[40] br[40] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_41 bl[41] br[41] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_42 bl[42] br[42] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_43 bl[43] br[43] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_44 bl[44] br[44] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_45 bl[45] br[45] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_46 bl[46] br[46] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_47 bl[47] br[47] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_48 bl[48] br[48] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_49 bl[49] br[49] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_50 bl[50] br[50] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_51 bl[51] br[51] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_52 bl[52] br[52] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_53 bl[53] br[53] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_54 bl[54] br[54] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_55 bl[55] br[55] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_56 bl[56] br[56] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_57 bl[57] br[57] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_58 bl[58] br[58] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_59 bl[59] br[59] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_60 bl[60] br[60] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_61 bl[61] br[61] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_62 bl[62] br[62] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_63 bl[63] br[63] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_8_0 bl[0] br[0] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_1 bl[1] br[1] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_2 bl[2] br[2] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_3 bl[3] br[3] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_4 bl[4] br[4] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_5 bl[5] br[5] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_6 bl[6] br[6] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_7 bl[7] br[7] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_8 bl[8] br[8] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_9 bl[9] br[9] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_10 bl[10] br[10] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_11 bl[11] br[11] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_12 bl[12] br[12] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_13 bl[13] br[13] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_14 bl[14] br[14] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_15 bl[15] br[15] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_16 bl[16] br[16] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_17 bl[17] br[17] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_18 bl[18] br[18] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_19 bl[19] br[19] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_20 bl[20] br[20] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_21 bl[21] br[21] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_22 bl[22] br[22] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_23 bl[23] br[23] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_24 bl[24] br[24] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_25 bl[25] br[25] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_26 bl[26] br[26] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_27 bl[27] br[27] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_28 bl[28] br[28] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_29 bl[29] br[29] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_30 bl[30] br[30] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_31 bl[31] br[31] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_32 bl[32] br[32] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_33 bl[33] br[33] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_34 bl[34] br[34] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_35 bl[35] br[35] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_36 bl[36] br[36] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_37 bl[37] br[37] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_38 bl[38] br[38] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_39 bl[39] br[39] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_40 bl[40] br[40] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_41 bl[41] br[41] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_42 bl[42] br[42] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_43 bl[43] br[43] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_44 bl[44] br[44] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_45 bl[45] br[45] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_46 bl[46] br[46] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_47 bl[47] br[47] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_48 bl[48] br[48] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_49 bl[49] br[49] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_50 bl[50] br[50] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_51 bl[51] br[51] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_52 bl[52] br[52] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_53 bl[53] br[53] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_54 bl[54] br[54] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_55 bl[55] br[55] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_56 bl[56] br[56] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_57 bl[57] br[57] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_58 bl[58] br[58] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_59 bl[59] br[59] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_60 bl[60] br[60] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_61 bl[61] br[61] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_62 bl[62] br[62] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_63 bl[63] br[63] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_9_0 bl[0] br[0] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_1 bl[1] br[1] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_2 bl[2] br[2] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_3 bl[3] br[3] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_4 bl[4] br[4] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_5 bl[5] br[5] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_6 bl[6] br[6] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_7 bl[7] br[7] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_8 bl[8] br[8] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_9 bl[9] br[9] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_10 bl[10] br[10] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_11 bl[11] br[11] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_12 bl[12] br[12] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_13 bl[13] br[13] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_14 bl[14] br[14] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_15 bl[15] br[15] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_16 bl[16] br[16] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_17 bl[17] br[17] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_18 bl[18] br[18] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_19 bl[19] br[19] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_20 bl[20] br[20] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_21 bl[21] br[21] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_22 bl[22] br[22] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_23 bl[23] br[23] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_24 bl[24] br[24] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_25 bl[25] br[25] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_26 bl[26] br[26] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_27 bl[27] br[27] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_28 bl[28] br[28] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_29 bl[29] br[29] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_30 bl[30] br[30] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_31 bl[31] br[31] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_32 bl[32] br[32] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_33 bl[33] br[33] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_34 bl[34] br[34] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_35 bl[35] br[35] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_36 bl[36] br[36] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_37 bl[37] br[37] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_38 bl[38] br[38] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_39 bl[39] br[39] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_40 bl[40] br[40] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_41 bl[41] br[41] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_42 bl[42] br[42] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_43 bl[43] br[43] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_44 bl[44] br[44] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_45 bl[45] br[45] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_46 bl[46] br[46] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_47 bl[47] br[47] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_48 bl[48] br[48] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_49 bl[49] br[49] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_50 bl[50] br[50] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_51 bl[51] br[51] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_52 bl[52] br[52] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_53 bl[53] br[53] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_54 bl[54] br[54] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_55 bl[55] br[55] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_56 bl[56] br[56] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_57 bl[57] br[57] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_58 bl[58] br[58] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_59 bl[59] br[59] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_60 bl[60] br[60] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_61 bl[61] br[61] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_62 bl[62] br[62] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_63 bl[63] br[63] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_10_0 bl[0] br[0] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_1 bl[1] br[1] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_2 bl[2] br[2] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_3 bl[3] br[3] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_4 bl[4] br[4] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_5 bl[5] br[5] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_6 bl[6] br[6] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_7 bl[7] br[7] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_8 bl[8] br[8] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_9 bl[9] br[9] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_10 bl[10] br[10] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_11 bl[11] br[11] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_12 bl[12] br[12] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_13 bl[13] br[13] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_14 bl[14] br[14] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_15 bl[15] br[15] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_16 bl[16] br[16] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_17 bl[17] br[17] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_18 bl[18] br[18] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_19 bl[19] br[19] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_20 bl[20] br[20] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_21 bl[21] br[21] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_22 bl[22] br[22] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_23 bl[23] br[23] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_24 bl[24] br[24] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_25 bl[25] br[25] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_26 bl[26] br[26] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_27 bl[27] br[27] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_28 bl[28] br[28] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_29 bl[29] br[29] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_30 bl[30] br[30] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_31 bl[31] br[31] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_32 bl[32] br[32] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_33 bl[33] br[33] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_34 bl[34] br[34] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_35 bl[35] br[35] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_36 bl[36] br[36] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_37 bl[37] br[37] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_38 bl[38] br[38] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_39 bl[39] br[39] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_40 bl[40] br[40] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_41 bl[41] br[41] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_42 bl[42] br[42] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_43 bl[43] br[43] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_44 bl[44] br[44] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_45 bl[45] br[45] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_46 bl[46] br[46] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_47 bl[47] br[47] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_48 bl[48] br[48] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_49 bl[49] br[49] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_50 bl[50] br[50] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_51 bl[51] br[51] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_52 bl[52] br[52] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_53 bl[53] br[53] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_54 bl[54] br[54] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_55 bl[55] br[55] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_56 bl[56] br[56] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_57 bl[57] br[57] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_58 bl[58] br[58] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_59 bl[59] br[59] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_60 bl[60] br[60] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_61 bl[61] br[61] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_62 bl[62] br[62] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_63 bl[63] br[63] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_11_0 bl[0] br[0] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_1 bl[1] br[1] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_2 bl[2] br[2] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_3 bl[3] br[3] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_4 bl[4] br[4] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_5 bl[5] br[5] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_6 bl[6] br[6] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_7 bl[7] br[7] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_8 bl[8] br[8] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_9 bl[9] br[9] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_10 bl[10] br[10] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_11 bl[11] br[11] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_12 bl[12] br[12] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_13 bl[13] br[13] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_14 bl[14] br[14] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_15 bl[15] br[15] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_16 bl[16] br[16] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_17 bl[17] br[17] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_18 bl[18] br[18] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_19 bl[19] br[19] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_20 bl[20] br[20] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_21 bl[21] br[21] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_22 bl[22] br[22] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_23 bl[23] br[23] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_24 bl[24] br[24] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_25 bl[25] br[25] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_26 bl[26] br[26] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_27 bl[27] br[27] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_28 bl[28] br[28] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_29 bl[29] br[29] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_30 bl[30] br[30] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_31 bl[31] br[31] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_32 bl[32] br[32] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_33 bl[33] br[33] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_34 bl[34] br[34] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_35 bl[35] br[35] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_36 bl[36] br[36] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_37 bl[37] br[37] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_38 bl[38] br[38] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_39 bl[39] br[39] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_40 bl[40] br[40] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_41 bl[41] br[41] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_42 bl[42] br[42] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_43 bl[43] br[43] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_44 bl[44] br[44] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_45 bl[45] br[45] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_46 bl[46] br[46] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_47 bl[47] br[47] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_48 bl[48] br[48] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_49 bl[49] br[49] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_50 bl[50] br[50] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_51 bl[51] br[51] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_52 bl[52] br[52] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_53 bl[53] br[53] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_54 bl[54] br[54] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_55 bl[55] br[55] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_56 bl[56] br[56] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_57 bl[57] br[57] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_58 bl[58] br[58] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_59 bl[59] br[59] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_60 bl[60] br[60] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_61 bl[61] br[61] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_62 bl[62] br[62] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_63 bl[63] br[63] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_12_0 bl[0] br[0] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_1 bl[1] br[1] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_2 bl[2] br[2] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_3 bl[3] br[3] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_4 bl[4] br[4] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_5 bl[5] br[5] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_6 bl[6] br[6] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_7 bl[7] br[7] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_8 bl[8] br[8] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_9 bl[9] br[9] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_10 bl[10] br[10] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_11 bl[11] br[11] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_12 bl[12] br[12] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_13 bl[13] br[13] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_14 bl[14] br[14] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_15 bl[15] br[15] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_16 bl[16] br[16] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_17 bl[17] br[17] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_18 bl[18] br[18] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_19 bl[19] br[19] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_20 bl[20] br[20] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_21 bl[21] br[21] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_22 bl[22] br[22] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_23 bl[23] br[23] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_24 bl[24] br[24] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_25 bl[25] br[25] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_26 bl[26] br[26] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_27 bl[27] br[27] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_28 bl[28] br[28] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_29 bl[29] br[29] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_30 bl[30] br[30] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_31 bl[31] br[31] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_32 bl[32] br[32] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_33 bl[33] br[33] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_34 bl[34] br[34] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_35 bl[35] br[35] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_36 bl[36] br[36] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_37 bl[37] br[37] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_38 bl[38] br[38] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_39 bl[39] br[39] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_40 bl[40] br[40] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_41 bl[41] br[41] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_42 bl[42] br[42] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_43 bl[43] br[43] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_44 bl[44] br[44] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_45 bl[45] br[45] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_46 bl[46] br[46] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_47 bl[47] br[47] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_48 bl[48] br[48] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_49 bl[49] br[49] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_50 bl[50] br[50] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_51 bl[51] br[51] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_52 bl[52] br[52] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_53 bl[53] br[53] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_54 bl[54] br[54] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_55 bl[55] br[55] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_56 bl[56] br[56] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_57 bl[57] br[57] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_58 bl[58] br[58] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_59 bl[59] br[59] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_60 bl[60] br[60] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_61 bl[61] br[61] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_62 bl[62] br[62] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_63 bl[63] br[63] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_13_0 bl[0] br[0] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_1 bl[1] br[1] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_2 bl[2] br[2] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_3 bl[3] br[3] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_4 bl[4] br[4] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_5 bl[5] br[5] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_6 bl[6] br[6] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_7 bl[7] br[7] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_8 bl[8] br[8] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_9 bl[9] br[9] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_10 bl[10] br[10] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_11 bl[11] br[11] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_12 bl[12] br[12] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_13 bl[13] br[13] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_14 bl[14] br[14] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_15 bl[15] br[15] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_16 bl[16] br[16] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_17 bl[17] br[17] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_18 bl[18] br[18] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_19 bl[19] br[19] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_20 bl[20] br[20] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_21 bl[21] br[21] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_22 bl[22] br[22] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_23 bl[23] br[23] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_24 bl[24] br[24] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_25 bl[25] br[25] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_26 bl[26] br[26] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_27 bl[27] br[27] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_28 bl[28] br[28] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_29 bl[29] br[29] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_30 bl[30] br[30] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_31 bl[31] br[31] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_32 bl[32] br[32] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_33 bl[33] br[33] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_34 bl[34] br[34] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_35 bl[35] br[35] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_36 bl[36] br[36] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_37 bl[37] br[37] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_38 bl[38] br[38] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_39 bl[39] br[39] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_40 bl[40] br[40] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_41 bl[41] br[41] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_42 bl[42] br[42] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_43 bl[43] br[43] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_44 bl[44] br[44] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_45 bl[45] br[45] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_46 bl[46] br[46] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_47 bl[47] br[47] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_48 bl[48] br[48] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_49 bl[49] br[49] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_50 bl[50] br[50] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_51 bl[51] br[51] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_52 bl[52] br[52] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_53 bl[53] br[53] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_54 bl[54] br[54] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_55 bl[55] br[55] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_56 bl[56] br[56] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_57 bl[57] br[57] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_58 bl[58] br[58] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_59 bl[59] br[59] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_60 bl[60] br[60] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_61 bl[61] br[61] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_62 bl[62] br[62] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_63 bl[63] br[63] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_14_0 bl[0] br[0] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_1 bl[1] br[1] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_2 bl[2] br[2] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_3 bl[3] br[3] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_4 bl[4] br[4] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_5 bl[5] br[5] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_6 bl[6] br[6] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_7 bl[7] br[7] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_8 bl[8] br[8] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_9 bl[9] br[9] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_10 bl[10] br[10] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_11 bl[11] br[11] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_12 bl[12] br[12] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_13 bl[13] br[13] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_14 bl[14] br[14] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_15 bl[15] br[15] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_16 bl[16] br[16] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_17 bl[17] br[17] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_18 bl[18] br[18] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_19 bl[19] br[19] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_20 bl[20] br[20] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_21 bl[21] br[21] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_22 bl[22] br[22] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_23 bl[23] br[23] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_24 bl[24] br[24] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_25 bl[25] br[25] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_26 bl[26] br[26] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_27 bl[27] br[27] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_28 bl[28] br[28] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_29 bl[29] br[29] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_30 bl[30] br[30] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_31 bl[31] br[31] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_32 bl[32] br[32] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_33 bl[33] br[33] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_34 bl[34] br[34] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_35 bl[35] br[35] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_36 bl[36] br[36] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_37 bl[37] br[37] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_38 bl[38] br[38] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_39 bl[39] br[39] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_40 bl[40] br[40] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_41 bl[41] br[41] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_42 bl[42] br[42] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_43 bl[43] br[43] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_44 bl[44] br[44] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_45 bl[45] br[45] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_46 bl[46] br[46] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_47 bl[47] br[47] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_48 bl[48] br[48] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_49 bl[49] br[49] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_50 bl[50] br[50] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_51 bl[51] br[51] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_52 bl[52] br[52] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_53 bl[53] br[53] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_54 bl[54] br[54] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_55 bl[55] br[55] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_56 bl[56] br[56] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_57 bl[57] br[57] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_58 bl[58] br[58] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_59 bl[59] br[59] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_60 bl[60] br[60] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_61 bl[61] br[61] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_62 bl[62] br[62] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_63 bl[63] br[63] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_15_0 bl[0] br[0] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_1 bl[1] br[1] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_2 bl[2] br[2] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_3 bl[3] br[3] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_4 bl[4] br[4] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_5 bl[5] br[5] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_6 bl[6] br[6] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_7 bl[7] br[7] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_8 bl[8] br[8] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_9 bl[9] br[9] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_10 bl[10] br[10] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_11 bl[11] br[11] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_12 bl[12] br[12] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_13 bl[13] br[13] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_14 bl[14] br[14] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_15 bl[15] br[15] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_16 bl[16] br[16] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_17 bl[17] br[17] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_18 bl[18] br[18] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_19 bl[19] br[19] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_20 bl[20] br[20] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_21 bl[21] br[21] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_22 bl[22] br[22] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_23 bl[23] br[23] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_24 bl[24] br[24] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_25 bl[25] br[25] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_26 bl[26] br[26] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_27 bl[27] br[27] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_28 bl[28] br[28] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_29 bl[29] br[29] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_30 bl[30] br[30] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_31 bl[31] br[31] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_32 bl[32] br[32] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_33 bl[33] br[33] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_34 bl[34] br[34] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_35 bl[35] br[35] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_36 bl[36] br[36] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_37 bl[37] br[37] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_38 bl[38] br[38] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_39 bl[39] br[39] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_40 bl[40] br[40] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_41 bl[41] br[41] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_42 bl[42] br[42] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_43 bl[43] br[43] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_44 bl[44] br[44] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_45 bl[45] br[45] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_46 bl[46] br[46] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_47 bl[47] br[47] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_48 bl[48] br[48] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_49 bl[49] br[49] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_50 bl[50] br[50] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_51 bl[51] br[51] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_52 bl[52] br[52] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_53 bl[53] br[53] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_54 bl[54] br[54] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_55 bl[55] br[55] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_56 bl[56] br[56] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_57 bl[57] br[57] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_58 bl[58] br[58] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_59 bl[59] br[59] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_60 bl[60] br[60] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_61 bl[61] br[61] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_62 bl[62] br[62] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_63 bl[63] br[63] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_16_0 bl[0] br[0] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_1 bl[1] br[1] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_2 bl[2] br[2] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_3 bl[3] br[3] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_4 bl[4] br[4] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_5 bl[5] br[5] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_6 bl[6] br[6] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_7 bl[7] br[7] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_8 bl[8] br[8] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_9 bl[9] br[9] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_10 bl[10] br[10] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_11 bl[11] br[11] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_12 bl[12] br[12] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_13 bl[13] br[13] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_14 bl[14] br[14] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_15 bl[15] br[15] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_16 bl[16] br[16] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_17 bl[17] br[17] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_18 bl[18] br[18] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_19 bl[19] br[19] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_20 bl[20] br[20] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_21 bl[21] br[21] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_22 bl[22] br[22] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_23 bl[23] br[23] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_24 bl[24] br[24] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_25 bl[25] br[25] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_26 bl[26] br[26] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_27 bl[27] br[27] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_28 bl[28] br[28] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_29 bl[29] br[29] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_30 bl[30] br[30] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_31 bl[31] br[31] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_32 bl[32] br[32] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_33 bl[33] br[33] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_34 bl[34] br[34] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_35 bl[35] br[35] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_36 bl[36] br[36] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_37 bl[37] br[37] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_38 bl[38] br[38] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_39 bl[39] br[39] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_40 bl[40] br[40] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_41 bl[41] br[41] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_42 bl[42] br[42] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_43 bl[43] br[43] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_44 bl[44] br[44] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_45 bl[45] br[45] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_46 bl[46] br[46] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_47 bl[47] br[47] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_48 bl[48] br[48] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_49 bl[49] br[49] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_50 bl[50] br[50] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_51 bl[51] br[51] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_52 bl[52] br[52] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_53 bl[53] br[53] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_54 bl[54] br[54] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_55 bl[55] br[55] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_56 bl[56] br[56] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_57 bl[57] br[57] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_58 bl[58] br[58] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_59 bl[59] br[59] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_60 bl[60] br[60] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_61 bl[61] br[61] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_62 bl[62] br[62] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_63 bl[63] br[63] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_17_0 bl[0] br[0] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_1 bl[1] br[1] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_2 bl[2] br[2] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_3 bl[3] br[3] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_4 bl[4] br[4] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_5 bl[5] br[5] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_6 bl[6] br[6] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_7 bl[7] br[7] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_8 bl[8] br[8] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_9 bl[9] br[9] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_10 bl[10] br[10] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_11 bl[11] br[11] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_12 bl[12] br[12] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_13 bl[13] br[13] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_14 bl[14] br[14] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_15 bl[15] br[15] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_16 bl[16] br[16] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_17 bl[17] br[17] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_18 bl[18] br[18] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_19 bl[19] br[19] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_20 bl[20] br[20] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_21 bl[21] br[21] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_22 bl[22] br[22] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_23 bl[23] br[23] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_24 bl[24] br[24] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_25 bl[25] br[25] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_26 bl[26] br[26] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_27 bl[27] br[27] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_28 bl[28] br[28] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_29 bl[29] br[29] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_30 bl[30] br[30] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_31 bl[31] br[31] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_32 bl[32] br[32] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_33 bl[33] br[33] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_34 bl[34] br[34] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_35 bl[35] br[35] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_36 bl[36] br[36] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_37 bl[37] br[37] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_38 bl[38] br[38] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_39 bl[39] br[39] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_40 bl[40] br[40] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_41 bl[41] br[41] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_42 bl[42] br[42] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_43 bl[43] br[43] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_44 bl[44] br[44] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_45 bl[45] br[45] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_46 bl[46] br[46] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_47 bl[47] br[47] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_48 bl[48] br[48] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_49 bl[49] br[49] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_50 bl[50] br[50] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_51 bl[51] br[51] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_52 bl[52] br[52] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_53 bl[53] br[53] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_54 bl[54] br[54] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_55 bl[55] br[55] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_56 bl[56] br[56] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_57 bl[57] br[57] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_58 bl[58] br[58] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_59 bl[59] br[59] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_60 bl[60] br[60] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_61 bl[61] br[61] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_62 bl[62] br[62] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_63 bl[63] br[63] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_18_0 bl[0] br[0] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_1 bl[1] br[1] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_2 bl[2] br[2] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_3 bl[3] br[3] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_4 bl[4] br[4] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_5 bl[5] br[5] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_6 bl[6] br[6] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_7 bl[7] br[7] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_8 bl[8] br[8] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_9 bl[9] br[9] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_10 bl[10] br[10] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_11 bl[11] br[11] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_12 bl[12] br[12] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_13 bl[13] br[13] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_14 bl[14] br[14] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_15 bl[15] br[15] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_16 bl[16] br[16] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_17 bl[17] br[17] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_18 bl[18] br[18] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_19 bl[19] br[19] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_20 bl[20] br[20] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_21 bl[21] br[21] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_22 bl[22] br[22] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_23 bl[23] br[23] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_24 bl[24] br[24] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_25 bl[25] br[25] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_26 bl[26] br[26] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_27 bl[27] br[27] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_28 bl[28] br[28] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_29 bl[29] br[29] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_30 bl[30] br[30] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_31 bl[31] br[31] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_32 bl[32] br[32] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_33 bl[33] br[33] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_34 bl[34] br[34] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_35 bl[35] br[35] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_36 bl[36] br[36] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_37 bl[37] br[37] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_38 bl[38] br[38] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_39 bl[39] br[39] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_40 bl[40] br[40] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_41 bl[41] br[41] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_42 bl[42] br[42] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_43 bl[43] br[43] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_44 bl[44] br[44] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_45 bl[45] br[45] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_46 bl[46] br[46] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_47 bl[47] br[47] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_48 bl[48] br[48] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_49 bl[49] br[49] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_50 bl[50] br[50] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_51 bl[51] br[51] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_52 bl[52] br[52] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_53 bl[53] br[53] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_54 bl[54] br[54] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_55 bl[55] br[55] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_56 bl[56] br[56] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_57 bl[57] br[57] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_58 bl[58] br[58] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_59 bl[59] br[59] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_60 bl[60] br[60] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_61 bl[61] br[61] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_62 bl[62] br[62] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_63 bl[63] br[63] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_19_0 bl[0] br[0] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_1 bl[1] br[1] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_2 bl[2] br[2] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_3 bl[3] br[3] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_4 bl[4] br[4] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_5 bl[5] br[5] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_6 bl[6] br[6] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_7 bl[7] br[7] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_8 bl[8] br[8] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_9 bl[9] br[9] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_10 bl[10] br[10] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_11 bl[11] br[11] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_12 bl[12] br[12] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_13 bl[13] br[13] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_14 bl[14] br[14] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_15 bl[15] br[15] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_16 bl[16] br[16] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_17 bl[17] br[17] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_18 bl[18] br[18] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_19 bl[19] br[19] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_20 bl[20] br[20] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_21 bl[21] br[21] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_22 bl[22] br[22] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_23 bl[23] br[23] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_24 bl[24] br[24] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_25 bl[25] br[25] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_26 bl[26] br[26] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_27 bl[27] br[27] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_28 bl[28] br[28] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_29 bl[29] br[29] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_30 bl[30] br[30] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_31 bl[31] br[31] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_32 bl[32] br[32] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_33 bl[33] br[33] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_34 bl[34] br[34] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_35 bl[35] br[35] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_36 bl[36] br[36] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_37 bl[37] br[37] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_38 bl[38] br[38] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_39 bl[39] br[39] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_40 bl[40] br[40] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_41 bl[41] br[41] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_42 bl[42] br[42] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_43 bl[43] br[43] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_44 bl[44] br[44] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_45 bl[45] br[45] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_46 bl[46] br[46] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_47 bl[47] br[47] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_48 bl[48] br[48] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_49 bl[49] br[49] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_50 bl[50] br[50] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_51 bl[51] br[51] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_52 bl[52] br[52] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_53 bl[53] br[53] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_54 bl[54] br[54] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_55 bl[55] br[55] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_56 bl[56] br[56] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_57 bl[57] br[57] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_58 bl[58] br[58] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_59 bl[59] br[59] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_60 bl[60] br[60] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_61 bl[61] br[61] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_62 bl[62] br[62] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_63 bl[63] br[63] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_20_0 bl[0] br[0] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_1 bl[1] br[1] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_2 bl[2] br[2] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_3 bl[3] br[3] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_4 bl[4] br[4] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_5 bl[5] br[5] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_6 bl[6] br[6] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_7 bl[7] br[7] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_8 bl[8] br[8] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_9 bl[9] br[9] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_10 bl[10] br[10] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_11 bl[11] br[11] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_12 bl[12] br[12] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_13 bl[13] br[13] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_14 bl[14] br[14] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_15 bl[15] br[15] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_16 bl[16] br[16] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_17 bl[17] br[17] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_18 bl[18] br[18] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_19 bl[19] br[19] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_20 bl[20] br[20] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_21 bl[21] br[21] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_22 bl[22] br[22] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_23 bl[23] br[23] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_24 bl[24] br[24] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_25 bl[25] br[25] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_26 bl[26] br[26] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_27 bl[27] br[27] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_28 bl[28] br[28] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_29 bl[29] br[29] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_30 bl[30] br[30] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_31 bl[31] br[31] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_32 bl[32] br[32] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_33 bl[33] br[33] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_34 bl[34] br[34] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_35 bl[35] br[35] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_36 bl[36] br[36] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_37 bl[37] br[37] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_38 bl[38] br[38] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_39 bl[39] br[39] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_40 bl[40] br[40] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_41 bl[41] br[41] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_42 bl[42] br[42] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_43 bl[43] br[43] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_44 bl[44] br[44] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_45 bl[45] br[45] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_46 bl[46] br[46] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_47 bl[47] br[47] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_48 bl[48] br[48] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_49 bl[49] br[49] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_50 bl[50] br[50] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_51 bl[51] br[51] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_52 bl[52] br[52] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_53 bl[53] br[53] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_54 bl[54] br[54] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_55 bl[55] br[55] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_56 bl[56] br[56] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_57 bl[57] br[57] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_58 bl[58] br[58] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_59 bl[59] br[59] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_60 bl[60] br[60] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_61 bl[61] br[61] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_62 bl[62] br[62] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_63 bl[63] br[63] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_21_0 bl[0] br[0] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_1 bl[1] br[1] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_2 bl[2] br[2] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_3 bl[3] br[3] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_4 bl[4] br[4] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_5 bl[5] br[5] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_6 bl[6] br[6] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_7 bl[7] br[7] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_8 bl[8] br[8] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_9 bl[9] br[9] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_10 bl[10] br[10] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_11 bl[11] br[11] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_12 bl[12] br[12] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_13 bl[13] br[13] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_14 bl[14] br[14] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_15 bl[15] br[15] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_16 bl[16] br[16] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_17 bl[17] br[17] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_18 bl[18] br[18] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_19 bl[19] br[19] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_20 bl[20] br[20] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_21 bl[21] br[21] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_22 bl[22] br[22] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_23 bl[23] br[23] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_24 bl[24] br[24] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_25 bl[25] br[25] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_26 bl[26] br[26] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_27 bl[27] br[27] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_28 bl[28] br[28] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_29 bl[29] br[29] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_30 bl[30] br[30] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_31 bl[31] br[31] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_32 bl[32] br[32] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_33 bl[33] br[33] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_34 bl[34] br[34] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_35 bl[35] br[35] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_36 bl[36] br[36] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_37 bl[37] br[37] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_38 bl[38] br[38] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_39 bl[39] br[39] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_40 bl[40] br[40] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_41 bl[41] br[41] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_42 bl[42] br[42] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_43 bl[43] br[43] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_44 bl[44] br[44] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_45 bl[45] br[45] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_46 bl[46] br[46] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_47 bl[47] br[47] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_48 bl[48] br[48] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_49 bl[49] br[49] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_50 bl[50] br[50] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_51 bl[51] br[51] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_52 bl[52] br[52] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_53 bl[53] br[53] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_54 bl[54] br[54] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_55 bl[55] br[55] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_56 bl[56] br[56] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_57 bl[57] br[57] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_58 bl[58] br[58] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_59 bl[59] br[59] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_60 bl[60] br[60] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_61 bl[61] br[61] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_62 bl[62] br[62] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_63 bl[63] br[63] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_22_0 bl[0] br[0] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_1 bl[1] br[1] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_2 bl[2] br[2] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_3 bl[3] br[3] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_4 bl[4] br[4] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_5 bl[5] br[5] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_6 bl[6] br[6] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_7 bl[7] br[7] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_8 bl[8] br[8] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_9 bl[9] br[9] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_10 bl[10] br[10] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_11 bl[11] br[11] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_12 bl[12] br[12] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_13 bl[13] br[13] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_14 bl[14] br[14] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_15 bl[15] br[15] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_16 bl[16] br[16] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_17 bl[17] br[17] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_18 bl[18] br[18] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_19 bl[19] br[19] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_20 bl[20] br[20] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_21 bl[21] br[21] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_22 bl[22] br[22] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_23 bl[23] br[23] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_24 bl[24] br[24] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_25 bl[25] br[25] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_26 bl[26] br[26] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_27 bl[27] br[27] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_28 bl[28] br[28] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_29 bl[29] br[29] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_30 bl[30] br[30] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_31 bl[31] br[31] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_32 bl[32] br[32] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_33 bl[33] br[33] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_34 bl[34] br[34] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_35 bl[35] br[35] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_36 bl[36] br[36] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_37 bl[37] br[37] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_38 bl[38] br[38] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_39 bl[39] br[39] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_40 bl[40] br[40] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_41 bl[41] br[41] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_42 bl[42] br[42] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_43 bl[43] br[43] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_44 bl[44] br[44] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_45 bl[45] br[45] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_46 bl[46] br[46] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_47 bl[47] br[47] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_48 bl[48] br[48] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_49 bl[49] br[49] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_50 bl[50] br[50] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_51 bl[51] br[51] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_52 bl[52] br[52] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_53 bl[53] br[53] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_54 bl[54] br[54] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_55 bl[55] br[55] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_56 bl[56] br[56] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_57 bl[57] br[57] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_58 bl[58] br[58] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_59 bl[59] br[59] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_60 bl[60] br[60] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_61 bl[61] br[61] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_62 bl[62] br[62] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_63 bl[63] br[63] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_23_0 bl[0] br[0] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_1 bl[1] br[1] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_2 bl[2] br[2] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_3 bl[3] br[3] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_4 bl[4] br[4] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_5 bl[5] br[5] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_6 bl[6] br[6] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_7 bl[7] br[7] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_8 bl[8] br[8] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_9 bl[9] br[9] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_10 bl[10] br[10] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_11 bl[11] br[11] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_12 bl[12] br[12] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_13 bl[13] br[13] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_14 bl[14] br[14] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_15 bl[15] br[15] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_16 bl[16] br[16] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_17 bl[17] br[17] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_18 bl[18] br[18] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_19 bl[19] br[19] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_20 bl[20] br[20] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_21 bl[21] br[21] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_22 bl[22] br[22] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_23 bl[23] br[23] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_24 bl[24] br[24] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_25 bl[25] br[25] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_26 bl[26] br[26] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_27 bl[27] br[27] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_28 bl[28] br[28] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_29 bl[29] br[29] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_30 bl[30] br[30] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_31 bl[31] br[31] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_32 bl[32] br[32] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_33 bl[33] br[33] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_34 bl[34] br[34] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_35 bl[35] br[35] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_36 bl[36] br[36] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_37 bl[37] br[37] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_38 bl[38] br[38] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_39 bl[39] br[39] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_40 bl[40] br[40] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_41 bl[41] br[41] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_42 bl[42] br[42] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_43 bl[43] br[43] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_44 bl[44] br[44] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_45 bl[45] br[45] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_46 bl[46] br[46] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_47 bl[47] br[47] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_48 bl[48] br[48] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_49 bl[49] br[49] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_50 bl[50] br[50] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_51 bl[51] br[51] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_52 bl[52] br[52] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_53 bl[53] br[53] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_54 bl[54] br[54] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_55 bl[55] br[55] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_56 bl[56] br[56] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_57 bl[57] br[57] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_58 bl[58] br[58] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_59 bl[59] br[59] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_60 bl[60] br[60] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_61 bl[61] br[61] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_62 bl[62] br[62] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_63 bl[63] br[63] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_24_0 bl[0] br[0] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_1 bl[1] br[1] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_2 bl[2] br[2] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_3 bl[3] br[3] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_4 bl[4] br[4] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_5 bl[5] br[5] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_6 bl[6] br[6] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_7 bl[7] br[7] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_8 bl[8] br[8] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_9 bl[9] br[9] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_10 bl[10] br[10] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_11 bl[11] br[11] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_12 bl[12] br[12] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_13 bl[13] br[13] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_14 bl[14] br[14] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_15 bl[15] br[15] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_16 bl[16] br[16] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_17 bl[17] br[17] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_18 bl[18] br[18] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_19 bl[19] br[19] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_20 bl[20] br[20] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_21 bl[21] br[21] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_22 bl[22] br[22] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_23 bl[23] br[23] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_24 bl[24] br[24] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_25 bl[25] br[25] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_26 bl[26] br[26] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_27 bl[27] br[27] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_28 bl[28] br[28] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_29 bl[29] br[29] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_30 bl[30] br[30] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_31 bl[31] br[31] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_32 bl[32] br[32] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_33 bl[33] br[33] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_34 bl[34] br[34] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_35 bl[35] br[35] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_36 bl[36] br[36] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_37 bl[37] br[37] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_38 bl[38] br[38] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_39 bl[39] br[39] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_40 bl[40] br[40] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_41 bl[41] br[41] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_42 bl[42] br[42] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_43 bl[43] br[43] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_44 bl[44] br[44] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_45 bl[45] br[45] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_46 bl[46] br[46] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_47 bl[47] br[47] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_48 bl[48] br[48] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_49 bl[49] br[49] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_50 bl[50] br[50] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_51 bl[51] br[51] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_52 bl[52] br[52] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_53 bl[53] br[53] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_54 bl[54] br[54] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_55 bl[55] br[55] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_56 bl[56] br[56] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_57 bl[57] br[57] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_58 bl[58] br[58] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_59 bl[59] br[59] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_60 bl[60] br[60] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_61 bl[61] br[61] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_62 bl[62] br[62] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_63 bl[63] br[63] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_25_0 bl[0] br[0] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_1 bl[1] br[1] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_2 bl[2] br[2] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_3 bl[3] br[3] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_4 bl[4] br[4] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_5 bl[5] br[5] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_6 bl[6] br[6] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_7 bl[7] br[7] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_8 bl[8] br[8] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_9 bl[9] br[9] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_10 bl[10] br[10] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_11 bl[11] br[11] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_12 bl[12] br[12] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_13 bl[13] br[13] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_14 bl[14] br[14] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_15 bl[15] br[15] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_16 bl[16] br[16] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_17 bl[17] br[17] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_18 bl[18] br[18] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_19 bl[19] br[19] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_20 bl[20] br[20] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_21 bl[21] br[21] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_22 bl[22] br[22] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_23 bl[23] br[23] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_24 bl[24] br[24] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_25 bl[25] br[25] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_26 bl[26] br[26] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_27 bl[27] br[27] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_28 bl[28] br[28] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_29 bl[29] br[29] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_30 bl[30] br[30] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_31 bl[31] br[31] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_32 bl[32] br[32] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_33 bl[33] br[33] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_34 bl[34] br[34] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_35 bl[35] br[35] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_36 bl[36] br[36] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_37 bl[37] br[37] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_38 bl[38] br[38] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_39 bl[39] br[39] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_40 bl[40] br[40] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_41 bl[41] br[41] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_42 bl[42] br[42] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_43 bl[43] br[43] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_44 bl[44] br[44] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_45 bl[45] br[45] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_46 bl[46] br[46] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_47 bl[47] br[47] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_48 bl[48] br[48] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_49 bl[49] br[49] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_50 bl[50] br[50] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_51 bl[51] br[51] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_52 bl[52] br[52] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_53 bl[53] br[53] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_54 bl[54] br[54] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_55 bl[55] br[55] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_56 bl[56] br[56] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_57 bl[57] br[57] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_58 bl[58] br[58] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_59 bl[59] br[59] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_60 bl[60] br[60] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_61 bl[61] br[61] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_62 bl[62] br[62] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_63 bl[63] br[63] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_26_0 bl[0] br[0] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_1 bl[1] br[1] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_2 bl[2] br[2] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_3 bl[3] br[3] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_4 bl[4] br[4] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_5 bl[5] br[5] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_6 bl[6] br[6] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_7 bl[7] br[7] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_8 bl[8] br[8] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_9 bl[9] br[9] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_10 bl[10] br[10] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_11 bl[11] br[11] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_12 bl[12] br[12] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_13 bl[13] br[13] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_14 bl[14] br[14] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_15 bl[15] br[15] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_16 bl[16] br[16] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_17 bl[17] br[17] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_18 bl[18] br[18] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_19 bl[19] br[19] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_20 bl[20] br[20] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_21 bl[21] br[21] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_22 bl[22] br[22] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_23 bl[23] br[23] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_24 bl[24] br[24] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_25 bl[25] br[25] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_26 bl[26] br[26] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_27 bl[27] br[27] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_28 bl[28] br[28] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_29 bl[29] br[29] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_30 bl[30] br[30] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_31 bl[31] br[31] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_32 bl[32] br[32] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_33 bl[33] br[33] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_34 bl[34] br[34] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_35 bl[35] br[35] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_36 bl[36] br[36] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_37 bl[37] br[37] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_38 bl[38] br[38] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_39 bl[39] br[39] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_40 bl[40] br[40] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_41 bl[41] br[41] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_42 bl[42] br[42] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_43 bl[43] br[43] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_44 bl[44] br[44] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_45 bl[45] br[45] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_46 bl[46] br[46] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_47 bl[47] br[47] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_48 bl[48] br[48] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_49 bl[49] br[49] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_50 bl[50] br[50] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_51 bl[51] br[51] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_52 bl[52] br[52] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_53 bl[53] br[53] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_54 bl[54] br[54] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_55 bl[55] br[55] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_56 bl[56] br[56] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_57 bl[57] br[57] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_58 bl[58] br[58] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_59 bl[59] br[59] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_60 bl[60] br[60] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_61 bl[61] br[61] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_62 bl[62] br[62] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_63 bl[63] br[63] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_27_0 bl[0] br[0] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_1 bl[1] br[1] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_2 bl[2] br[2] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_3 bl[3] br[3] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_4 bl[4] br[4] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_5 bl[5] br[5] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_6 bl[6] br[6] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_7 bl[7] br[7] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_8 bl[8] br[8] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_9 bl[9] br[9] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_10 bl[10] br[10] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_11 bl[11] br[11] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_12 bl[12] br[12] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_13 bl[13] br[13] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_14 bl[14] br[14] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_15 bl[15] br[15] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_16 bl[16] br[16] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_17 bl[17] br[17] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_18 bl[18] br[18] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_19 bl[19] br[19] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_20 bl[20] br[20] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_21 bl[21] br[21] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_22 bl[22] br[22] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_23 bl[23] br[23] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_24 bl[24] br[24] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_25 bl[25] br[25] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_26 bl[26] br[26] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_27 bl[27] br[27] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_28 bl[28] br[28] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_29 bl[29] br[29] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_30 bl[30] br[30] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_31 bl[31] br[31] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_32 bl[32] br[32] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_33 bl[33] br[33] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_34 bl[34] br[34] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_35 bl[35] br[35] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_36 bl[36] br[36] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_37 bl[37] br[37] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_38 bl[38] br[38] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_39 bl[39] br[39] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_40 bl[40] br[40] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_41 bl[41] br[41] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_42 bl[42] br[42] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_43 bl[43] br[43] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_44 bl[44] br[44] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_45 bl[45] br[45] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_46 bl[46] br[46] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_47 bl[47] br[47] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_48 bl[48] br[48] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_49 bl[49] br[49] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_50 bl[50] br[50] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_51 bl[51] br[51] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_52 bl[52] br[52] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_53 bl[53] br[53] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_54 bl[54] br[54] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_55 bl[55] br[55] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_56 bl[56] br[56] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_57 bl[57] br[57] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_58 bl[58] br[58] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_59 bl[59] br[59] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_60 bl[60] br[60] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_61 bl[61] br[61] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_62 bl[62] br[62] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_63 bl[63] br[63] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_28_0 bl[0] br[0] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_1 bl[1] br[1] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_2 bl[2] br[2] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_3 bl[3] br[3] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_4 bl[4] br[4] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_5 bl[5] br[5] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_6 bl[6] br[6] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_7 bl[7] br[7] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_8 bl[8] br[8] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_9 bl[9] br[9] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_10 bl[10] br[10] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_11 bl[11] br[11] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_12 bl[12] br[12] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_13 bl[13] br[13] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_14 bl[14] br[14] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_15 bl[15] br[15] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_16 bl[16] br[16] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_17 bl[17] br[17] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_18 bl[18] br[18] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_19 bl[19] br[19] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_20 bl[20] br[20] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_21 bl[21] br[21] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_22 bl[22] br[22] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_23 bl[23] br[23] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_24 bl[24] br[24] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_25 bl[25] br[25] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_26 bl[26] br[26] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_27 bl[27] br[27] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_28 bl[28] br[28] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_29 bl[29] br[29] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_30 bl[30] br[30] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_31 bl[31] br[31] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_32 bl[32] br[32] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_33 bl[33] br[33] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_34 bl[34] br[34] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_35 bl[35] br[35] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_36 bl[36] br[36] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_37 bl[37] br[37] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_38 bl[38] br[38] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_39 bl[39] br[39] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_40 bl[40] br[40] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_41 bl[41] br[41] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_42 bl[42] br[42] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_43 bl[43] br[43] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_44 bl[44] br[44] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_45 bl[45] br[45] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_46 bl[46] br[46] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_47 bl[47] br[47] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_48 bl[48] br[48] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_49 bl[49] br[49] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_50 bl[50] br[50] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_51 bl[51] br[51] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_52 bl[52] br[52] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_53 bl[53] br[53] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_54 bl[54] br[54] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_55 bl[55] br[55] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_56 bl[56] br[56] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_57 bl[57] br[57] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_58 bl[58] br[58] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_59 bl[59] br[59] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_60 bl[60] br[60] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_61 bl[61] br[61] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_62 bl[62] br[62] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_63 bl[63] br[63] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_29_0 bl[0] br[0] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_1 bl[1] br[1] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_2 bl[2] br[2] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_3 bl[3] br[3] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_4 bl[4] br[4] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_5 bl[5] br[5] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_6 bl[6] br[6] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_7 bl[7] br[7] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_8 bl[8] br[8] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_9 bl[9] br[9] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_10 bl[10] br[10] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_11 bl[11] br[11] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_12 bl[12] br[12] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_13 bl[13] br[13] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_14 bl[14] br[14] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_15 bl[15] br[15] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_16 bl[16] br[16] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_17 bl[17] br[17] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_18 bl[18] br[18] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_19 bl[19] br[19] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_20 bl[20] br[20] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_21 bl[21] br[21] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_22 bl[22] br[22] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_23 bl[23] br[23] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_24 bl[24] br[24] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_25 bl[25] br[25] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_26 bl[26] br[26] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_27 bl[27] br[27] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_28 bl[28] br[28] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_29 bl[29] br[29] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_30 bl[30] br[30] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_31 bl[31] br[31] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_32 bl[32] br[32] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_33 bl[33] br[33] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_34 bl[34] br[34] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_35 bl[35] br[35] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_36 bl[36] br[36] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_37 bl[37] br[37] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_38 bl[38] br[38] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_39 bl[39] br[39] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_40 bl[40] br[40] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_41 bl[41] br[41] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_42 bl[42] br[42] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_43 bl[43] br[43] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_44 bl[44] br[44] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_45 bl[45] br[45] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_46 bl[46] br[46] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_47 bl[47] br[47] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_48 bl[48] br[48] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_49 bl[49] br[49] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_50 bl[50] br[50] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_51 bl[51] br[51] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_52 bl[52] br[52] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_53 bl[53] br[53] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_54 bl[54] br[54] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_55 bl[55] br[55] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_56 bl[56] br[56] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_57 bl[57] br[57] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_58 bl[58] br[58] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_59 bl[59] br[59] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_60 bl[60] br[60] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_61 bl[61] br[61] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_62 bl[62] br[62] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_63 bl[63] br[63] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_30_0 bl[0] br[0] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_1 bl[1] br[1] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_2 bl[2] br[2] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_3 bl[3] br[3] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_4 bl[4] br[4] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_5 bl[5] br[5] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_6 bl[6] br[6] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_7 bl[7] br[7] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_8 bl[8] br[8] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_9 bl[9] br[9] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_10 bl[10] br[10] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_11 bl[11] br[11] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_12 bl[12] br[12] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_13 bl[13] br[13] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_14 bl[14] br[14] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_15 bl[15] br[15] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_16 bl[16] br[16] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_17 bl[17] br[17] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_18 bl[18] br[18] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_19 bl[19] br[19] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_20 bl[20] br[20] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_21 bl[21] br[21] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_22 bl[22] br[22] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_23 bl[23] br[23] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_24 bl[24] br[24] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_25 bl[25] br[25] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_26 bl[26] br[26] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_27 bl[27] br[27] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_28 bl[28] br[28] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_29 bl[29] br[29] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_30 bl[30] br[30] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_31 bl[31] br[31] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_32 bl[32] br[32] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_33 bl[33] br[33] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_34 bl[34] br[34] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_35 bl[35] br[35] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_36 bl[36] br[36] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_37 bl[37] br[37] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_38 bl[38] br[38] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_39 bl[39] br[39] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_40 bl[40] br[40] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_41 bl[41] br[41] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_42 bl[42] br[42] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_43 bl[43] br[43] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_44 bl[44] br[44] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_45 bl[45] br[45] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_46 bl[46] br[46] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_47 bl[47] br[47] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_48 bl[48] br[48] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_49 bl[49] br[49] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_50 bl[50] br[50] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_51 bl[51] br[51] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_52 bl[52] br[52] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_53 bl[53] br[53] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_54 bl[54] br[54] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_55 bl[55] br[55] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_56 bl[56] br[56] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_57 bl[57] br[57] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_58 bl[58] br[58] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_59 bl[59] br[59] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_60 bl[60] br[60] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_61 bl[61] br[61] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_62 bl[62] br[62] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_63 bl[63] br[63] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_31_0 bl[0] br[0] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_1 bl[1] br[1] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_2 bl[2] br[2] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_3 bl[3] br[3] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_4 bl[4] br[4] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_5 bl[5] br[5] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_6 bl[6] br[6] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_7 bl[7] br[7] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_8 bl[8] br[8] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_9 bl[9] br[9] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_10 bl[10] br[10] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_11 bl[11] br[11] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_12 bl[12] br[12] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_13 bl[13] br[13] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_14 bl[14] br[14] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_15 bl[15] br[15] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_16 bl[16] br[16] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_17 bl[17] br[17] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_18 bl[18] br[18] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_19 bl[19] br[19] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_20 bl[20] br[20] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_21 bl[21] br[21] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_22 bl[22] br[22] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_23 bl[23] br[23] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_24 bl[24] br[24] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_25 bl[25] br[25] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_26 bl[26] br[26] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_27 bl[27] br[27] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_28 bl[28] br[28] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_29 bl[29] br[29] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_30 bl[30] br[30] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_31 bl[31] br[31] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_32 bl[32] br[32] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_33 bl[33] br[33] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_34 bl[34] br[34] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_35 bl[35] br[35] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_36 bl[36] br[36] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_37 bl[37] br[37] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_38 bl[38] br[38] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_39 bl[39] br[39] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_40 bl[40] br[40] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_41 bl[41] br[41] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_42 bl[42] br[42] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_43 bl[43] br[43] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_44 bl[44] br[44] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_45 bl[45] br[45] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_46 bl[46] br[46] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_47 bl[47] br[47] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_48 bl[48] br[48] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_49 bl[49] br[49] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_50 bl[50] br[50] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_51 bl[51] br[51] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_52 bl[52] br[52] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_53 bl[53] br[53] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_54 bl[54] br[54] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_55 bl[55] br[55] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_56 bl[56] br[56] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_57 bl[57] br[57] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_58 bl[58] br[58] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_59 bl[59] br[59] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_60 bl[60] br[60] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_61 bl[61] br[61] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_62 bl[62] br[62] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_63 bl[63] br[63] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_32_0 bl[0] br[0] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_1 bl[1] br[1] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_2 bl[2] br[2] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_3 bl[3] br[3] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_4 bl[4] br[4] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_5 bl[5] br[5] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_6 bl[6] br[6] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_7 bl[7] br[7] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_8 bl[8] br[8] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_9 bl[9] br[9] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_10 bl[10] br[10] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_11 bl[11] br[11] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_12 bl[12] br[12] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_13 bl[13] br[13] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_14 bl[14] br[14] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_15 bl[15] br[15] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_16 bl[16] br[16] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_17 bl[17] br[17] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_18 bl[18] br[18] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_19 bl[19] br[19] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_20 bl[20] br[20] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_21 bl[21] br[21] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_22 bl[22] br[22] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_23 bl[23] br[23] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_24 bl[24] br[24] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_25 bl[25] br[25] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_26 bl[26] br[26] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_27 bl[27] br[27] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_28 bl[28] br[28] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_29 bl[29] br[29] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_30 bl[30] br[30] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_31 bl[31] br[31] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_32 bl[32] br[32] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_33 bl[33] br[33] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_34 bl[34] br[34] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_35 bl[35] br[35] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_36 bl[36] br[36] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_37 bl[37] br[37] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_38 bl[38] br[38] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_39 bl[39] br[39] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_40 bl[40] br[40] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_41 bl[41] br[41] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_42 bl[42] br[42] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_43 bl[43] br[43] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_44 bl[44] br[44] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_45 bl[45] br[45] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_46 bl[46] br[46] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_47 bl[47] br[47] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_48 bl[48] br[48] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_49 bl[49] br[49] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_50 bl[50] br[50] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_51 bl[51] br[51] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_52 bl[52] br[52] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_53 bl[53] br[53] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_54 bl[54] br[54] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_55 bl[55] br[55] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_56 bl[56] br[56] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_57 bl[57] br[57] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_58 bl[58] br[58] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_59 bl[59] br[59] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_60 bl[60] br[60] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_61 bl[61] br[61] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_62 bl[62] br[62] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_63 bl[63] br[63] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_33_0 bl[0] br[0] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_1 bl[1] br[1] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_2 bl[2] br[2] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_3 bl[3] br[3] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_4 bl[4] br[4] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_5 bl[5] br[5] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_6 bl[6] br[6] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_7 bl[7] br[7] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_8 bl[8] br[8] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_9 bl[9] br[9] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_10 bl[10] br[10] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_11 bl[11] br[11] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_12 bl[12] br[12] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_13 bl[13] br[13] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_14 bl[14] br[14] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_15 bl[15] br[15] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_16 bl[16] br[16] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_17 bl[17] br[17] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_18 bl[18] br[18] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_19 bl[19] br[19] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_20 bl[20] br[20] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_21 bl[21] br[21] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_22 bl[22] br[22] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_23 bl[23] br[23] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_24 bl[24] br[24] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_25 bl[25] br[25] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_26 bl[26] br[26] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_27 bl[27] br[27] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_28 bl[28] br[28] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_29 bl[29] br[29] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_30 bl[30] br[30] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_31 bl[31] br[31] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_32 bl[32] br[32] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_33 bl[33] br[33] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_34 bl[34] br[34] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_35 bl[35] br[35] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_36 bl[36] br[36] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_37 bl[37] br[37] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_38 bl[38] br[38] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_39 bl[39] br[39] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_40 bl[40] br[40] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_41 bl[41] br[41] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_42 bl[42] br[42] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_43 bl[43] br[43] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_44 bl[44] br[44] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_45 bl[45] br[45] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_46 bl[46] br[46] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_47 bl[47] br[47] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_48 bl[48] br[48] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_49 bl[49] br[49] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_50 bl[50] br[50] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_51 bl[51] br[51] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_52 bl[52] br[52] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_53 bl[53] br[53] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_54 bl[54] br[54] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_55 bl[55] br[55] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_56 bl[56] br[56] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_57 bl[57] br[57] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_58 bl[58] br[58] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_59 bl[59] br[59] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_60 bl[60] br[60] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_61 bl[61] br[61] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_62 bl[62] br[62] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_63 bl[63] br[63] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_34_0 bl[0] br[0] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_1 bl[1] br[1] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_2 bl[2] br[2] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_3 bl[3] br[3] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_4 bl[4] br[4] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_5 bl[5] br[5] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_6 bl[6] br[6] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_7 bl[7] br[7] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_8 bl[8] br[8] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_9 bl[9] br[9] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_10 bl[10] br[10] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_11 bl[11] br[11] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_12 bl[12] br[12] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_13 bl[13] br[13] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_14 bl[14] br[14] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_15 bl[15] br[15] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_16 bl[16] br[16] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_17 bl[17] br[17] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_18 bl[18] br[18] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_19 bl[19] br[19] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_20 bl[20] br[20] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_21 bl[21] br[21] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_22 bl[22] br[22] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_23 bl[23] br[23] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_24 bl[24] br[24] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_25 bl[25] br[25] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_26 bl[26] br[26] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_27 bl[27] br[27] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_28 bl[28] br[28] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_29 bl[29] br[29] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_30 bl[30] br[30] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_31 bl[31] br[31] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_32 bl[32] br[32] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_33 bl[33] br[33] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_34 bl[34] br[34] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_35 bl[35] br[35] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_36 bl[36] br[36] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_37 bl[37] br[37] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_38 bl[38] br[38] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_39 bl[39] br[39] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_40 bl[40] br[40] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_41 bl[41] br[41] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_42 bl[42] br[42] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_43 bl[43] br[43] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_44 bl[44] br[44] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_45 bl[45] br[45] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_46 bl[46] br[46] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_47 bl[47] br[47] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_48 bl[48] br[48] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_49 bl[49] br[49] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_50 bl[50] br[50] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_51 bl[51] br[51] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_52 bl[52] br[52] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_53 bl[53] br[53] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_54 bl[54] br[54] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_55 bl[55] br[55] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_56 bl[56] br[56] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_57 bl[57] br[57] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_58 bl[58] br[58] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_59 bl[59] br[59] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_60 bl[60] br[60] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_61 bl[61] br[61] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_62 bl[62] br[62] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_63 bl[63] br[63] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_35_0 bl[0] br[0] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_1 bl[1] br[1] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_2 bl[2] br[2] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_3 bl[3] br[3] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_4 bl[4] br[4] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_5 bl[5] br[5] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_6 bl[6] br[6] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_7 bl[7] br[7] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_8 bl[8] br[8] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_9 bl[9] br[9] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_10 bl[10] br[10] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_11 bl[11] br[11] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_12 bl[12] br[12] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_13 bl[13] br[13] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_14 bl[14] br[14] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_15 bl[15] br[15] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_16 bl[16] br[16] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_17 bl[17] br[17] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_18 bl[18] br[18] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_19 bl[19] br[19] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_20 bl[20] br[20] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_21 bl[21] br[21] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_22 bl[22] br[22] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_23 bl[23] br[23] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_24 bl[24] br[24] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_25 bl[25] br[25] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_26 bl[26] br[26] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_27 bl[27] br[27] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_28 bl[28] br[28] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_29 bl[29] br[29] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_30 bl[30] br[30] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_31 bl[31] br[31] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_32 bl[32] br[32] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_33 bl[33] br[33] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_34 bl[34] br[34] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_35 bl[35] br[35] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_36 bl[36] br[36] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_37 bl[37] br[37] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_38 bl[38] br[38] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_39 bl[39] br[39] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_40 bl[40] br[40] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_41 bl[41] br[41] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_42 bl[42] br[42] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_43 bl[43] br[43] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_44 bl[44] br[44] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_45 bl[45] br[45] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_46 bl[46] br[46] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_47 bl[47] br[47] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_48 bl[48] br[48] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_49 bl[49] br[49] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_50 bl[50] br[50] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_51 bl[51] br[51] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_52 bl[52] br[52] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_53 bl[53] br[53] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_54 bl[54] br[54] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_55 bl[55] br[55] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_56 bl[56] br[56] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_57 bl[57] br[57] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_58 bl[58] br[58] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_59 bl[59] br[59] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_60 bl[60] br[60] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_61 bl[61] br[61] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_62 bl[62] br[62] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_63 bl[63] br[63] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_36_0 bl[0] br[0] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_1 bl[1] br[1] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_2 bl[2] br[2] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_3 bl[3] br[3] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_4 bl[4] br[4] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_5 bl[5] br[5] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_6 bl[6] br[6] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_7 bl[7] br[7] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_8 bl[8] br[8] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_9 bl[9] br[9] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_10 bl[10] br[10] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_11 bl[11] br[11] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_12 bl[12] br[12] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_13 bl[13] br[13] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_14 bl[14] br[14] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_15 bl[15] br[15] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_16 bl[16] br[16] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_17 bl[17] br[17] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_18 bl[18] br[18] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_19 bl[19] br[19] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_20 bl[20] br[20] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_21 bl[21] br[21] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_22 bl[22] br[22] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_23 bl[23] br[23] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_24 bl[24] br[24] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_25 bl[25] br[25] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_26 bl[26] br[26] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_27 bl[27] br[27] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_28 bl[28] br[28] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_29 bl[29] br[29] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_30 bl[30] br[30] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_31 bl[31] br[31] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_32 bl[32] br[32] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_33 bl[33] br[33] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_34 bl[34] br[34] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_35 bl[35] br[35] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_36 bl[36] br[36] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_37 bl[37] br[37] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_38 bl[38] br[38] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_39 bl[39] br[39] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_40 bl[40] br[40] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_41 bl[41] br[41] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_42 bl[42] br[42] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_43 bl[43] br[43] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_44 bl[44] br[44] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_45 bl[45] br[45] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_46 bl[46] br[46] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_47 bl[47] br[47] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_48 bl[48] br[48] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_49 bl[49] br[49] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_50 bl[50] br[50] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_51 bl[51] br[51] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_52 bl[52] br[52] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_53 bl[53] br[53] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_54 bl[54] br[54] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_55 bl[55] br[55] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_56 bl[56] br[56] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_57 bl[57] br[57] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_58 bl[58] br[58] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_59 bl[59] br[59] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_60 bl[60] br[60] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_61 bl[61] br[61] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_62 bl[62] br[62] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_63 bl[63] br[63] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_37_0 bl[0] br[0] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_1 bl[1] br[1] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_2 bl[2] br[2] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_3 bl[3] br[3] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_4 bl[4] br[4] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_5 bl[5] br[5] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_6 bl[6] br[6] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_7 bl[7] br[7] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_8 bl[8] br[8] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_9 bl[9] br[9] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_10 bl[10] br[10] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_11 bl[11] br[11] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_12 bl[12] br[12] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_13 bl[13] br[13] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_14 bl[14] br[14] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_15 bl[15] br[15] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_16 bl[16] br[16] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_17 bl[17] br[17] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_18 bl[18] br[18] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_19 bl[19] br[19] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_20 bl[20] br[20] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_21 bl[21] br[21] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_22 bl[22] br[22] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_23 bl[23] br[23] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_24 bl[24] br[24] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_25 bl[25] br[25] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_26 bl[26] br[26] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_27 bl[27] br[27] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_28 bl[28] br[28] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_29 bl[29] br[29] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_30 bl[30] br[30] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_31 bl[31] br[31] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_32 bl[32] br[32] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_33 bl[33] br[33] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_34 bl[34] br[34] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_35 bl[35] br[35] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_36 bl[36] br[36] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_37 bl[37] br[37] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_38 bl[38] br[38] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_39 bl[39] br[39] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_40 bl[40] br[40] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_41 bl[41] br[41] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_42 bl[42] br[42] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_43 bl[43] br[43] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_44 bl[44] br[44] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_45 bl[45] br[45] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_46 bl[46] br[46] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_47 bl[47] br[47] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_48 bl[48] br[48] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_49 bl[49] br[49] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_50 bl[50] br[50] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_51 bl[51] br[51] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_52 bl[52] br[52] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_53 bl[53] br[53] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_54 bl[54] br[54] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_55 bl[55] br[55] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_56 bl[56] br[56] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_57 bl[57] br[57] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_58 bl[58] br[58] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_59 bl[59] br[59] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_60 bl[60] br[60] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_61 bl[61] br[61] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_62 bl[62] br[62] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_63 bl[63] br[63] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_38_0 bl[0] br[0] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_1 bl[1] br[1] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_2 bl[2] br[2] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_3 bl[3] br[3] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_4 bl[4] br[4] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_5 bl[5] br[5] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_6 bl[6] br[6] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_7 bl[7] br[7] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_8 bl[8] br[8] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_9 bl[9] br[9] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_10 bl[10] br[10] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_11 bl[11] br[11] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_12 bl[12] br[12] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_13 bl[13] br[13] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_14 bl[14] br[14] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_15 bl[15] br[15] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_16 bl[16] br[16] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_17 bl[17] br[17] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_18 bl[18] br[18] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_19 bl[19] br[19] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_20 bl[20] br[20] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_21 bl[21] br[21] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_22 bl[22] br[22] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_23 bl[23] br[23] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_24 bl[24] br[24] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_25 bl[25] br[25] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_26 bl[26] br[26] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_27 bl[27] br[27] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_28 bl[28] br[28] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_29 bl[29] br[29] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_30 bl[30] br[30] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_31 bl[31] br[31] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_32 bl[32] br[32] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_33 bl[33] br[33] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_34 bl[34] br[34] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_35 bl[35] br[35] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_36 bl[36] br[36] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_37 bl[37] br[37] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_38 bl[38] br[38] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_39 bl[39] br[39] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_40 bl[40] br[40] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_41 bl[41] br[41] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_42 bl[42] br[42] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_43 bl[43] br[43] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_44 bl[44] br[44] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_45 bl[45] br[45] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_46 bl[46] br[46] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_47 bl[47] br[47] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_48 bl[48] br[48] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_49 bl[49] br[49] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_50 bl[50] br[50] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_51 bl[51] br[51] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_52 bl[52] br[52] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_53 bl[53] br[53] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_54 bl[54] br[54] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_55 bl[55] br[55] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_56 bl[56] br[56] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_57 bl[57] br[57] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_58 bl[58] br[58] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_59 bl[59] br[59] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_60 bl[60] br[60] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_61 bl[61] br[61] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_62 bl[62] br[62] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_63 bl[63] br[63] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_39_0 bl[0] br[0] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_1 bl[1] br[1] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_2 bl[2] br[2] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_3 bl[3] br[3] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_4 bl[4] br[4] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_5 bl[5] br[5] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_6 bl[6] br[6] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_7 bl[7] br[7] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_8 bl[8] br[8] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_9 bl[9] br[9] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_10 bl[10] br[10] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_11 bl[11] br[11] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_12 bl[12] br[12] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_13 bl[13] br[13] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_14 bl[14] br[14] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_15 bl[15] br[15] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_16 bl[16] br[16] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_17 bl[17] br[17] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_18 bl[18] br[18] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_19 bl[19] br[19] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_20 bl[20] br[20] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_21 bl[21] br[21] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_22 bl[22] br[22] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_23 bl[23] br[23] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_24 bl[24] br[24] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_25 bl[25] br[25] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_26 bl[26] br[26] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_27 bl[27] br[27] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_28 bl[28] br[28] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_29 bl[29] br[29] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_30 bl[30] br[30] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_31 bl[31] br[31] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_32 bl[32] br[32] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_33 bl[33] br[33] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_34 bl[34] br[34] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_35 bl[35] br[35] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_36 bl[36] br[36] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_37 bl[37] br[37] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_38 bl[38] br[38] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_39 bl[39] br[39] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_40 bl[40] br[40] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_41 bl[41] br[41] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_42 bl[42] br[42] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_43 bl[43] br[43] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_44 bl[44] br[44] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_45 bl[45] br[45] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_46 bl[46] br[46] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_47 bl[47] br[47] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_48 bl[48] br[48] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_49 bl[49] br[49] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_50 bl[50] br[50] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_51 bl[51] br[51] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_52 bl[52] br[52] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_53 bl[53] br[53] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_54 bl[54] br[54] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_55 bl[55] br[55] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_56 bl[56] br[56] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_57 bl[57] br[57] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_58 bl[58] br[58] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_59 bl[59] br[59] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_60 bl[60] br[60] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_61 bl[61] br[61] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_62 bl[62] br[62] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_63 bl[63] br[63] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_40_0 bl[0] br[0] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_1 bl[1] br[1] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_2 bl[2] br[2] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_3 bl[3] br[3] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_4 bl[4] br[4] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_5 bl[5] br[5] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_6 bl[6] br[6] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_7 bl[7] br[7] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_8 bl[8] br[8] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_9 bl[9] br[9] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_10 bl[10] br[10] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_11 bl[11] br[11] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_12 bl[12] br[12] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_13 bl[13] br[13] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_14 bl[14] br[14] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_15 bl[15] br[15] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_16 bl[16] br[16] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_17 bl[17] br[17] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_18 bl[18] br[18] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_19 bl[19] br[19] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_20 bl[20] br[20] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_21 bl[21] br[21] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_22 bl[22] br[22] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_23 bl[23] br[23] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_24 bl[24] br[24] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_25 bl[25] br[25] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_26 bl[26] br[26] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_27 bl[27] br[27] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_28 bl[28] br[28] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_29 bl[29] br[29] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_30 bl[30] br[30] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_31 bl[31] br[31] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_32 bl[32] br[32] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_33 bl[33] br[33] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_34 bl[34] br[34] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_35 bl[35] br[35] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_36 bl[36] br[36] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_37 bl[37] br[37] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_38 bl[38] br[38] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_39 bl[39] br[39] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_40 bl[40] br[40] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_41 bl[41] br[41] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_42 bl[42] br[42] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_43 bl[43] br[43] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_44 bl[44] br[44] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_45 bl[45] br[45] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_46 bl[46] br[46] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_47 bl[47] br[47] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_48 bl[48] br[48] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_49 bl[49] br[49] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_50 bl[50] br[50] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_51 bl[51] br[51] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_52 bl[52] br[52] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_53 bl[53] br[53] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_54 bl[54] br[54] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_55 bl[55] br[55] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_56 bl[56] br[56] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_57 bl[57] br[57] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_58 bl[58] br[58] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_59 bl[59] br[59] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_60 bl[60] br[60] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_61 bl[61] br[61] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_62 bl[62] br[62] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_63 bl[63] br[63] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_41_0 bl[0] br[0] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_1 bl[1] br[1] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_2 bl[2] br[2] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_3 bl[3] br[3] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_4 bl[4] br[4] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_5 bl[5] br[5] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_6 bl[6] br[6] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_7 bl[7] br[7] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_8 bl[8] br[8] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_9 bl[9] br[9] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_10 bl[10] br[10] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_11 bl[11] br[11] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_12 bl[12] br[12] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_13 bl[13] br[13] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_14 bl[14] br[14] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_15 bl[15] br[15] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_16 bl[16] br[16] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_17 bl[17] br[17] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_18 bl[18] br[18] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_19 bl[19] br[19] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_20 bl[20] br[20] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_21 bl[21] br[21] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_22 bl[22] br[22] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_23 bl[23] br[23] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_24 bl[24] br[24] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_25 bl[25] br[25] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_26 bl[26] br[26] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_27 bl[27] br[27] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_28 bl[28] br[28] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_29 bl[29] br[29] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_30 bl[30] br[30] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_31 bl[31] br[31] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_32 bl[32] br[32] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_33 bl[33] br[33] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_34 bl[34] br[34] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_35 bl[35] br[35] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_36 bl[36] br[36] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_37 bl[37] br[37] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_38 bl[38] br[38] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_39 bl[39] br[39] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_40 bl[40] br[40] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_41 bl[41] br[41] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_42 bl[42] br[42] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_43 bl[43] br[43] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_44 bl[44] br[44] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_45 bl[45] br[45] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_46 bl[46] br[46] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_47 bl[47] br[47] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_48 bl[48] br[48] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_49 bl[49] br[49] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_50 bl[50] br[50] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_51 bl[51] br[51] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_52 bl[52] br[52] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_53 bl[53] br[53] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_54 bl[54] br[54] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_55 bl[55] br[55] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_56 bl[56] br[56] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_57 bl[57] br[57] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_58 bl[58] br[58] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_59 bl[59] br[59] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_60 bl[60] br[60] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_61 bl[61] br[61] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_62 bl[62] br[62] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_63 bl[63] br[63] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_42_0 bl[0] br[0] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_1 bl[1] br[1] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_2 bl[2] br[2] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_3 bl[3] br[3] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_4 bl[4] br[4] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_5 bl[5] br[5] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_6 bl[6] br[6] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_7 bl[7] br[7] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_8 bl[8] br[8] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_9 bl[9] br[9] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_10 bl[10] br[10] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_11 bl[11] br[11] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_12 bl[12] br[12] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_13 bl[13] br[13] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_14 bl[14] br[14] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_15 bl[15] br[15] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_16 bl[16] br[16] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_17 bl[17] br[17] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_18 bl[18] br[18] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_19 bl[19] br[19] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_20 bl[20] br[20] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_21 bl[21] br[21] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_22 bl[22] br[22] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_23 bl[23] br[23] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_24 bl[24] br[24] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_25 bl[25] br[25] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_26 bl[26] br[26] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_27 bl[27] br[27] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_28 bl[28] br[28] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_29 bl[29] br[29] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_30 bl[30] br[30] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_31 bl[31] br[31] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_32 bl[32] br[32] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_33 bl[33] br[33] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_34 bl[34] br[34] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_35 bl[35] br[35] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_36 bl[36] br[36] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_37 bl[37] br[37] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_38 bl[38] br[38] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_39 bl[39] br[39] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_40 bl[40] br[40] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_41 bl[41] br[41] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_42 bl[42] br[42] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_43 bl[43] br[43] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_44 bl[44] br[44] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_45 bl[45] br[45] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_46 bl[46] br[46] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_47 bl[47] br[47] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_48 bl[48] br[48] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_49 bl[49] br[49] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_50 bl[50] br[50] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_51 bl[51] br[51] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_52 bl[52] br[52] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_53 bl[53] br[53] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_54 bl[54] br[54] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_55 bl[55] br[55] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_56 bl[56] br[56] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_57 bl[57] br[57] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_58 bl[58] br[58] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_59 bl[59] br[59] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_60 bl[60] br[60] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_61 bl[61] br[61] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_62 bl[62] br[62] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_63 bl[63] br[63] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_43_0 bl[0] br[0] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_1 bl[1] br[1] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_2 bl[2] br[2] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_3 bl[3] br[3] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_4 bl[4] br[4] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_5 bl[5] br[5] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_6 bl[6] br[6] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_7 bl[7] br[7] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_8 bl[8] br[8] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_9 bl[9] br[9] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_10 bl[10] br[10] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_11 bl[11] br[11] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_12 bl[12] br[12] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_13 bl[13] br[13] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_14 bl[14] br[14] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_15 bl[15] br[15] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_16 bl[16] br[16] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_17 bl[17] br[17] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_18 bl[18] br[18] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_19 bl[19] br[19] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_20 bl[20] br[20] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_21 bl[21] br[21] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_22 bl[22] br[22] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_23 bl[23] br[23] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_24 bl[24] br[24] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_25 bl[25] br[25] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_26 bl[26] br[26] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_27 bl[27] br[27] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_28 bl[28] br[28] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_29 bl[29] br[29] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_30 bl[30] br[30] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_31 bl[31] br[31] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_32 bl[32] br[32] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_33 bl[33] br[33] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_34 bl[34] br[34] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_35 bl[35] br[35] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_36 bl[36] br[36] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_37 bl[37] br[37] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_38 bl[38] br[38] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_39 bl[39] br[39] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_40 bl[40] br[40] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_41 bl[41] br[41] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_42 bl[42] br[42] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_43 bl[43] br[43] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_44 bl[44] br[44] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_45 bl[45] br[45] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_46 bl[46] br[46] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_47 bl[47] br[47] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_48 bl[48] br[48] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_49 bl[49] br[49] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_50 bl[50] br[50] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_51 bl[51] br[51] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_52 bl[52] br[52] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_53 bl[53] br[53] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_54 bl[54] br[54] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_55 bl[55] br[55] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_56 bl[56] br[56] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_57 bl[57] br[57] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_58 bl[58] br[58] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_59 bl[59] br[59] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_60 bl[60] br[60] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_61 bl[61] br[61] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_62 bl[62] br[62] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_63 bl[63] br[63] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_44_0 bl[0] br[0] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_1 bl[1] br[1] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_2 bl[2] br[2] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_3 bl[3] br[3] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_4 bl[4] br[4] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_5 bl[5] br[5] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_6 bl[6] br[6] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_7 bl[7] br[7] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_8 bl[8] br[8] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_9 bl[9] br[9] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_10 bl[10] br[10] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_11 bl[11] br[11] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_12 bl[12] br[12] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_13 bl[13] br[13] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_14 bl[14] br[14] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_15 bl[15] br[15] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_16 bl[16] br[16] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_17 bl[17] br[17] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_18 bl[18] br[18] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_19 bl[19] br[19] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_20 bl[20] br[20] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_21 bl[21] br[21] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_22 bl[22] br[22] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_23 bl[23] br[23] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_24 bl[24] br[24] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_25 bl[25] br[25] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_26 bl[26] br[26] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_27 bl[27] br[27] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_28 bl[28] br[28] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_29 bl[29] br[29] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_30 bl[30] br[30] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_31 bl[31] br[31] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_32 bl[32] br[32] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_33 bl[33] br[33] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_34 bl[34] br[34] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_35 bl[35] br[35] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_36 bl[36] br[36] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_37 bl[37] br[37] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_38 bl[38] br[38] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_39 bl[39] br[39] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_40 bl[40] br[40] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_41 bl[41] br[41] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_42 bl[42] br[42] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_43 bl[43] br[43] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_44 bl[44] br[44] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_45 bl[45] br[45] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_46 bl[46] br[46] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_47 bl[47] br[47] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_48 bl[48] br[48] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_49 bl[49] br[49] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_50 bl[50] br[50] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_51 bl[51] br[51] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_52 bl[52] br[52] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_53 bl[53] br[53] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_54 bl[54] br[54] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_55 bl[55] br[55] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_56 bl[56] br[56] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_57 bl[57] br[57] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_58 bl[58] br[58] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_59 bl[59] br[59] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_60 bl[60] br[60] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_61 bl[61] br[61] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_62 bl[62] br[62] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_63 bl[63] br[63] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_45_0 bl[0] br[0] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_1 bl[1] br[1] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_2 bl[2] br[2] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_3 bl[3] br[3] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_4 bl[4] br[4] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_5 bl[5] br[5] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_6 bl[6] br[6] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_7 bl[7] br[7] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_8 bl[8] br[8] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_9 bl[9] br[9] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_10 bl[10] br[10] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_11 bl[11] br[11] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_12 bl[12] br[12] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_13 bl[13] br[13] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_14 bl[14] br[14] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_15 bl[15] br[15] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_16 bl[16] br[16] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_17 bl[17] br[17] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_18 bl[18] br[18] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_19 bl[19] br[19] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_20 bl[20] br[20] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_21 bl[21] br[21] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_22 bl[22] br[22] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_23 bl[23] br[23] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_24 bl[24] br[24] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_25 bl[25] br[25] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_26 bl[26] br[26] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_27 bl[27] br[27] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_28 bl[28] br[28] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_29 bl[29] br[29] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_30 bl[30] br[30] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_31 bl[31] br[31] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_32 bl[32] br[32] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_33 bl[33] br[33] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_34 bl[34] br[34] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_35 bl[35] br[35] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_36 bl[36] br[36] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_37 bl[37] br[37] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_38 bl[38] br[38] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_39 bl[39] br[39] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_40 bl[40] br[40] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_41 bl[41] br[41] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_42 bl[42] br[42] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_43 bl[43] br[43] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_44 bl[44] br[44] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_45 bl[45] br[45] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_46 bl[46] br[46] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_47 bl[47] br[47] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_48 bl[48] br[48] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_49 bl[49] br[49] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_50 bl[50] br[50] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_51 bl[51] br[51] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_52 bl[52] br[52] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_53 bl[53] br[53] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_54 bl[54] br[54] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_55 bl[55] br[55] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_56 bl[56] br[56] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_57 bl[57] br[57] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_58 bl[58] br[58] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_59 bl[59] br[59] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_60 bl[60] br[60] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_61 bl[61] br[61] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_62 bl[62] br[62] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_63 bl[63] br[63] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_46_0 bl[0] br[0] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_1 bl[1] br[1] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_2 bl[2] br[2] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_3 bl[3] br[3] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_4 bl[4] br[4] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_5 bl[5] br[5] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_6 bl[6] br[6] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_7 bl[7] br[7] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_8 bl[8] br[8] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_9 bl[9] br[9] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_10 bl[10] br[10] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_11 bl[11] br[11] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_12 bl[12] br[12] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_13 bl[13] br[13] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_14 bl[14] br[14] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_15 bl[15] br[15] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_16 bl[16] br[16] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_17 bl[17] br[17] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_18 bl[18] br[18] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_19 bl[19] br[19] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_20 bl[20] br[20] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_21 bl[21] br[21] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_22 bl[22] br[22] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_23 bl[23] br[23] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_24 bl[24] br[24] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_25 bl[25] br[25] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_26 bl[26] br[26] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_27 bl[27] br[27] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_28 bl[28] br[28] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_29 bl[29] br[29] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_30 bl[30] br[30] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_31 bl[31] br[31] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_32 bl[32] br[32] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_33 bl[33] br[33] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_34 bl[34] br[34] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_35 bl[35] br[35] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_36 bl[36] br[36] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_37 bl[37] br[37] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_38 bl[38] br[38] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_39 bl[39] br[39] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_40 bl[40] br[40] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_41 bl[41] br[41] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_42 bl[42] br[42] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_43 bl[43] br[43] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_44 bl[44] br[44] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_45 bl[45] br[45] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_46 bl[46] br[46] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_47 bl[47] br[47] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_48 bl[48] br[48] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_49 bl[49] br[49] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_50 bl[50] br[50] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_51 bl[51] br[51] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_52 bl[52] br[52] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_53 bl[53] br[53] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_54 bl[54] br[54] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_55 bl[55] br[55] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_56 bl[56] br[56] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_57 bl[57] br[57] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_58 bl[58] br[58] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_59 bl[59] br[59] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_60 bl[60] br[60] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_61 bl[61] br[61] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_62 bl[62] br[62] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_63 bl[63] br[63] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_47_0 bl[0] br[0] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_1 bl[1] br[1] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_2 bl[2] br[2] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_3 bl[3] br[3] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_4 bl[4] br[4] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_5 bl[5] br[5] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_6 bl[6] br[6] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_7 bl[7] br[7] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_8 bl[8] br[8] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_9 bl[9] br[9] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_10 bl[10] br[10] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_11 bl[11] br[11] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_12 bl[12] br[12] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_13 bl[13] br[13] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_14 bl[14] br[14] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_15 bl[15] br[15] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_16 bl[16] br[16] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_17 bl[17] br[17] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_18 bl[18] br[18] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_19 bl[19] br[19] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_20 bl[20] br[20] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_21 bl[21] br[21] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_22 bl[22] br[22] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_23 bl[23] br[23] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_24 bl[24] br[24] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_25 bl[25] br[25] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_26 bl[26] br[26] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_27 bl[27] br[27] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_28 bl[28] br[28] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_29 bl[29] br[29] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_30 bl[30] br[30] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_31 bl[31] br[31] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_32 bl[32] br[32] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_33 bl[33] br[33] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_34 bl[34] br[34] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_35 bl[35] br[35] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_36 bl[36] br[36] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_37 bl[37] br[37] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_38 bl[38] br[38] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_39 bl[39] br[39] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_40 bl[40] br[40] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_41 bl[41] br[41] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_42 bl[42] br[42] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_43 bl[43] br[43] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_44 bl[44] br[44] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_45 bl[45] br[45] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_46 bl[46] br[46] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_47 bl[47] br[47] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_48 bl[48] br[48] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_49 bl[49] br[49] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_50 bl[50] br[50] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_51 bl[51] br[51] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_52 bl[52] br[52] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_53 bl[53] br[53] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_54 bl[54] br[54] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_55 bl[55] br[55] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_56 bl[56] br[56] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_57 bl[57] br[57] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_58 bl[58] br[58] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_59 bl[59] br[59] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_60 bl[60] br[60] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_61 bl[61] br[61] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_62 bl[62] br[62] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_63 bl[63] br[63] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_48_0 bl[0] br[0] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_1 bl[1] br[1] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_2 bl[2] br[2] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_3 bl[3] br[3] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_4 bl[4] br[4] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_5 bl[5] br[5] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_6 bl[6] br[6] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_7 bl[7] br[7] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_8 bl[8] br[8] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_9 bl[9] br[9] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_10 bl[10] br[10] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_11 bl[11] br[11] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_12 bl[12] br[12] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_13 bl[13] br[13] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_14 bl[14] br[14] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_15 bl[15] br[15] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_16 bl[16] br[16] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_17 bl[17] br[17] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_18 bl[18] br[18] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_19 bl[19] br[19] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_20 bl[20] br[20] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_21 bl[21] br[21] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_22 bl[22] br[22] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_23 bl[23] br[23] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_24 bl[24] br[24] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_25 bl[25] br[25] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_26 bl[26] br[26] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_27 bl[27] br[27] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_28 bl[28] br[28] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_29 bl[29] br[29] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_30 bl[30] br[30] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_31 bl[31] br[31] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_32 bl[32] br[32] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_33 bl[33] br[33] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_34 bl[34] br[34] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_35 bl[35] br[35] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_36 bl[36] br[36] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_37 bl[37] br[37] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_38 bl[38] br[38] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_39 bl[39] br[39] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_40 bl[40] br[40] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_41 bl[41] br[41] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_42 bl[42] br[42] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_43 bl[43] br[43] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_44 bl[44] br[44] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_45 bl[45] br[45] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_46 bl[46] br[46] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_47 bl[47] br[47] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_48 bl[48] br[48] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_49 bl[49] br[49] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_50 bl[50] br[50] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_51 bl[51] br[51] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_52 bl[52] br[52] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_53 bl[53] br[53] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_54 bl[54] br[54] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_55 bl[55] br[55] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_56 bl[56] br[56] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_57 bl[57] br[57] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_58 bl[58] br[58] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_59 bl[59] br[59] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_60 bl[60] br[60] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_61 bl[61] br[61] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_62 bl[62] br[62] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_63 bl[63] br[63] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_49_0 bl[0] br[0] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_1 bl[1] br[1] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_2 bl[2] br[2] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_3 bl[3] br[3] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_4 bl[4] br[4] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_5 bl[5] br[5] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_6 bl[6] br[6] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_7 bl[7] br[7] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_8 bl[8] br[8] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_9 bl[9] br[9] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_10 bl[10] br[10] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_11 bl[11] br[11] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_12 bl[12] br[12] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_13 bl[13] br[13] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_14 bl[14] br[14] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_15 bl[15] br[15] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_16 bl[16] br[16] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_17 bl[17] br[17] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_18 bl[18] br[18] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_19 bl[19] br[19] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_20 bl[20] br[20] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_21 bl[21] br[21] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_22 bl[22] br[22] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_23 bl[23] br[23] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_24 bl[24] br[24] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_25 bl[25] br[25] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_26 bl[26] br[26] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_27 bl[27] br[27] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_28 bl[28] br[28] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_29 bl[29] br[29] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_30 bl[30] br[30] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_31 bl[31] br[31] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_32 bl[32] br[32] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_33 bl[33] br[33] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_34 bl[34] br[34] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_35 bl[35] br[35] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_36 bl[36] br[36] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_37 bl[37] br[37] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_38 bl[38] br[38] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_39 bl[39] br[39] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_40 bl[40] br[40] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_41 bl[41] br[41] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_42 bl[42] br[42] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_43 bl[43] br[43] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_44 bl[44] br[44] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_45 bl[45] br[45] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_46 bl[46] br[46] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_47 bl[47] br[47] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_48 bl[48] br[48] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_49 bl[49] br[49] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_50 bl[50] br[50] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_51 bl[51] br[51] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_52 bl[52] br[52] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_53 bl[53] br[53] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_54 bl[54] br[54] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_55 bl[55] br[55] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_56 bl[56] br[56] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_57 bl[57] br[57] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_58 bl[58] br[58] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_59 bl[59] br[59] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_60 bl[60] br[60] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_61 bl[61] br[61] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_62 bl[62] br[62] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_63 bl[63] br[63] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_50_0 bl[0] br[0] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_1 bl[1] br[1] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_2 bl[2] br[2] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_3 bl[3] br[3] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_4 bl[4] br[4] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_5 bl[5] br[5] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_6 bl[6] br[6] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_7 bl[7] br[7] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_8 bl[8] br[8] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_9 bl[9] br[9] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_10 bl[10] br[10] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_11 bl[11] br[11] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_12 bl[12] br[12] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_13 bl[13] br[13] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_14 bl[14] br[14] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_15 bl[15] br[15] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_16 bl[16] br[16] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_17 bl[17] br[17] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_18 bl[18] br[18] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_19 bl[19] br[19] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_20 bl[20] br[20] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_21 bl[21] br[21] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_22 bl[22] br[22] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_23 bl[23] br[23] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_24 bl[24] br[24] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_25 bl[25] br[25] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_26 bl[26] br[26] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_27 bl[27] br[27] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_28 bl[28] br[28] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_29 bl[29] br[29] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_30 bl[30] br[30] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_31 bl[31] br[31] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_32 bl[32] br[32] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_33 bl[33] br[33] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_34 bl[34] br[34] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_35 bl[35] br[35] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_36 bl[36] br[36] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_37 bl[37] br[37] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_38 bl[38] br[38] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_39 bl[39] br[39] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_40 bl[40] br[40] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_41 bl[41] br[41] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_42 bl[42] br[42] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_43 bl[43] br[43] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_44 bl[44] br[44] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_45 bl[45] br[45] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_46 bl[46] br[46] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_47 bl[47] br[47] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_48 bl[48] br[48] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_49 bl[49] br[49] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_50 bl[50] br[50] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_51 bl[51] br[51] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_52 bl[52] br[52] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_53 bl[53] br[53] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_54 bl[54] br[54] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_55 bl[55] br[55] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_56 bl[56] br[56] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_57 bl[57] br[57] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_58 bl[58] br[58] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_59 bl[59] br[59] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_60 bl[60] br[60] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_61 bl[61] br[61] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_62 bl[62] br[62] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_63 bl[63] br[63] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_51_0 bl[0] br[0] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_1 bl[1] br[1] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_2 bl[2] br[2] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_3 bl[3] br[3] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_4 bl[4] br[4] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_5 bl[5] br[5] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_6 bl[6] br[6] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_7 bl[7] br[7] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_8 bl[8] br[8] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_9 bl[9] br[9] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_10 bl[10] br[10] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_11 bl[11] br[11] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_12 bl[12] br[12] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_13 bl[13] br[13] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_14 bl[14] br[14] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_15 bl[15] br[15] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_16 bl[16] br[16] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_17 bl[17] br[17] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_18 bl[18] br[18] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_19 bl[19] br[19] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_20 bl[20] br[20] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_21 bl[21] br[21] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_22 bl[22] br[22] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_23 bl[23] br[23] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_24 bl[24] br[24] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_25 bl[25] br[25] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_26 bl[26] br[26] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_27 bl[27] br[27] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_28 bl[28] br[28] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_29 bl[29] br[29] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_30 bl[30] br[30] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_31 bl[31] br[31] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_32 bl[32] br[32] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_33 bl[33] br[33] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_34 bl[34] br[34] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_35 bl[35] br[35] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_36 bl[36] br[36] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_37 bl[37] br[37] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_38 bl[38] br[38] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_39 bl[39] br[39] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_40 bl[40] br[40] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_41 bl[41] br[41] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_42 bl[42] br[42] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_43 bl[43] br[43] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_44 bl[44] br[44] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_45 bl[45] br[45] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_46 bl[46] br[46] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_47 bl[47] br[47] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_48 bl[48] br[48] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_49 bl[49] br[49] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_50 bl[50] br[50] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_51 bl[51] br[51] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_52 bl[52] br[52] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_53 bl[53] br[53] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_54 bl[54] br[54] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_55 bl[55] br[55] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_56 bl[56] br[56] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_57 bl[57] br[57] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_58 bl[58] br[58] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_59 bl[59] br[59] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_60 bl[60] br[60] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_61 bl[61] br[61] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_62 bl[62] br[62] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_63 bl[63] br[63] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_52_0 bl[0] br[0] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_1 bl[1] br[1] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_2 bl[2] br[2] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_3 bl[3] br[3] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_4 bl[4] br[4] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_5 bl[5] br[5] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_6 bl[6] br[6] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_7 bl[7] br[7] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_8 bl[8] br[8] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_9 bl[9] br[9] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_10 bl[10] br[10] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_11 bl[11] br[11] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_12 bl[12] br[12] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_13 bl[13] br[13] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_14 bl[14] br[14] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_15 bl[15] br[15] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_16 bl[16] br[16] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_17 bl[17] br[17] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_18 bl[18] br[18] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_19 bl[19] br[19] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_20 bl[20] br[20] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_21 bl[21] br[21] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_22 bl[22] br[22] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_23 bl[23] br[23] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_24 bl[24] br[24] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_25 bl[25] br[25] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_26 bl[26] br[26] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_27 bl[27] br[27] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_28 bl[28] br[28] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_29 bl[29] br[29] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_30 bl[30] br[30] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_31 bl[31] br[31] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_32 bl[32] br[32] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_33 bl[33] br[33] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_34 bl[34] br[34] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_35 bl[35] br[35] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_36 bl[36] br[36] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_37 bl[37] br[37] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_38 bl[38] br[38] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_39 bl[39] br[39] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_40 bl[40] br[40] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_41 bl[41] br[41] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_42 bl[42] br[42] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_43 bl[43] br[43] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_44 bl[44] br[44] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_45 bl[45] br[45] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_46 bl[46] br[46] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_47 bl[47] br[47] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_48 bl[48] br[48] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_49 bl[49] br[49] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_50 bl[50] br[50] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_51 bl[51] br[51] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_52 bl[52] br[52] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_53 bl[53] br[53] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_54 bl[54] br[54] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_55 bl[55] br[55] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_56 bl[56] br[56] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_57 bl[57] br[57] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_58 bl[58] br[58] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_59 bl[59] br[59] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_60 bl[60] br[60] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_61 bl[61] br[61] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_62 bl[62] br[62] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_63 bl[63] br[63] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_53_0 bl[0] br[0] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_1 bl[1] br[1] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_2 bl[2] br[2] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_3 bl[3] br[3] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_4 bl[4] br[4] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_5 bl[5] br[5] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_6 bl[6] br[6] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_7 bl[7] br[7] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_8 bl[8] br[8] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_9 bl[9] br[9] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_10 bl[10] br[10] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_11 bl[11] br[11] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_12 bl[12] br[12] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_13 bl[13] br[13] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_14 bl[14] br[14] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_15 bl[15] br[15] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_16 bl[16] br[16] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_17 bl[17] br[17] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_18 bl[18] br[18] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_19 bl[19] br[19] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_20 bl[20] br[20] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_21 bl[21] br[21] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_22 bl[22] br[22] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_23 bl[23] br[23] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_24 bl[24] br[24] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_25 bl[25] br[25] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_26 bl[26] br[26] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_27 bl[27] br[27] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_28 bl[28] br[28] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_29 bl[29] br[29] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_30 bl[30] br[30] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_31 bl[31] br[31] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_32 bl[32] br[32] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_33 bl[33] br[33] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_34 bl[34] br[34] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_35 bl[35] br[35] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_36 bl[36] br[36] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_37 bl[37] br[37] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_38 bl[38] br[38] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_39 bl[39] br[39] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_40 bl[40] br[40] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_41 bl[41] br[41] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_42 bl[42] br[42] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_43 bl[43] br[43] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_44 bl[44] br[44] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_45 bl[45] br[45] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_46 bl[46] br[46] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_47 bl[47] br[47] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_48 bl[48] br[48] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_49 bl[49] br[49] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_50 bl[50] br[50] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_51 bl[51] br[51] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_52 bl[52] br[52] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_53 bl[53] br[53] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_54 bl[54] br[54] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_55 bl[55] br[55] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_56 bl[56] br[56] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_57 bl[57] br[57] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_58 bl[58] br[58] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_59 bl[59] br[59] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_60 bl[60] br[60] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_61 bl[61] br[61] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_62 bl[62] br[62] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_63 bl[63] br[63] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_54_0 bl[0] br[0] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_1 bl[1] br[1] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_2 bl[2] br[2] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_3 bl[3] br[3] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_4 bl[4] br[4] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_5 bl[5] br[5] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_6 bl[6] br[6] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_7 bl[7] br[7] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_8 bl[8] br[8] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_9 bl[9] br[9] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_10 bl[10] br[10] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_11 bl[11] br[11] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_12 bl[12] br[12] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_13 bl[13] br[13] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_14 bl[14] br[14] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_15 bl[15] br[15] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_16 bl[16] br[16] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_17 bl[17] br[17] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_18 bl[18] br[18] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_19 bl[19] br[19] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_20 bl[20] br[20] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_21 bl[21] br[21] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_22 bl[22] br[22] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_23 bl[23] br[23] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_24 bl[24] br[24] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_25 bl[25] br[25] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_26 bl[26] br[26] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_27 bl[27] br[27] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_28 bl[28] br[28] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_29 bl[29] br[29] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_30 bl[30] br[30] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_31 bl[31] br[31] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_32 bl[32] br[32] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_33 bl[33] br[33] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_34 bl[34] br[34] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_35 bl[35] br[35] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_36 bl[36] br[36] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_37 bl[37] br[37] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_38 bl[38] br[38] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_39 bl[39] br[39] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_40 bl[40] br[40] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_41 bl[41] br[41] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_42 bl[42] br[42] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_43 bl[43] br[43] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_44 bl[44] br[44] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_45 bl[45] br[45] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_46 bl[46] br[46] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_47 bl[47] br[47] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_48 bl[48] br[48] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_49 bl[49] br[49] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_50 bl[50] br[50] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_51 bl[51] br[51] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_52 bl[52] br[52] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_53 bl[53] br[53] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_54 bl[54] br[54] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_55 bl[55] br[55] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_56 bl[56] br[56] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_57 bl[57] br[57] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_58 bl[58] br[58] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_59 bl[59] br[59] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_60 bl[60] br[60] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_61 bl[61] br[61] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_62 bl[62] br[62] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_63 bl[63] br[63] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_55_0 bl[0] br[0] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_1 bl[1] br[1] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_2 bl[2] br[2] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_3 bl[3] br[3] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_4 bl[4] br[4] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_5 bl[5] br[5] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_6 bl[6] br[6] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_7 bl[7] br[7] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_8 bl[8] br[8] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_9 bl[9] br[9] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_10 bl[10] br[10] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_11 bl[11] br[11] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_12 bl[12] br[12] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_13 bl[13] br[13] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_14 bl[14] br[14] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_15 bl[15] br[15] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_16 bl[16] br[16] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_17 bl[17] br[17] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_18 bl[18] br[18] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_19 bl[19] br[19] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_20 bl[20] br[20] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_21 bl[21] br[21] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_22 bl[22] br[22] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_23 bl[23] br[23] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_24 bl[24] br[24] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_25 bl[25] br[25] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_26 bl[26] br[26] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_27 bl[27] br[27] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_28 bl[28] br[28] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_29 bl[29] br[29] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_30 bl[30] br[30] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_31 bl[31] br[31] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_32 bl[32] br[32] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_33 bl[33] br[33] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_34 bl[34] br[34] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_35 bl[35] br[35] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_36 bl[36] br[36] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_37 bl[37] br[37] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_38 bl[38] br[38] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_39 bl[39] br[39] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_40 bl[40] br[40] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_41 bl[41] br[41] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_42 bl[42] br[42] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_43 bl[43] br[43] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_44 bl[44] br[44] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_45 bl[45] br[45] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_46 bl[46] br[46] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_47 bl[47] br[47] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_48 bl[48] br[48] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_49 bl[49] br[49] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_50 bl[50] br[50] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_51 bl[51] br[51] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_52 bl[52] br[52] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_53 bl[53] br[53] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_54 bl[54] br[54] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_55 bl[55] br[55] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_56 bl[56] br[56] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_57 bl[57] br[57] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_58 bl[58] br[58] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_59 bl[59] br[59] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_60 bl[60] br[60] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_61 bl[61] br[61] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_62 bl[62] br[62] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_63 bl[63] br[63] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_56_0 bl[0] br[0] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_1 bl[1] br[1] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_2 bl[2] br[2] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_3 bl[3] br[3] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_4 bl[4] br[4] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_5 bl[5] br[5] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_6 bl[6] br[6] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_7 bl[7] br[7] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_8 bl[8] br[8] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_9 bl[9] br[9] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_10 bl[10] br[10] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_11 bl[11] br[11] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_12 bl[12] br[12] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_13 bl[13] br[13] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_14 bl[14] br[14] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_15 bl[15] br[15] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_16 bl[16] br[16] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_17 bl[17] br[17] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_18 bl[18] br[18] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_19 bl[19] br[19] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_20 bl[20] br[20] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_21 bl[21] br[21] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_22 bl[22] br[22] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_23 bl[23] br[23] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_24 bl[24] br[24] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_25 bl[25] br[25] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_26 bl[26] br[26] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_27 bl[27] br[27] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_28 bl[28] br[28] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_29 bl[29] br[29] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_30 bl[30] br[30] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_31 bl[31] br[31] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_32 bl[32] br[32] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_33 bl[33] br[33] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_34 bl[34] br[34] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_35 bl[35] br[35] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_36 bl[36] br[36] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_37 bl[37] br[37] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_38 bl[38] br[38] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_39 bl[39] br[39] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_40 bl[40] br[40] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_41 bl[41] br[41] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_42 bl[42] br[42] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_43 bl[43] br[43] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_44 bl[44] br[44] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_45 bl[45] br[45] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_46 bl[46] br[46] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_47 bl[47] br[47] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_48 bl[48] br[48] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_49 bl[49] br[49] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_50 bl[50] br[50] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_51 bl[51] br[51] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_52 bl[52] br[52] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_53 bl[53] br[53] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_54 bl[54] br[54] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_55 bl[55] br[55] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_56 bl[56] br[56] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_57 bl[57] br[57] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_58 bl[58] br[58] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_59 bl[59] br[59] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_60 bl[60] br[60] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_61 bl[61] br[61] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_62 bl[62] br[62] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_63 bl[63] br[63] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_57_0 bl[0] br[0] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_1 bl[1] br[1] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_2 bl[2] br[2] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_3 bl[3] br[3] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_4 bl[4] br[4] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_5 bl[5] br[5] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_6 bl[6] br[6] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_7 bl[7] br[7] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_8 bl[8] br[8] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_9 bl[9] br[9] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_10 bl[10] br[10] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_11 bl[11] br[11] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_12 bl[12] br[12] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_13 bl[13] br[13] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_14 bl[14] br[14] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_15 bl[15] br[15] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_16 bl[16] br[16] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_17 bl[17] br[17] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_18 bl[18] br[18] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_19 bl[19] br[19] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_20 bl[20] br[20] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_21 bl[21] br[21] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_22 bl[22] br[22] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_23 bl[23] br[23] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_24 bl[24] br[24] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_25 bl[25] br[25] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_26 bl[26] br[26] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_27 bl[27] br[27] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_28 bl[28] br[28] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_29 bl[29] br[29] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_30 bl[30] br[30] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_31 bl[31] br[31] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_32 bl[32] br[32] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_33 bl[33] br[33] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_34 bl[34] br[34] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_35 bl[35] br[35] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_36 bl[36] br[36] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_37 bl[37] br[37] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_38 bl[38] br[38] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_39 bl[39] br[39] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_40 bl[40] br[40] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_41 bl[41] br[41] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_42 bl[42] br[42] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_43 bl[43] br[43] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_44 bl[44] br[44] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_45 bl[45] br[45] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_46 bl[46] br[46] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_47 bl[47] br[47] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_48 bl[48] br[48] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_49 bl[49] br[49] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_50 bl[50] br[50] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_51 bl[51] br[51] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_52 bl[52] br[52] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_53 bl[53] br[53] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_54 bl[54] br[54] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_55 bl[55] br[55] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_56 bl[56] br[56] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_57 bl[57] br[57] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_58 bl[58] br[58] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_59 bl[59] br[59] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_60 bl[60] br[60] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_61 bl[61] br[61] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_62 bl[62] br[62] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_63 bl[63] br[63] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_58_0 bl[0] br[0] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_1 bl[1] br[1] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_2 bl[2] br[2] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_3 bl[3] br[3] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_4 bl[4] br[4] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_5 bl[5] br[5] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_6 bl[6] br[6] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_7 bl[7] br[7] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_8 bl[8] br[8] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_9 bl[9] br[9] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_10 bl[10] br[10] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_11 bl[11] br[11] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_12 bl[12] br[12] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_13 bl[13] br[13] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_14 bl[14] br[14] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_15 bl[15] br[15] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_16 bl[16] br[16] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_17 bl[17] br[17] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_18 bl[18] br[18] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_19 bl[19] br[19] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_20 bl[20] br[20] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_21 bl[21] br[21] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_22 bl[22] br[22] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_23 bl[23] br[23] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_24 bl[24] br[24] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_25 bl[25] br[25] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_26 bl[26] br[26] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_27 bl[27] br[27] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_28 bl[28] br[28] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_29 bl[29] br[29] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_30 bl[30] br[30] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_31 bl[31] br[31] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_32 bl[32] br[32] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_33 bl[33] br[33] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_34 bl[34] br[34] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_35 bl[35] br[35] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_36 bl[36] br[36] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_37 bl[37] br[37] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_38 bl[38] br[38] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_39 bl[39] br[39] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_40 bl[40] br[40] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_41 bl[41] br[41] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_42 bl[42] br[42] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_43 bl[43] br[43] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_44 bl[44] br[44] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_45 bl[45] br[45] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_46 bl[46] br[46] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_47 bl[47] br[47] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_48 bl[48] br[48] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_49 bl[49] br[49] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_50 bl[50] br[50] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_51 bl[51] br[51] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_52 bl[52] br[52] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_53 bl[53] br[53] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_54 bl[54] br[54] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_55 bl[55] br[55] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_56 bl[56] br[56] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_57 bl[57] br[57] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_58 bl[58] br[58] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_59 bl[59] br[59] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_60 bl[60] br[60] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_61 bl[61] br[61] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_62 bl[62] br[62] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_63 bl[63] br[63] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_59_0 bl[0] br[0] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_1 bl[1] br[1] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_2 bl[2] br[2] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_3 bl[3] br[3] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_4 bl[4] br[4] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_5 bl[5] br[5] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_6 bl[6] br[6] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_7 bl[7] br[7] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_8 bl[8] br[8] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_9 bl[9] br[9] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_10 bl[10] br[10] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_11 bl[11] br[11] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_12 bl[12] br[12] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_13 bl[13] br[13] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_14 bl[14] br[14] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_15 bl[15] br[15] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_16 bl[16] br[16] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_17 bl[17] br[17] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_18 bl[18] br[18] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_19 bl[19] br[19] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_20 bl[20] br[20] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_21 bl[21] br[21] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_22 bl[22] br[22] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_23 bl[23] br[23] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_24 bl[24] br[24] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_25 bl[25] br[25] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_26 bl[26] br[26] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_27 bl[27] br[27] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_28 bl[28] br[28] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_29 bl[29] br[29] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_30 bl[30] br[30] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_31 bl[31] br[31] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_32 bl[32] br[32] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_33 bl[33] br[33] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_34 bl[34] br[34] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_35 bl[35] br[35] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_36 bl[36] br[36] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_37 bl[37] br[37] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_38 bl[38] br[38] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_39 bl[39] br[39] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_40 bl[40] br[40] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_41 bl[41] br[41] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_42 bl[42] br[42] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_43 bl[43] br[43] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_44 bl[44] br[44] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_45 bl[45] br[45] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_46 bl[46] br[46] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_47 bl[47] br[47] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_48 bl[48] br[48] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_49 bl[49] br[49] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_50 bl[50] br[50] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_51 bl[51] br[51] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_52 bl[52] br[52] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_53 bl[53] br[53] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_54 bl[54] br[54] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_55 bl[55] br[55] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_56 bl[56] br[56] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_57 bl[57] br[57] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_58 bl[58] br[58] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_59 bl[59] br[59] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_60 bl[60] br[60] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_61 bl[61] br[61] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_62 bl[62] br[62] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_63 bl[63] br[63] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_60_0 bl[0] br[0] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_1 bl[1] br[1] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_2 bl[2] br[2] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_3 bl[3] br[3] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_4 bl[4] br[4] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_5 bl[5] br[5] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_6 bl[6] br[6] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_7 bl[7] br[7] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_8 bl[8] br[8] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_9 bl[9] br[9] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_10 bl[10] br[10] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_11 bl[11] br[11] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_12 bl[12] br[12] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_13 bl[13] br[13] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_14 bl[14] br[14] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_15 bl[15] br[15] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_16 bl[16] br[16] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_17 bl[17] br[17] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_18 bl[18] br[18] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_19 bl[19] br[19] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_20 bl[20] br[20] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_21 bl[21] br[21] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_22 bl[22] br[22] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_23 bl[23] br[23] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_24 bl[24] br[24] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_25 bl[25] br[25] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_26 bl[26] br[26] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_27 bl[27] br[27] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_28 bl[28] br[28] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_29 bl[29] br[29] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_30 bl[30] br[30] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_31 bl[31] br[31] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_32 bl[32] br[32] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_33 bl[33] br[33] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_34 bl[34] br[34] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_35 bl[35] br[35] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_36 bl[36] br[36] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_37 bl[37] br[37] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_38 bl[38] br[38] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_39 bl[39] br[39] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_40 bl[40] br[40] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_41 bl[41] br[41] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_42 bl[42] br[42] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_43 bl[43] br[43] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_44 bl[44] br[44] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_45 bl[45] br[45] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_46 bl[46] br[46] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_47 bl[47] br[47] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_48 bl[48] br[48] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_49 bl[49] br[49] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_50 bl[50] br[50] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_51 bl[51] br[51] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_52 bl[52] br[52] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_53 bl[53] br[53] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_54 bl[54] br[54] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_55 bl[55] br[55] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_56 bl[56] br[56] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_57 bl[57] br[57] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_58 bl[58] br[58] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_59 bl[59] br[59] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_60 bl[60] br[60] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_61 bl[61] br[61] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_62 bl[62] br[62] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_63 bl[63] br[63] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_61_0 bl[0] br[0] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_1 bl[1] br[1] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_2 bl[2] br[2] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_3 bl[3] br[3] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_4 bl[4] br[4] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_5 bl[5] br[5] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_6 bl[6] br[6] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_7 bl[7] br[7] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_8 bl[8] br[8] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_9 bl[9] br[9] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_10 bl[10] br[10] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_11 bl[11] br[11] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_12 bl[12] br[12] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_13 bl[13] br[13] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_14 bl[14] br[14] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_15 bl[15] br[15] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_16 bl[16] br[16] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_17 bl[17] br[17] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_18 bl[18] br[18] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_19 bl[19] br[19] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_20 bl[20] br[20] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_21 bl[21] br[21] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_22 bl[22] br[22] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_23 bl[23] br[23] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_24 bl[24] br[24] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_25 bl[25] br[25] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_26 bl[26] br[26] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_27 bl[27] br[27] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_28 bl[28] br[28] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_29 bl[29] br[29] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_30 bl[30] br[30] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_31 bl[31] br[31] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_32 bl[32] br[32] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_33 bl[33] br[33] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_34 bl[34] br[34] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_35 bl[35] br[35] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_36 bl[36] br[36] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_37 bl[37] br[37] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_38 bl[38] br[38] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_39 bl[39] br[39] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_40 bl[40] br[40] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_41 bl[41] br[41] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_42 bl[42] br[42] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_43 bl[43] br[43] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_44 bl[44] br[44] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_45 bl[45] br[45] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_46 bl[46] br[46] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_47 bl[47] br[47] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_48 bl[48] br[48] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_49 bl[49] br[49] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_50 bl[50] br[50] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_51 bl[51] br[51] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_52 bl[52] br[52] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_53 bl[53] br[53] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_54 bl[54] br[54] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_55 bl[55] br[55] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_56 bl[56] br[56] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_57 bl[57] br[57] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_58 bl[58] br[58] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_59 bl[59] br[59] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_60 bl[60] br[60] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_61 bl[61] br[61] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_62 bl[62] br[62] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_63 bl[63] br[63] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_62_0 bl[0] br[0] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_1 bl[1] br[1] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_2 bl[2] br[2] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_3 bl[3] br[3] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_4 bl[4] br[4] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_5 bl[5] br[5] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_6 bl[6] br[6] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_7 bl[7] br[7] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_8 bl[8] br[8] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_9 bl[9] br[9] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_10 bl[10] br[10] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_11 bl[11] br[11] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_12 bl[12] br[12] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_13 bl[13] br[13] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_14 bl[14] br[14] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_15 bl[15] br[15] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_16 bl[16] br[16] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_17 bl[17] br[17] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_18 bl[18] br[18] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_19 bl[19] br[19] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_20 bl[20] br[20] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_21 bl[21] br[21] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_22 bl[22] br[22] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_23 bl[23] br[23] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_24 bl[24] br[24] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_25 bl[25] br[25] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_26 bl[26] br[26] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_27 bl[27] br[27] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_28 bl[28] br[28] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_29 bl[29] br[29] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_30 bl[30] br[30] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_31 bl[31] br[31] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_32 bl[32] br[32] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_33 bl[33] br[33] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_34 bl[34] br[34] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_35 bl[35] br[35] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_36 bl[36] br[36] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_37 bl[37] br[37] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_38 bl[38] br[38] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_39 bl[39] br[39] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_40 bl[40] br[40] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_41 bl[41] br[41] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_42 bl[42] br[42] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_43 bl[43] br[43] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_44 bl[44] br[44] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_45 bl[45] br[45] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_46 bl[46] br[46] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_47 bl[47] br[47] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_48 bl[48] br[48] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_49 bl[49] br[49] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_50 bl[50] br[50] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_51 bl[51] br[51] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_52 bl[52] br[52] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_53 bl[53] br[53] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_54 bl[54] br[54] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_55 bl[55] br[55] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_56 bl[56] br[56] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_57 bl[57] br[57] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_58 bl[58] br[58] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_59 bl[59] br[59] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_60 bl[60] br[60] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_61 bl[61] br[61] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_62 bl[62] br[62] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_63 bl[63] br[63] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_63_0 bl[0] br[0] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_1 bl[1] br[1] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_2 bl[2] br[2] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_3 bl[3] br[3] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_4 bl[4] br[4] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_5 bl[5] br[5] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_6 bl[6] br[6] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_7 bl[7] br[7] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_8 bl[8] br[8] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_9 bl[9] br[9] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_10 bl[10] br[10] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_11 bl[11] br[11] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_12 bl[12] br[12] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_13 bl[13] br[13] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_14 bl[14] br[14] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_15 bl[15] br[15] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_16 bl[16] br[16] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_17 bl[17] br[17] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_18 bl[18] br[18] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_19 bl[19] br[19] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_20 bl[20] br[20] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_21 bl[21] br[21] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_22 bl[22] br[22] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_23 bl[23] br[23] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_24 bl[24] br[24] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_25 bl[25] br[25] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_26 bl[26] br[26] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_27 bl[27] br[27] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_28 bl[28] br[28] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_29 bl[29] br[29] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_30 bl[30] br[30] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_31 bl[31] br[31] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_32 bl[32] br[32] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_33 bl[33] br[33] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_34 bl[34] br[34] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_35 bl[35] br[35] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_36 bl[36] br[36] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_37 bl[37] br[37] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_38 bl[38] br[38] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_39 bl[39] br[39] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_40 bl[40] br[40] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_41 bl[41] br[41] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_42 bl[42] br[42] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_43 bl[43] br[43] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_44 bl[44] br[44] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_45 bl[45] br[45] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_46 bl[46] br[46] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_47 bl[47] br[47] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_48 bl[48] br[48] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_49 bl[49] br[49] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_50 bl[50] br[50] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_51 bl[51] br[51] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_52 bl[52] br[52] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_53 bl[53] br[53] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_54 bl[54] br[54] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_55 bl[55] br[55] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_56 bl[56] br[56] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_57 bl[57] br[57] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_58 bl[58] br[58] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_59 bl[59] br[59] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_60 bl[60] br[60] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_61 bl[61] br[61] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_62 bl[62] br[62] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_63 bl[63] br[63] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_64_0 bl[0] br[0] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_1 bl[1] br[1] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_2 bl[2] br[2] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_3 bl[3] br[3] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_4 bl[4] br[4] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_5 bl[5] br[5] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_6 bl[6] br[6] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_7 bl[7] br[7] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_8 bl[8] br[8] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_9 bl[9] br[9] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_10 bl[10] br[10] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_11 bl[11] br[11] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_12 bl[12] br[12] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_13 bl[13] br[13] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_14 bl[14] br[14] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_15 bl[15] br[15] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_16 bl[16] br[16] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_17 bl[17] br[17] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_18 bl[18] br[18] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_19 bl[19] br[19] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_20 bl[20] br[20] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_21 bl[21] br[21] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_22 bl[22] br[22] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_23 bl[23] br[23] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_24 bl[24] br[24] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_25 bl[25] br[25] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_26 bl[26] br[26] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_27 bl[27] br[27] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_28 bl[28] br[28] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_29 bl[29] br[29] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_30 bl[30] br[30] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_31 bl[31] br[31] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_32 bl[32] br[32] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_33 bl[33] br[33] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_34 bl[34] br[34] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_35 bl[35] br[35] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_36 bl[36] br[36] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_37 bl[37] br[37] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_38 bl[38] br[38] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_39 bl[39] br[39] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_40 bl[40] br[40] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_41 bl[41] br[41] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_42 bl[42] br[42] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_43 bl[43] br[43] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_44 bl[44] br[44] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_45 bl[45] br[45] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_46 bl[46] br[46] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_47 bl[47] br[47] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_48 bl[48] br[48] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_49 bl[49] br[49] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_50 bl[50] br[50] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_51 bl[51] br[51] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_52 bl[52] br[52] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_53 bl[53] br[53] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_54 bl[54] br[54] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_55 bl[55] br[55] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_56 bl[56] br[56] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_57 bl[57] br[57] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_58 bl[58] br[58] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_59 bl[59] br[59] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_60 bl[60] br[60] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_61 bl[61] br[61] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_62 bl[62] br[62] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_64_63 bl[63] br[63] vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xcell_65_0 bl[0] br[0] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_1 bl[1] br[1] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_2 bl[2] br[2] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_3 bl[3] br[3] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_4 bl[4] br[4] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_5 bl[5] br[5] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_6 bl[6] br[6] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_7 bl[7] br[7] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_8 bl[8] br[8] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_9 bl[9] br[9] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_10 bl[10] br[10] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_11 bl[11] br[11] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_12 bl[12] br[12] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_13 bl[13] br[13] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_14 bl[14] br[14] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_15 bl[15] br[15] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_16 bl[16] br[16] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_17 bl[17] br[17] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_18 bl[18] br[18] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_19 bl[19] br[19] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_20 bl[20] br[20] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_21 bl[21] br[21] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_22 bl[22] br[22] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_23 bl[23] br[23] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_24 bl[24] br[24] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_25 bl[25] br[25] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_26 bl[26] br[26] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_27 bl[27] br[27] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_28 bl[28] br[28] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_29 bl[29] br[29] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_30 bl[30] br[30] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_31 bl[31] br[31] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_32 bl[32] br[32] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_33 bl[33] br[33] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_34 bl[34] br[34] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_35 bl[35] br[35] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_36 bl[36] br[36] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_37 bl[37] br[37] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_38 bl[38] br[38] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_39 bl[39] br[39] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_40 bl[40] br[40] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_41 bl[41] br[41] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_42 bl[42] br[42] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_43 bl[43] br[43] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_44 bl[44] br[44] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_45 bl[45] br[45] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_46 bl[46] br[46] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_47 bl[47] br[47] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_48 bl[48] br[48] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_49 bl[49] br[49] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_50 bl[50] br[50] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_51 bl[51] br[51] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_52 bl[52] br[52] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_53 bl[53] br[53] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_54 bl[54] br[54] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_55 bl[55] br[55] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_56 bl[56] br[56] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_57 bl[57] br[57] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_58 bl[58] br[58] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_59 bl[59] br[59] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_60 bl[60] br[60] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_61 bl[61] br[61] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_62 bl[62] br[62] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_65_63 bl[63] br[63] vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xcell_66_0 bl[0] br[0] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_1 bl[1] br[1] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_2 bl[2] br[2] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_3 bl[3] br[3] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_4 bl[4] br[4] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_5 bl[5] br[5] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_6 bl[6] br[6] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_7 bl[7] br[7] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_8 bl[8] br[8] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_9 bl[9] br[9] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_10 bl[10] br[10] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_11 bl[11] br[11] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_12 bl[12] br[12] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_13 bl[13] br[13] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_14 bl[14] br[14] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_15 bl[15] br[15] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_16 bl[16] br[16] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_17 bl[17] br[17] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_18 bl[18] br[18] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_19 bl[19] br[19] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_20 bl[20] br[20] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_21 bl[21] br[21] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_22 bl[22] br[22] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_23 bl[23] br[23] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_24 bl[24] br[24] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_25 bl[25] br[25] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_26 bl[26] br[26] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_27 bl[27] br[27] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_28 bl[28] br[28] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_29 bl[29] br[29] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_30 bl[30] br[30] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_31 bl[31] br[31] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_32 bl[32] br[32] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_33 bl[33] br[33] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_34 bl[34] br[34] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_35 bl[35] br[35] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_36 bl[36] br[36] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_37 bl[37] br[37] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_38 bl[38] br[38] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_39 bl[39] br[39] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_40 bl[40] br[40] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_41 bl[41] br[41] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_42 bl[42] br[42] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_43 bl[43] br[43] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_44 bl[44] br[44] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_45 bl[45] br[45] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_46 bl[46] br[46] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_47 bl[47] br[47] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_48 bl[48] br[48] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_49 bl[49] br[49] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_50 bl[50] br[50] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_51 bl[51] br[51] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_52 bl[52] br[52] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_53 bl[53] br[53] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_54 bl[54] br[54] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_55 bl[55] br[55] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_56 bl[56] br[56] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_57 bl[57] br[57] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_58 bl[58] br[58] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_59 bl[59] br[59] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_60 bl[60] br[60] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_61 bl[61] br[61] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_62 bl[62] br[62] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_66_63 bl[63] br[63] vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xcell_67_0 bl[0] br[0] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_1 bl[1] br[1] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_2 bl[2] br[2] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_3 bl[3] br[3] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_4 bl[4] br[4] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_5 bl[5] br[5] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_6 bl[6] br[6] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_7 bl[7] br[7] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_8 bl[8] br[8] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_9 bl[9] br[9] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_10 bl[10] br[10] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_11 bl[11] br[11] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_12 bl[12] br[12] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_13 bl[13] br[13] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_14 bl[14] br[14] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_15 bl[15] br[15] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_16 bl[16] br[16] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_17 bl[17] br[17] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_18 bl[18] br[18] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_19 bl[19] br[19] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_20 bl[20] br[20] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_21 bl[21] br[21] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_22 bl[22] br[22] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_23 bl[23] br[23] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_24 bl[24] br[24] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_25 bl[25] br[25] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_26 bl[26] br[26] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_27 bl[27] br[27] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_28 bl[28] br[28] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_29 bl[29] br[29] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_30 bl[30] br[30] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_31 bl[31] br[31] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_32 bl[32] br[32] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_33 bl[33] br[33] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_34 bl[34] br[34] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_35 bl[35] br[35] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_36 bl[36] br[36] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_37 bl[37] br[37] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_38 bl[38] br[38] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_39 bl[39] br[39] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_40 bl[40] br[40] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_41 bl[41] br[41] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_42 bl[42] br[42] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_43 bl[43] br[43] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_44 bl[44] br[44] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_45 bl[45] br[45] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_46 bl[46] br[46] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_47 bl[47] br[47] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_48 bl[48] br[48] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_49 bl[49] br[49] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_50 bl[50] br[50] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_51 bl[51] br[51] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_52 bl[52] br[52] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_53 bl[53] br[53] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_54 bl[54] br[54] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_55 bl[55] br[55] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_56 bl[56] br[56] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_57 bl[57] br[57] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_58 bl[58] br[58] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_59 bl[59] br[59] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_60 bl[60] br[60] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_61 bl[61] br[61] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_62 bl[62] br[62] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_67_63 bl[63] br[63] vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xcell_68_0 bl[0] br[0] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_1 bl[1] br[1] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_2 bl[2] br[2] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_3 bl[3] br[3] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_4 bl[4] br[4] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_5 bl[5] br[5] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_6 bl[6] br[6] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_7 bl[7] br[7] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_8 bl[8] br[8] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_9 bl[9] br[9] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_10 bl[10] br[10] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_11 bl[11] br[11] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_12 bl[12] br[12] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_13 bl[13] br[13] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_14 bl[14] br[14] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_15 bl[15] br[15] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_16 bl[16] br[16] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_17 bl[17] br[17] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_18 bl[18] br[18] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_19 bl[19] br[19] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_20 bl[20] br[20] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_21 bl[21] br[21] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_22 bl[22] br[22] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_23 bl[23] br[23] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_24 bl[24] br[24] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_25 bl[25] br[25] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_26 bl[26] br[26] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_27 bl[27] br[27] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_28 bl[28] br[28] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_29 bl[29] br[29] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_30 bl[30] br[30] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_31 bl[31] br[31] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_32 bl[32] br[32] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_33 bl[33] br[33] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_34 bl[34] br[34] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_35 bl[35] br[35] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_36 bl[36] br[36] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_37 bl[37] br[37] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_38 bl[38] br[38] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_39 bl[39] br[39] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_40 bl[40] br[40] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_41 bl[41] br[41] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_42 bl[42] br[42] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_43 bl[43] br[43] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_44 bl[44] br[44] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_45 bl[45] br[45] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_46 bl[46] br[46] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_47 bl[47] br[47] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_48 bl[48] br[48] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_49 bl[49] br[49] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_50 bl[50] br[50] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_51 bl[51] br[51] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_52 bl[52] br[52] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_53 bl[53] br[53] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_54 bl[54] br[54] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_55 bl[55] br[55] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_56 bl[56] br[56] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_57 bl[57] br[57] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_58 bl[58] br[58] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_59 bl[59] br[59] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_60 bl[60] br[60] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_61 bl[61] br[61] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_62 bl[62] br[62] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_68_63 bl[63] br[63] vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xcell_69_0 bl[0] br[0] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_1 bl[1] br[1] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_2 bl[2] br[2] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_3 bl[3] br[3] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_4 bl[4] br[4] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_5 bl[5] br[5] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_6 bl[6] br[6] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_7 bl[7] br[7] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_8 bl[8] br[8] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_9 bl[9] br[9] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_10 bl[10] br[10] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_11 bl[11] br[11] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_12 bl[12] br[12] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_13 bl[13] br[13] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_14 bl[14] br[14] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_15 bl[15] br[15] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_16 bl[16] br[16] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_17 bl[17] br[17] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_18 bl[18] br[18] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_19 bl[19] br[19] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_20 bl[20] br[20] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_21 bl[21] br[21] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_22 bl[22] br[22] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_23 bl[23] br[23] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_24 bl[24] br[24] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_25 bl[25] br[25] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_26 bl[26] br[26] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_27 bl[27] br[27] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_28 bl[28] br[28] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_29 bl[29] br[29] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_30 bl[30] br[30] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_31 bl[31] br[31] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_32 bl[32] br[32] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_33 bl[33] br[33] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_34 bl[34] br[34] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_35 bl[35] br[35] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_36 bl[36] br[36] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_37 bl[37] br[37] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_38 bl[38] br[38] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_39 bl[39] br[39] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_40 bl[40] br[40] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_41 bl[41] br[41] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_42 bl[42] br[42] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_43 bl[43] br[43] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_44 bl[44] br[44] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_45 bl[45] br[45] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_46 bl[46] br[46] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_47 bl[47] br[47] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_48 bl[48] br[48] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_49 bl[49] br[49] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_50 bl[50] br[50] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_51 bl[51] br[51] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_52 bl[52] br[52] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_53 bl[53] br[53] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_54 bl[54] br[54] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_55 bl[55] br[55] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_56 bl[56] br[56] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_57 bl[57] br[57] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_58 bl[58] br[58] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_59 bl[59] br[59] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_60 bl[60] br[60] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_61 bl[61] br[61] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_62 bl[62] br[62] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_69_63 bl[63] br[63] vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xcell_70_0 bl[0] br[0] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_1 bl[1] br[1] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_2 bl[2] br[2] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_3 bl[3] br[3] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_4 bl[4] br[4] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_5 bl[5] br[5] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_6 bl[6] br[6] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_7 bl[7] br[7] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_8 bl[8] br[8] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_9 bl[9] br[9] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_10 bl[10] br[10] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_11 bl[11] br[11] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_12 bl[12] br[12] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_13 bl[13] br[13] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_14 bl[14] br[14] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_15 bl[15] br[15] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_16 bl[16] br[16] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_17 bl[17] br[17] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_18 bl[18] br[18] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_19 bl[19] br[19] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_20 bl[20] br[20] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_21 bl[21] br[21] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_22 bl[22] br[22] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_23 bl[23] br[23] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_24 bl[24] br[24] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_25 bl[25] br[25] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_26 bl[26] br[26] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_27 bl[27] br[27] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_28 bl[28] br[28] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_29 bl[29] br[29] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_30 bl[30] br[30] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_31 bl[31] br[31] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_32 bl[32] br[32] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_33 bl[33] br[33] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_34 bl[34] br[34] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_35 bl[35] br[35] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_36 bl[36] br[36] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_37 bl[37] br[37] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_38 bl[38] br[38] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_39 bl[39] br[39] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_40 bl[40] br[40] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_41 bl[41] br[41] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_42 bl[42] br[42] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_43 bl[43] br[43] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_44 bl[44] br[44] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_45 bl[45] br[45] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_46 bl[46] br[46] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_47 bl[47] br[47] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_48 bl[48] br[48] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_49 bl[49] br[49] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_50 bl[50] br[50] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_51 bl[51] br[51] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_52 bl[52] br[52] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_53 bl[53] br[53] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_54 bl[54] br[54] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_55 bl[55] br[55] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_56 bl[56] br[56] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_57 bl[57] br[57] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_58 bl[58] br[58] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_59 bl[59] br[59] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_60 bl[60] br[60] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_61 bl[61] br[61] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_62 bl[62] br[62] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_70_63 bl[63] br[63] vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xcell_71_0 bl[0] br[0] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_1 bl[1] br[1] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_2 bl[2] br[2] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_3 bl[3] br[3] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_4 bl[4] br[4] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_5 bl[5] br[5] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_6 bl[6] br[6] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_7 bl[7] br[7] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_8 bl[8] br[8] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_9 bl[9] br[9] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_10 bl[10] br[10] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_11 bl[11] br[11] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_12 bl[12] br[12] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_13 bl[13] br[13] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_14 bl[14] br[14] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_15 bl[15] br[15] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_16 bl[16] br[16] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_17 bl[17] br[17] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_18 bl[18] br[18] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_19 bl[19] br[19] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_20 bl[20] br[20] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_21 bl[21] br[21] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_22 bl[22] br[22] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_23 bl[23] br[23] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_24 bl[24] br[24] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_25 bl[25] br[25] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_26 bl[26] br[26] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_27 bl[27] br[27] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_28 bl[28] br[28] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_29 bl[29] br[29] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_30 bl[30] br[30] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_31 bl[31] br[31] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_32 bl[32] br[32] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_33 bl[33] br[33] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_34 bl[34] br[34] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_35 bl[35] br[35] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_36 bl[36] br[36] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_37 bl[37] br[37] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_38 bl[38] br[38] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_39 bl[39] br[39] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_40 bl[40] br[40] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_41 bl[41] br[41] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_42 bl[42] br[42] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_43 bl[43] br[43] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_44 bl[44] br[44] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_45 bl[45] br[45] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_46 bl[46] br[46] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_47 bl[47] br[47] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_48 bl[48] br[48] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_49 bl[49] br[49] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_50 bl[50] br[50] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_51 bl[51] br[51] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_52 bl[52] br[52] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_53 bl[53] br[53] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_54 bl[54] br[54] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_55 bl[55] br[55] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_56 bl[56] br[56] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_57 bl[57] br[57] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_58 bl[58] br[58] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_59 bl[59] br[59] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_60 bl[60] br[60] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_61 bl[61] br[61] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_62 bl[62] br[62] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_71_63 bl[63] br[63] vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xcell_72_0 bl[0] br[0] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_1 bl[1] br[1] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_2 bl[2] br[2] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_3 bl[3] br[3] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_4 bl[4] br[4] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_5 bl[5] br[5] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_6 bl[6] br[6] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_7 bl[7] br[7] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_8 bl[8] br[8] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_9 bl[9] br[9] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_10 bl[10] br[10] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_11 bl[11] br[11] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_12 bl[12] br[12] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_13 bl[13] br[13] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_14 bl[14] br[14] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_15 bl[15] br[15] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_16 bl[16] br[16] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_17 bl[17] br[17] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_18 bl[18] br[18] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_19 bl[19] br[19] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_20 bl[20] br[20] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_21 bl[21] br[21] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_22 bl[22] br[22] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_23 bl[23] br[23] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_24 bl[24] br[24] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_25 bl[25] br[25] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_26 bl[26] br[26] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_27 bl[27] br[27] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_28 bl[28] br[28] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_29 bl[29] br[29] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_30 bl[30] br[30] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_31 bl[31] br[31] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_32 bl[32] br[32] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_33 bl[33] br[33] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_34 bl[34] br[34] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_35 bl[35] br[35] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_36 bl[36] br[36] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_37 bl[37] br[37] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_38 bl[38] br[38] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_39 bl[39] br[39] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_40 bl[40] br[40] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_41 bl[41] br[41] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_42 bl[42] br[42] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_43 bl[43] br[43] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_44 bl[44] br[44] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_45 bl[45] br[45] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_46 bl[46] br[46] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_47 bl[47] br[47] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_48 bl[48] br[48] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_49 bl[49] br[49] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_50 bl[50] br[50] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_51 bl[51] br[51] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_52 bl[52] br[52] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_53 bl[53] br[53] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_54 bl[54] br[54] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_55 bl[55] br[55] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_56 bl[56] br[56] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_57 bl[57] br[57] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_58 bl[58] br[58] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_59 bl[59] br[59] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_60 bl[60] br[60] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_61 bl[61] br[61] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_62 bl[62] br[62] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_72_63 bl[63] br[63] vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xcell_73_0 bl[0] br[0] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_1 bl[1] br[1] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_2 bl[2] br[2] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_3 bl[3] br[3] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_4 bl[4] br[4] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_5 bl[5] br[5] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_6 bl[6] br[6] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_7 bl[7] br[7] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_8 bl[8] br[8] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_9 bl[9] br[9] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_10 bl[10] br[10] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_11 bl[11] br[11] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_12 bl[12] br[12] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_13 bl[13] br[13] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_14 bl[14] br[14] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_15 bl[15] br[15] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_16 bl[16] br[16] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_17 bl[17] br[17] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_18 bl[18] br[18] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_19 bl[19] br[19] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_20 bl[20] br[20] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_21 bl[21] br[21] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_22 bl[22] br[22] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_23 bl[23] br[23] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_24 bl[24] br[24] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_25 bl[25] br[25] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_26 bl[26] br[26] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_27 bl[27] br[27] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_28 bl[28] br[28] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_29 bl[29] br[29] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_30 bl[30] br[30] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_31 bl[31] br[31] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_32 bl[32] br[32] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_33 bl[33] br[33] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_34 bl[34] br[34] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_35 bl[35] br[35] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_36 bl[36] br[36] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_37 bl[37] br[37] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_38 bl[38] br[38] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_39 bl[39] br[39] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_40 bl[40] br[40] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_41 bl[41] br[41] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_42 bl[42] br[42] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_43 bl[43] br[43] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_44 bl[44] br[44] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_45 bl[45] br[45] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_46 bl[46] br[46] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_47 bl[47] br[47] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_48 bl[48] br[48] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_49 bl[49] br[49] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_50 bl[50] br[50] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_51 bl[51] br[51] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_52 bl[52] br[52] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_53 bl[53] br[53] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_54 bl[54] br[54] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_55 bl[55] br[55] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_56 bl[56] br[56] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_57 bl[57] br[57] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_58 bl[58] br[58] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_59 bl[59] br[59] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_60 bl[60] br[60] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_61 bl[61] br[61] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_62 bl[62] br[62] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_73_63 bl[63] br[63] vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xcell_74_0 bl[0] br[0] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_1 bl[1] br[1] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_2 bl[2] br[2] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_3 bl[3] br[3] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_4 bl[4] br[4] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_5 bl[5] br[5] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_6 bl[6] br[6] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_7 bl[7] br[7] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_8 bl[8] br[8] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_9 bl[9] br[9] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_10 bl[10] br[10] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_11 bl[11] br[11] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_12 bl[12] br[12] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_13 bl[13] br[13] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_14 bl[14] br[14] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_15 bl[15] br[15] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_16 bl[16] br[16] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_17 bl[17] br[17] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_18 bl[18] br[18] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_19 bl[19] br[19] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_20 bl[20] br[20] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_21 bl[21] br[21] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_22 bl[22] br[22] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_23 bl[23] br[23] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_24 bl[24] br[24] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_25 bl[25] br[25] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_26 bl[26] br[26] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_27 bl[27] br[27] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_28 bl[28] br[28] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_29 bl[29] br[29] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_30 bl[30] br[30] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_31 bl[31] br[31] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_32 bl[32] br[32] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_33 bl[33] br[33] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_34 bl[34] br[34] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_35 bl[35] br[35] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_36 bl[36] br[36] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_37 bl[37] br[37] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_38 bl[38] br[38] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_39 bl[39] br[39] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_40 bl[40] br[40] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_41 bl[41] br[41] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_42 bl[42] br[42] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_43 bl[43] br[43] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_44 bl[44] br[44] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_45 bl[45] br[45] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_46 bl[46] br[46] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_47 bl[47] br[47] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_48 bl[48] br[48] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_49 bl[49] br[49] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_50 bl[50] br[50] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_51 bl[51] br[51] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_52 bl[52] br[52] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_53 bl[53] br[53] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_54 bl[54] br[54] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_55 bl[55] br[55] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_56 bl[56] br[56] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_57 bl[57] br[57] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_58 bl[58] br[58] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_59 bl[59] br[59] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_60 bl[60] br[60] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_61 bl[61] br[61] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_62 bl[62] br[62] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_74_63 bl[63] br[63] vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xcell_75_0 bl[0] br[0] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_1 bl[1] br[1] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_2 bl[2] br[2] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_3 bl[3] br[3] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_4 bl[4] br[4] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_5 bl[5] br[5] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_6 bl[6] br[6] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_7 bl[7] br[7] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_8 bl[8] br[8] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_9 bl[9] br[9] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_10 bl[10] br[10] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_11 bl[11] br[11] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_12 bl[12] br[12] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_13 bl[13] br[13] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_14 bl[14] br[14] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_15 bl[15] br[15] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_16 bl[16] br[16] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_17 bl[17] br[17] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_18 bl[18] br[18] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_19 bl[19] br[19] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_20 bl[20] br[20] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_21 bl[21] br[21] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_22 bl[22] br[22] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_23 bl[23] br[23] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_24 bl[24] br[24] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_25 bl[25] br[25] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_26 bl[26] br[26] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_27 bl[27] br[27] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_28 bl[28] br[28] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_29 bl[29] br[29] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_30 bl[30] br[30] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_31 bl[31] br[31] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_32 bl[32] br[32] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_33 bl[33] br[33] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_34 bl[34] br[34] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_35 bl[35] br[35] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_36 bl[36] br[36] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_37 bl[37] br[37] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_38 bl[38] br[38] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_39 bl[39] br[39] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_40 bl[40] br[40] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_41 bl[41] br[41] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_42 bl[42] br[42] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_43 bl[43] br[43] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_44 bl[44] br[44] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_45 bl[45] br[45] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_46 bl[46] br[46] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_47 bl[47] br[47] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_48 bl[48] br[48] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_49 bl[49] br[49] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_50 bl[50] br[50] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_51 bl[51] br[51] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_52 bl[52] br[52] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_53 bl[53] br[53] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_54 bl[54] br[54] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_55 bl[55] br[55] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_56 bl[56] br[56] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_57 bl[57] br[57] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_58 bl[58] br[58] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_59 bl[59] br[59] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_60 bl[60] br[60] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_61 bl[61] br[61] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_62 bl[62] br[62] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_75_63 bl[63] br[63] vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xcell_76_0 bl[0] br[0] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_1 bl[1] br[1] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_2 bl[2] br[2] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_3 bl[3] br[3] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_4 bl[4] br[4] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_5 bl[5] br[5] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_6 bl[6] br[6] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_7 bl[7] br[7] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_8 bl[8] br[8] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_9 bl[9] br[9] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_10 bl[10] br[10] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_11 bl[11] br[11] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_12 bl[12] br[12] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_13 bl[13] br[13] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_14 bl[14] br[14] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_15 bl[15] br[15] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_16 bl[16] br[16] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_17 bl[17] br[17] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_18 bl[18] br[18] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_19 bl[19] br[19] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_20 bl[20] br[20] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_21 bl[21] br[21] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_22 bl[22] br[22] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_23 bl[23] br[23] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_24 bl[24] br[24] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_25 bl[25] br[25] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_26 bl[26] br[26] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_27 bl[27] br[27] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_28 bl[28] br[28] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_29 bl[29] br[29] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_30 bl[30] br[30] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_31 bl[31] br[31] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_32 bl[32] br[32] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_33 bl[33] br[33] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_34 bl[34] br[34] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_35 bl[35] br[35] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_36 bl[36] br[36] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_37 bl[37] br[37] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_38 bl[38] br[38] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_39 bl[39] br[39] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_40 bl[40] br[40] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_41 bl[41] br[41] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_42 bl[42] br[42] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_43 bl[43] br[43] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_44 bl[44] br[44] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_45 bl[45] br[45] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_46 bl[46] br[46] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_47 bl[47] br[47] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_48 bl[48] br[48] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_49 bl[49] br[49] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_50 bl[50] br[50] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_51 bl[51] br[51] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_52 bl[52] br[52] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_53 bl[53] br[53] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_54 bl[54] br[54] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_55 bl[55] br[55] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_56 bl[56] br[56] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_57 bl[57] br[57] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_58 bl[58] br[58] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_59 bl[59] br[59] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_60 bl[60] br[60] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_61 bl[61] br[61] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_62 bl[62] br[62] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_76_63 bl[63] br[63] vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xcell_77_0 bl[0] br[0] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_1 bl[1] br[1] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_2 bl[2] br[2] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_3 bl[3] br[3] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_4 bl[4] br[4] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_5 bl[5] br[5] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_6 bl[6] br[6] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_7 bl[7] br[7] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_8 bl[8] br[8] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_9 bl[9] br[9] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_10 bl[10] br[10] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_11 bl[11] br[11] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_12 bl[12] br[12] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_13 bl[13] br[13] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_14 bl[14] br[14] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_15 bl[15] br[15] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_16 bl[16] br[16] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_17 bl[17] br[17] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_18 bl[18] br[18] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_19 bl[19] br[19] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_20 bl[20] br[20] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_21 bl[21] br[21] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_22 bl[22] br[22] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_23 bl[23] br[23] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_24 bl[24] br[24] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_25 bl[25] br[25] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_26 bl[26] br[26] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_27 bl[27] br[27] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_28 bl[28] br[28] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_29 bl[29] br[29] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_30 bl[30] br[30] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_31 bl[31] br[31] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_32 bl[32] br[32] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_33 bl[33] br[33] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_34 bl[34] br[34] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_35 bl[35] br[35] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_36 bl[36] br[36] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_37 bl[37] br[37] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_38 bl[38] br[38] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_39 bl[39] br[39] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_40 bl[40] br[40] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_41 bl[41] br[41] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_42 bl[42] br[42] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_43 bl[43] br[43] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_44 bl[44] br[44] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_45 bl[45] br[45] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_46 bl[46] br[46] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_47 bl[47] br[47] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_48 bl[48] br[48] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_49 bl[49] br[49] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_50 bl[50] br[50] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_51 bl[51] br[51] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_52 bl[52] br[52] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_53 bl[53] br[53] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_54 bl[54] br[54] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_55 bl[55] br[55] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_56 bl[56] br[56] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_57 bl[57] br[57] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_58 bl[58] br[58] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_59 bl[59] br[59] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_60 bl[60] br[60] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_61 bl[61] br[61] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_62 bl[62] br[62] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_77_63 bl[63] br[63] vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xcell_78_0 bl[0] br[0] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_1 bl[1] br[1] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_2 bl[2] br[2] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_3 bl[3] br[3] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_4 bl[4] br[4] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_5 bl[5] br[5] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_6 bl[6] br[6] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_7 bl[7] br[7] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_8 bl[8] br[8] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_9 bl[9] br[9] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_10 bl[10] br[10] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_11 bl[11] br[11] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_12 bl[12] br[12] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_13 bl[13] br[13] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_14 bl[14] br[14] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_15 bl[15] br[15] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_16 bl[16] br[16] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_17 bl[17] br[17] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_18 bl[18] br[18] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_19 bl[19] br[19] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_20 bl[20] br[20] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_21 bl[21] br[21] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_22 bl[22] br[22] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_23 bl[23] br[23] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_24 bl[24] br[24] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_25 bl[25] br[25] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_26 bl[26] br[26] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_27 bl[27] br[27] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_28 bl[28] br[28] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_29 bl[29] br[29] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_30 bl[30] br[30] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_31 bl[31] br[31] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_32 bl[32] br[32] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_33 bl[33] br[33] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_34 bl[34] br[34] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_35 bl[35] br[35] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_36 bl[36] br[36] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_37 bl[37] br[37] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_38 bl[38] br[38] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_39 bl[39] br[39] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_40 bl[40] br[40] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_41 bl[41] br[41] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_42 bl[42] br[42] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_43 bl[43] br[43] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_44 bl[44] br[44] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_45 bl[45] br[45] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_46 bl[46] br[46] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_47 bl[47] br[47] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_48 bl[48] br[48] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_49 bl[49] br[49] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_50 bl[50] br[50] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_51 bl[51] br[51] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_52 bl[52] br[52] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_53 bl[53] br[53] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_54 bl[54] br[54] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_55 bl[55] br[55] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_56 bl[56] br[56] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_57 bl[57] br[57] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_58 bl[58] br[58] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_59 bl[59] br[59] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_60 bl[60] br[60] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_61 bl[61] br[61] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_62 bl[62] br[62] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_78_63 bl[63] br[63] vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xcell_79_0 bl[0] br[0] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_1 bl[1] br[1] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_2 bl[2] br[2] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_3 bl[3] br[3] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_4 bl[4] br[4] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_5 bl[5] br[5] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_6 bl[6] br[6] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_7 bl[7] br[7] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_8 bl[8] br[8] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_9 bl[9] br[9] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_10 bl[10] br[10] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_11 bl[11] br[11] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_12 bl[12] br[12] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_13 bl[13] br[13] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_14 bl[14] br[14] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_15 bl[15] br[15] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_16 bl[16] br[16] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_17 bl[17] br[17] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_18 bl[18] br[18] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_19 bl[19] br[19] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_20 bl[20] br[20] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_21 bl[21] br[21] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_22 bl[22] br[22] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_23 bl[23] br[23] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_24 bl[24] br[24] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_25 bl[25] br[25] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_26 bl[26] br[26] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_27 bl[27] br[27] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_28 bl[28] br[28] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_29 bl[29] br[29] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_30 bl[30] br[30] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_31 bl[31] br[31] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_32 bl[32] br[32] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_33 bl[33] br[33] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_34 bl[34] br[34] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_35 bl[35] br[35] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_36 bl[36] br[36] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_37 bl[37] br[37] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_38 bl[38] br[38] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_39 bl[39] br[39] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_40 bl[40] br[40] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_41 bl[41] br[41] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_42 bl[42] br[42] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_43 bl[43] br[43] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_44 bl[44] br[44] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_45 bl[45] br[45] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_46 bl[46] br[46] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_47 bl[47] br[47] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_48 bl[48] br[48] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_49 bl[49] br[49] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_50 bl[50] br[50] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_51 bl[51] br[51] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_52 bl[52] br[52] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_53 bl[53] br[53] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_54 bl[54] br[54] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_55 bl[55] br[55] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_56 bl[56] br[56] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_57 bl[57] br[57] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_58 bl[58] br[58] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_59 bl[59] br[59] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_60 bl[60] br[60] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_61 bl[61] br[61] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_62 bl[62] br[62] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_79_63 bl[63] br[63] vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xcell_80_0 bl[0] br[0] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_1 bl[1] br[1] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_2 bl[2] br[2] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_3 bl[3] br[3] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_4 bl[4] br[4] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_5 bl[5] br[5] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_6 bl[6] br[6] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_7 bl[7] br[7] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_8 bl[8] br[8] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_9 bl[9] br[9] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_10 bl[10] br[10] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_11 bl[11] br[11] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_12 bl[12] br[12] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_13 bl[13] br[13] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_14 bl[14] br[14] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_15 bl[15] br[15] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_16 bl[16] br[16] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_17 bl[17] br[17] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_18 bl[18] br[18] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_19 bl[19] br[19] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_20 bl[20] br[20] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_21 bl[21] br[21] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_22 bl[22] br[22] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_23 bl[23] br[23] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_24 bl[24] br[24] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_25 bl[25] br[25] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_26 bl[26] br[26] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_27 bl[27] br[27] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_28 bl[28] br[28] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_29 bl[29] br[29] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_30 bl[30] br[30] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_31 bl[31] br[31] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_32 bl[32] br[32] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_33 bl[33] br[33] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_34 bl[34] br[34] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_35 bl[35] br[35] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_36 bl[36] br[36] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_37 bl[37] br[37] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_38 bl[38] br[38] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_39 bl[39] br[39] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_40 bl[40] br[40] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_41 bl[41] br[41] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_42 bl[42] br[42] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_43 bl[43] br[43] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_44 bl[44] br[44] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_45 bl[45] br[45] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_46 bl[46] br[46] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_47 bl[47] br[47] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_48 bl[48] br[48] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_49 bl[49] br[49] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_50 bl[50] br[50] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_51 bl[51] br[51] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_52 bl[52] br[52] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_53 bl[53] br[53] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_54 bl[54] br[54] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_55 bl[55] br[55] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_56 bl[56] br[56] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_57 bl[57] br[57] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_58 bl[58] br[58] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_59 bl[59] br[59] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_60 bl[60] br[60] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_61 bl[61] br[61] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_62 bl[62] br[62] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_80_63 bl[63] br[63] vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xcell_81_0 bl[0] br[0] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_1 bl[1] br[1] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_2 bl[2] br[2] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_3 bl[3] br[3] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_4 bl[4] br[4] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_5 bl[5] br[5] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_6 bl[6] br[6] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_7 bl[7] br[7] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_8 bl[8] br[8] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_9 bl[9] br[9] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_10 bl[10] br[10] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_11 bl[11] br[11] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_12 bl[12] br[12] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_13 bl[13] br[13] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_14 bl[14] br[14] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_15 bl[15] br[15] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_16 bl[16] br[16] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_17 bl[17] br[17] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_18 bl[18] br[18] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_19 bl[19] br[19] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_20 bl[20] br[20] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_21 bl[21] br[21] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_22 bl[22] br[22] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_23 bl[23] br[23] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_24 bl[24] br[24] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_25 bl[25] br[25] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_26 bl[26] br[26] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_27 bl[27] br[27] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_28 bl[28] br[28] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_29 bl[29] br[29] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_30 bl[30] br[30] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_31 bl[31] br[31] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_32 bl[32] br[32] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_33 bl[33] br[33] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_34 bl[34] br[34] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_35 bl[35] br[35] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_36 bl[36] br[36] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_37 bl[37] br[37] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_38 bl[38] br[38] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_39 bl[39] br[39] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_40 bl[40] br[40] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_41 bl[41] br[41] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_42 bl[42] br[42] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_43 bl[43] br[43] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_44 bl[44] br[44] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_45 bl[45] br[45] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_46 bl[46] br[46] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_47 bl[47] br[47] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_48 bl[48] br[48] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_49 bl[49] br[49] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_50 bl[50] br[50] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_51 bl[51] br[51] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_52 bl[52] br[52] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_53 bl[53] br[53] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_54 bl[54] br[54] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_55 bl[55] br[55] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_56 bl[56] br[56] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_57 bl[57] br[57] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_58 bl[58] br[58] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_59 bl[59] br[59] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_60 bl[60] br[60] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_61 bl[61] br[61] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_62 bl[62] br[62] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_81_63 bl[63] br[63] vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xcell_82_0 bl[0] br[0] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_1 bl[1] br[1] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_2 bl[2] br[2] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_3 bl[3] br[3] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_4 bl[4] br[4] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_5 bl[5] br[5] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_6 bl[6] br[6] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_7 bl[7] br[7] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_8 bl[8] br[8] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_9 bl[9] br[9] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_10 bl[10] br[10] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_11 bl[11] br[11] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_12 bl[12] br[12] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_13 bl[13] br[13] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_14 bl[14] br[14] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_15 bl[15] br[15] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_16 bl[16] br[16] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_17 bl[17] br[17] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_18 bl[18] br[18] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_19 bl[19] br[19] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_20 bl[20] br[20] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_21 bl[21] br[21] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_22 bl[22] br[22] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_23 bl[23] br[23] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_24 bl[24] br[24] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_25 bl[25] br[25] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_26 bl[26] br[26] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_27 bl[27] br[27] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_28 bl[28] br[28] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_29 bl[29] br[29] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_30 bl[30] br[30] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_31 bl[31] br[31] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_32 bl[32] br[32] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_33 bl[33] br[33] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_34 bl[34] br[34] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_35 bl[35] br[35] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_36 bl[36] br[36] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_37 bl[37] br[37] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_38 bl[38] br[38] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_39 bl[39] br[39] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_40 bl[40] br[40] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_41 bl[41] br[41] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_42 bl[42] br[42] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_43 bl[43] br[43] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_44 bl[44] br[44] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_45 bl[45] br[45] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_46 bl[46] br[46] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_47 bl[47] br[47] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_48 bl[48] br[48] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_49 bl[49] br[49] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_50 bl[50] br[50] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_51 bl[51] br[51] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_52 bl[52] br[52] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_53 bl[53] br[53] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_54 bl[54] br[54] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_55 bl[55] br[55] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_56 bl[56] br[56] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_57 bl[57] br[57] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_58 bl[58] br[58] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_59 bl[59] br[59] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_60 bl[60] br[60] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_61 bl[61] br[61] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_62 bl[62] br[62] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_82_63 bl[63] br[63] vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xcell_83_0 bl[0] br[0] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_1 bl[1] br[1] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_2 bl[2] br[2] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_3 bl[3] br[3] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_4 bl[4] br[4] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_5 bl[5] br[5] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_6 bl[6] br[6] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_7 bl[7] br[7] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_8 bl[8] br[8] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_9 bl[9] br[9] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_10 bl[10] br[10] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_11 bl[11] br[11] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_12 bl[12] br[12] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_13 bl[13] br[13] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_14 bl[14] br[14] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_15 bl[15] br[15] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_16 bl[16] br[16] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_17 bl[17] br[17] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_18 bl[18] br[18] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_19 bl[19] br[19] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_20 bl[20] br[20] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_21 bl[21] br[21] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_22 bl[22] br[22] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_23 bl[23] br[23] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_24 bl[24] br[24] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_25 bl[25] br[25] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_26 bl[26] br[26] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_27 bl[27] br[27] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_28 bl[28] br[28] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_29 bl[29] br[29] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_30 bl[30] br[30] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_31 bl[31] br[31] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_32 bl[32] br[32] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_33 bl[33] br[33] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_34 bl[34] br[34] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_35 bl[35] br[35] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_36 bl[36] br[36] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_37 bl[37] br[37] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_38 bl[38] br[38] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_39 bl[39] br[39] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_40 bl[40] br[40] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_41 bl[41] br[41] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_42 bl[42] br[42] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_43 bl[43] br[43] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_44 bl[44] br[44] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_45 bl[45] br[45] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_46 bl[46] br[46] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_47 bl[47] br[47] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_48 bl[48] br[48] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_49 bl[49] br[49] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_50 bl[50] br[50] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_51 bl[51] br[51] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_52 bl[52] br[52] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_53 bl[53] br[53] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_54 bl[54] br[54] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_55 bl[55] br[55] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_56 bl[56] br[56] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_57 bl[57] br[57] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_58 bl[58] br[58] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_59 bl[59] br[59] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_60 bl[60] br[60] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_61 bl[61] br[61] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_62 bl[62] br[62] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_83_63 bl[63] br[63] vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xcell_84_0 bl[0] br[0] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_1 bl[1] br[1] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_2 bl[2] br[2] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_3 bl[3] br[3] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_4 bl[4] br[4] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_5 bl[5] br[5] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_6 bl[6] br[6] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_7 bl[7] br[7] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_8 bl[8] br[8] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_9 bl[9] br[9] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_10 bl[10] br[10] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_11 bl[11] br[11] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_12 bl[12] br[12] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_13 bl[13] br[13] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_14 bl[14] br[14] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_15 bl[15] br[15] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_16 bl[16] br[16] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_17 bl[17] br[17] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_18 bl[18] br[18] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_19 bl[19] br[19] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_20 bl[20] br[20] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_21 bl[21] br[21] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_22 bl[22] br[22] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_23 bl[23] br[23] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_24 bl[24] br[24] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_25 bl[25] br[25] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_26 bl[26] br[26] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_27 bl[27] br[27] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_28 bl[28] br[28] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_29 bl[29] br[29] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_30 bl[30] br[30] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_31 bl[31] br[31] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_32 bl[32] br[32] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_33 bl[33] br[33] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_34 bl[34] br[34] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_35 bl[35] br[35] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_36 bl[36] br[36] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_37 bl[37] br[37] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_38 bl[38] br[38] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_39 bl[39] br[39] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_40 bl[40] br[40] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_41 bl[41] br[41] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_42 bl[42] br[42] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_43 bl[43] br[43] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_44 bl[44] br[44] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_45 bl[45] br[45] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_46 bl[46] br[46] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_47 bl[47] br[47] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_48 bl[48] br[48] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_49 bl[49] br[49] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_50 bl[50] br[50] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_51 bl[51] br[51] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_52 bl[52] br[52] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_53 bl[53] br[53] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_54 bl[54] br[54] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_55 bl[55] br[55] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_56 bl[56] br[56] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_57 bl[57] br[57] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_58 bl[58] br[58] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_59 bl[59] br[59] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_60 bl[60] br[60] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_61 bl[61] br[61] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_62 bl[62] br[62] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_84_63 bl[63] br[63] vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xcell_85_0 bl[0] br[0] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_1 bl[1] br[1] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_2 bl[2] br[2] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_3 bl[3] br[3] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_4 bl[4] br[4] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_5 bl[5] br[5] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_6 bl[6] br[6] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_7 bl[7] br[7] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_8 bl[8] br[8] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_9 bl[9] br[9] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_10 bl[10] br[10] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_11 bl[11] br[11] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_12 bl[12] br[12] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_13 bl[13] br[13] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_14 bl[14] br[14] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_15 bl[15] br[15] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_16 bl[16] br[16] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_17 bl[17] br[17] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_18 bl[18] br[18] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_19 bl[19] br[19] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_20 bl[20] br[20] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_21 bl[21] br[21] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_22 bl[22] br[22] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_23 bl[23] br[23] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_24 bl[24] br[24] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_25 bl[25] br[25] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_26 bl[26] br[26] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_27 bl[27] br[27] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_28 bl[28] br[28] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_29 bl[29] br[29] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_30 bl[30] br[30] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_31 bl[31] br[31] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_32 bl[32] br[32] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_33 bl[33] br[33] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_34 bl[34] br[34] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_35 bl[35] br[35] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_36 bl[36] br[36] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_37 bl[37] br[37] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_38 bl[38] br[38] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_39 bl[39] br[39] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_40 bl[40] br[40] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_41 bl[41] br[41] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_42 bl[42] br[42] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_43 bl[43] br[43] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_44 bl[44] br[44] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_45 bl[45] br[45] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_46 bl[46] br[46] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_47 bl[47] br[47] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_48 bl[48] br[48] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_49 bl[49] br[49] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_50 bl[50] br[50] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_51 bl[51] br[51] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_52 bl[52] br[52] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_53 bl[53] br[53] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_54 bl[54] br[54] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_55 bl[55] br[55] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_56 bl[56] br[56] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_57 bl[57] br[57] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_58 bl[58] br[58] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_59 bl[59] br[59] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_60 bl[60] br[60] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_61 bl[61] br[61] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_62 bl[62] br[62] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_85_63 bl[63] br[63] vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xcell_86_0 bl[0] br[0] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_1 bl[1] br[1] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_2 bl[2] br[2] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_3 bl[3] br[3] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_4 bl[4] br[4] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_5 bl[5] br[5] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_6 bl[6] br[6] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_7 bl[7] br[7] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_8 bl[8] br[8] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_9 bl[9] br[9] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_10 bl[10] br[10] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_11 bl[11] br[11] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_12 bl[12] br[12] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_13 bl[13] br[13] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_14 bl[14] br[14] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_15 bl[15] br[15] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_16 bl[16] br[16] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_17 bl[17] br[17] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_18 bl[18] br[18] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_19 bl[19] br[19] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_20 bl[20] br[20] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_21 bl[21] br[21] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_22 bl[22] br[22] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_23 bl[23] br[23] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_24 bl[24] br[24] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_25 bl[25] br[25] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_26 bl[26] br[26] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_27 bl[27] br[27] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_28 bl[28] br[28] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_29 bl[29] br[29] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_30 bl[30] br[30] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_31 bl[31] br[31] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_32 bl[32] br[32] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_33 bl[33] br[33] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_34 bl[34] br[34] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_35 bl[35] br[35] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_36 bl[36] br[36] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_37 bl[37] br[37] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_38 bl[38] br[38] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_39 bl[39] br[39] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_40 bl[40] br[40] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_41 bl[41] br[41] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_42 bl[42] br[42] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_43 bl[43] br[43] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_44 bl[44] br[44] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_45 bl[45] br[45] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_46 bl[46] br[46] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_47 bl[47] br[47] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_48 bl[48] br[48] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_49 bl[49] br[49] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_50 bl[50] br[50] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_51 bl[51] br[51] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_52 bl[52] br[52] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_53 bl[53] br[53] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_54 bl[54] br[54] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_55 bl[55] br[55] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_56 bl[56] br[56] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_57 bl[57] br[57] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_58 bl[58] br[58] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_59 bl[59] br[59] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_60 bl[60] br[60] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_61 bl[61] br[61] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_62 bl[62] br[62] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_86_63 bl[63] br[63] vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xcell_87_0 bl[0] br[0] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_1 bl[1] br[1] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_2 bl[2] br[2] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_3 bl[3] br[3] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_4 bl[4] br[4] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_5 bl[5] br[5] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_6 bl[6] br[6] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_7 bl[7] br[7] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_8 bl[8] br[8] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_9 bl[9] br[9] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_10 bl[10] br[10] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_11 bl[11] br[11] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_12 bl[12] br[12] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_13 bl[13] br[13] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_14 bl[14] br[14] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_15 bl[15] br[15] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_16 bl[16] br[16] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_17 bl[17] br[17] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_18 bl[18] br[18] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_19 bl[19] br[19] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_20 bl[20] br[20] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_21 bl[21] br[21] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_22 bl[22] br[22] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_23 bl[23] br[23] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_24 bl[24] br[24] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_25 bl[25] br[25] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_26 bl[26] br[26] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_27 bl[27] br[27] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_28 bl[28] br[28] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_29 bl[29] br[29] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_30 bl[30] br[30] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_31 bl[31] br[31] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_32 bl[32] br[32] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_33 bl[33] br[33] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_34 bl[34] br[34] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_35 bl[35] br[35] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_36 bl[36] br[36] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_37 bl[37] br[37] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_38 bl[38] br[38] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_39 bl[39] br[39] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_40 bl[40] br[40] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_41 bl[41] br[41] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_42 bl[42] br[42] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_43 bl[43] br[43] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_44 bl[44] br[44] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_45 bl[45] br[45] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_46 bl[46] br[46] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_47 bl[47] br[47] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_48 bl[48] br[48] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_49 bl[49] br[49] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_50 bl[50] br[50] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_51 bl[51] br[51] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_52 bl[52] br[52] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_53 bl[53] br[53] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_54 bl[54] br[54] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_55 bl[55] br[55] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_56 bl[56] br[56] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_57 bl[57] br[57] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_58 bl[58] br[58] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_59 bl[59] br[59] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_60 bl[60] br[60] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_61 bl[61] br[61] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_62 bl[62] br[62] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_87_63 bl[63] br[63] vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xcell_88_0 bl[0] br[0] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_1 bl[1] br[1] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_2 bl[2] br[2] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_3 bl[3] br[3] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_4 bl[4] br[4] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_5 bl[5] br[5] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_6 bl[6] br[6] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_7 bl[7] br[7] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_8 bl[8] br[8] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_9 bl[9] br[9] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_10 bl[10] br[10] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_11 bl[11] br[11] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_12 bl[12] br[12] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_13 bl[13] br[13] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_14 bl[14] br[14] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_15 bl[15] br[15] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_16 bl[16] br[16] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_17 bl[17] br[17] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_18 bl[18] br[18] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_19 bl[19] br[19] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_20 bl[20] br[20] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_21 bl[21] br[21] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_22 bl[22] br[22] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_23 bl[23] br[23] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_24 bl[24] br[24] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_25 bl[25] br[25] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_26 bl[26] br[26] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_27 bl[27] br[27] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_28 bl[28] br[28] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_29 bl[29] br[29] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_30 bl[30] br[30] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_31 bl[31] br[31] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_32 bl[32] br[32] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_33 bl[33] br[33] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_34 bl[34] br[34] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_35 bl[35] br[35] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_36 bl[36] br[36] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_37 bl[37] br[37] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_38 bl[38] br[38] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_39 bl[39] br[39] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_40 bl[40] br[40] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_41 bl[41] br[41] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_42 bl[42] br[42] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_43 bl[43] br[43] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_44 bl[44] br[44] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_45 bl[45] br[45] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_46 bl[46] br[46] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_47 bl[47] br[47] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_48 bl[48] br[48] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_49 bl[49] br[49] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_50 bl[50] br[50] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_51 bl[51] br[51] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_52 bl[52] br[52] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_53 bl[53] br[53] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_54 bl[54] br[54] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_55 bl[55] br[55] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_56 bl[56] br[56] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_57 bl[57] br[57] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_58 bl[58] br[58] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_59 bl[59] br[59] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_60 bl[60] br[60] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_61 bl[61] br[61] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_62 bl[62] br[62] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_88_63 bl[63] br[63] vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xcell_89_0 bl[0] br[0] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_1 bl[1] br[1] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_2 bl[2] br[2] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_3 bl[3] br[3] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_4 bl[4] br[4] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_5 bl[5] br[5] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_6 bl[6] br[6] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_7 bl[7] br[7] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_8 bl[8] br[8] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_9 bl[9] br[9] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_10 bl[10] br[10] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_11 bl[11] br[11] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_12 bl[12] br[12] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_13 bl[13] br[13] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_14 bl[14] br[14] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_15 bl[15] br[15] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_16 bl[16] br[16] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_17 bl[17] br[17] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_18 bl[18] br[18] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_19 bl[19] br[19] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_20 bl[20] br[20] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_21 bl[21] br[21] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_22 bl[22] br[22] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_23 bl[23] br[23] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_24 bl[24] br[24] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_25 bl[25] br[25] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_26 bl[26] br[26] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_27 bl[27] br[27] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_28 bl[28] br[28] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_29 bl[29] br[29] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_30 bl[30] br[30] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_31 bl[31] br[31] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_32 bl[32] br[32] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_33 bl[33] br[33] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_34 bl[34] br[34] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_35 bl[35] br[35] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_36 bl[36] br[36] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_37 bl[37] br[37] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_38 bl[38] br[38] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_39 bl[39] br[39] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_40 bl[40] br[40] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_41 bl[41] br[41] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_42 bl[42] br[42] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_43 bl[43] br[43] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_44 bl[44] br[44] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_45 bl[45] br[45] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_46 bl[46] br[46] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_47 bl[47] br[47] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_48 bl[48] br[48] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_49 bl[49] br[49] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_50 bl[50] br[50] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_51 bl[51] br[51] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_52 bl[52] br[52] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_53 bl[53] br[53] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_54 bl[54] br[54] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_55 bl[55] br[55] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_56 bl[56] br[56] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_57 bl[57] br[57] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_58 bl[58] br[58] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_59 bl[59] br[59] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_60 bl[60] br[60] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_61 bl[61] br[61] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_62 bl[62] br[62] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_89_63 bl[63] br[63] vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xcell_90_0 bl[0] br[0] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_1 bl[1] br[1] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_2 bl[2] br[2] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_3 bl[3] br[3] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_4 bl[4] br[4] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_5 bl[5] br[5] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_6 bl[6] br[6] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_7 bl[7] br[7] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_8 bl[8] br[8] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_9 bl[9] br[9] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_10 bl[10] br[10] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_11 bl[11] br[11] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_12 bl[12] br[12] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_13 bl[13] br[13] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_14 bl[14] br[14] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_15 bl[15] br[15] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_16 bl[16] br[16] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_17 bl[17] br[17] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_18 bl[18] br[18] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_19 bl[19] br[19] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_20 bl[20] br[20] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_21 bl[21] br[21] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_22 bl[22] br[22] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_23 bl[23] br[23] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_24 bl[24] br[24] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_25 bl[25] br[25] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_26 bl[26] br[26] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_27 bl[27] br[27] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_28 bl[28] br[28] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_29 bl[29] br[29] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_30 bl[30] br[30] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_31 bl[31] br[31] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_32 bl[32] br[32] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_33 bl[33] br[33] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_34 bl[34] br[34] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_35 bl[35] br[35] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_36 bl[36] br[36] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_37 bl[37] br[37] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_38 bl[38] br[38] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_39 bl[39] br[39] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_40 bl[40] br[40] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_41 bl[41] br[41] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_42 bl[42] br[42] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_43 bl[43] br[43] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_44 bl[44] br[44] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_45 bl[45] br[45] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_46 bl[46] br[46] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_47 bl[47] br[47] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_48 bl[48] br[48] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_49 bl[49] br[49] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_50 bl[50] br[50] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_51 bl[51] br[51] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_52 bl[52] br[52] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_53 bl[53] br[53] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_54 bl[54] br[54] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_55 bl[55] br[55] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_56 bl[56] br[56] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_57 bl[57] br[57] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_58 bl[58] br[58] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_59 bl[59] br[59] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_60 bl[60] br[60] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_61 bl[61] br[61] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_62 bl[62] br[62] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_90_63 bl[63] br[63] vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xcell_91_0 bl[0] br[0] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_1 bl[1] br[1] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_2 bl[2] br[2] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_3 bl[3] br[3] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_4 bl[4] br[4] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_5 bl[5] br[5] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_6 bl[6] br[6] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_7 bl[7] br[7] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_8 bl[8] br[8] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_9 bl[9] br[9] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_10 bl[10] br[10] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_11 bl[11] br[11] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_12 bl[12] br[12] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_13 bl[13] br[13] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_14 bl[14] br[14] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_15 bl[15] br[15] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_16 bl[16] br[16] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_17 bl[17] br[17] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_18 bl[18] br[18] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_19 bl[19] br[19] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_20 bl[20] br[20] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_21 bl[21] br[21] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_22 bl[22] br[22] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_23 bl[23] br[23] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_24 bl[24] br[24] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_25 bl[25] br[25] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_26 bl[26] br[26] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_27 bl[27] br[27] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_28 bl[28] br[28] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_29 bl[29] br[29] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_30 bl[30] br[30] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_31 bl[31] br[31] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_32 bl[32] br[32] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_33 bl[33] br[33] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_34 bl[34] br[34] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_35 bl[35] br[35] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_36 bl[36] br[36] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_37 bl[37] br[37] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_38 bl[38] br[38] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_39 bl[39] br[39] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_40 bl[40] br[40] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_41 bl[41] br[41] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_42 bl[42] br[42] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_43 bl[43] br[43] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_44 bl[44] br[44] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_45 bl[45] br[45] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_46 bl[46] br[46] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_47 bl[47] br[47] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_48 bl[48] br[48] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_49 bl[49] br[49] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_50 bl[50] br[50] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_51 bl[51] br[51] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_52 bl[52] br[52] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_53 bl[53] br[53] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_54 bl[54] br[54] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_55 bl[55] br[55] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_56 bl[56] br[56] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_57 bl[57] br[57] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_58 bl[58] br[58] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_59 bl[59] br[59] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_60 bl[60] br[60] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_61 bl[61] br[61] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_62 bl[62] br[62] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_91_63 bl[63] br[63] vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xcell_92_0 bl[0] br[0] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_1 bl[1] br[1] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_2 bl[2] br[2] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_3 bl[3] br[3] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_4 bl[4] br[4] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_5 bl[5] br[5] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_6 bl[6] br[6] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_7 bl[7] br[7] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_8 bl[8] br[8] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_9 bl[9] br[9] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_10 bl[10] br[10] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_11 bl[11] br[11] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_12 bl[12] br[12] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_13 bl[13] br[13] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_14 bl[14] br[14] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_15 bl[15] br[15] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_16 bl[16] br[16] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_17 bl[17] br[17] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_18 bl[18] br[18] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_19 bl[19] br[19] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_20 bl[20] br[20] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_21 bl[21] br[21] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_22 bl[22] br[22] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_23 bl[23] br[23] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_24 bl[24] br[24] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_25 bl[25] br[25] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_26 bl[26] br[26] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_27 bl[27] br[27] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_28 bl[28] br[28] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_29 bl[29] br[29] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_30 bl[30] br[30] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_31 bl[31] br[31] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_32 bl[32] br[32] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_33 bl[33] br[33] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_34 bl[34] br[34] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_35 bl[35] br[35] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_36 bl[36] br[36] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_37 bl[37] br[37] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_38 bl[38] br[38] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_39 bl[39] br[39] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_40 bl[40] br[40] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_41 bl[41] br[41] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_42 bl[42] br[42] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_43 bl[43] br[43] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_44 bl[44] br[44] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_45 bl[45] br[45] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_46 bl[46] br[46] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_47 bl[47] br[47] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_48 bl[48] br[48] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_49 bl[49] br[49] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_50 bl[50] br[50] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_51 bl[51] br[51] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_52 bl[52] br[52] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_53 bl[53] br[53] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_54 bl[54] br[54] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_55 bl[55] br[55] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_56 bl[56] br[56] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_57 bl[57] br[57] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_58 bl[58] br[58] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_59 bl[59] br[59] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_60 bl[60] br[60] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_61 bl[61] br[61] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_62 bl[62] br[62] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_92_63 bl[63] br[63] vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xcell_93_0 bl[0] br[0] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_1 bl[1] br[1] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_2 bl[2] br[2] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_3 bl[3] br[3] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_4 bl[4] br[4] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_5 bl[5] br[5] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_6 bl[6] br[6] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_7 bl[7] br[7] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_8 bl[8] br[8] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_9 bl[9] br[9] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_10 bl[10] br[10] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_11 bl[11] br[11] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_12 bl[12] br[12] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_13 bl[13] br[13] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_14 bl[14] br[14] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_15 bl[15] br[15] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_16 bl[16] br[16] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_17 bl[17] br[17] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_18 bl[18] br[18] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_19 bl[19] br[19] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_20 bl[20] br[20] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_21 bl[21] br[21] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_22 bl[22] br[22] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_23 bl[23] br[23] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_24 bl[24] br[24] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_25 bl[25] br[25] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_26 bl[26] br[26] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_27 bl[27] br[27] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_28 bl[28] br[28] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_29 bl[29] br[29] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_30 bl[30] br[30] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_31 bl[31] br[31] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_32 bl[32] br[32] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_33 bl[33] br[33] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_34 bl[34] br[34] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_35 bl[35] br[35] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_36 bl[36] br[36] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_37 bl[37] br[37] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_38 bl[38] br[38] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_39 bl[39] br[39] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_40 bl[40] br[40] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_41 bl[41] br[41] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_42 bl[42] br[42] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_43 bl[43] br[43] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_44 bl[44] br[44] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_45 bl[45] br[45] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_46 bl[46] br[46] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_47 bl[47] br[47] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_48 bl[48] br[48] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_49 bl[49] br[49] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_50 bl[50] br[50] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_51 bl[51] br[51] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_52 bl[52] br[52] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_53 bl[53] br[53] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_54 bl[54] br[54] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_55 bl[55] br[55] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_56 bl[56] br[56] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_57 bl[57] br[57] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_58 bl[58] br[58] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_59 bl[59] br[59] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_60 bl[60] br[60] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_61 bl[61] br[61] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_62 bl[62] br[62] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_93_63 bl[63] br[63] vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xcell_94_0 bl[0] br[0] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_1 bl[1] br[1] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_2 bl[2] br[2] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_3 bl[3] br[3] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_4 bl[4] br[4] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_5 bl[5] br[5] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_6 bl[6] br[6] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_7 bl[7] br[7] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_8 bl[8] br[8] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_9 bl[9] br[9] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_10 bl[10] br[10] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_11 bl[11] br[11] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_12 bl[12] br[12] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_13 bl[13] br[13] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_14 bl[14] br[14] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_15 bl[15] br[15] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_16 bl[16] br[16] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_17 bl[17] br[17] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_18 bl[18] br[18] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_19 bl[19] br[19] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_20 bl[20] br[20] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_21 bl[21] br[21] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_22 bl[22] br[22] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_23 bl[23] br[23] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_24 bl[24] br[24] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_25 bl[25] br[25] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_26 bl[26] br[26] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_27 bl[27] br[27] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_28 bl[28] br[28] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_29 bl[29] br[29] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_30 bl[30] br[30] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_31 bl[31] br[31] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_32 bl[32] br[32] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_33 bl[33] br[33] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_34 bl[34] br[34] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_35 bl[35] br[35] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_36 bl[36] br[36] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_37 bl[37] br[37] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_38 bl[38] br[38] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_39 bl[39] br[39] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_40 bl[40] br[40] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_41 bl[41] br[41] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_42 bl[42] br[42] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_43 bl[43] br[43] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_44 bl[44] br[44] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_45 bl[45] br[45] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_46 bl[46] br[46] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_47 bl[47] br[47] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_48 bl[48] br[48] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_49 bl[49] br[49] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_50 bl[50] br[50] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_51 bl[51] br[51] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_52 bl[52] br[52] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_53 bl[53] br[53] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_54 bl[54] br[54] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_55 bl[55] br[55] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_56 bl[56] br[56] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_57 bl[57] br[57] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_58 bl[58] br[58] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_59 bl[59] br[59] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_60 bl[60] br[60] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_61 bl[61] br[61] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_62 bl[62] br[62] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_94_63 bl[63] br[63] vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xcell_95_0 bl[0] br[0] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_1 bl[1] br[1] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_2 bl[2] br[2] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_3 bl[3] br[3] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_4 bl[4] br[4] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_5 bl[5] br[5] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_6 bl[6] br[6] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_7 bl[7] br[7] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_8 bl[8] br[8] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_9 bl[9] br[9] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_10 bl[10] br[10] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_11 bl[11] br[11] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_12 bl[12] br[12] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_13 bl[13] br[13] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_14 bl[14] br[14] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_15 bl[15] br[15] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_16 bl[16] br[16] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_17 bl[17] br[17] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_18 bl[18] br[18] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_19 bl[19] br[19] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_20 bl[20] br[20] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_21 bl[21] br[21] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_22 bl[22] br[22] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_23 bl[23] br[23] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_24 bl[24] br[24] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_25 bl[25] br[25] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_26 bl[26] br[26] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_27 bl[27] br[27] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_28 bl[28] br[28] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_29 bl[29] br[29] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_30 bl[30] br[30] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_31 bl[31] br[31] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_32 bl[32] br[32] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_33 bl[33] br[33] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_34 bl[34] br[34] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_35 bl[35] br[35] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_36 bl[36] br[36] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_37 bl[37] br[37] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_38 bl[38] br[38] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_39 bl[39] br[39] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_40 bl[40] br[40] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_41 bl[41] br[41] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_42 bl[42] br[42] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_43 bl[43] br[43] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_44 bl[44] br[44] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_45 bl[45] br[45] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_46 bl[46] br[46] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_47 bl[47] br[47] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_48 bl[48] br[48] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_49 bl[49] br[49] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_50 bl[50] br[50] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_51 bl[51] br[51] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_52 bl[52] br[52] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_53 bl[53] br[53] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_54 bl[54] br[54] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_55 bl[55] br[55] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_56 bl[56] br[56] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_57 bl[57] br[57] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_58 bl[58] br[58] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_59 bl[59] br[59] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_60 bl[60] br[60] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_61 bl[61] br[61] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_62 bl[62] br[62] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_95_63 bl[63] br[63] vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xcell_96_0 bl[0] br[0] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_1 bl[1] br[1] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_2 bl[2] br[2] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_3 bl[3] br[3] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_4 bl[4] br[4] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_5 bl[5] br[5] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_6 bl[6] br[6] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_7 bl[7] br[7] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_8 bl[8] br[8] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_9 bl[9] br[9] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_10 bl[10] br[10] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_11 bl[11] br[11] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_12 bl[12] br[12] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_13 bl[13] br[13] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_14 bl[14] br[14] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_15 bl[15] br[15] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_16 bl[16] br[16] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_17 bl[17] br[17] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_18 bl[18] br[18] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_19 bl[19] br[19] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_20 bl[20] br[20] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_21 bl[21] br[21] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_22 bl[22] br[22] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_23 bl[23] br[23] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_24 bl[24] br[24] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_25 bl[25] br[25] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_26 bl[26] br[26] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_27 bl[27] br[27] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_28 bl[28] br[28] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_29 bl[29] br[29] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_30 bl[30] br[30] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_31 bl[31] br[31] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_32 bl[32] br[32] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_33 bl[33] br[33] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_34 bl[34] br[34] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_35 bl[35] br[35] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_36 bl[36] br[36] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_37 bl[37] br[37] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_38 bl[38] br[38] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_39 bl[39] br[39] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_40 bl[40] br[40] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_41 bl[41] br[41] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_42 bl[42] br[42] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_43 bl[43] br[43] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_44 bl[44] br[44] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_45 bl[45] br[45] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_46 bl[46] br[46] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_47 bl[47] br[47] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_48 bl[48] br[48] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_49 bl[49] br[49] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_50 bl[50] br[50] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_51 bl[51] br[51] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_52 bl[52] br[52] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_53 bl[53] br[53] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_54 bl[54] br[54] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_55 bl[55] br[55] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_56 bl[56] br[56] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_57 bl[57] br[57] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_58 bl[58] br[58] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_59 bl[59] br[59] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_60 bl[60] br[60] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_61 bl[61] br[61] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_62 bl[62] br[62] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_96_63 bl[63] br[63] vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xcell_97_0 bl[0] br[0] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_1 bl[1] br[1] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_2 bl[2] br[2] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_3 bl[3] br[3] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_4 bl[4] br[4] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_5 bl[5] br[5] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_6 bl[6] br[6] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_7 bl[7] br[7] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_8 bl[8] br[8] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_9 bl[9] br[9] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_10 bl[10] br[10] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_11 bl[11] br[11] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_12 bl[12] br[12] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_13 bl[13] br[13] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_14 bl[14] br[14] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_15 bl[15] br[15] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_16 bl[16] br[16] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_17 bl[17] br[17] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_18 bl[18] br[18] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_19 bl[19] br[19] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_20 bl[20] br[20] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_21 bl[21] br[21] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_22 bl[22] br[22] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_23 bl[23] br[23] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_24 bl[24] br[24] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_25 bl[25] br[25] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_26 bl[26] br[26] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_27 bl[27] br[27] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_28 bl[28] br[28] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_29 bl[29] br[29] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_30 bl[30] br[30] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_31 bl[31] br[31] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_32 bl[32] br[32] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_33 bl[33] br[33] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_34 bl[34] br[34] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_35 bl[35] br[35] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_36 bl[36] br[36] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_37 bl[37] br[37] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_38 bl[38] br[38] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_39 bl[39] br[39] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_40 bl[40] br[40] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_41 bl[41] br[41] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_42 bl[42] br[42] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_43 bl[43] br[43] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_44 bl[44] br[44] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_45 bl[45] br[45] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_46 bl[46] br[46] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_47 bl[47] br[47] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_48 bl[48] br[48] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_49 bl[49] br[49] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_50 bl[50] br[50] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_51 bl[51] br[51] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_52 bl[52] br[52] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_53 bl[53] br[53] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_54 bl[54] br[54] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_55 bl[55] br[55] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_56 bl[56] br[56] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_57 bl[57] br[57] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_58 bl[58] br[58] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_59 bl[59] br[59] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_60 bl[60] br[60] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_61 bl[61] br[61] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_62 bl[62] br[62] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_97_63 bl[63] br[63] vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xcell_98_0 bl[0] br[0] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_1 bl[1] br[1] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_2 bl[2] br[2] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_3 bl[3] br[3] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_4 bl[4] br[4] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_5 bl[5] br[5] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_6 bl[6] br[6] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_7 bl[7] br[7] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_8 bl[8] br[8] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_9 bl[9] br[9] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_10 bl[10] br[10] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_11 bl[11] br[11] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_12 bl[12] br[12] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_13 bl[13] br[13] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_14 bl[14] br[14] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_15 bl[15] br[15] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_16 bl[16] br[16] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_17 bl[17] br[17] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_18 bl[18] br[18] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_19 bl[19] br[19] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_20 bl[20] br[20] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_21 bl[21] br[21] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_22 bl[22] br[22] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_23 bl[23] br[23] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_24 bl[24] br[24] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_25 bl[25] br[25] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_26 bl[26] br[26] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_27 bl[27] br[27] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_28 bl[28] br[28] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_29 bl[29] br[29] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_30 bl[30] br[30] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_31 bl[31] br[31] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_32 bl[32] br[32] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_33 bl[33] br[33] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_34 bl[34] br[34] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_35 bl[35] br[35] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_36 bl[36] br[36] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_37 bl[37] br[37] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_38 bl[38] br[38] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_39 bl[39] br[39] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_40 bl[40] br[40] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_41 bl[41] br[41] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_42 bl[42] br[42] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_43 bl[43] br[43] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_44 bl[44] br[44] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_45 bl[45] br[45] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_46 bl[46] br[46] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_47 bl[47] br[47] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_48 bl[48] br[48] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_49 bl[49] br[49] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_50 bl[50] br[50] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_51 bl[51] br[51] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_52 bl[52] br[52] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_53 bl[53] br[53] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_54 bl[54] br[54] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_55 bl[55] br[55] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_56 bl[56] br[56] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_57 bl[57] br[57] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_58 bl[58] br[58] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_59 bl[59] br[59] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_60 bl[60] br[60] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_61 bl[61] br[61] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_62 bl[62] br[62] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_98_63 bl[63] br[63] vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xcell_99_0 bl[0] br[0] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_1 bl[1] br[1] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_2 bl[2] br[2] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_3 bl[3] br[3] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_4 bl[4] br[4] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_5 bl[5] br[5] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_6 bl[6] br[6] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_7 bl[7] br[7] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_8 bl[8] br[8] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_9 bl[9] br[9] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_10 bl[10] br[10] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_11 bl[11] br[11] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_12 bl[12] br[12] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_13 bl[13] br[13] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_14 bl[14] br[14] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_15 bl[15] br[15] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_16 bl[16] br[16] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_17 bl[17] br[17] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_18 bl[18] br[18] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_19 bl[19] br[19] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_20 bl[20] br[20] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_21 bl[21] br[21] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_22 bl[22] br[22] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_23 bl[23] br[23] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_24 bl[24] br[24] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_25 bl[25] br[25] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_26 bl[26] br[26] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_27 bl[27] br[27] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_28 bl[28] br[28] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_29 bl[29] br[29] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_30 bl[30] br[30] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_31 bl[31] br[31] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_32 bl[32] br[32] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_33 bl[33] br[33] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_34 bl[34] br[34] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_35 bl[35] br[35] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_36 bl[36] br[36] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_37 bl[37] br[37] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_38 bl[38] br[38] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_39 bl[39] br[39] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_40 bl[40] br[40] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_41 bl[41] br[41] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_42 bl[42] br[42] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_43 bl[43] br[43] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_44 bl[44] br[44] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_45 bl[45] br[45] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_46 bl[46] br[46] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_47 bl[47] br[47] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_48 bl[48] br[48] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_49 bl[49] br[49] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_50 bl[50] br[50] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_51 bl[51] br[51] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_52 bl[52] br[52] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_53 bl[53] br[53] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_54 bl[54] br[54] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_55 bl[55] br[55] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_56 bl[56] br[56] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_57 bl[57] br[57] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_58 bl[58] br[58] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_59 bl[59] br[59] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_60 bl[60] br[60] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_61 bl[61] br[61] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_62 bl[62] br[62] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_99_63 bl[63] br[63] vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xcell_100_0 bl[0] br[0] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_1 bl[1] br[1] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_2 bl[2] br[2] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_3 bl[3] br[3] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_4 bl[4] br[4] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_5 bl[5] br[5] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_6 bl[6] br[6] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_7 bl[7] br[7] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_8 bl[8] br[8] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_9 bl[9] br[9] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_10 bl[10] br[10] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_11 bl[11] br[11] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_12 bl[12] br[12] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_13 bl[13] br[13] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_14 bl[14] br[14] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_15 bl[15] br[15] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_16 bl[16] br[16] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_17 bl[17] br[17] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_18 bl[18] br[18] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_19 bl[19] br[19] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_20 bl[20] br[20] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_21 bl[21] br[21] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_22 bl[22] br[22] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_23 bl[23] br[23] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_24 bl[24] br[24] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_25 bl[25] br[25] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_26 bl[26] br[26] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_27 bl[27] br[27] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_28 bl[28] br[28] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_29 bl[29] br[29] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_30 bl[30] br[30] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_31 bl[31] br[31] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_32 bl[32] br[32] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_33 bl[33] br[33] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_34 bl[34] br[34] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_35 bl[35] br[35] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_36 bl[36] br[36] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_37 bl[37] br[37] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_38 bl[38] br[38] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_39 bl[39] br[39] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_40 bl[40] br[40] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_41 bl[41] br[41] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_42 bl[42] br[42] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_43 bl[43] br[43] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_44 bl[44] br[44] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_45 bl[45] br[45] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_46 bl[46] br[46] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_47 bl[47] br[47] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_48 bl[48] br[48] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_49 bl[49] br[49] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_50 bl[50] br[50] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_51 bl[51] br[51] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_52 bl[52] br[52] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_53 bl[53] br[53] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_54 bl[54] br[54] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_55 bl[55] br[55] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_56 bl[56] br[56] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_57 bl[57] br[57] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_58 bl[58] br[58] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_59 bl[59] br[59] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_60 bl[60] br[60] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_61 bl[61] br[61] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_62 bl[62] br[62] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_100_63 bl[63] br[63] vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xcell_101_0 bl[0] br[0] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_1 bl[1] br[1] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_2 bl[2] br[2] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_3 bl[3] br[3] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_4 bl[4] br[4] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_5 bl[5] br[5] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_6 bl[6] br[6] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_7 bl[7] br[7] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_8 bl[8] br[8] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_9 bl[9] br[9] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_10 bl[10] br[10] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_11 bl[11] br[11] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_12 bl[12] br[12] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_13 bl[13] br[13] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_14 bl[14] br[14] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_15 bl[15] br[15] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_16 bl[16] br[16] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_17 bl[17] br[17] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_18 bl[18] br[18] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_19 bl[19] br[19] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_20 bl[20] br[20] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_21 bl[21] br[21] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_22 bl[22] br[22] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_23 bl[23] br[23] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_24 bl[24] br[24] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_25 bl[25] br[25] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_26 bl[26] br[26] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_27 bl[27] br[27] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_28 bl[28] br[28] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_29 bl[29] br[29] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_30 bl[30] br[30] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_31 bl[31] br[31] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_32 bl[32] br[32] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_33 bl[33] br[33] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_34 bl[34] br[34] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_35 bl[35] br[35] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_36 bl[36] br[36] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_37 bl[37] br[37] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_38 bl[38] br[38] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_39 bl[39] br[39] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_40 bl[40] br[40] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_41 bl[41] br[41] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_42 bl[42] br[42] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_43 bl[43] br[43] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_44 bl[44] br[44] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_45 bl[45] br[45] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_46 bl[46] br[46] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_47 bl[47] br[47] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_48 bl[48] br[48] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_49 bl[49] br[49] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_50 bl[50] br[50] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_51 bl[51] br[51] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_52 bl[52] br[52] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_53 bl[53] br[53] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_54 bl[54] br[54] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_55 bl[55] br[55] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_56 bl[56] br[56] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_57 bl[57] br[57] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_58 bl[58] br[58] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_59 bl[59] br[59] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_60 bl[60] br[60] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_61 bl[61] br[61] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_62 bl[62] br[62] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_101_63 bl[63] br[63] vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xcell_102_0 bl[0] br[0] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_1 bl[1] br[1] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_2 bl[2] br[2] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_3 bl[3] br[3] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_4 bl[4] br[4] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_5 bl[5] br[5] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_6 bl[6] br[6] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_7 bl[7] br[7] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_8 bl[8] br[8] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_9 bl[9] br[9] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_10 bl[10] br[10] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_11 bl[11] br[11] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_12 bl[12] br[12] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_13 bl[13] br[13] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_14 bl[14] br[14] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_15 bl[15] br[15] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_16 bl[16] br[16] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_17 bl[17] br[17] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_18 bl[18] br[18] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_19 bl[19] br[19] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_20 bl[20] br[20] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_21 bl[21] br[21] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_22 bl[22] br[22] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_23 bl[23] br[23] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_24 bl[24] br[24] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_25 bl[25] br[25] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_26 bl[26] br[26] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_27 bl[27] br[27] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_28 bl[28] br[28] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_29 bl[29] br[29] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_30 bl[30] br[30] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_31 bl[31] br[31] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_32 bl[32] br[32] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_33 bl[33] br[33] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_34 bl[34] br[34] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_35 bl[35] br[35] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_36 bl[36] br[36] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_37 bl[37] br[37] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_38 bl[38] br[38] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_39 bl[39] br[39] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_40 bl[40] br[40] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_41 bl[41] br[41] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_42 bl[42] br[42] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_43 bl[43] br[43] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_44 bl[44] br[44] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_45 bl[45] br[45] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_46 bl[46] br[46] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_47 bl[47] br[47] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_48 bl[48] br[48] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_49 bl[49] br[49] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_50 bl[50] br[50] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_51 bl[51] br[51] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_52 bl[52] br[52] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_53 bl[53] br[53] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_54 bl[54] br[54] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_55 bl[55] br[55] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_56 bl[56] br[56] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_57 bl[57] br[57] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_58 bl[58] br[58] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_59 bl[59] br[59] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_60 bl[60] br[60] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_61 bl[61] br[61] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_62 bl[62] br[62] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_102_63 bl[63] br[63] vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xcell_103_0 bl[0] br[0] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_1 bl[1] br[1] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_2 bl[2] br[2] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_3 bl[3] br[3] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_4 bl[4] br[4] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_5 bl[5] br[5] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_6 bl[6] br[6] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_7 bl[7] br[7] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_8 bl[8] br[8] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_9 bl[9] br[9] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_10 bl[10] br[10] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_11 bl[11] br[11] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_12 bl[12] br[12] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_13 bl[13] br[13] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_14 bl[14] br[14] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_15 bl[15] br[15] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_16 bl[16] br[16] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_17 bl[17] br[17] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_18 bl[18] br[18] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_19 bl[19] br[19] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_20 bl[20] br[20] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_21 bl[21] br[21] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_22 bl[22] br[22] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_23 bl[23] br[23] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_24 bl[24] br[24] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_25 bl[25] br[25] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_26 bl[26] br[26] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_27 bl[27] br[27] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_28 bl[28] br[28] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_29 bl[29] br[29] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_30 bl[30] br[30] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_31 bl[31] br[31] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_32 bl[32] br[32] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_33 bl[33] br[33] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_34 bl[34] br[34] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_35 bl[35] br[35] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_36 bl[36] br[36] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_37 bl[37] br[37] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_38 bl[38] br[38] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_39 bl[39] br[39] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_40 bl[40] br[40] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_41 bl[41] br[41] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_42 bl[42] br[42] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_43 bl[43] br[43] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_44 bl[44] br[44] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_45 bl[45] br[45] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_46 bl[46] br[46] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_47 bl[47] br[47] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_48 bl[48] br[48] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_49 bl[49] br[49] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_50 bl[50] br[50] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_51 bl[51] br[51] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_52 bl[52] br[52] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_53 bl[53] br[53] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_54 bl[54] br[54] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_55 bl[55] br[55] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_56 bl[56] br[56] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_57 bl[57] br[57] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_58 bl[58] br[58] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_59 bl[59] br[59] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_60 bl[60] br[60] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_61 bl[61] br[61] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_62 bl[62] br[62] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_103_63 bl[63] br[63] vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xcell_104_0 bl[0] br[0] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_1 bl[1] br[1] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_2 bl[2] br[2] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_3 bl[3] br[3] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_4 bl[4] br[4] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_5 bl[5] br[5] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_6 bl[6] br[6] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_7 bl[7] br[7] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_8 bl[8] br[8] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_9 bl[9] br[9] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_10 bl[10] br[10] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_11 bl[11] br[11] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_12 bl[12] br[12] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_13 bl[13] br[13] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_14 bl[14] br[14] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_15 bl[15] br[15] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_16 bl[16] br[16] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_17 bl[17] br[17] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_18 bl[18] br[18] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_19 bl[19] br[19] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_20 bl[20] br[20] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_21 bl[21] br[21] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_22 bl[22] br[22] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_23 bl[23] br[23] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_24 bl[24] br[24] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_25 bl[25] br[25] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_26 bl[26] br[26] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_27 bl[27] br[27] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_28 bl[28] br[28] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_29 bl[29] br[29] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_30 bl[30] br[30] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_31 bl[31] br[31] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_32 bl[32] br[32] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_33 bl[33] br[33] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_34 bl[34] br[34] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_35 bl[35] br[35] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_36 bl[36] br[36] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_37 bl[37] br[37] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_38 bl[38] br[38] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_39 bl[39] br[39] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_40 bl[40] br[40] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_41 bl[41] br[41] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_42 bl[42] br[42] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_43 bl[43] br[43] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_44 bl[44] br[44] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_45 bl[45] br[45] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_46 bl[46] br[46] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_47 bl[47] br[47] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_48 bl[48] br[48] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_49 bl[49] br[49] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_50 bl[50] br[50] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_51 bl[51] br[51] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_52 bl[52] br[52] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_53 bl[53] br[53] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_54 bl[54] br[54] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_55 bl[55] br[55] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_56 bl[56] br[56] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_57 bl[57] br[57] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_58 bl[58] br[58] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_59 bl[59] br[59] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_60 bl[60] br[60] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_61 bl[61] br[61] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_62 bl[62] br[62] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_104_63 bl[63] br[63] vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xcell_105_0 bl[0] br[0] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_1 bl[1] br[1] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_2 bl[2] br[2] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_3 bl[3] br[3] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_4 bl[4] br[4] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_5 bl[5] br[5] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_6 bl[6] br[6] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_7 bl[7] br[7] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_8 bl[8] br[8] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_9 bl[9] br[9] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_10 bl[10] br[10] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_11 bl[11] br[11] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_12 bl[12] br[12] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_13 bl[13] br[13] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_14 bl[14] br[14] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_15 bl[15] br[15] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_16 bl[16] br[16] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_17 bl[17] br[17] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_18 bl[18] br[18] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_19 bl[19] br[19] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_20 bl[20] br[20] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_21 bl[21] br[21] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_22 bl[22] br[22] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_23 bl[23] br[23] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_24 bl[24] br[24] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_25 bl[25] br[25] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_26 bl[26] br[26] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_27 bl[27] br[27] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_28 bl[28] br[28] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_29 bl[29] br[29] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_30 bl[30] br[30] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_31 bl[31] br[31] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_32 bl[32] br[32] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_33 bl[33] br[33] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_34 bl[34] br[34] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_35 bl[35] br[35] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_36 bl[36] br[36] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_37 bl[37] br[37] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_38 bl[38] br[38] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_39 bl[39] br[39] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_40 bl[40] br[40] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_41 bl[41] br[41] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_42 bl[42] br[42] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_43 bl[43] br[43] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_44 bl[44] br[44] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_45 bl[45] br[45] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_46 bl[46] br[46] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_47 bl[47] br[47] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_48 bl[48] br[48] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_49 bl[49] br[49] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_50 bl[50] br[50] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_51 bl[51] br[51] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_52 bl[52] br[52] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_53 bl[53] br[53] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_54 bl[54] br[54] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_55 bl[55] br[55] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_56 bl[56] br[56] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_57 bl[57] br[57] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_58 bl[58] br[58] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_59 bl[59] br[59] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_60 bl[60] br[60] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_61 bl[61] br[61] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_62 bl[62] br[62] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_105_63 bl[63] br[63] vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xcell_106_0 bl[0] br[0] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_1 bl[1] br[1] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_2 bl[2] br[2] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_3 bl[3] br[3] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_4 bl[4] br[4] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_5 bl[5] br[5] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_6 bl[6] br[6] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_7 bl[7] br[7] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_8 bl[8] br[8] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_9 bl[9] br[9] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_10 bl[10] br[10] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_11 bl[11] br[11] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_12 bl[12] br[12] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_13 bl[13] br[13] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_14 bl[14] br[14] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_15 bl[15] br[15] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_16 bl[16] br[16] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_17 bl[17] br[17] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_18 bl[18] br[18] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_19 bl[19] br[19] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_20 bl[20] br[20] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_21 bl[21] br[21] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_22 bl[22] br[22] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_23 bl[23] br[23] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_24 bl[24] br[24] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_25 bl[25] br[25] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_26 bl[26] br[26] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_27 bl[27] br[27] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_28 bl[28] br[28] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_29 bl[29] br[29] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_30 bl[30] br[30] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_31 bl[31] br[31] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_32 bl[32] br[32] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_33 bl[33] br[33] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_34 bl[34] br[34] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_35 bl[35] br[35] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_36 bl[36] br[36] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_37 bl[37] br[37] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_38 bl[38] br[38] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_39 bl[39] br[39] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_40 bl[40] br[40] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_41 bl[41] br[41] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_42 bl[42] br[42] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_43 bl[43] br[43] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_44 bl[44] br[44] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_45 bl[45] br[45] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_46 bl[46] br[46] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_47 bl[47] br[47] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_48 bl[48] br[48] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_49 bl[49] br[49] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_50 bl[50] br[50] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_51 bl[51] br[51] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_52 bl[52] br[52] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_53 bl[53] br[53] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_54 bl[54] br[54] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_55 bl[55] br[55] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_56 bl[56] br[56] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_57 bl[57] br[57] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_58 bl[58] br[58] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_59 bl[59] br[59] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_60 bl[60] br[60] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_61 bl[61] br[61] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_62 bl[62] br[62] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_106_63 bl[63] br[63] vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xcell_107_0 bl[0] br[0] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_1 bl[1] br[1] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_2 bl[2] br[2] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_3 bl[3] br[3] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_4 bl[4] br[4] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_5 bl[5] br[5] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_6 bl[6] br[6] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_7 bl[7] br[7] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_8 bl[8] br[8] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_9 bl[9] br[9] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_10 bl[10] br[10] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_11 bl[11] br[11] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_12 bl[12] br[12] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_13 bl[13] br[13] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_14 bl[14] br[14] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_15 bl[15] br[15] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_16 bl[16] br[16] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_17 bl[17] br[17] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_18 bl[18] br[18] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_19 bl[19] br[19] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_20 bl[20] br[20] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_21 bl[21] br[21] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_22 bl[22] br[22] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_23 bl[23] br[23] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_24 bl[24] br[24] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_25 bl[25] br[25] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_26 bl[26] br[26] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_27 bl[27] br[27] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_28 bl[28] br[28] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_29 bl[29] br[29] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_30 bl[30] br[30] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_31 bl[31] br[31] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_32 bl[32] br[32] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_33 bl[33] br[33] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_34 bl[34] br[34] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_35 bl[35] br[35] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_36 bl[36] br[36] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_37 bl[37] br[37] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_38 bl[38] br[38] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_39 bl[39] br[39] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_40 bl[40] br[40] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_41 bl[41] br[41] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_42 bl[42] br[42] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_43 bl[43] br[43] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_44 bl[44] br[44] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_45 bl[45] br[45] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_46 bl[46] br[46] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_47 bl[47] br[47] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_48 bl[48] br[48] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_49 bl[49] br[49] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_50 bl[50] br[50] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_51 bl[51] br[51] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_52 bl[52] br[52] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_53 bl[53] br[53] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_54 bl[54] br[54] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_55 bl[55] br[55] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_56 bl[56] br[56] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_57 bl[57] br[57] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_58 bl[58] br[58] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_59 bl[59] br[59] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_60 bl[60] br[60] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_61 bl[61] br[61] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_62 bl[62] br[62] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_107_63 bl[63] br[63] vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xcell_108_0 bl[0] br[0] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_1 bl[1] br[1] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_2 bl[2] br[2] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_3 bl[3] br[3] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_4 bl[4] br[4] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_5 bl[5] br[5] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_6 bl[6] br[6] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_7 bl[7] br[7] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_8 bl[8] br[8] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_9 bl[9] br[9] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_10 bl[10] br[10] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_11 bl[11] br[11] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_12 bl[12] br[12] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_13 bl[13] br[13] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_14 bl[14] br[14] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_15 bl[15] br[15] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_16 bl[16] br[16] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_17 bl[17] br[17] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_18 bl[18] br[18] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_19 bl[19] br[19] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_20 bl[20] br[20] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_21 bl[21] br[21] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_22 bl[22] br[22] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_23 bl[23] br[23] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_24 bl[24] br[24] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_25 bl[25] br[25] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_26 bl[26] br[26] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_27 bl[27] br[27] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_28 bl[28] br[28] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_29 bl[29] br[29] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_30 bl[30] br[30] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_31 bl[31] br[31] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_32 bl[32] br[32] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_33 bl[33] br[33] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_34 bl[34] br[34] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_35 bl[35] br[35] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_36 bl[36] br[36] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_37 bl[37] br[37] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_38 bl[38] br[38] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_39 bl[39] br[39] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_40 bl[40] br[40] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_41 bl[41] br[41] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_42 bl[42] br[42] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_43 bl[43] br[43] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_44 bl[44] br[44] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_45 bl[45] br[45] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_46 bl[46] br[46] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_47 bl[47] br[47] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_48 bl[48] br[48] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_49 bl[49] br[49] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_50 bl[50] br[50] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_51 bl[51] br[51] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_52 bl[52] br[52] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_53 bl[53] br[53] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_54 bl[54] br[54] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_55 bl[55] br[55] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_56 bl[56] br[56] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_57 bl[57] br[57] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_58 bl[58] br[58] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_59 bl[59] br[59] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_60 bl[60] br[60] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_61 bl[61] br[61] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_62 bl[62] br[62] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_108_63 bl[63] br[63] vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xcell_109_0 bl[0] br[0] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_1 bl[1] br[1] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_2 bl[2] br[2] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_3 bl[3] br[3] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_4 bl[4] br[4] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_5 bl[5] br[5] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_6 bl[6] br[6] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_7 bl[7] br[7] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_8 bl[8] br[8] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_9 bl[9] br[9] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_10 bl[10] br[10] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_11 bl[11] br[11] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_12 bl[12] br[12] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_13 bl[13] br[13] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_14 bl[14] br[14] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_15 bl[15] br[15] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_16 bl[16] br[16] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_17 bl[17] br[17] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_18 bl[18] br[18] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_19 bl[19] br[19] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_20 bl[20] br[20] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_21 bl[21] br[21] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_22 bl[22] br[22] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_23 bl[23] br[23] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_24 bl[24] br[24] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_25 bl[25] br[25] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_26 bl[26] br[26] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_27 bl[27] br[27] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_28 bl[28] br[28] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_29 bl[29] br[29] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_30 bl[30] br[30] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_31 bl[31] br[31] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_32 bl[32] br[32] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_33 bl[33] br[33] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_34 bl[34] br[34] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_35 bl[35] br[35] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_36 bl[36] br[36] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_37 bl[37] br[37] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_38 bl[38] br[38] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_39 bl[39] br[39] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_40 bl[40] br[40] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_41 bl[41] br[41] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_42 bl[42] br[42] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_43 bl[43] br[43] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_44 bl[44] br[44] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_45 bl[45] br[45] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_46 bl[46] br[46] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_47 bl[47] br[47] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_48 bl[48] br[48] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_49 bl[49] br[49] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_50 bl[50] br[50] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_51 bl[51] br[51] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_52 bl[52] br[52] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_53 bl[53] br[53] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_54 bl[54] br[54] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_55 bl[55] br[55] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_56 bl[56] br[56] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_57 bl[57] br[57] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_58 bl[58] br[58] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_59 bl[59] br[59] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_60 bl[60] br[60] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_61 bl[61] br[61] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_62 bl[62] br[62] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_109_63 bl[63] br[63] vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xcell_110_0 bl[0] br[0] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_1 bl[1] br[1] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_2 bl[2] br[2] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_3 bl[3] br[3] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_4 bl[4] br[4] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_5 bl[5] br[5] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_6 bl[6] br[6] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_7 bl[7] br[7] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_8 bl[8] br[8] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_9 bl[9] br[9] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_10 bl[10] br[10] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_11 bl[11] br[11] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_12 bl[12] br[12] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_13 bl[13] br[13] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_14 bl[14] br[14] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_15 bl[15] br[15] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_16 bl[16] br[16] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_17 bl[17] br[17] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_18 bl[18] br[18] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_19 bl[19] br[19] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_20 bl[20] br[20] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_21 bl[21] br[21] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_22 bl[22] br[22] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_23 bl[23] br[23] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_24 bl[24] br[24] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_25 bl[25] br[25] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_26 bl[26] br[26] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_27 bl[27] br[27] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_28 bl[28] br[28] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_29 bl[29] br[29] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_30 bl[30] br[30] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_31 bl[31] br[31] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_32 bl[32] br[32] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_33 bl[33] br[33] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_34 bl[34] br[34] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_35 bl[35] br[35] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_36 bl[36] br[36] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_37 bl[37] br[37] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_38 bl[38] br[38] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_39 bl[39] br[39] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_40 bl[40] br[40] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_41 bl[41] br[41] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_42 bl[42] br[42] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_43 bl[43] br[43] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_44 bl[44] br[44] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_45 bl[45] br[45] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_46 bl[46] br[46] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_47 bl[47] br[47] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_48 bl[48] br[48] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_49 bl[49] br[49] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_50 bl[50] br[50] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_51 bl[51] br[51] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_52 bl[52] br[52] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_53 bl[53] br[53] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_54 bl[54] br[54] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_55 bl[55] br[55] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_56 bl[56] br[56] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_57 bl[57] br[57] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_58 bl[58] br[58] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_59 bl[59] br[59] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_60 bl[60] br[60] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_61 bl[61] br[61] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_62 bl[62] br[62] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_110_63 bl[63] br[63] vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xcell_111_0 bl[0] br[0] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_1 bl[1] br[1] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_2 bl[2] br[2] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_3 bl[3] br[3] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_4 bl[4] br[4] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_5 bl[5] br[5] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_6 bl[6] br[6] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_7 bl[7] br[7] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_8 bl[8] br[8] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_9 bl[9] br[9] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_10 bl[10] br[10] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_11 bl[11] br[11] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_12 bl[12] br[12] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_13 bl[13] br[13] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_14 bl[14] br[14] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_15 bl[15] br[15] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_16 bl[16] br[16] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_17 bl[17] br[17] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_18 bl[18] br[18] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_19 bl[19] br[19] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_20 bl[20] br[20] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_21 bl[21] br[21] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_22 bl[22] br[22] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_23 bl[23] br[23] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_24 bl[24] br[24] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_25 bl[25] br[25] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_26 bl[26] br[26] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_27 bl[27] br[27] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_28 bl[28] br[28] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_29 bl[29] br[29] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_30 bl[30] br[30] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_31 bl[31] br[31] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_32 bl[32] br[32] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_33 bl[33] br[33] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_34 bl[34] br[34] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_35 bl[35] br[35] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_36 bl[36] br[36] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_37 bl[37] br[37] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_38 bl[38] br[38] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_39 bl[39] br[39] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_40 bl[40] br[40] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_41 bl[41] br[41] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_42 bl[42] br[42] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_43 bl[43] br[43] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_44 bl[44] br[44] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_45 bl[45] br[45] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_46 bl[46] br[46] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_47 bl[47] br[47] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_48 bl[48] br[48] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_49 bl[49] br[49] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_50 bl[50] br[50] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_51 bl[51] br[51] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_52 bl[52] br[52] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_53 bl[53] br[53] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_54 bl[54] br[54] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_55 bl[55] br[55] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_56 bl[56] br[56] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_57 bl[57] br[57] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_58 bl[58] br[58] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_59 bl[59] br[59] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_60 bl[60] br[60] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_61 bl[61] br[61] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_62 bl[62] br[62] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_111_63 bl[63] br[63] vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xcell_112_0 bl[0] br[0] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_1 bl[1] br[1] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_2 bl[2] br[2] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_3 bl[3] br[3] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_4 bl[4] br[4] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_5 bl[5] br[5] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_6 bl[6] br[6] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_7 bl[7] br[7] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_8 bl[8] br[8] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_9 bl[9] br[9] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_10 bl[10] br[10] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_11 bl[11] br[11] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_12 bl[12] br[12] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_13 bl[13] br[13] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_14 bl[14] br[14] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_15 bl[15] br[15] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_16 bl[16] br[16] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_17 bl[17] br[17] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_18 bl[18] br[18] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_19 bl[19] br[19] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_20 bl[20] br[20] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_21 bl[21] br[21] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_22 bl[22] br[22] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_23 bl[23] br[23] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_24 bl[24] br[24] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_25 bl[25] br[25] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_26 bl[26] br[26] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_27 bl[27] br[27] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_28 bl[28] br[28] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_29 bl[29] br[29] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_30 bl[30] br[30] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_31 bl[31] br[31] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_32 bl[32] br[32] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_33 bl[33] br[33] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_34 bl[34] br[34] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_35 bl[35] br[35] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_36 bl[36] br[36] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_37 bl[37] br[37] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_38 bl[38] br[38] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_39 bl[39] br[39] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_40 bl[40] br[40] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_41 bl[41] br[41] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_42 bl[42] br[42] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_43 bl[43] br[43] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_44 bl[44] br[44] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_45 bl[45] br[45] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_46 bl[46] br[46] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_47 bl[47] br[47] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_48 bl[48] br[48] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_49 bl[49] br[49] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_50 bl[50] br[50] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_51 bl[51] br[51] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_52 bl[52] br[52] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_53 bl[53] br[53] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_54 bl[54] br[54] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_55 bl[55] br[55] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_56 bl[56] br[56] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_57 bl[57] br[57] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_58 bl[58] br[58] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_59 bl[59] br[59] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_60 bl[60] br[60] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_61 bl[61] br[61] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_62 bl[62] br[62] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_112_63 bl[63] br[63] vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xcell_113_0 bl[0] br[0] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_1 bl[1] br[1] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_2 bl[2] br[2] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_3 bl[3] br[3] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_4 bl[4] br[4] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_5 bl[5] br[5] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_6 bl[6] br[6] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_7 bl[7] br[7] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_8 bl[8] br[8] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_9 bl[9] br[9] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_10 bl[10] br[10] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_11 bl[11] br[11] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_12 bl[12] br[12] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_13 bl[13] br[13] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_14 bl[14] br[14] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_15 bl[15] br[15] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_16 bl[16] br[16] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_17 bl[17] br[17] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_18 bl[18] br[18] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_19 bl[19] br[19] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_20 bl[20] br[20] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_21 bl[21] br[21] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_22 bl[22] br[22] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_23 bl[23] br[23] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_24 bl[24] br[24] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_25 bl[25] br[25] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_26 bl[26] br[26] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_27 bl[27] br[27] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_28 bl[28] br[28] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_29 bl[29] br[29] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_30 bl[30] br[30] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_31 bl[31] br[31] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_32 bl[32] br[32] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_33 bl[33] br[33] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_34 bl[34] br[34] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_35 bl[35] br[35] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_36 bl[36] br[36] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_37 bl[37] br[37] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_38 bl[38] br[38] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_39 bl[39] br[39] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_40 bl[40] br[40] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_41 bl[41] br[41] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_42 bl[42] br[42] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_43 bl[43] br[43] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_44 bl[44] br[44] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_45 bl[45] br[45] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_46 bl[46] br[46] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_47 bl[47] br[47] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_48 bl[48] br[48] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_49 bl[49] br[49] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_50 bl[50] br[50] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_51 bl[51] br[51] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_52 bl[52] br[52] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_53 bl[53] br[53] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_54 bl[54] br[54] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_55 bl[55] br[55] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_56 bl[56] br[56] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_57 bl[57] br[57] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_58 bl[58] br[58] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_59 bl[59] br[59] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_60 bl[60] br[60] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_61 bl[61] br[61] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_62 bl[62] br[62] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_113_63 bl[63] br[63] vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xcell_114_0 bl[0] br[0] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_1 bl[1] br[1] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_2 bl[2] br[2] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_3 bl[3] br[3] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_4 bl[4] br[4] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_5 bl[5] br[5] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_6 bl[6] br[6] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_7 bl[7] br[7] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_8 bl[8] br[8] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_9 bl[9] br[9] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_10 bl[10] br[10] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_11 bl[11] br[11] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_12 bl[12] br[12] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_13 bl[13] br[13] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_14 bl[14] br[14] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_15 bl[15] br[15] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_16 bl[16] br[16] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_17 bl[17] br[17] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_18 bl[18] br[18] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_19 bl[19] br[19] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_20 bl[20] br[20] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_21 bl[21] br[21] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_22 bl[22] br[22] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_23 bl[23] br[23] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_24 bl[24] br[24] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_25 bl[25] br[25] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_26 bl[26] br[26] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_27 bl[27] br[27] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_28 bl[28] br[28] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_29 bl[29] br[29] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_30 bl[30] br[30] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_31 bl[31] br[31] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_32 bl[32] br[32] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_33 bl[33] br[33] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_34 bl[34] br[34] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_35 bl[35] br[35] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_36 bl[36] br[36] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_37 bl[37] br[37] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_38 bl[38] br[38] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_39 bl[39] br[39] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_40 bl[40] br[40] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_41 bl[41] br[41] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_42 bl[42] br[42] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_43 bl[43] br[43] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_44 bl[44] br[44] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_45 bl[45] br[45] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_46 bl[46] br[46] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_47 bl[47] br[47] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_48 bl[48] br[48] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_49 bl[49] br[49] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_50 bl[50] br[50] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_51 bl[51] br[51] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_52 bl[52] br[52] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_53 bl[53] br[53] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_54 bl[54] br[54] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_55 bl[55] br[55] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_56 bl[56] br[56] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_57 bl[57] br[57] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_58 bl[58] br[58] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_59 bl[59] br[59] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_60 bl[60] br[60] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_61 bl[61] br[61] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_62 bl[62] br[62] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_114_63 bl[63] br[63] vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xcell_115_0 bl[0] br[0] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_1 bl[1] br[1] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_2 bl[2] br[2] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_3 bl[3] br[3] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_4 bl[4] br[4] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_5 bl[5] br[5] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_6 bl[6] br[6] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_7 bl[7] br[7] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_8 bl[8] br[8] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_9 bl[9] br[9] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_10 bl[10] br[10] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_11 bl[11] br[11] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_12 bl[12] br[12] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_13 bl[13] br[13] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_14 bl[14] br[14] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_15 bl[15] br[15] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_16 bl[16] br[16] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_17 bl[17] br[17] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_18 bl[18] br[18] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_19 bl[19] br[19] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_20 bl[20] br[20] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_21 bl[21] br[21] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_22 bl[22] br[22] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_23 bl[23] br[23] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_24 bl[24] br[24] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_25 bl[25] br[25] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_26 bl[26] br[26] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_27 bl[27] br[27] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_28 bl[28] br[28] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_29 bl[29] br[29] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_30 bl[30] br[30] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_31 bl[31] br[31] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_32 bl[32] br[32] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_33 bl[33] br[33] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_34 bl[34] br[34] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_35 bl[35] br[35] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_36 bl[36] br[36] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_37 bl[37] br[37] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_38 bl[38] br[38] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_39 bl[39] br[39] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_40 bl[40] br[40] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_41 bl[41] br[41] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_42 bl[42] br[42] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_43 bl[43] br[43] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_44 bl[44] br[44] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_45 bl[45] br[45] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_46 bl[46] br[46] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_47 bl[47] br[47] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_48 bl[48] br[48] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_49 bl[49] br[49] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_50 bl[50] br[50] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_51 bl[51] br[51] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_52 bl[52] br[52] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_53 bl[53] br[53] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_54 bl[54] br[54] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_55 bl[55] br[55] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_56 bl[56] br[56] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_57 bl[57] br[57] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_58 bl[58] br[58] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_59 bl[59] br[59] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_60 bl[60] br[60] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_61 bl[61] br[61] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_62 bl[62] br[62] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_115_63 bl[63] br[63] vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xcell_116_0 bl[0] br[0] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_1 bl[1] br[1] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_2 bl[2] br[2] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_3 bl[3] br[3] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_4 bl[4] br[4] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_5 bl[5] br[5] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_6 bl[6] br[6] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_7 bl[7] br[7] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_8 bl[8] br[8] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_9 bl[9] br[9] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_10 bl[10] br[10] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_11 bl[11] br[11] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_12 bl[12] br[12] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_13 bl[13] br[13] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_14 bl[14] br[14] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_15 bl[15] br[15] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_16 bl[16] br[16] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_17 bl[17] br[17] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_18 bl[18] br[18] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_19 bl[19] br[19] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_20 bl[20] br[20] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_21 bl[21] br[21] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_22 bl[22] br[22] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_23 bl[23] br[23] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_24 bl[24] br[24] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_25 bl[25] br[25] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_26 bl[26] br[26] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_27 bl[27] br[27] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_28 bl[28] br[28] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_29 bl[29] br[29] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_30 bl[30] br[30] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_31 bl[31] br[31] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_32 bl[32] br[32] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_33 bl[33] br[33] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_34 bl[34] br[34] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_35 bl[35] br[35] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_36 bl[36] br[36] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_37 bl[37] br[37] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_38 bl[38] br[38] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_39 bl[39] br[39] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_40 bl[40] br[40] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_41 bl[41] br[41] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_42 bl[42] br[42] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_43 bl[43] br[43] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_44 bl[44] br[44] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_45 bl[45] br[45] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_46 bl[46] br[46] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_47 bl[47] br[47] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_48 bl[48] br[48] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_49 bl[49] br[49] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_50 bl[50] br[50] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_51 bl[51] br[51] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_52 bl[52] br[52] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_53 bl[53] br[53] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_54 bl[54] br[54] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_55 bl[55] br[55] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_56 bl[56] br[56] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_57 bl[57] br[57] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_58 bl[58] br[58] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_59 bl[59] br[59] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_60 bl[60] br[60] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_61 bl[61] br[61] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_62 bl[62] br[62] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_116_63 bl[63] br[63] vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xcell_117_0 bl[0] br[0] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_1 bl[1] br[1] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_2 bl[2] br[2] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_3 bl[3] br[3] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_4 bl[4] br[4] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_5 bl[5] br[5] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_6 bl[6] br[6] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_7 bl[7] br[7] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_8 bl[8] br[8] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_9 bl[9] br[9] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_10 bl[10] br[10] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_11 bl[11] br[11] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_12 bl[12] br[12] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_13 bl[13] br[13] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_14 bl[14] br[14] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_15 bl[15] br[15] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_16 bl[16] br[16] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_17 bl[17] br[17] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_18 bl[18] br[18] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_19 bl[19] br[19] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_20 bl[20] br[20] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_21 bl[21] br[21] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_22 bl[22] br[22] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_23 bl[23] br[23] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_24 bl[24] br[24] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_25 bl[25] br[25] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_26 bl[26] br[26] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_27 bl[27] br[27] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_28 bl[28] br[28] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_29 bl[29] br[29] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_30 bl[30] br[30] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_31 bl[31] br[31] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_32 bl[32] br[32] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_33 bl[33] br[33] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_34 bl[34] br[34] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_35 bl[35] br[35] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_36 bl[36] br[36] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_37 bl[37] br[37] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_38 bl[38] br[38] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_39 bl[39] br[39] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_40 bl[40] br[40] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_41 bl[41] br[41] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_42 bl[42] br[42] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_43 bl[43] br[43] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_44 bl[44] br[44] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_45 bl[45] br[45] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_46 bl[46] br[46] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_47 bl[47] br[47] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_48 bl[48] br[48] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_49 bl[49] br[49] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_50 bl[50] br[50] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_51 bl[51] br[51] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_52 bl[52] br[52] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_53 bl[53] br[53] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_54 bl[54] br[54] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_55 bl[55] br[55] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_56 bl[56] br[56] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_57 bl[57] br[57] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_58 bl[58] br[58] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_59 bl[59] br[59] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_60 bl[60] br[60] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_61 bl[61] br[61] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_62 bl[62] br[62] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_117_63 bl[63] br[63] vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xcell_118_0 bl[0] br[0] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_1 bl[1] br[1] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_2 bl[2] br[2] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_3 bl[3] br[3] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_4 bl[4] br[4] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_5 bl[5] br[5] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_6 bl[6] br[6] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_7 bl[7] br[7] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_8 bl[8] br[8] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_9 bl[9] br[9] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_10 bl[10] br[10] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_11 bl[11] br[11] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_12 bl[12] br[12] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_13 bl[13] br[13] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_14 bl[14] br[14] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_15 bl[15] br[15] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_16 bl[16] br[16] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_17 bl[17] br[17] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_18 bl[18] br[18] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_19 bl[19] br[19] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_20 bl[20] br[20] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_21 bl[21] br[21] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_22 bl[22] br[22] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_23 bl[23] br[23] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_24 bl[24] br[24] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_25 bl[25] br[25] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_26 bl[26] br[26] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_27 bl[27] br[27] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_28 bl[28] br[28] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_29 bl[29] br[29] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_30 bl[30] br[30] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_31 bl[31] br[31] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_32 bl[32] br[32] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_33 bl[33] br[33] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_34 bl[34] br[34] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_35 bl[35] br[35] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_36 bl[36] br[36] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_37 bl[37] br[37] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_38 bl[38] br[38] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_39 bl[39] br[39] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_40 bl[40] br[40] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_41 bl[41] br[41] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_42 bl[42] br[42] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_43 bl[43] br[43] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_44 bl[44] br[44] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_45 bl[45] br[45] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_46 bl[46] br[46] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_47 bl[47] br[47] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_48 bl[48] br[48] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_49 bl[49] br[49] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_50 bl[50] br[50] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_51 bl[51] br[51] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_52 bl[52] br[52] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_53 bl[53] br[53] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_54 bl[54] br[54] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_55 bl[55] br[55] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_56 bl[56] br[56] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_57 bl[57] br[57] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_58 bl[58] br[58] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_59 bl[59] br[59] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_60 bl[60] br[60] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_61 bl[61] br[61] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_62 bl[62] br[62] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_118_63 bl[63] br[63] vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xcell_119_0 bl[0] br[0] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_1 bl[1] br[1] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_2 bl[2] br[2] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_3 bl[3] br[3] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_4 bl[4] br[4] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_5 bl[5] br[5] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_6 bl[6] br[6] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_7 bl[7] br[7] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_8 bl[8] br[8] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_9 bl[9] br[9] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_10 bl[10] br[10] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_11 bl[11] br[11] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_12 bl[12] br[12] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_13 bl[13] br[13] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_14 bl[14] br[14] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_15 bl[15] br[15] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_16 bl[16] br[16] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_17 bl[17] br[17] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_18 bl[18] br[18] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_19 bl[19] br[19] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_20 bl[20] br[20] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_21 bl[21] br[21] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_22 bl[22] br[22] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_23 bl[23] br[23] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_24 bl[24] br[24] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_25 bl[25] br[25] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_26 bl[26] br[26] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_27 bl[27] br[27] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_28 bl[28] br[28] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_29 bl[29] br[29] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_30 bl[30] br[30] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_31 bl[31] br[31] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_32 bl[32] br[32] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_33 bl[33] br[33] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_34 bl[34] br[34] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_35 bl[35] br[35] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_36 bl[36] br[36] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_37 bl[37] br[37] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_38 bl[38] br[38] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_39 bl[39] br[39] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_40 bl[40] br[40] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_41 bl[41] br[41] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_42 bl[42] br[42] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_43 bl[43] br[43] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_44 bl[44] br[44] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_45 bl[45] br[45] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_46 bl[46] br[46] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_47 bl[47] br[47] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_48 bl[48] br[48] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_49 bl[49] br[49] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_50 bl[50] br[50] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_51 bl[51] br[51] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_52 bl[52] br[52] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_53 bl[53] br[53] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_54 bl[54] br[54] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_55 bl[55] br[55] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_56 bl[56] br[56] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_57 bl[57] br[57] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_58 bl[58] br[58] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_59 bl[59] br[59] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_60 bl[60] br[60] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_61 bl[61] br[61] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_62 bl[62] br[62] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_119_63 bl[63] br[63] vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xcell_120_0 bl[0] br[0] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_1 bl[1] br[1] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_2 bl[2] br[2] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_3 bl[3] br[3] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_4 bl[4] br[4] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_5 bl[5] br[5] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_6 bl[6] br[6] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_7 bl[7] br[7] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_8 bl[8] br[8] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_9 bl[9] br[9] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_10 bl[10] br[10] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_11 bl[11] br[11] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_12 bl[12] br[12] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_13 bl[13] br[13] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_14 bl[14] br[14] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_15 bl[15] br[15] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_16 bl[16] br[16] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_17 bl[17] br[17] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_18 bl[18] br[18] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_19 bl[19] br[19] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_20 bl[20] br[20] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_21 bl[21] br[21] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_22 bl[22] br[22] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_23 bl[23] br[23] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_24 bl[24] br[24] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_25 bl[25] br[25] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_26 bl[26] br[26] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_27 bl[27] br[27] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_28 bl[28] br[28] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_29 bl[29] br[29] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_30 bl[30] br[30] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_31 bl[31] br[31] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_32 bl[32] br[32] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_33 bl[33] br[33] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_34 bl[34] br[34] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_35 bl[35] br[35] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_36 bl[36] br[36] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_37 bl[37] br[37] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_38 bl[38] br[38] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_39 bl[39] br[39] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_40 bl[40] br[40] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_41 bl[41] br[41] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_42 bl[42] br[42] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_43 bl[43] br[43] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_44 bl[44] br[44] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_45 bl[45] br[45] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_46 bl[46] br[46] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_47 bl[47] br[47] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_48 bl[48] br[48] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_49 bl[49] br[49] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_50 bl[50] br[50] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_51 bl[51] br[51] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_52 bl[52] br[52] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_53 bl[53] br[53] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_54 bl[54] br[54] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_55 bl[55] br[55] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_56 bl[56] br[56] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_57 bl[57] br[57] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_58 bl[58] br[58] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_59 bl[59] br[59] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_60 bl[60] br[60] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_61 bl[61] br[61] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_62 bl[62] br[62] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_120_63 bl[63] br[63] vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xcell_121_0 bl[0] br[0] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_1 bl[1] br[1] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_2 bl[2] br[2] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_3 bl[3] br[3] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_4 bl[4] br[4] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_5 bl[5] br[5] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_6 bl[6] br[6] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_7 bl[7] br[7] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_8 bl[8] br[8] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_9 bl[9] br[9] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_10 bl[10] br[10] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_11 bl[11] br[11] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_12 bl[12] br[12] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_13 bl[13] br[13] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_14 bl[14] br[14] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_15 bl[15] br[15] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_16 bl[16] br[16] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_17 bl[17] br[17] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_18 bl[18] br[18] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_19 bl[19] br[19] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_20 bl[20] br[20] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_21 bl[21] br[21] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_22 bl[22] br[22] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_23 bl[23] br[23] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_24 bl[24] br[24] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_25 bl[25] br[25] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_26 bl[26] br[26] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_27 bl[27] br[27] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_28 bl[28] br[28] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_29 bl[29] br[29] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_30 bl[30] br[30] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_31 bl[31] br[31] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_32 bl[32] br[32] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_33 bl[33] br[33] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_34 bl[34] br[34] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_35 bl[35] br[35] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_36 bl[36] br[36] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_37 bl[37] br[37] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_38 bl[38] br[38] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_39 bl[39] br[39] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_40 bl[40] br[40] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_41 bl[41] br[41] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_42 bl[42] br[42] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_43 bl[43] br[43] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_44 bl[44] br[44] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_45 bl[45] br[45] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_46 bl[46] br[46] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_47 bl[47] br[47] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_48 bl[48] br[48] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_49 bl[49] br[49] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_50 bl[50] br[50] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_51 bl[51] br[51] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_52 bl[52] br[52] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_53 bl[53] br[53] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_54 bl[54] br[54] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_55 bl[55] br[55] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_56 bl[56] br[56] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_57 bl[57] br[57] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_58 bl[58] br[58] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_59 bl[59] br[59] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_60 bl[60] br[60] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_61 bl[61] br[61] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_62 bl[62] br[62] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_121_63 bl[63] br[63] vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xcell_122_0 bl[0] br[0] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_1 bl[1] br[1] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_2 bl[2] br[2] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_3 bl[3] br[3] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_4 bl[4] br[4] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_5 bl[5] br[5] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_6 bl[6] br[6] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_7 bl[7] br[7] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_8 bl[8] br[8] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_9 bl[9] br[9] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_10 bl[10] br[10] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_11 bl[11] br[11] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_12 bl[12] br[12] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_13 bl[13] br[13] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_14 bl[14] br[14] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_15 bl[15] br[15] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_16 bl[16] br[16] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_17 bl[17] br[17] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_18 bl[18] br[18] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_19 bl[19] br[19] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_20 bl[20] br[20] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_21 bl[21] br[21] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_22 bl[22] br[22] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_23 bl[23] br[23] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_24 bl[24] br[24] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_25 bl[25] br[25] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_26 bl[26] br[26] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_27 bl[27] br[27] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_28 bl[28] br[28] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_29 bl[29] br[29] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_30 bl[30] br[30] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_31 bl[31] br[31] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_32 bl[32] br[32] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_33 bl[33] br[33] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_34 bl[34] br[34] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_35 bl[35] br[35] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_36 bl[36] br[36] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_37 bl[37] br[37] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_38 bl[38] br[38] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_39 bl[39] br[39] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_40 bl[40] br[40] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_41 bl[41] br[41] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_42 bl[42] br[42] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_43 bl[43] br[43] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_44 bl[44] br[44] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_45 bl[45] br[45] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_46 bl[46] br[46] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_47 bl[47] br[47] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_48 bl[48] br[48] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_49 bl[49] br[49] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_50 bl[50] br[50] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_51 bl[51] br[51] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_52 bl[52] br[52] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_53 bl[53] br[53] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_54 bl[54] br[54] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_55 bl[55] br[55] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_56 bl[56] br[56] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_57 bl[57] br[57] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_58 bl[58] br[58] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_59 bl[59] br[59] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_60 bl[60] br[60] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_61 bl[61] br[61] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_62 bl[62] br[62] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_122_63 bl[63] br[63] vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xcell_123_0 bl[0] br[0] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_1 bl[1] br[1] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_2 bl[2] br[2] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_3 bl[3] br[3] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_4 bl[4] br[4] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_5 bl[5] br[5] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_6 bl[6] br[6] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_7 bl[7] br[7] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_8 bl[8] br[8] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_9 bl[9] br[9] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_10 bl[10] br[10] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_11 bl[11] br[11] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_12 bl[12] br[12] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_13 bl[13] br[13] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_14 bl[14] br[14] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_15 bl[15] br[15] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_16 bl[16] br[16] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_17 bl[17] br[17] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_18 bl[18] br[18] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_19 bl[19] br[19] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_20 bl[20] br[20] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_21 bl[21] br[21] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_22 bl[22] br[22] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_23 bl[23] br[23] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_24 bl[24] br[24] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_25 bl[25] br[25] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_26 bl[26] br[26] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_27 bl[27] br[27] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_28 bl[28] br[28] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_29 bl[29] br[29] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_30 bl[30] br[30] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_31 bl[31] br[31] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_32 bl[32] br[32] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_33 bl[33] br[33] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_34 bl[34] br[34] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_35 bl[35] br[35] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_36 bl[36] br[36] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_37 bl[37] br[37] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_38 bl[38] br[38] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_39 bl[39] br[39] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_40 bl[40] br[40] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_41 bl[41] br[41] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_42 bl[42] br[42] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_43 bl[43] br[43] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_44 bl[44] br[44] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_45 bl[45] br[45] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_46 bl[46] br[46] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_47 bl[47] br[47] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_48 bl[48] br[48] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_49 bl[49] br[49] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_50 bl[50] br[50] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_51 bl[51] br[51] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_52 bl[52] br[52] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_53 bl[53] br[53] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_54 bl[54] br[54] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_55 bl[55] br[55] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_56 bl[56] br[56] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_57 bl[57] br[57] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_58 bl[58] br[58] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_59 bl[59] br[59] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_60 bl[60] br[60] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_61 bl[61] br[61] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_62 bl[62] br[62] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_123_63 bl[63] br[63] vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xcell_124_0 bl[0] br[0] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_1 bl[1] br[1] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_2 bl[2] br[2] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_3 bl[3] br[3] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_4 bl[4] br[4] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_5 bl[5] br[5] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_6 bl[6] br[6] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_7 bl[7] br[7] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_8 bl[8] br[8] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_9 bl[9] br[9] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_10 bl[10] br[10] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_11 bl[11] br[11] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_12 bl[12] br[12] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_13 bl[13] br[13] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_14 bl[14] br[14] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_15 bl[15] br[15] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_16 bl[16] br[16] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_17 bl[17] br[17] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_18 bl[18] br[18] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_19 bl[19] br[19] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_20 bl[20] br[20] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_21 bl[21] br[21] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_22 bl[22] br[22] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_23 bl[23] br[23] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_24 bl[24] br[24] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_25 bl[25] br[25] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_26 bl[26] br[26] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_27 bl[27] br[27] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_28 bl[28] br[28] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_29 bl[29] br[29] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_30 bl[30] br[30] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_31 bl[31] br[31] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_32 bl[32] br[32] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_33 bl[33] br[33] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_34 bl[34] br[34] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_35 bl[35] br[35] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_36 bl[36] br[36] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_37 bl[37] br[37] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_38 bl[38] br[38] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_39 bl[39] br[39] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_40 bl[40] br[40] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_41 bl[41] br[41] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_42 bl[42] br[42] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_43 bl[43] br[43] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_44 bl[44] br[44] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_45 bl[45] br[45] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_46 bl[46] br[46] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_47 bl[47] br[47] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_48 bl[48] br[48] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_49 bl[49] br[49] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_50 bl[50] br[50] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_51 bl[51] br[51] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_52 bl[52] br[52] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_53 bl[53] br[53] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_54 bl[54] br[54] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_55 bl[55] br[55] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_56 bl[56] br[56] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_57 bl[57] br[57] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_58 bl[58] br[58] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_59 bl[59] br[59] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_60 bl[60] br[60] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_61 bl[61] br[61] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_62 bl[62] br[62] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_124_63 bl[63] br[63] vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xcell_125_0 bl[0] br[0] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_1 bl[1] br[1] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_2 bl[2] br[2] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_3 bl[3] br[3] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_4 bl[4] br[4] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_5 bl[5] br[5] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_6 bl[6] br[6] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_7 bl[7] br[7] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_8 bl[8] br[8] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_9 bl[9] br[9] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_10 bl[10] br[10] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_11 bl[11] br[11] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_12 bl[12] br[12] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_13 bl[13] br[13] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_14 bl[14] br[14] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_15 bl[15] br[15] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_16 bl[16] br[16] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_17 bl[17] br[17] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_18 bl[18] br[18] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_19 bl[19] br[19] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_20 bl[20] br[20] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_21 bl[21] br[21] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_22 bl[22] br[22] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_23 bl[23] br[23] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_24 bl[24] br[24] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_25 bl[25] br[25] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_26 bl[26] br[26] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_27 bl[27] br[27] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_28 bl[28] br[28] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_29 bl[29] br[29] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_30 bl[30] br[30] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_31 bl[31] br[31] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_32 bl[32] br[32] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_33 bl[33] br[33] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_34 bl[34] br[34] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_35 bl[35] br[35] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_36 bl[36] br[36] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_37 bl[37] br[37] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_38 bl[38] br[38] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_39 bl[39] br[39] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_40 bl[40] br[40] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_41 bl[41] br[41] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_42 bl[42] br[42] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_43 bl[43] br[43] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_44 bl[44] br[44] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_45 bl[45] br[45] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_46 bl[46] br[46] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_47 bl[47] br[47] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_48 bl[48] br[48] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_49 bl[49] br[49] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_50 bl[50] br[50] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_51 bl[51] br[51] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_52 bl[52] br[52] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_53 bl[53] br[53] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_54 bl[54] br[54] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_55 bl[55] br[55] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_56 bl[56] br[56] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_57 bl[57] br[57] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_58 bl[58] br[58] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_59 bl[59] br[59] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_60 bl[60] br[60] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_61 bl[61] br[61] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_62 bl[62] br[62] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_125_63 bl[63] br[63] vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xcell_126_0 bl[0] br[0] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_1 bl[1] br[1] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_2 bl[2] br[2] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_3 bl[3] br[3] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_4 bl[4] br[4] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_5 bl[5] br[5] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_6 bl[6] br[6] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_7 bl[7] br[7] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_8 bl[8] br[8] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_9 bl[9] br[9] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_10 bl[10] br[10] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_11 bl[11] br[11] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_12 bl[12] br[12] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_13 bl[13] br[13] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_14 bl[14] br[14] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_15 bl[15] br[15] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_16 bl[16] br[16] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_17 bl[17] br[17] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_18 bl[18] br[18] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_19 bl[19] br[19] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_20 bl[20] br[20] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_21 bl[21] br[21] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_22 bl[22] br[22] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_23 bl[23] br[23] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_24 bl[24] br[24] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_25 bl[25] br[25] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_26 bl[26] br[26] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_27 bl[27] br[27] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_28 bl[28] br[28] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_29 bl[29] br[29] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_30 bl[30] br[30] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_31 bl[31] br[31] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_32 bl[32] br[32] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_33 bl[33] br[33] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_34 bl[34] br[34] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_35 bl[35] br[35] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_36 bl[36] br[36] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_37 bl[37] br[37] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_38 bl[38] br[38] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_39 bl[39] br[39] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_40 bl[40] br[40] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_41 bl[41] br[41] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_42 bl[42] br[42] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_43 bl[43] br[43] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_44 bl[44] br[44] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_45 bl[45] br[45] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_46 bl[46] br[46] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_47 bl[47] br[47] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_48 bl[48] br[48] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_49 bl[49] br[49] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_50 bl[50] br[50] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_51 bl[51] br[51] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_52 bl[52] br[52] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_53 bl[53] br[53] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_54 bl[54] br[54] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_55 bl[55] br[55] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_56 bl[56] br[56] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_57 bl[57] br[57] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_58 bl[58] br[58] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_59 bl[59] br[59] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_60 bl[60] br[60] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_61 bl[61] br[61] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_62 bl[62] br[62] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_126_63 bl[63] br[63] vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xcell_127_0 bl[0] br[0] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_1 bl[1] br[1] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_2 bl[2] br[2] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_3 bl[3] br[3] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_4 bl[4] br[4] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_5 bl[5] br[5] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_6 bl[6] br[6] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_7 bl[7] br[7] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_8 bl[8] br[8] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_9 bl[9] br[9] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_10 bl[10] br[10] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_11 bl[11] br[11] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_12 bl[12] br[12] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_13 bl[13] br[13] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_14 bl[14] br[14] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_15 bl[15] br[15] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_16 bl[16] br[16] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_17 bl[17] br[17] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_18 bl[18] br[18] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_19 bl[19] br[19] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_20 bl[20] br[20] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_21 bl[21] br[21] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_22 bl[22] br[22] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_23 bl[23] br[23] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_24 bl[24] br[24] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_25 bl[25] br[25] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_26 bl[26] br[26] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_27 bl[27] br[27] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_28 bl[28] br[28] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_29 bl[29] br[29] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_30 bl[30] br[30] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_31 bl[31] br[31] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_32 bl[32] br[32] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_33 bl[33] br[33] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_34 bl[34] br[34] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_35 bl[35] br[35] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_36 bl[36] br[36] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_37 bl[37] br[37] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_38 bl[38] br[38] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_39 bl[39] br[39] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_40 bl[40] br[40] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_41 bl[41] br[41] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_42 bl[42] br[42] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_43 bl[43] br[43] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_44 bl[44] br[44] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_45 bl[45] br[45] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_46 bl[46] br[46] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_47 bl[47] br[47] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_48 bl[48] br[48] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_49 bl[49] br[49] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_50 bl[50] br[50] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_51 bl[51] br[51] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_52 bl[52] br[52] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_53 bl[53] br[53] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_54 bl[54] br[54] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_55 bl[55] br[55] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_56 bl[56] br[56] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_57 bl[57] br[57] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_58 bl[58] br[58] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_59 bl[59] br[59] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_60 bl[60] br[60] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_61 bl[61] br[61] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_62 bl[62] br[62] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_127_63 bl[63] br[63] vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xcell_128_0 bl[0] br[0] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_1 bl[1] br[1] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_2 bl[2] br[2] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_3 bl[3] br[3] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_4 bl[4] br[4] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_5 bl[5] br[5] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_6 bl[6] br[6] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_7 bl[7] br[7] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_8 bl[8] br[8] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_9 bl[9] br[9] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_10 bl[10] br[10] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_11 bl[11] br[11] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_12 bl[12] br[12] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_13 bl[13] br[13] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_14 bl[14] br[14] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_15 bl[15] br[15] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_16 bl[16] br[16] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_17 bl[17] br[17] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_18 bl[18] br[18] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_19 bl[19] br[19] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_20 bl[20] br[20] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_21 bl[21] br[21] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_22 bl[22] br[22] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_23 bl[23] br[23] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_24 bl[24] br[24] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_25 bl[25] br[25] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_26 bl[26] br[26] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_27 bl[27] br[27] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_28 bl[28] br[28] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_29 bl[29] br[29] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_30 bl[30] br[30] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_31 bl[31] br[31] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_32 bl[32] br[32] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_33 bl[33] br[33] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_34 bl[34] br[34] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_35 bl[35] br[35] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_36 bl[36] br[36] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_37 bl[37] br[37] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_38 bl[38] br[38] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_39 bl[39] br[39] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_40 bl[40] br[40] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_41 bl[41] br[41] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_42 bl[42] br[42] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_43 bl[43] br[43] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_44 bl[44] br[44] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_45 bl[45] br[45] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_46 bl[46] br[46] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_47 bl[47] br[47] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_48 bl[48] br[48] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_49 bl[49] br[49] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_50 bl[50] br[50] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_51 bl[51] br[51] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_52 bl[52] br[52] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_53 bl[53] br[53] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_54 bl[54] br[54] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_55 bl[55] br[55] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_56 bl[56] br[56] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_57 bl[57] br[57] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_58 bl[58] br[58] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_59 bl[59] br[59] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_60 bl[60] br[60] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_61 bl[61] br[61] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_62 bl[62] br[62] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_128_63 bl[63] br[63] vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xcell_129_0 bl[0] br[0] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_1 bl[1] br[1] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_2 bl[2] br[2] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_3 bl[3] br[3] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_4 bl[4] br[4] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_5 bl[5] br[5] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_6 bl[6] br[6] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_7 bl[7] br[7] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_8 bl[8] br[8] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_9 bl[9] br[9] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_10 bl[10] br[10] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_11 bl[11] br[11] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_12 bl[12] br[12] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_13 bl[13] br[13] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_14 bl[14] br[14] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_15 bl[15] br[15] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_16 bl[16] br[16] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_17 bl[17] br[17] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_18 bl[18] br[18] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_19 bl[19] br[19] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_20 bl[20] br[20] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_21 bl[21] br[21] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_22 bl[22] br[22] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_23 bl[23] br[23] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_24 bl[24] br[24] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_25 bl[25] br[25] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_26 bl[26] br[26] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_27 bl[27] br[27] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_28 bl[28] br[28] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_29 bl[29] br[29] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_30 bl[30] br[30] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_31 bl[31] br[31] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_32 bl[32] br[32] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_33 bl[33] br[33] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_34 bl[34] br[34] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_35 bl[35] br[35] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_36 bl[36] br[36] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_37 bl[37] br[37] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_38 bl[38] br[38] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_39 bl[39] br[39] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_40 bl[40] br[40] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_41 bl[41] br[41] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_42 bl[42] br[42] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_43 bl[43] br[43] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_44 bl[44] br[44] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_45 bl[45] br[45] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_46 bl[46] br[46] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_47 bl[47] br[47] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_48 bl[48] br[48] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_49 bl[49] br[49] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_50 bl[50] br[50] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_51 bl[51] br[51] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_52 bl[52] br[52] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_53 bl[53] br[53] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_54 bl[54] br[54] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_55 bl[55] br[55] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_56 bl[56] br[56] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_57 bl[57] br[57] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_58 bl[58] br[58] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_59 bl[59] br[59] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_60 bl[60] br[60] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_61 bl[61] br[61] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_62 bl[62] br[62] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_129_63 bl[63] br[63] vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xcell_130_0 bl[0] br[0] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_1 bl[1] br[1] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_2 bl[2] br[2] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_3 bl[3] br[3] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_4 bl[4] br[4] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_5 bl[5] br[5] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_6 bl[6] br[6] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_7 bl[7] br[7] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_8 bl[8] br[8] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_9 bl[9] br[9] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_10 bl[10] br[10] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_11 bl[11] br[11] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_12 bl[12] br[12] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_13 bl[13] br[13] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_14 bl[14] br[14] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_15 bl[15] br[15] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_16 bl[16] br[16] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_17 bl[17] br[17] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_18 bl[18] br[18] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_19 bl[19] br[19] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_20 bl[20] br[20] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_21 bl[21] br[21] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_22 bl[22] br[22] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_23 bl[23] br[23] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_24 bl[24] br[24] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_25 bl[25] br[25] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_26 bl[26] br[26] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_27 bl[27] br[27] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_28 bl[28] br[28] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_29 bl[29] br[29] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_30 bl[30] br[30] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_31 bl[31] br[31] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_32 bl[32] br[32] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_33 bl[33] br[33] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_34 bl[34] br[34] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_35 bl[35] br[35] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_36 bl[36] br[36] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_37 bl[37] br[37] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_38 bl[38] br[38] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_39 bl[39] br[39] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_40 bl[40] br[40] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_41 bl[41] br[41] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_42 bl[42] br[42] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_43 bl[43] br[43] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_44 bl[44] br[44] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_45 bl[45] br[45] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_46 bl[46] br[46] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_47 bl[47] br[47] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_48 bl[48] br[48] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_49 bl[49] br[49] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_50 bl[50] br[50] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_51 bl[51] br[51] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_52 bl[52] br[52] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_53 bl[53] br[53] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_54 bl[54] br[54] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_55 bl[55] br[55] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_56 bl[56] br[56] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_57 bl[57] br[57] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_58 bl[58] br[58] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_59 bl[59] br[59] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_60 bl[60] br[60] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_61 bl[61] br[61] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_62 bl[62] br[62] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_130_63 bl[63] br[63] vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xcell_131_0 bl[0] br[0] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_1 bl[1] br[1] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_2 bl[2] br[2] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_3 bl[3] br[3] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_4 bl[4] br[4] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_5 bl[5] br[5] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_6 bl[6] br[6] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_7 bl[7] br[7] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_8 bl[8] br[8] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_9 bl[9] br[9] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_10 bl[10] br[10] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_11 bl[11] br[11] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_12 bl[12] br[12] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_13 bl[13] br[13] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_14 bl[14] br[14] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_15 bl[15] br[15] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_16 bl[16] br[16] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_17 bl[17] br[17] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_18 bl[18] br[18] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_19 bl[19] br[19] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_20 bl[20] br[20] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_21 bl[21] br[21] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_22 bl[22] br[22] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_23 bl[23] br[23] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_24 bl[24] br[24] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_25 bl[25] br[25] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_26 bl[26] br[26] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_27 bl[27] br[27] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_28 bl[28] br[28] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_29 bl[29] br[29] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_30 bl[30] br[30] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_31 bl[31] br[31] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_32 bl[32] br[32] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_33 bl[33] br[33] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_34 bl[34] br[34] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_35 bl[35] br[35] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_36 bl[36] br[36] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_37 bl[37] br[37] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_38 bl[38] br[38] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_39 bl[39] br[39] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_40 bl[40] br[40] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_41 bl[41] br[41] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_42 bl[42] br[42] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_43 bl[43] br[43] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_44 bl[44] br[44] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_45 bl[45] br[45] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_46 bl[46] br[46] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_47 bl[47] br[47] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_48 bl[48] br[48] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_49 bl[49] br[49] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_50 bl[50] br[50] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_51 bl[51] br[51] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_52 bl[52] br[52] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_53 bl[53] br[53] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_54 bl[54] br[54] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_55 bl[55] br[55] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_56 bl[56] br[56] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_57 bl[57] br[57] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_58 bl[58] br[58] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_59 bl[59] br[59] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_60 bl[60] br[60] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_61 bl[61] br[61] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_62 bl[62] br[62] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_131_63 bl[63] br[63] vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xcell_132_0 bl[0] br[0] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_1 bl[1] br[1] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_2 bl[2] br[2] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_3 bl[3] br[3] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_4 bl[4] br[4] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_5 bl[5] br[5] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_6 bl[6] br[6] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_7 bl[7] br[7] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_8 bl[8] br[8] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_9 bl[9] br[9] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_10 bl[10] br[10] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_11 bl[11] br[11] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_12 bl[12] br[12] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_13 bl[13] br[13] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_14 bl[14] br[14] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_15 bl[15] br[15] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_16 bl[16] br[16] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_17 bl[17] br[17] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_18 bl[18] br[18] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_19 bl[19] br[19] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_20 bl[20] br[20] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_21 bl[21] br[21] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_22 bl[22] br[22] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_23 bl[23] br[23] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_24 bl[24] br[24] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_25 bl[25] br[25] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_26 bl[26] br[26] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_27 bl[27] br[27] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_28 bl[28] br[28] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_29 bl[29] br[29] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_30 bl[30] br[30] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_31 bl[31] br[31] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_32 bl[32] br[32] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_33 bl[33] br[33] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_34 bl[34] br[34] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_35 bl[35] br[35] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_36 bl[36] br[36] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_37 bl[37] br[37] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_38 bl[38] br[38] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_39 bl[39] br[39] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_40 bl[40] br[40] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_41 bl[41] br[41] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_42 bl[42] br[42] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_43 bl[43] br[43] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_44 bl[44] br[44] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_45 bl[45] br[45] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_46 bl[46] br[46] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_47 bl[47] br[47] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_48 bl[48] br[48] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_49 bl[49] br[49] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_50 bl[50] br[50] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_51 bl[51] br[51] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_52 bl[52] br[52] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_53 bl[53] br[53] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_54 bl[54] br[54] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_55 bl[55] br[55] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_56 bl[56] br[56] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_57 bl[57] br[57] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_58 bl[58] br[58] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_59 bl[59] br[59] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_60 bl[60] br[60] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_61 bl[61] br[61] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_62 bl[62] br[62] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_132_63 bl[63] br[63] vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xcell_133_0 bl[0] br[0] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_1 bl[1] br[1] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_2 bl[2] br[2] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_3 bl[3] br[3] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_4 bl[4] br[4] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_5 bl[5] br[5] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_6 bl[6] br[6] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_7 bl[7] br[7] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_8 bl[8] br[8] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_9 bl[9] br[9] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_10 bl[10] br[10] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_11 bl[11] br[11] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_12 bl[12] br[12] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_13 bl[13] br[13] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_14 bl[14] br[14] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_15 bl[15] br[15] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_16 bl[16] br[16] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_17 bl[17] br[17] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_18 bl[18] br[18] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_19 bl[19] br[19] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_20 bl[20] br[20] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_21 bl[21] br[21] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_22 bl[22] br[22] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_23 bl[23] br[23] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_24 bl[24] br[24] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_25 bl[25] br[25] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_26 bl[26] br[26] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_27 bl[27] br[27] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_28 bl[28] br[28] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_29 bl[29] br[29] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_30 bl[30] br[30] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_31 bl[31] br[31] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_32 bl[32] br[32] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_33 bl[33] br[33] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_34 bl[34] br[34] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_35 bl[35] br[35] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_36 bl[36] br[36] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_37 bl[37] br[37] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_38 bl[38] br[38] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_39 bl[39] br[39] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_40 bl[40] br[40] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_41 bl[41] br[41] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_42 bl[42] br[42] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_43 bl[43] br[43] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_44 bl[44] br[44] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_45 bl[45] br[45] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_46 bl[46] br[46] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_47 bl[47] br[47] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_48 bl[48] br[48] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_49 bl[49] br[49] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_50 bl[50] br[50] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_51 bl[51] br[51] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_52 bl[52] br[52] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_53 bl[53] br[53] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_54 bl[54] br[54] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_55 bl[55] br[55] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_56 bl[56] br[56] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_57 bl[57] br[57] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_58 bl[58] br[58] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_59 bl[59] br[59] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_60 bl[60] br[60] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_61 bl[61] br[61] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_62 bl[62] br[62] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_133_63 bl[63] br[63] vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xcell_134_0 bl[0] br[0] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_1 bl[1] br[1] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_2 bl[2] br[2] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_3 bl[3] br[3] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_4 bl[4] br[4] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_5 bl[5] br[5] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_6 bl[6] br[6] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_7 bl[7] br[7] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_8 bl[8] br[8] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_9 bl[9] br[9] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_10 bl[10] br[10] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_11 bl[11] br[11] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_12 bl[12] br[12] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_13 bl[13] br[13] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_14 bl[14] br[14] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_15 bl[15] br[15] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_16 bl[16] br[16] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_17 bl[17] br[17] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_18 bl[18] br[18] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_19 bl[19] br[19] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_20 bl[20] br[20] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_21 bl[21] br[21] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_22 bl[22] br[22] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_23 bl[23] br[23] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_24 bl[24] br[24] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_25 bl[25] br[25] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_26 bl[26] br[26] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_27 bl[27] br[27] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_28 bl[28] br[28] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_29 bl[29] br[29] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_30 bl[30] br[30] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_31 bl[31] br[31] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_32 bl[32] br[32] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_33 bl[33] br[33] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_34 bl[34] br[34] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_35 bl[35] br[35] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_36 bl[36] br[36] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_37 bl[37] br[37] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_38 bl[38] br[38] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_39 bl[39] br[39] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_40 bl[40] br[40] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_41 bl[41] br[41] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_42 bl[42] br[42] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_43 bl[43] br[43] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_44 bl[44] br[44] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_45 bl[45] br[45] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_46 bl[46] br[46] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_47 bl[47] br[47] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_48 bl[48] br[48] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_49 bl[49] br[49] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_50 bl[50] br[50] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_51 bl[51] br[51] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_52 bl[52] br[52] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_53 bl[53] br[53] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_54 bl[54] br[54] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_55 bl[55] br[55] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_56 bl[56] br[56] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_57 bl[57] br[57] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_58 bl[58] br[58] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_59 bl[59] br[59] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_60 bl[60] br[60] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_61 bl[61] br[61] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_62 bl[62] br[62] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_134_63 bl[63] br[63] vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xcell_135_0 bl[0] br[0] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_1 bl[1] br[1] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_2 bl[2] br[2] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_3 bl[3] br[3] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_4 bl[4] br[4] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_5 bl[5] br[5] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_6 bl[6] br[6] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_7 bl[7] br[7] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_8 bl[8] br[8] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_9 bl[9] br[9] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_10 bl[10] br[10] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_11 bl[11] br[11] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_12 bl[12] br[12] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_13 bl[13] br[13] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_14 bl[14] br[14] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_15 bl[15] br[15] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_16 bl[16] br[16] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_17 bl[17] br[17] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_18 bl[18] br[18] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_19 bl[19] br[19] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_20 bl[20] br[20] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_21 bl[21] br[21] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_22 bl[22] br[22] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_23 bl[23] br[23] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_24 bl[24] br[24] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_25 bl[25] br[25] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_26 bl[26] br[26] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_27 bl[27] br[27] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_28 bl[28] br[28] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_29 bl[29] br[29] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_30 bl[30] br[30] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_31 bl[31] br[31] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_32 bl[32] br[32] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_33 bl[33] br[33] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_34 bl[34] br[34] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_35 bl[35] br[35] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_36 bl[36] br[36] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_37 bl[37] br[37] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_38 bl[38] br[38] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_39 bl[39] br[39] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_40 bl[40] br[40] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_41 bl[41] br[41] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_42 bl[42] br[42] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_43 bl[43] br[43] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_44 bl[44] br[44] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_45 bl[45] br[45] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_46 bl[46] br[46] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_47 bl[47] br[47] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_48 bl[48] br[48] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_49 bl[49] br[49] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_50 bl[50] br[50] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_51 bl[51] br[51] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_52 bl[52] br[52] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_53 bl[53] br[53] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_54 bl[54] br[54] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_55 bl[55] br[55] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_56 bl[56] br[56] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_57 bl[57] br[57] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_58 bl[58] br[58] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_59 bl[59] br[59] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_60 bl[60] br[60] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_61 bl[61] br[61] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_62 bl[62] br[62] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_135_63 bl[63] br[63] vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xcell_136_0 bl[0] br[0] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_1 bl[1] br[1] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_2 bl[2] br[2] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_3 bl[3] br[3] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_4 bl[4] br[4] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_5 bl[5] br[5] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_6 bl[6] br[6] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_7 bl[7] br[7] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_8 bl[8] br[8] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_9 bl[9] br[9] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_10 bl[10] br[10] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_11 bl[11] br[11] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_12 bl[12] br[12] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_13 bl[13] br[13] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_14 bl[14] br[14] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_15 bl[15] br[15] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_16 bl[16] br[16] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_17 bl[17] br[17] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_18 bl[18] br[18] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_19 bl[19] br[19] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_20 bl[20] br[20] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_21 bl[21] br[21] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_22 bl[22] br[22] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_23 bl[23] br[23] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_24 bl[24] br[24] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_25 bl[25] br[25] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_26 bl[26] br[26] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_27 bl[27] br[27] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_28 bl[28] br[28] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_29 bl[29] br[29] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_30 bl[30] br[30] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_31 bl[31] br[31] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_32 bl[32] br[32] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_33 bl[33] br[33] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_34 bl[34] br[34] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_35 bl[35] br[35] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_36 bl[36] br[36] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_37 bl[37] br[37] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_38 bl[38] br[38] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_39 bl[39] br[39] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_40 bl[40] br[40] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_41 bl[41] br[41] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_42 bl[42] br[42] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_43 bl[43] br[43] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_44 bl[44] br[44] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_45 bl[45] br[45] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_46 bl[46] br[46] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_47 bl[47] br[47] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_48 bl[48] br[48] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_49 bl[49] br[49] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_50 bl[50] br[50] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_51 bl[51] br[51] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_52 bl[52] br[52] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_53 bl[53] br[53] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_54 bl[54] br[54] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_55 bl[55] br[55] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_56 bl[56] br[56] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_57 bl[57] br[57] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_58 bl[58] br[58] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_59 bl[59] br[59] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_60 bl[60] br[60] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_61 bl[61] br[61] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_62 bl[62] br[62] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_136_63 bl[63] br[63] vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xcell_137_0 bl[0] br[0] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_1 bl[1] br[1] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_2 bl[2] br[2] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_3 bl[3] br[3] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_4 bl[4] br[4] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_5 bl[5] br[5] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_6 bl[6] br[6] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_7 bl[7] br[7] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_8 bl[8] br[8] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_9 bl[9] br[9] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_10 bl[10] br[10] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_11 bl[11] br[11] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_12 bl[12] br[12] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_13 bl[13] br[13] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_14 bl[14] br[14] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_15 bl[15] br[15] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_16 bl[16] br[16] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_17 bl[17] br[17] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_18 bl[18] br[18] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_19 bl[19] br[19] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_20 bl[20] br[20] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_21 bl[21] br[21] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_22 bl[22] br[22] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_23 bl[23] br[23] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_24 bl[24] br[24] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_25 bl[25] br[25] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_26 bl[26] br[26] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_27 bl[27] br[27] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_28 bl[28] br[28] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_29 bl[29] br[29] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_30 bl[30] br[30] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_31 bl[31] br[31] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_32 bl[32] br[32] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_33 bl[33] br[33] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_34 bl[34] br[34] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_35 bl[35] br[35] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_36 bl[36] br[36] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_37 bl[37] br[37] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_38 bl[38] br[38] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_39 bl[39] br[39] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_40 bl[40] br[40] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_41 bl[41] br[41] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_42 bl[42] br[42] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_43 bl[43] br[43] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_44 bl[44] br[44] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_45 bl[45] br[45] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_46 bl[46] br[46] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_47 bl[47] br[47] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_48 bl[48] br[48] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_49 bl[49] br[49] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_50 bl[50] br[50] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_51 bl[51] br[51] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_52 bl[52] br[52] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_53 bl[53] br[53] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_54 bl[54] br[54] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_55 bl[55] br[55] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_56 bl[56] br[56] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_57 bl[57] br[57] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_58 bl[58] br[58] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_59 bl[59] br[59] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_60 bl[60] br[60] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_61 bl[61] br[61] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_62 bl[62] br[62] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_137_63 bl[63] br[63] vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xcell_138_0 bl[0] br[0] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_1 bl[1] br[1] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_2 bl[2] br[2] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_3 bl[3] br[3] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_4 bl[4] br[4] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_5 bl[5] br[5] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_6 bl[6] br[6] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_7 bl[7] br[7] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_8 bl[8] br[8] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_9 bl[9] br[9] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_10 bl[10] br[10] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_11 bl[11] br[11] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_12 bl[12] br[12] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_13 bl[13] br[13] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_14 bl[14] br[14] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_15 bl[15] br[15] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_16 bl[16] br[16] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_17 bl[17] br[17] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_18 bl[18] br[18] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_19 bl[19] br[19] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_20 bl[20] br[20] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_21 bl[21] br[21] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_22 bl[22] br[22] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_23 bl[23] br[23] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_24 bl[24] br[24] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_25 bl[25] br[25] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_26 bl[26] br[26] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_27 bl[27] br[27] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_28 bl[28] br[28] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_29 bl[29] br[29] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_30 bl[30] br[30] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_31 bl[31] br[31] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_32 bl[32] br[32] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_33 bl[33] br[33] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_34 bl[34] br[34] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_35 bl[35] br[35] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_36 bl[36] br[36] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_37 bl[37] br[37] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_38 bl[38] br[38] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_39 bl[39] br[39] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_40 bl[40] br[40] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_41 bl[41] br[41] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_42 bl[42] br[42] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_43 bl[43] br[43] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_44 bl[44] br[44] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_45 bl[45] br[45] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_46 bl[46] br[46] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_47 bl[47] br[47] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_48 bl[48] br[48] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_49 bl[49] br[49] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_50 bl[50] br[50] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_51 bl[51] br[51] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_52 bl[52] br[52] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_53 bl[53] br[53] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_54 bl[54] br[54] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_55 bl[55] br[55] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_56 bl[56] br[56] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_57 bl[57] br[57] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_58 bl[58] br[58] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_59 bl[59] br[59] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_60 bl[60] br[60] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_61 bl[61] br[61] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_62 bl[62] br[62] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_138_63 bl[63] br[63] vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xcell_139_0 bl[0] br[0] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_1 bl[1] br[1] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_2 bl[2] br[2] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_3 bl[3] br[3] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_4 bl[4] br[4] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_5 bl[5] br[5] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_6 bl[6] br[6] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_7 bl[7] br[7] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_8 bl[8] br[8] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_9 bl[9] br[9] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_10 bl[10] br[10] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_11 bl[11] br[11] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_12 bl[12] br[12] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_13 bl[13] br[13] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_14 bl[14] br[14] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_15 bl[15] br[15] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_16 bl[16] br[16] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_17 bl[17] br[17] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_18 bl[18] br[18] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_19 bl[19] br[19] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_20 bl[20] br[20] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_21 bl[21] br[21] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_22 bl[22] br[22] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_23 bl[23] br[23] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_24 bl[24] br[24] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_25 bl[25] br[25] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_26 bl[26] br[26] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_27 bl[27] br[27] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_28 bl[28] br[28] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_29 bl[29] br[29] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_30 bl[30] br[30] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_31 bl[31] br[31] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_32 bl[32] br[32] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_33 bl[33] br[33] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_34 bl[34] br[34] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_35 bl[35] br[35] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_36 bl[36] br[36] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_37 bl[37] br[37] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_38 bl[38] br[38] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_39 bl[39] br[39] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_40 bl[40] br[40] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_41 bl[41] br[41] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_42 bl[42] br[42] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_43 bl[43] br[43] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_44 bl[44] br[44] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_45 bl[45] br[45] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_46 bl[46] br[46] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_47 bl[47] br[47] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_48 bl[48] br[48] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_49 bl[49] br[49] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_50 bl[50] br[50] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_51 bl[51] br[51] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_52 bl[52] br[52] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_53 bl[53] br[53] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_54 bl[54] br[54] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_55 bl[55] br[55] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_56 bl[56] br[56] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_57 bl[57] br[57] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_58 bl[58] br[58] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_59 bl[59] br[59] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_60 bl[60] br[60] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_61 bl[61] br[61] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_62 bl[62] br[62] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_139_63 bl[63] br[63] vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xcell_140_0 bl[0] br[0] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_1 bl[1] br[1] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_2 bl[2] br[2] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_3 bl[3] br[3] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_4 bl[4] br[4] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_5 bl[5] br[5] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_6 bl[6] br[6] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_7 bl[7] br[7] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_8 bl[8] br[8] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_9 bl[9] br[9] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_10 bl[10] br[10] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_11 bl[11] br[11] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_12 bl[12] br[12] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_13 bl[13] br[13] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_14 bl[14] br[14] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_15 bl[15] br[15] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_16 bl[16] br[16] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_17 bl[17] br[17] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_18 bl[18] br[18] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_19 bl[19] br[19] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_20 bl[20] br[20] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_21 bl[21] br[21] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_22 bl[22] br[22] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_23 bl[23] br[23] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_24 bl[24] br[24] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_25 bl[25] br[25] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_26 bl[26] br[26] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_27 bl[27] br[27] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_28 bl[28] br[28] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_29 bl[29] br[29] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_30 bl[30] br[30] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_31 bl[31] br[31] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_32 bl[32] br[32] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_33 bl[33] br[33] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_34 bl[34] br[34] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_35 bl[35] br[35] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_36 bl[36] br[36] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_37 bl[37] br[37] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_38 bl[38] br[38] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_39 bl[39] br[39] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_40 bl[40] br[40] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_41 bl[41] br[41] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_42 bl[42] br[42] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_43 bl[43] br[43] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_44 bl[44] br[44] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_45 bl[45] br[45] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_46 bl[46] br[46] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_47 bl[47] br[47] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_48 bl[48] br[48] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_49 bl[49] br[49] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_50 bl[50] br[50] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_51 bl[51] br[51] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_52 bl[52] br[52] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_53 bl[53] br[53] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_54 bl[54] br[54] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_55 bl[55] br[55] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_56 bl[56] br[56] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_57 bl[57] br[57] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_58 bl[58] br[58] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_59 bl[59] br[59] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_60 bl[60] br[60] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_61 bl[61] br[61] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_62 bl[62] br[62] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_140_63 bl[63] br[63] vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xcell_141_0 bl[0] br[0] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_1 bl[1] br[1] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_2 bl[2] br[2] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_3 bl[3] br[3] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_4 bl[4] br[4] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_5 bl[5] br[5] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_6 bl[6] br[6] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_7 bl[7] br[7] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_8 bl[8] br[8] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_9 bl[9] br[9] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_10 bl[10] br[10] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_11 bl[11] br[11] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_12 bl[12] br[12] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_13 bl[13] br[13] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_14 bl[14] br[14] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_15 bl[15] br[15] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_16 bl[16] br[16] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_17 bl[17] br[17] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_18 bl[18] br[18] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_19 bl[19] br[19] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_20 bl[20] br[20] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_21 bl[21] br[21] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_22 bl[22] br[22] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_23 bl[23] br[23] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_24 bl[24] br[24] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_25 bl[25] br[25] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_26 bl[26] br[26] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_27 bl[27] br[27] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_28 bl[28] br[28] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_29 bl[29] br[29] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_30 bl[30] br[30] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_31 bl[31] br[31] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_32 bl[32] br[32] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_33 bl[33] br[33] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_34 bl[34] br[34] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_35 bl[35] br[35] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_36 bl[36] br[36] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_37 bl[37] br[37] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_38 bl[38] br[38] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_39 bl[39] br[39] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_40 bl[40] br[40] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_41 bl[41] br[41] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_42 bl[42] br[42] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_43 bl[43] br[43] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_44 bl[44] br[44] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_45 bl[45] br[45] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_46 bl[46] br[46] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_47 bl[47] br[47] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_48 bl[48] br[48] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_49 bl[49] br[49] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_50 bl[50] br[50] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_51 bl[51] br[51] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_52 bl[52] br[52] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_53 bl[53] br[53] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_54 bl[54] br[54] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_55 bl[55] br[55] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_56 bl[56] br[56] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_57 bl[57] br[57] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_58 bl[58] br[58] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_59 bl[59] br[59] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_60 bl[60] br[60] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_61 bl[61] br[61] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_62 bl[62] br[62] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_141_63 bl[63] br[63] vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xcell_142_0 bl[0] br[0] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_1 bl[1] br[1] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_2 bl[2] br[2] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_3 bl[3] br[3] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_4 bl[4] br[4] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_5 bl[5] br[5] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_6 bl[6] br[6] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_7 bl[7] br[7] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_8 bl[8] br[8] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_9 bl[9] br[9] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_10 bl[10] br[10] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_11 bl[11] br[11] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_12 bl[12] br[12] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_13 bl[13] br[13] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_14 bl[14] br[14] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_15 bl[15] br[15] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_16 bl[16] br[16] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_17 bl[17] br[17] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_18 bl[18] br[18] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_19 bl[19] br[19] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_20 bl[20] br[20] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_21 bl[21] br[21] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_22 bl[22] br[22] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_23 bl[23] br[23] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_24 bl[24] br[24] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_25 bl[25] br[25] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_26 bl[26] br[26] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_27 bl[27] br[27] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_28 bl[28] br[28] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_29 bl[29] br[29] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_30 bl[30] br[30] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_31 bl[31] br[31] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_32 bl[32] br[32] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_33 bl[33] br[33] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_34 bl[34] br[34] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_35 bl[35] br[35] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_36 bl[36] br[36] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_37 bl[37] br[37] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_38 bl[38] br[38] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_39 bl[39] br[39] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_40 bl[40] br[40] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_41 bl[41] br[41] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_42 bl[42] br[42] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_43 bl[43] br[43] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_44 bl[44] br[44] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_45 bl[45] br[45] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_46 bl[46] br[46] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_47 bl[47] br[47] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_48 bl[48] br[48] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_49 bl[49] br[49] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_50 bl[50] br[50] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_51 bl[51] br[51] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_52 bl[52] br[52] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_53 bl[53] br[53] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_54 bl[54] br[54] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_55 bl[55] br[55] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_56 bl[56] br[56] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_57 bl[57] br[57] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_58 bl[58] br[58] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_59 bl[59] br[59] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_60 bl[60] br[60] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_61 bl[61] br[61] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_62 bl[62] br[62] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_142_63 bl[63] br[63] vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xcell_143_0 bl[0] br[0] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_1 bl[1] br[1] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_2 bl[2] br[2] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_3 bl[3] br[3] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_4 bl[4] br[4] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_5 bl[5] br[5] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_6 bl[6] br[6] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_7 bl[7] br[7] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_8 bl[8] br[8] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_9 bl[9] br[9] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_10 bl[10] br[10] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_11 bl[11] br[11] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_12 bl[12] br[12] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_13 bl[13] br[13] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_14 bl[14] br[14] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_15 bl[15] br[15] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_16 bl[16] br[16] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_17 bl[17] br[17] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_18 bl[18] br[18] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_19 bl[19] br[19] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_20 bl[20] br[20] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_21 bl[21] br[21] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_22 bl[22] br[22] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_23 bl[23] br[23] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_24 bl[24] br[24] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_25 bl[25] br[25] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_26 bl[26] br[26] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_27 bl[27] br[27] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_28 bl[28] br[28] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_29 bl[29] br[29] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_30 bl[30] br[30] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_31 bl[31] br[31] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_32 bl[32] br[32] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_33 bl[33] br[33] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_34 bl[34] br[34] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_35 bl[35] br[35] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_36 bl[36] br[36] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_37 bl[37] br[37] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_38 bl[38] br[38] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_39 bl[39] br[39] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_40 bl[40] br[40] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_41 bl[41] br[41] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_42 bl[42] br[42] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_43 bl[43] br[43] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_44 bl[44] br[44] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_45 bl[45] br[45] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_46 bl[46] br[46] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_47 bl[47] br[47] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_48 bl[48] br[48] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_49 bl[49] br[49] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_50 bl[50] br[50] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_51 bl[51] br[51] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_52 bl[52] br[52] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_53 bl[53] br[53] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_54 bl[54] br[54] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_55 bl[55] br[55] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_56 bl[56] br[56] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_57 bl[57] br[57] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_58 bl[58] br[58] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_59 bl[59] br[59] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_60 bl[60] br[60] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_61 bl[61] br[61] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_62 bl[62] br[62] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_143_63 bl[63] br[63] vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xcell_144_0 bl[0] br[0] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_1 bl[1] br[1] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_2 bl[2] br[2] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_3 bl[3] br[3] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_4 bl[4] br[4] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_5 bl[5] br[5] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_6 bl[6] br[6] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_7 bl[7] br[7] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_8 bl[8] br[8] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_9 bl[9] br[9] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_10 bl[10] br[10] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_11 bl[11] br[11] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_12 bl[12] br[12] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_13 bl[13] br[13] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_14 bl[14] br[14] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_15 bl[15] br[15] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_16 bl[16] br[16] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_17 bl[17] br[17] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_18 bl[18] br[18] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_19 bl[19] br[19] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_20 bl[20] br[20] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_21 bl[21] br[21] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_22 bl[22] br[22] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_23 bl[23] br[23] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_24 bl[24] br[24] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_25 bl[25] br[25] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_26 bl[26] br[26] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_27 bl[27] br[27] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_28 bl[28] br[28] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_29 bl[29] br[29] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_30 bl[30] br[30] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_31 bl[31] br[31] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_32 bl[32] br[32] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_33 bl[33] br[33] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_34 bl[34] br[34] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_35 bl[35] br[35] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_36 bl[36] br[36] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_37 bl[37] br[37] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_38 bl[38] br[38] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_39 bl[39] br[39] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_40 bl[40] br[40] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_41 bl[41] br[41] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_42 bl[42] br[42] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_43 bl[43] br[43] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_44 bl[44] br[44] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_45 bl[45] br[45] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_46 bl[46] br[46] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_47 bl[47] br[47] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_48 bl[48] br[48] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_49 bl[49] br[49] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_50 bl[50] br[50] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_51 bl[51] br[51] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_52 bl[52] br[52] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_53 bl[53] br[53] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_54 bl[54] br[54] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_55 bl[55] br[55] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_56 bl[56] br[56] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_57 bl[57] br[57] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_58 bl[58] br[58] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_59 bl[59] br[59] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_60 bl[60] br[60] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_61 bl[61] br[61] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_62 bl[62] br[62] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_144_63 bl[63] br[63] vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xcell_145_0 bl[0] br[0] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_1 bl[1] br[1] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_2 bl[2] br[2] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_3 bl[3] br[3] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_4 bl[4] br[4] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_5 bl[5] br[5] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_6 bl[6] br[6] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_7 bl[7] br[7] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_8 bl[8] br[8] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_9 bl[9] br[9] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_10 bl[10] br[10] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_11 bl[11] br[11] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_12 bl[12] br[12] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_13 bl[13] br[13] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_14 bl[14] br[14] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_15 bl[15] br[15] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_16 bl[16] br[16] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_17 bl[17] br[17] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_18 bl[18] br[18] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_19 bl[19] br[19] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_20 bl[20] br[20] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_21 bl[21] br[21] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_22 bl[22] br[22] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_23 bl[23] br[23] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_24 bl[24] br[24] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_25 bl[25] br[25] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_26 bl[26] br[26] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_27 bl[27] br[27] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_28 bl[28] br[28] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_29 bl[29] br[29] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_30 bl[30] br[30] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_31 bl[31] br[31] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_32 bl[32] br[32] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_33 bl[33] br[33] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_34 bl[34] br[34] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_35 bl[35] br[35] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_36 bl[36] br[36] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_37 bl[37] br[37] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_38 bl[38] br[38] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_39 bl[39] br[39] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_40 bl[40] br[40] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_41 bl[41] br[41] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_42 bl[42] br[42] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_43 bl[43] br[43] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_44 bl[44] br[44] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_45 bl[45] br[45] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_46 bl[46] br[46] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_47 bl[47] br[47] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_48 bl[48] br[48] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_49 bl[49] br[49] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_50 bl[50] br[50] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_51 bl[51] br[51] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_52 bl[52] br[52] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_53 bl[53] br[53] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_54 bl[54] br[54] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_55 bl[55] br[55] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_56 bl[56] br[56] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_57 bl[57] br[57] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_58 bl[58] br[58] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_59 bl[59] br[59] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_60 bl[60] br[60] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_61 bl[61] br[61] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_62 bl[62] br[62] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_145_63 bl[63] br[63] vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xcell_146_0 bl[0] br[0] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_1 bl[1] br[1] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_2 bl[2] br[2] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_3 bl[3] br[3] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_4 bl[4] br[4] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_5 bl[5] br[5] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_6 bl[6] br[6] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_7 bl[7] br[7] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_8 bl[8] br[8] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_9 bl[9] br[9] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_10 bl[10] br[10] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_11 bl[11] br[11] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_12 bl[12] br[12] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_13 bl[13] br[13] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_14 bl[14] br[14] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_15 bl[15] br[15] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_16 bl[16] br[16] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_17 bl[17] br[17] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_18 bl[18] br[18] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_19 bl[19] br[19] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_20 bl[20] br[20] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_21 bl[21] br[21] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_22 bl[22] br[22] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_23 bl[23] br[23] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_24 bl[24] br[24] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_25 bl[25] br[25] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_26 bl[26] br[26] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_27 bl[27] br[27] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_28 bl[28] br[28] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_29 bl[29] br[29] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_30 bl[30] br[30] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_31 bl[31] br[31] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_32 bl[32] br[32] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_33 bl[33] br[33] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_34 bl[34] br[34] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_35 bl[35] br[35] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_36 bl[36] br[36] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_37 bl[37] br[37] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_38 bl[38] br[38] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_39 bl[39] br[39] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_40 bl[40] br[40] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_41 bl[41] br[41] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_42 bl[42] br[42] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_43 bl[43] br[43] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_44 bl[44] br[44] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_45 bl[45] br[45] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_46 bl[46] br[46] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_47 bl[47] br[47] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_48 bl[48] br[48] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_49 bl[49] br[49] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_50 bl[50] br[50] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_51 bl[51] br[51] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_52 bl[52] br[52] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_53 bl[53] br[53] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_54 bl[54] br[54] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_55 bl[55] br[55] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_56 bl[56] br[56] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_57 bl[57] br[57] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_58 bl[58] br[58] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_59 bl[59] br[59] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_60 bl[60] br[60] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_61 bl[61] br[61] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_62 bl[62] br[62] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_146_63 bl[63] br[63] vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xcell_147_0 bl[0] br[0] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_1 bl[1] br[1] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_2 bl[2] br[2] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_3 bl[3] br[3] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_4 bl[4] br[4] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_5 bl[5] br[5] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_6 bl[6] br[6] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_7 bl[7] br[7] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_8 bl[8] br[8] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_9 bl[9] br[9] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_10 bl[10] br[10] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_11 bl[11] br[11] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_12 bl[12] br[12] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_13 bl[13] br[13] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_14 bl[14] br[14] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_15 bl[15] br[15] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_16 bl[16] br[16] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_17 bl[17] br[17] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_18 bl[18] br[18] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_19 bl[19] br[19] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_20 bl[20] br[20] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_21 bl[21] br[21] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_22 bl[22] br[22] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_23 bl[23] br[23] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_24 bl[24] br[24] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_25 bl[25] br[25] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_26 bl[26] br[26] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_27 bl[27] br[27] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_28 bl[28] br[28] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_29 bl[29] br[29] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_30 bl[30] br[30] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_31 bl[31] br[31] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_32 bl[32] br[32] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_33 bl[33] br[33] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_34 bl[34] br[34] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_35 bl[35] br[35] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_36 bl[36] br[36] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_37 bl[37] br[37] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_38 bl[38] br[38] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_39 bl[39] br[39] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_40 bl[40] br[40] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_41 bl[41] br[41] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_42 bl[42] br[42] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_43 bl[43] br[43] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_44 bl[44] br[44] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_45 bl[45] br[45] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_46 bl[46] br[46] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_47 bl[47] br[47] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_48 bl[48] br[48] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_49 bl[49] br[49] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_50 bl[50] br[50] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_51 bl[51] br[51] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_52 bl[52] br[52] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_53 bl[53] br[53] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_54 bl[54] br[54] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_55 bl[55] br[55] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_56 bl[56] br[56] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_57 bl[57] br[57] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_58 bl[58] br[58] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_59 bl[59] br[59] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_60 bl[60] br[60] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_61 bl[61] br[61] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_62 bl[62] br[62] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_147_63 bl[63] br[63] vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xcell_148_0 bl[0] br[0] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_1 bl[1] br[1] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_2 bl[2] br[2] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_3 bl[3] br[3] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_4 bl[4] br[4] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_5 bl[5] br[5] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_6 bl[6] br[6] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_7 bl[7] br[7] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_8 bl[8] br[8] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_9 bl[9] br[9] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_10 bl[10] br[10] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_11 bl[11] br[11] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_12 bl[12] br[12] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_13 bl[13] br[13] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_14 bl[14] br[14] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_15 bl[15] br[15] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_16 bl[16] br[16] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_17 bl[17] br[17] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_18 bl[18] br[18] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_19 bl[19] br[19] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_20 bl[20] br[20] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_21 bl[21] br[21] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_22 bl[22] br[22] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_23 bl[23] br[23] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_24 bl[24] br[24] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_25 bl[25] br[25] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_26 bl[26] br[26] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_27 bl[27] br[27] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_28 bl[28] br[28] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_29 bl[29] br[29] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_30 bl[30] br[30] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_31 bl[31] br[31] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_32 bl[32] br[32] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_33 bl[33] br[33] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_34 bl[34] br[34] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_35 bl[35] br[35] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_36 bl[36] br[36] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_37 bl[37] br[37] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_38 bl[38] br[38] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_39 bl[39] br[39] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_40 bl[40] br[40] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_41 bl[41] br[41] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_42 bl[42] br[42] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_43 bl[43] br[43] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_44 bl[44] br[44] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_45 bl[45] br[45] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_46 bl[46] br[46] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_47 bl[47] br[47] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_48 bl[48] br[48] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_49 bl[49] br[49] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_50 bl[50] br[50] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_51 bl[51] br[51] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_52 bl[52] br[52] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_53 bl[53] br[53] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_54 bl[54] br[54] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_55 bl[55] br[55] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_56 bl[56] br[56] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_57 bl[57] br[57] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_58 bl[58] br[58] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_59 bl[59] br[59] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_60 bl[60] br[60] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_61 bl[61] br[61] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_62 bl[62] br[62] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_148_63 bl[63] br[63] vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xcell_149_0 bl[0] br[0] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_1 bl[1] br[1] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_2 bl[2] br[2] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_3 bl[3] br[3] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_4 bl[4] br[4] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_5 bl[5] br[5] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_6 bl[6] br[6] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_7 bl[7] br[7] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_8 bl[8] br[8] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_9 bl[9] br[9] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_10 bl[10] br[10] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_11 bl[11] br[11] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_12 bl[12] br[12] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_13 bl[13] br[13] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_14 bl[14] br[14] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_15 bl[15] br[15] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_16 bl[16] br[16] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_17 bl[17] br[17] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_18 bl[18] br[18] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_19 bl[19] br[19] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_20 bl[20] br[20] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_21 bl[21] br[21] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_22 bl[22] br[22] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_23 bl[23] br[23] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_24 bl[24] br[24] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_25 bl[25] br[25] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_26 bl[26] br[26] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_27 bl[27] br[27] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_28 bl[28] br[28] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_29 bl[29] br[29] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_30 bl[30] br[30] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_31 bl[31] br[31] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_32 bl[32] br[32] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_33 bl[33] br[33] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_34 bl[34] br[34] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_35 bl[35] br[35] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_36 bl[36] br[36] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_37 bl[37] br[37] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_38 bl[38] br[38] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_39 bl[39] br[39] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_40 bl[40] br[40] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_41 bl[41] br[41] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_42 bl[42] br[42] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_43 bl[43] br[43] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_44 bl[44] br[44] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_45 bl[45] br[45] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_46 bl[46] br[46] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_47 bl[47] br[47] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_48 bl[48] br[48] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_49 bl[49] br[49] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_50 bl[50] br[50] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_51 bl[51] br[51] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_52 bl[52] br[52] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_53 bl[53] br[53] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_54 bl[54] br[54] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_55 bl[55] br[55] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_56 bl[56] br[56] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_57 bl[57] br[57] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_58 bl[58] br[58] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_59 bl[59] br[59] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_60 bl[60] br[60] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_61 bl[61] br[61] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_62 bl[62] br[62] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_149_63 bl[63] br[63] vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xcell_150_0 bl[0] br[0] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_1 bl[1] br[1] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_2 bl[2] br[2] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_3 bl[3] br[3] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_4 bl[4] br[4] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_5 bl[5] br[5] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_6 bl[6] br[6] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_7 bl[7] br[7] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_8 bl[8] br[8] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_9 bl[9] br[9] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_10 bl[10] br[10] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_11 bl[11] br[11] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_12 bl[12] br[12] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_13 bl[13] br[13] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_14 bl[14] br[14] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_15 bl[15] br[15] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_16 bl[16] br[16] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_17 bl[17] br[17] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_18 bl[18] br[18] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_19 bl[19] br[19] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_20 bl[20] br[20] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_21 bl[21] br[21] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_22 bl[22] br[22] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_23 bl[23] br[23] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_24 bl[24] br[24] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_25 bl[25] br[25] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_26 bl[26] br[26] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_27 bl[27] br[27] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_28 bl[28] br[28] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_29 bl[29] br[29] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_30 bl[30] br[30] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_31 bl[31] br[31] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_32 bl[32] br[32] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_33 bl[33] br[33] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_34 bl[34] br[34] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_35 bl[35] br[35] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_36 bl[36] br[36] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_37 bl[37] br[37] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_38 bl[38] br[38] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_39 bl[39] br[39] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_40 bl[40] br[40] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_41 bl[41] br[41] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_42 bl[42] br[42] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_43 bl[43] br[43] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_44 bl[44] br[44] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_45 bl[45] br[45] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_46 bl[46] br[46] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_47 bl[47] br[47] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_48 bl[48] br[48] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_49 bl[49] br[49] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_50 bl[50] br[50] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_51 bl[51] br[51] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_52 bl[52] br[52] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_53 bl[53] br[53] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_54 bl[54] br[54] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_55 bl[55] br[55] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_56 bl[56] br[56] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_57 bl[57] br[57] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_58 bl[58] br[58] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_59 bl[59] br[59] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_60 bl[60] br[60] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_61 bl[61] br[61] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_62 bl[62] br[62] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_150_63 bl[63] br[63] vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xcell_151_0 bl[0] br[0] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_1 bl[1] br[1] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_2 bl[2] br[2] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_3 bl[3] br[3] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_4 bl[4] br[4] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_5 bl[5] br[5] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_6 bl[6] br[6] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_7 bl[7] br[7] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_8 bl[8] br[8] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_9 bl[9] br[9] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_10 bl[10] br[10] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_11 bl[11] br[11] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_12 bl[12] br[12] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_13 bl[13] br[13] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_14 bl[14] br[14] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_15 bl[15] br[15] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_16 bl[16] br[16] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_17 bl[17] br[17] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_18 bl[18] br[18] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_19 bl[19] br[19] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_20 bl[20] br[20] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_21 bl[21] br[21] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_22 bl[22] br[22] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_23 bl[23] br[23] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_24 bl[24] br[24] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_25 bl[25] br[25] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_26 bl[26] br[26] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_27 bl[27] br[27] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_28 bl[28] br[28] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_29 bl[29] br[29] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_30 bl[30] br[30] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_31 bl[31] br[31] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_32 bl[32] br[32] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_33 bl[33] br[33] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_34 bl[34] br[34] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_35 bl[35] br[35] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_36 bl[36] br[36] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_37 bl[37] br[37] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_38 bl[38] br[38] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_39 bl[39] br[39] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_40 bl[40] br[40] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_41 bl[41] br[41] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_42 bl[42] br[42] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_43 bl[43] br[43] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_44 bl[44] br[44] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_45 bl[45] br[45] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_46 bl[46] br[46] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_47 bl[47] br[47] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_48 bl[48] br[48] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_49 bl[49] br[49] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_50 bl[50] br[50] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_51 bl[51] br[51] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_52 bl[52] br[52] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_53 bl[53] br[53] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_54 bl[54] br[54] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_55 bl[55] br[55] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_56 bl[56] br[56] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_57 bl[57] br[57] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_58 bl[58] br[58] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_59 bl[59] br[59] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_60 bl[60] br[60] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_61 bl[61] br[61] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_62 bl[62] br[62] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_151_63 bl[63] br[63] vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xcell_152_0 bl[0] br[0] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_1 bl[1] br[1] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_2 bl[2] br[2] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_3 bl[3] br[3] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_4 bl[4] br[4] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_5 bl[5] br[5] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_6 bl[6] br[6] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_7 bl[7] br[7] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_8 bl[8] br[8] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_9 bl[9] br[9] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_10 bl[10] br[10] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_11 bl[11] br[11] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_12 bl[12] br[12] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_13 bl[13] br[13] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_14 bl[14] br[14] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_15 bl[15] br[15] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_16 bl[16] br[16] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_17 bl[17] br[17] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_18 bl[18] br[18] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_19 bl[19] br[19] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_20 bl[20] br[20] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_21 bl[21] br[21] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_22 bl[22] br[22] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_23 bl[23] br[23] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_24 bl[24] br[24] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_25 bl[25] br[25] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_26 bl[26] br[26] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_27 bl[27] br[27] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_28 bl[28] br[28] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_29 bl[29] br[29] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_30 bl[30] br[30] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_31 bl[31] br[31] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_32 bl[32] br[32] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_33 bl[33] br[33] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_34 bl[34] br[34] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_35 bl[35] br[35] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_36 bl[36] br[36] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_37 bl[37] br[37] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_38 bl[38] br[38] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_39 bl[39] br[39] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_40 bl[40] br[40] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_41 bl[41] br[41] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_42 bl[42] br[42] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_43 bl[43] br[43] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_44 bl[44] br[44] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_45 bl[45] br[45] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_46 bl[46] br[46] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_47 bl[47] br[47] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_48 bl[48] br[48] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_49 bl[49] br[49] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_50 bl[50] br[50] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_51 bl[51] br[51] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_52 bl[52] br[52] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_53 bl[53] br[53] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_54 bl[54] br[54] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_55 bl[55] br[55] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_56 bl[56] br[56] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_57 bl[57] br[57] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_58 bl[58] br[58] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_59 bl[59] br[59] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_60 bl[60] br[60] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_61 bl[61] br[61] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_62 bl[62] br[62] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_152_63 bl[63] br[63] vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xcell_153_0 bl[0] br[0] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_1 bl[1] br[1] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_2 bl[2] br[2] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_3 bl[3] br[3] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_4 bl[4] br[4] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_5 bl[5] br[5] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_6 bl[6] br[6] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_7 bl[7] br[7] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_8 bl[8] br[8] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_9 bl[9] br[9] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_10 bl[10] br[10] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_11 bl[11] br[11] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_12 bl[12] br[12] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_13 bl[13] br[13] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_14 bl[14] br[14] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_15 bl[15] br[15] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_16 bl[16] br[16] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_17 bl[17] br[17] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_18 bl[18] br[18] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_19 bl[19] br[19] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_20 bl[20] br[20] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_21 bl[21] br[21] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_22 bl[22] br[22] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_23 bl[23] br[23] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_24 bl[24] br[24] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_25 bl[25] br[25] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_26 bl[26] br[26] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_27 bl[27] br[27] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_28 bl[28] br[28] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_29 bl[29] br[29] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_30 bl[30] br[30] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_31 bl[31] br[31] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_32 bl[32] br[32] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_33 bl[33] br[33] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_34 bl[34] br[34] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_35 bl[35] br[35] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_36 bl[36] br[36] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_37 bl[37] br[37] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_38 bl[38] br[38] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_39 bl[39] br[39] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_40 bl[40] br[40] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_41 bl[41] br[41] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_42 bl[42] br[42] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_43 bl[43] br[43] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_44 bl[44] br[44] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_45 bl[45] br[45] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_46 bl[46] br[46] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_47 bl[47] br[47] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_48 bl[48] br[48] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_49 bl[49] br[49] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_50 bl[50] br[50] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_51 bl[51] br[51] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_52 bl[52] br[52] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_53 bl[53] br[53] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_54 bl[54] br[54] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_55 bl[55] br[55] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_56 bl[56] br[56] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_57 bl[57] br[57] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_58 bl[58] br[58] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_59 bl[59] br[59] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_60 bl[60] br[60] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_61 bl[61] br[61] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_62 bl[62] br[62] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_153_63 bl[63] br[63] vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xcell_154_0 bl[0] br[0] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_1 bl[1] br[1] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_2 bl[2] br[2] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_3 bl[3] br[3] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_4 bl[4] br[4] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_5 bl[5] br[5] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_6 bl[6] br[6] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_7 bl[7] br[7] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_8 bl[8] br[8] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_9 bl[9] br[9] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_10 bl[10] br[10] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_11 bl[11] br[11] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_12 bl[12] br[12] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_13 bl[13] br[13] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_14 bl[14] br[14] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_15 bl[15] br[15] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_16 bl[16] br[16] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_17 bl[17] br[17] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_18 bl[18] br[18] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_19 bl[19] br[19] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_20 bl[20] br[20] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_21 bl[21] br[21] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_22 bl[22] br[22] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_23 bl[23] br[23] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_24 bl[24] br[24] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_25 bl[25] br[25] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_26 bl[26] br[26] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_27 bl[27] br[27] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_28 bl[28] br[28] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_29 bl[29] br[29] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_30 bl[30] br[30] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_31 bl[31] br[31] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_32 bl[32] br[32] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_33 bl[33] br[33] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_34 bl[34] br[34] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_35 bl[35] br[35] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_36 bl[36] br[36] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_37 bl[37] br[37] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_38 bl[38] br[38] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_39 bl[39] br[39] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_40 bl[40] br[40] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_41 bl[41] br[41] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_42 bl[42] br[42] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_43 bl[43] br[43] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_44 bl[44] br[44] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_45 bl[45] br[45] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_46 bl[46] br[46] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_47 bl[47] br[47] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_48 bl[48] br[48] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_49 bl[49] br[49] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_50 bl[50] br[50] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_51 bl[51] br[51] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_52 bl[52] br[52] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_53 bl[53] br[53] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_54 bl[54] br[54] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_55 bl[55] br[55] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_56 bl[56] br[56] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_57 bl[57] br[57] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_58 bl[58] br[58] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_59 bl[59] br[59] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_60 bl[60] br[60] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_61 bl[61] br[61] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_62 bl[62] br[62] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_154_63 bl[63] br[63] vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xcell_155_0 bl[0] br[0] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_1 bl[1] br[1] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_2 bl[2] br[2] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_3 bl[3] br[3] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_4 bl[4] br[4] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_5 bl[5] br[5] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_6 bl[6] br[6] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_7 bl[7] br[7] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_8 bl[8] br[8] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_9 bl[9] br[9] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_10 bl[10] br[10] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_11 bl[11] br[11] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_12 bl[12] br[12] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_13 bl[13] br[13] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_14 bl[14] br[14] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_15 bl[15] br[15] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_16 bl[16] br[16] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_17 bl[17] br[17] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_18 bl[18] br[18] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_19 bl[19] br[19] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_20 bl[20] br[20] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_21 bl[21] br[21] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_22 bl[22] br[22] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_23 bl[23] br[23] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_24 bl[24] br[24] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_25 bl[25] br[25] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_26 bl[26] br[26] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_27 bl[27] br[27] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_28 bl[28] br[28] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_29 bl[29] br[29] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_30 bl[30] br[30] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_31 bl[31] br[31] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_32 bl[32] br[32] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_33 bl[33] br[33] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_34 bl[34] br[34] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_35 bl[35] br[35] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_36 bl[36] br[36] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_37 bl[37] br[37] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_38 bl[38] br[38] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_39 bl[39] br[39] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_40 bl[40] br[40] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_41 bl[41] br[41] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_42 bl[42] br[42] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_43 bl[43] br[43] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_44 bl[44] br[44] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_45 bl[45] br[45] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_46 bl[46] br[46] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_47 bl[47] br[47] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_48 bl[48] br[48] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_49 bl[49] br[49] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_50 bl[50] br[50] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_51 bl[51] br[51] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_52 bl[52] br[52] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_53 bl[53] br[53] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_54 bl[54] br[54] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_55 bl[55] br[55] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_56 bl[56] br[56] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_57 bl[57] br[57] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_58 bl[58] br[58] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_59 bl[59] br[59] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_60 bl[60] br[60] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_61 bl[61] br[61] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_62 bl[62] br[62] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_155_63 bl[63] br[63] vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xcell_156_0 bl[0] br[0] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_1 bl[1] br[1] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_2 bl[2] br[2] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_3 bl[3] br[3] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_4 bl[4] br[4] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_5 bl[5] br[5] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_6 bl[6] br[6] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_7 bl[7] br[7] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_8 bl[8] br[8] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_9 bl[9] br[9] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_10 bl[10] br[10] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_11 bl[11] br[11] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_12 bl[12] br[12] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_13 bl[13] br[13] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_14 bl[14] br[14] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_15 bl[15] br[15] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_16 bl[16] br[16] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_17 bl[17] br[17] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_18 bl[18] br[18] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_19 bl[19] br[19] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_20 bl[20] br[20] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_21 bl[21] br[21] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_22 bl[22] br[22] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_23 bl[23] br[23] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_24 bl[24] br[24] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_25 bl[25] br[25] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_26 bl[26] br[26] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_27 bl[27] br[27] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_28 bl[28] br[28] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_29 bl[29] br[29] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_30 bl[30] br[30] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_31 bl[31] br[31] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_32 bl[32] br[32] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_33 bl[33] br[33] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_34 bl[34] br[34] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_35 bl[35] br[35] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_36 bl[36] br[36] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_37 bl[37] br[37] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_38 bl[38] br[38] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_39 bl[39] br[39] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_40 bl[40] br[40] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_41 bl[41] br[41] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_42 bl[42] br[42] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_43 bl[43] br[43] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_44 bl[44] br[44] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_45 bl[45] br[45] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_46 bl[46] br[46] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_47 bl[47] br[47] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_48 bl[48] br[48] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_49 bl[49] br[49] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_50 bl[50] br[50] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_51 bl[51] br[51] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_52 bl[52] br[52] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_53 bl[53] br[53] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_54 bl[54] br[54] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_55 bl[55] br[55] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_56 bl[56] br[56] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_57 bl[57] br[57] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_58 bl[58] br[58] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_59 bl[59] br[59] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_60 bl[60] br[60] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_61 bl[61] br[61] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_62 bl[62] br[62] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_156_63 bl[63] br[63] vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xcell_157_0 bl[0] br[0] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_1 bl[1] br[1] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_2 bl[2] br[2] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_3 bl[3] br[3] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_4 bl[4] br[4] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_5 bl[5] br[5] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_6 bl[6] br[6] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_7 bl[7] br[7] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_8 bl[8] br[8] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_9 bl[9] br[9] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_10 bl[10] br[10] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_11 bl[11] br[11] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_12 bl[12] br[12] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_13 bl[13] br[13] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_14 bl[14] br[14] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_15 bl[15] br[15] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_16 bl[16] br[16] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_17 bl[17] br[17] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_18 bl[18] br[18] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_19 bl[19] br[19] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_20 bl[20] br[20] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_21 bl[21] br[21] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_22 bl[22] br[22] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_23 bl[23] br[23] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_24 bl[24] br[24] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_25 bl[25] br[25] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_26 bl[26] br[26] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_27 bl[27] br[27] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_28 bl[28] br[28] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_29 bl[29] br[29] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_30 bl[30] br[30] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_31 bl[31] br[31] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_32 bl[32] br[32] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_33 bl[33] br[33] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_34 bl[34] br[34] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_35 bl[35] br[35] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_36 bl[36] br[36] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_37 bl[37] br[37] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_38 bl[38] br[38] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_39 bl[39] br[39] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_40 bl[40] br[40] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_41 bl[41] br[41] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_42 bl[42] br[42] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_43 bl[43] br[43] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_44 bl[44] br[44] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_45 bl[45] br[45] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_46 bl[46] br[46] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_47 bl[47] br[47] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_48 bl[48] br[48] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_49 bl[49] br[49] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_50 bl[50] br[50] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_51 bl[51] br[51] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_52 bl[52] br[52] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_53 bl[53] br[53] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_54 bl[54] br[54] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_55 bl[55] br[55] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_56 bl[56] br[56] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_57 bl[57] br[57] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_58 bl[58] br[58] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_59 bl[59] br[59] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_60 bl[60] br[60] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_61 bl[61] br[61] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_62 bl[62] br[62] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_157_63 bl[63] br[63] vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xcell_158_0 bl[0] br[0] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_1 bl[1] br[1] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_2 bl[2] br[2] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_3 bl[3] br[3] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_4 bl[4] br[4] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_5 bl[5] br[5] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_6 bl[6] br[6] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_7 bl[7] br[7] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_8 bl[8] br[8] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_9 bl[9] br[9] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_10 bl[10] br[10] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_11 bl[11] br[11] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_12 bl[12] br[12] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_13 bl[13] br[13] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_14 bl[14] br[14] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_15 bl[15] br[15] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_16 bl[16] br[16] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_17 bl[17] br[17] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_18 bl[18] br[18] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_19 bl[19] br[19] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_20 bl[20] br[20] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_21 bl[21] br[21] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_22 bl[22] br[22] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_23 bl[23] br[23] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_24 bl[24] br[24] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_25 bl[25] br[25] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_26 bl[26] br[26] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_27 bl[27] br[27] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_28 bl[28] br[28] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_29 bl[29] br[29] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_30 bl[30] br[30] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_31 bl[31] br[31] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_32 bl[32] br[32] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_33 bl[33] br[33] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_34 bl[34] br[34] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_35 bl[35] br[35] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_36 bl[36] br[36] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_37 bl[37] br[37] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_38 bl[38] br[38] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_39 bl[39] br[39] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_40 bl[40] br[40] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_41 bl[41] br[41] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_42 bl[42] br[42] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_43 bl[43] br[43] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_44 bl[44] br[44] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_45 bl[45] br[45] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_46 bl[46] br[46] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_47 bl[47] br[47] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_48 bl[48] br[48] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_49 bl[49] br[49] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_50 bl[50] br[50] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_51 bl[51] br[51] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_52 bl[52] br[52] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_53 bl[53] br[53] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_54 bl[54] br[54] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_55 bl[55] br[55] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_56 bl[56] br[56] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_57 bl[57] br[57] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_58 bl[58] br[58] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_59 bl[59] br[59] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_60 bl[60] br[60] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_61 bl[61] br[61] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_62 bl[62] br[62] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_158_63 bl[63] br[63] vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xcell_159_0 bl[0] br[0] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_1 bl[1] br[1] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_2 bl[2] br[2] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_3 bl[3] br[3] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_4 bl[4] br[4] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_5 bl[5] br[5] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_6 bl[6] br[6] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_7 bl[7] br[7] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_8 bl[8] br[8] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_9 bl[9] br[9] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_10 bl[10] br[10] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_11 bl[11] br[11] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_12 bl[12] br[12] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_13 bl[13] br[13] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_14 bl[14] br[14] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_15 bl[15] br[15] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_16 bl[16] br[16] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_17 bl[17] br[17] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_18 bl[18] br[18] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_19 bl[19] br[19] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_20 bl[20] br[20] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_21 bl[21] br[21] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_22 bl[22] br[22] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_23 bl[23] br[23] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_24 bl[24] br[24] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_25 bl[25] br[25] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_26 bl[26] br[26] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_27 bl[27] br[27] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_28 bl[28] br[28] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_29 bl[29] br[29] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_30 bl[30] br[30] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_31 bl[31] br[31] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_32 bl[32] br[32] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_33 bl[33] br[33] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_34 bl[34] br[34] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_35 bl[35] br[35] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_36 bl[36] br[36] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_37 bl[37] br[37] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_38 bl[38] br[38] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_39 bl[39] br[39] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_40 bl[40] br[40] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_41 bl[41] br[41] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_42 bl[42] br[42] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_43 bl[43] br[43] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_44 bl[44] br[44] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_45 bl[45] br[45] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_46 bl[46] br[46] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_47 bl[47] br[47] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_48 bl[48] br[48] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_49 bl[49] br[49] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_50 bl[50] br[50] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_51 bl[51] br[51] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_52 bl[52] br[52] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_53 bl[53] br[53] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_54 bl[54] br[54] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_55 bl[55] br[55] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_56 bl[56] br[56] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_57 bl[57] br[57] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_58 bl[58] br[58] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_59 bl[59] br[59] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_60 bl[60] br[60] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_61 bl[61] br[61] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_62 bl[62] br[62] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_159_63 bl[63] br[63] vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xcell_160_0 bl[0] br[0] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_1 bl[1] br[1] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_2 bl[2] br[2] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_3 bl[3] br[3] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_4 bl[4] br[4] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_5 bl[5] br[5] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_6 bl[6] br[6] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_7 bl[7] br[7] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_8 bl[8] br[8] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_9 bl[9] br[9] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_10 bl[10] br[10] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_11 bl[11] br[11] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_12 bl[12] br[12] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_13 bl[13] br[13] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_14 bl[14] br[14] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_15 bl[15] br[15] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_16 bl[16] br[16] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_17 bl[17] br[17] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_18 bl[18] br[18] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_19 bl[19] br[19] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_20 bl[20] br[20] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_21 bl[21] br[21] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_22 bl[22] br[22] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_23 bl[23] br[23] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_24 bl[24] br[24] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_25 bl[25] br[25] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_26 bl[26] br[26] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_27 bl[27] br[27] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_28 bl[28] br[28] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_29 bl[29] br[29] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_30 bl[30] br[30] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_31 bl[31] br[31] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_32 bl[32] br[32] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_33 bl[33] br[33] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_34 bl[34] br[34] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_35 bl[35] br[35] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_36 bl[36] br[36] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_37 bl[37] br[37] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_38 bl[38] br[38] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_39 bl[39] br[39] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_40 bl[40] br[40] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_41 bl[41] br[41] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_42 bl[42] br[42] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_43 bl[43] br[43] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_44 bl[44] br[44] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_45 bl[45] br[45] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_46 bl[46] br[46] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_47 bl[47] br[47] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_48 bl[48] br[48] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_49 bl[49] br[49] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_50 bl[50] br[50] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_51 bl[51] br[51] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_52 bl[52] br[52] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_53 bl[53] br[53] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_54 bl[54] br[54] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_55 bl[55] br[55] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_56 bl[56] br[56] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_57 bl[57] br[57] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_58 bl[58] br[58] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_59 bl[59] br[59] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_60 bl[60] br[60] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_61 bl[61] br[61] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_62 bl[62] br[62] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_160_63 bl[63] br[63] vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xcell_161_0 bl[0] br[0] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_1 bl[1] br[1] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_2 bl[2] br[2] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_3 bl[3] br[3] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_4 bl[4] br[4] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_5 bl[5] br[5] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_6 bl[6] br[6] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_7 bl[7] br[7] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_8 bl[8] br[8] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_9 bl[9] br[9] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_10 bl[10] br[10] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_11 bl[11] br[11] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_12 bl[12] br[12] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_13 bl[13] br[13] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_14 bl[14] br[14] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_15 bl[15] br[15] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_16 bl[16] br[16] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_17 bl[17] br[17] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_18 bl[18] br[18] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_19 bl[19] br[19] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_20 bl[20] br[20] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_21 bl[21] br[21] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_22 bl[22] br[22] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_23 bl[23] br[23] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_24 bl[24] br[24] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_25 bl[25] br[25] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_26 bl[26] br[26] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_27 bl[27] br[27] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_28 bl[28] br[28] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_29 bl[29] br[29] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_30 bl[30] br[30] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_31 bl[31] br[31] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_32 bl[32] br[32] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_33 bl[33] br[33] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_34 bl[34] br[34] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_35 bl[35] br[35] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_36 bl[36] br[36] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_37 bl[37] br[37] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_38 bl[38] br[38] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_39 bl[39] br[39] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_40 bl[40] br[40] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_41 bl[41] br[41] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_42 bl[42] br[42] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_43 bl[43] br[43] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_44 bl[44] br[44] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_45 bl[45] br[45] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_46 bl[46] br[46] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_47 bl[47] br[47] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_48 bl[48] br[48] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_49 bl[49] br[49] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_50 bl[50] br[50] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_51 bl[51] br[51] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_52 bl[52] br[52] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_53 bl[53] br[53] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_54 bl[54] br[54] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_55 bl[55] br[55] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_56 bl[56] br[56] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_57 bl[57] br[57] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_58 bl[58] br[58] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_59 bl[59] br[59] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_60 bl[60] br[60] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_61 bl[61] br[61] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_62 bl[62] br[62] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_161_63 bl[63] br[63] vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xcell_162_0 bl[0] br[0] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_1 bl[1] br[1] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_2 bl[2] br[2] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_3 bl[3] br[3] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_4 bl[4] br[4] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_5 bl[5] br[5] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_6 bl[6] br[6] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_7 bl[7] br[7] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_8 bl[8] br[8] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_9 bl[9] br[9] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_10 bl[10] br[10] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_11 bl[11] br[11] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_12 bl[12] br[12] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_13 bl[13] br[13] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_14 bl[14] br[14] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_15 bl[15] br[15] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_16 bl[16] br[16] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_17 bl[17] br[17] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_18 bl[18] br[18] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_19 bl[19] br[19] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_20 bl[20] br[20] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_21 bl[21] br[21] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_22 bl[22] br[22] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_23 bl[23] br[23] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_24 bl[24] br[24] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_25 bl[25] br[25] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_26 bl[26] br[26] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_27 bl[27] br[27] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_28 bl[28] br[28] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_29 bl[29] br[29] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_30 bl[30] br[30] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_31 bl[31] br[31] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_32 bl[32] br[32] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_33 bl[33] br[33] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_34 bl[34] br[34] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_35 bl[35] br[35] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_36 bl[36] br[36] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_37 bl[37] br[37] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_38 bl[38] br[38] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_39 bl[39] br[39] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_40 bl[40] br[40] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_41 bl[41] br[41] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_42 bl[42] br[42] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_43 bl[43] br[43] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_44 bl[44] br[44] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_45 bl[45] br[45] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_46 bl[46] br[46] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_47 bl[47] br[47] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_48 bl[48] br[48] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_49 bl[49] br[49] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_50 bl[50] br[50] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_51 bl[51] br[51] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_52 bl[52] br[52] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_53 bl[53] br[53] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_54 bl[54] br[54] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_55 bl[55] br[55] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_56 bl[56] br[56] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_57 bl[57] br[57] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_58 bl[58] br[58] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_59 bl[59] br[59] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_60 bl[60] br[60] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_61 bl[61] br[61] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_62 bl[62] br[62] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_162_63 bl[63] br[63] vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xcell_163_0 bl[0] br[0] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_1 bl[1] br[1] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_2 bl[2] br[2] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_3 bl[3] br[3] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_4 bl[4] br[4] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_5 bl[5] br[5] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_6 bl[6] br[6] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_7 bl[7] br[7] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_8 bl[8] br[8] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_9 bl[9] br[9] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_10 bl[10] br[10] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_11 bl[11] br[11] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_12 bl[12] br[12] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_13 bl[13] br[13] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_14 bl[14] br[14] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_15 bl[15] br[15] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_16 bl[16] br[16] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_17 bl[17] br[17] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_18 bl[18] br[18] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_19 bl[19] br[19] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_20 bl[20] br[20] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_21 bl[21] br[21] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_22 bl[22] br[22] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_23 bl[23] br[23] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_24 bl[24] br[24] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_25 bl[25] br[25] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_26 bl[26] br[26] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_27 bl[27] br[27] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_28 bl[28] br[28] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_29 bl[29] br[29] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_30 bl[30] br[30] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_31 bl[31] br[31] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_32 bl[32] br[32] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_33 bl[33] br[33] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_34 bl[34] br[34] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_35 bl[35] br[35] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_36 bl[36] br[36] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_37 bl[37] br[37] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_38 bl[38] br[38] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_39 bl[39] br[39] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_40 bl[40] br[40] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_41 bl[41] br[41] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_42 bl[42] br[42] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_43 bl[43] br[43] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_44 bl[44] br[44] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_45 bl[45] br[45] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_46 bl[46] br[46] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_47 bl[47] br[47] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_48 bl[48] br[48] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_49 bl[49] br[49] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_50 bl[50] br[50] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_51 bl[51] br[51] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_52 bl[52] br[52] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_53 bl[53] br[53] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_54 bl[54] br[54] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_55 bl[55] br[55] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_56 bl[56] br[56] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_57 bl[57] br[57] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_58 bl[58] br[58] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_59 bl[59] br[59] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_60 bl[60] br[60] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_61 bl[61] br[61] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_62 bl[62] br[62] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_163_63 bl[63] br[63] vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xcell_164_0 bl[0] br[0] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_1 bl[1] br[1] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_2 bl[2] br[2] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_3 bl[3] br[3] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_4 bl[4] br[4] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_5 bl[5] br[5] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_6 bl[6] br[6] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_7 bl[7] br[7] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_8 bl[8] br[8] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_9 bl[9] br[9] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_10 bl[10] br[10] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_11 bl[11] br[11] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_12 bl[12] br[12] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_13 bl[13] br[13] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_14 bl[14] br[14] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_15 bl[15] br[15] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_16 bl[16] br[16] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_17 bl[17] br[17] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_18 bl[18] br[18] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_19 bl[19] br[19] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_20 bl[20] br[20] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_21 bl[21] br[21] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_22 bl[22] br[22] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_23 bl[23] br[23] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_24 bl[24] br[24] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_25 bl[25] br[25] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_26 bl[26] br[26] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_27 bl[27] br[27] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_28 bl[28] br[28] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_29 bl[29] br[29] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_30 bl[30] br[30] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_31 bl[31] br[31] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_32 bl[32] br[32] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_33 bl[33] br[33] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_34 bl[34] br[34] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_35 bl[35] br[35] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_36 bl[36] br[36] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_37 bl[37] br[37] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_38 bl[38] br[38] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_39 bl[39] br[39] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_40 bl[40] br[40] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_41 bl[41] br[41] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_42 bl[42] br[42] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_43 bl[43] br[43] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_44 bl[44] br[44] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_45 bl[45] br[45] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_46 bl[46] br[46] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_47 bl[47] br[47] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_48 bl[48] br[48] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_49 bl[49] br[49] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_50 bl[50] br[50] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_51 bl[51] br[51] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_52 bl[52] br[52] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_53 bl[53] br[53] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_54 bl[54] br[54] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_55 bl[55] br[55] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_56 bl[56] br[56] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_57 bl[57] br[57] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_58 bl[58] br[58] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_59 bl[59] br[59] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_60 bl[60] br[60] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_61 bl[61] br[61] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_62 bl[62] br[62] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_164_63 bl[63] br[63] vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xcell_165_0 bl[0] br[0] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_1 bl[1] br[1] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_2 bl[2] br[2] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_3 bl[3] br[3] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_4 bl[4] br[4] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_5 bl[5] br[5] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_6 bl[6] br[6] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_7 bl[7] br[7] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_8 bl[8] br[8] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_9 bl[9] br[9] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_10 bl[10] br[10] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_11 bl[11] br[11] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_12 bl[12] br[12] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_13 bl[13] br[13] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_14 bl[14] br[14] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_15 bl[15] br[15] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_16 bl[16] br[16] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_17 bl[17] br[17] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_18 bl[18] br[18] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_19 bl[19] br[19] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_20 bl[20] br[20] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_21 bl[21] br[21] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_22 bl[22] br[22] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_23 bl[23] br[23] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_24 bl[24] br[24] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_25 bl[25] br[25] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_26 bl[26] br[26] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_27 bl[27] br[27] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_28 bl[28] br[28] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_29 bl[29] br[29] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_30 bl[30] br[30] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_31 bl[31] br[31] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_32 bl[32] br[32] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_33 bl[33] br[33] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_34 bl[34] br[34] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_35 bl[35] br[35] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_36 bl[36] br[36] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_37 bl[37] br[37] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_38 bl[38] br[38] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_39 bl[39] br[39] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_40 bl[40] br[40] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_41 bl[41] br[41] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_42 bl[42] br[42] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_43 bl[43] br[43] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_44 bl[44] br[44] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_45 bl[45] br[45] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_46 bl[46] br[46] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_47 bl[47] br[47] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_48 bl[48] br[48] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_49 bl[49] br[49] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_50 bl[50] br[50] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_51 bl[51] br[51] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_52 bl[52] br[52] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_53 bl[53] br[53] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_54 bl[54] br[54] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_55 bl[55] br[55] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_56 bl[56] br[56] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_57 bl[57] br[57] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_58 bl[58] br[58] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_59 bl[59] br[59] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_60 bl[60] br[60] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_61 bl[61] br[61] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_62 bl[62] br[62] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_165_63 bl[63] br[63] vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xcell_166_0 bl[0] br[0] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_1 bl[1] br[1] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_2 bl[2] br[2] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_3 bl[3] br[3] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_4 bl[4] br[4] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_5 bl[5] br[5] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_6 bl[6] br[6] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_7 bl[7] br[7] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_8 bl[8] br[8] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_9 bl[9] br[9] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_10 bl[10] br[10] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_11 bl[11] br[11] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_12 bl[12] br[12] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_13 bl[13] br[13] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_14 bl[14] br[14] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_15 bl[15] br[15] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_16 bl[16] br[16] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_17 bl[17] br[17] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_18 bl[18] br[18] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_19 bl[19] br[19] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_20 bl[20] br[20] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_21 bl[21] br[21] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_22 bl[22] br[22] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_23 bl[23] br[23] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_24 bl[24] br[24] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_25 bl[25] br[25] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_26 bl[26] br[26] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_27 bl[27] br[27] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_28 bl[28] br[28] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_29 bl[29] br[29] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_30 bl[30] br[30] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_31 bl[31] br[31] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_32 bl[32] br[32] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_33 bl[33] br[33] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_34 bl[34] br[34] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_35 bl[35] br[35] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_36 bl[36] br[36] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_37 bl[37] br[37] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_38 bl[38] br[38] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_39 bl[39] br[39] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_40 bl[40] br[40] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_41 bl[41] br[41] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_42 bl[42] br[42] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_43 bl[43] br[43] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_44 bl[44] br[44] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_45 bl[45] br[45] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_46 bl[46] br[46] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_47 bl[47] br[47] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_48 bl[48] br[48] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_49 bl[49] br[49] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_50 bl[50] br[50] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_51 bl[51] br[51] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_52 bl[52] br[52] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_53 bl[53] br[53] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_54 bl[54] br[54] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_55 bl[55] br[55] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_56 bl[56] br[56] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_57 bl[57] br[57] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_58 bl[58] br[58] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_59 bl[59] br[59] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_60 bl[60] br[60] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_61 bl[61] br[61] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_62 bl[62] br[62] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_166_63 bl[63] br[63] vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xcell_167_0 bl[0] br[0] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_1 bl[1] br[1] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_2 bl[2] br[2] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_3 bl[3] br[3] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_4 bl[4] br[4] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_5 bl[5] br[5] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_6 bl[6] br[6] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_7 bl[7] br[7] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_8 bl[8] br[8] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_9 bl[9] br[9] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_10 bl[10] br[10] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_11 bl[11] br[11] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_12 bl[12] br[12] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_13 bl[13] br[13] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_14 bl[14] br[14] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_15 bl[15] br[15] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_16 bl[16] br[16] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_17 bl[17] br[17] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_18 bl[18] br[18] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_19 bl[19] br[19] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_20 bl[20] br[20] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_21 bl[21] br[21] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_22 bl[22] br[22] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_23 bl[23] br[23] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_24 bl[24] br[24] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_25 bl[25] br[25] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_26 bl[26] br[26] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_27 bl[27] br[27] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_28 bl[28] br[28] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_29 bl[29] br[29] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_30 bl[30] br[30] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_31 bl[31] br[31] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_32 bl[32] br[32] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_33 bl[33] br[33] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_34 bl[34] br[34] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_35 bl[35] br[35] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_36 bl[36] br[36] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_37 bl[37] br[37] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_38 bl[38] br[38] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_39 bl[39] br[39] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_40 bl[40] br[40] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_41 bl[41] br[41] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_42 bl[42] br[42] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_43 bl[43] br[43] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_44 bl[44] br[44] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_45 bl[45] br[45] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_46 bl[46] br[46] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_47 bl[47] br[47] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_48 bl[48] br[48] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_49 bl[49] br[49] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_50 bl[50] br[50] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_51 bl[51] br[51] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_52 bl[52] br[52] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_53 bl[53] br[53] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_54 bl[54] br[54] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_55 bl[55] br[55] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_56 bl[56] br[56] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_57 bl[57] br[57] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_58 bl[58] br[58] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_59 bl[59] br[59] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_60 bl[60] br[60] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_61 bl[61] br[61] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_62 bl[62] br[62] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_167_63 bl[63] br[63] vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xcell_168_0 bl[0] br[0] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_1 bl[1] br[1] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_2 bl[2] br[2] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_3 bl[3] br[3] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_4 bl[4] br[4] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_5 bl[5] br[5] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_6 bl[6] br[6] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_7 bl[7] br[7] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_8 bl[8] br[8] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_9 bl[9] br[9] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_10 bl[10] br[10] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_11 bl[11] br[11] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_12 bl[12] br[12] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_13 bl[13] br[13] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_14 bl[14] br[14] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_15 bl[15] br[15] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_16 bl[16] br[16] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_17 bl[17] br[17] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_18 bl[18] br[18] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_19 bl[19] br[19] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_20 bl[20] br[20] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_21 bl[21] br[21] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_22 bl[22] br[22] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_23 bl[23] br[23] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_24 bl[24] br[24] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_25 bl[25] br[25] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_26 bl[26] br[26] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_27 bl[27] br[27] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_28 bl[28] br[28] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_29 bl[29] br[29] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_30 bl[30] br[30] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_31 bl[31] br[31] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_32 bl[32] br[32] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_33 bl[33] br[33] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_34 bl[34] br[34] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_35 bl[35] br[35] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_36 bl[36] br[36] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_37 bl[37] br[37] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_38 bl[38] br[38] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_39 bl[39] br[39] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_40 bl[40] br[40] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_41 bl[41] br[41] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_42 bl[42] br[42] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_43 bl[43] br[43] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_44 bl[44] br[44] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_45 bl[45] br[45] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_46 bl[46] br[46] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_47 bl[47] br[47] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_48 bl[48] br[48] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_49 bl[49] br[49] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_50 bl[50] br[50] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_51 bl[51] br[51] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_52 bl[52] br[52] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_53 bl[53] br[53] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_54 bl[54] br[54] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_55 bl[55] br[55] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_56 bl[56] br[56] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_57 bl[57] br[57] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_58 bl[58] br[58] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_59 bl[59] br[59] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_60 bl[60] br[60] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_61 bl[61] br[61] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_62 bl[62] br[62] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_168_63 bl[63] br[63] vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xcell_169_0 bl[0] br[0] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_1 bl[1] br[1] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_2 bl[2] br[2] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_3 bl[3] br[3] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_4 bl[4] br[4] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_5 bl[5] br[5] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_6 bl[6] br[6] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_7 bl[7] br[7] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_8 bl[8] br[8] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_9 bl[9] br[9] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_10 bl[10] br[10] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_11 bl[11] br[11] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_12 bl[12] br[12] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_13 bl[13] br[13] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_14 bl[14] br[14] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_15 bl[15] br[15] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_16 bl[16] br[16] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_17 bl[17] br[17] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_18 bl[18] br[18] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_19 bl[19] br[19] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_20 bl[20] br[20] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_21 bl[21] br[21] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_22 bl[22] br[22] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_23 bl[23] br[23] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_24 bl[24] br[24] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_25 bl[25] br[25] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_26 bl[26] br[26] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_27 bl[27] br[27] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_28 bl[28] br[28] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_29 bl[29] br[29] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_30 bl[30] br[30] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_31 bl[31] br[31] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_32 bl[32] br[32] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_33 bl[33] br[33] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_34 bl[34] br[34] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_35 bl[35] br[35] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_36 bl[36] br[36] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_37 bl[37] br[37] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_38 bl[38] br[38] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_39 bl[39] br[39] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_40 bl[40] br[40] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_41 bl[41] br[41] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_42 bl[42] br[42] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_43 bl[43] br[43] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_44 bl[44] br[44] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_45 bl[45] br[45] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_46 bl[46] br[46] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_47 bl[47] br[47] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_48 bl[48] br[48] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_49 bl[49] br[49] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_50 bl[50] br[50] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_51 bl[51] br[51] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_52 bl[52] br[52] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_53 bl[53] br[53] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_54 bl[54] br[54] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_55 bl[55] br[55] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_56 bl[56] br[56] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_57 bl[57] br[57] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_58 bl[58] br[58] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_59 bl[59] br[59] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_60 bl[60] br[60] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_61 bl[61] br[61] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_62 bl[62] br[62] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_169_63 bl[63] br[63] vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xcell_170_0 bl[0] br[0] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_1 bl[1] br[1] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_2 bl[2] br[2] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_3 bl[3] br[3] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_4 bl[4] br[4] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_5 bl[5] br[5] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_6 bl[6] br[6] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_7 bl[7] br[7] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_8 bl[8] br[8] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_9 bl[9] br[9] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_10 bl[10] br[10] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_11 bl[11] br[11] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_12 bl[12] br[12] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_13 bl[13] br[13] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_14 bl[14] br[14] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_15 bl[15] br[15] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_16 bl[16] br[16] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_17 bl[17] br[17] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_18 bl[18] br[18] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_19 bl[19] br[19] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_20 bl[20] br[20] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_21 bl[21] br[21] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_22 bl[22] br[22] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_23 bl[23] br[23] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_24 bl[24] br[24] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_25 bl[25] br[25] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_26 bl[26] br[26] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_27 bl[27] br[27] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_28 bl[28] br[28] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_29 bl[29] br[29] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_30 bl[30] br[30] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_31 bl[31] br[31] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_32 bl[32] br[32] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_33 bl[33] br[33] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_34 bl[34] br[34] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_35 bl[35] br[35] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_36 bl[36] br[36] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_37 bl[37] br[37] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_38 bl[38] br[38] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_39 bl[39] br[39] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_40 bl[40] br[40] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_41 bl[41] br[41] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_42 bl[42] br[42] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_43 bl[43] br[43] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_44 bl[44] br[44] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_45 bl[45] br[45] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_46 bl[46] br[46] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_47 bl[47] br[47] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_48 bl[48] br[48] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_49 bl[49] br[49] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_50 bl[50] br[50] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_51 bl[51] br[51] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_52 bl[52] br[52] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_53 bl[53] br[53] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_54 bl[54] br[54] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_55 bl[55] br[55] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_56 bl[56] br[56] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_57 bl[57] br[57] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_58 bl[58] br[58] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_59 bl[59] br[59] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_60 bl[60] br[60] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_61 bl[61] br[61] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_62 bl[62] br[62] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_170_63 bl[63] br[63] vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xcell_171_0 bl[0] br[0] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_1 bl[1] br[1] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_2 bl[2] br[2] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_3 bl[3] br[3] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_4 bl[4] br[4] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_5 bl[5] br[5] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_6 bl[6] br[6] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_7 bl[7] br[7] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_8 bl[8] br[8] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_9 bl[9] br[9] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_10 bl[10] br[10] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_11 bl[11] br[11] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_12 bl[12] br[12] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_13 bl[13] br[13] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_14 bl[14] br[14] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_15 bl[15] br[15] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_16 bl[16] br[16] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_17 bl[17] br[17] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_18 bl[18] br[18] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_19 bl[19] br[19] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_20 bl[20] br[20] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_21 bl[21] br[21] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_22 bl[22] br[22] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_23 bl[23] br[23] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_24 bl[24] br[24] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_25 bl[25] br[25] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_26 bl[26] br[26] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_27 bl[27] br[27] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_28 bl[28] br[28] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_29 bl[29] br[29] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_30 bl[30] br[30] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_31 bl[31] br[31] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_32 bl[32] br[32] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_33 bl[33] br[33] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_34 bl[34] br[34] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_35 bl[35] br[35] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_36 bl[36] br[36] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_37 bl[37] br[37] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_38 bl[38] br[38] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_39 bl[39] br[39] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_40 bl[40] br[40] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_41 bl[41] br[41] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_42 bl[42] br[42] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_43 bl[43] br[43] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_44 bl[44] br[44] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_45 bl[45] br[45] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_46 bl[46] br[46] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_47 bl[47] br[47] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_48 bl[48] br[48] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_49 bl[49] br[49] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_50 bl[50] br[50] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_51 bl[51] br[51] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_52 bl[52] br[52] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_53 bl[53] br[53] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_54 bl[54] br[54] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_55 bl[55] br[55] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_56 bl[56] br[56] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_57 bl[57] br[57] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_58 bl[58] br[58] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_59 bl[59] br[59] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_60 bl[60] br[60] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_61 bl[61] br[61] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_62 bl[62] br[62] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_171_63 bl[63] br[63] vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xcell_172_0 bl[0] br[0] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_1 bl[1] br[1] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_2 bl[2] br[2] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_3 bl[3] br[3] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_4 bl[4] br[4] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_5 bl[5] br[5] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_6 bl[6] br[6] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_7 bl[7] br[7] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_8 bl[8] br[8] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_9 bl[9] br[9] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_10 bl[10] br[10] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_11 bl[11] br[11] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_12 bl[12] br[12] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_13 bl[13] br[13] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_14 bl[14] br[14] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_15 bl[15] br[15] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_16 bl[16] br[16] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_17 bl[17] br[17] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_18 bl[18] br[18] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_19 bl[19] br[19] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_20 bl[20] br[20] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_21 bl[21] br[21] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_22 bl[22] br[22] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_23 bl[23] br[23] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_24 bl[24] br[24] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_25 bl[25] br[25] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_26 bl[26] br[26] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_27 bl[27] br[27] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_28 bl[28] br[28] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_29 bl[29] br[29] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_30 bl[30] br[30] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_31 bl[31] br[31] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_32 bl[32] br[32] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_33 bl[33] br[33] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_34 bl[34] br[34] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_35 bl[35] br[35] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_36 bl[36] br[36] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_37 bl[37] br[37] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_38 bl[38] br[38] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_39 bl[39] br[39] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_40 bl[40] br[40] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_41 bl[41] br[41] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_42 bl[42] br[42] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_43 bl[43] br[43] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_44 bl[44] br[44] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_45 bl[45] br[45] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_46 bl[46] br[46] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_47 bl[47] br[47] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_48 bl[48] br[48] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_49 bl[49] br[49] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_50 bl[50] br[50] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_51 bl[51] br[51] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_52 bl[52] br[52] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_53 bl[53] br[53] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_54 bl[54] br[54] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_55 bl[55] br[55] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_56 bl[56] br[56] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_57 bl[57] br[57] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_58 bl[58] br[58] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_59 bl[59] br[59] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_60 bl[60] br[60] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_61 bl[61] br[61] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_62 bl[62] br[62] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_172_63 bl[63] br[63] vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xcell_173_0 bl[0] br[0] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_1 bl[1] br[1] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_2 bl[2] br[2] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_3 bl[3] br[3] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_4 bl[4] br[4] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_5 bl[5] br[5] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_6 bl[6] br[6] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_7 bl[7] br[7] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_8 bl[8] br[8] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_9 bl[9] br[9] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_10 bl[10] br[10] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_11 bl[11] br[11] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_12 bl[12] br[12] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_13 bl[13] br[13] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_14 bl[14] br[14] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_15 bl[15] br[15] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_16 bl[16] br[16] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_17 bl[17] br[17] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_18 bl[18] br[18] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_19 bl[19] br[19] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_20 bl[20] br[20] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_21 bl[21] br[21] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_22 bl[22] br[22] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_23 bl[23] br[23] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_24 bl[24] br[24] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_25 bl[25] br[25] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_26 bl[26] br[26] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_27 bl[27] br[27] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_28 bl[28] br[28] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_29 bl[29] br[29] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_30 bl[30] br[30] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_31 bl[31] br[31] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_32 bl[32] br[32] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_33 bl[33] br[33] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_34 bl[34] br[34] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_35 bl[35] br[35] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_36 bl[36] br[36] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_37 bl[37] br[37] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_38 bl[38] br[38] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_39 bl[39] br[39] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_40 bl[40] br[40] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_41 bl[41] br[41] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_42 bl[42] br[42] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_43 bl[43] br[43] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_44 bl[44] br[44] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_45 bl[45] br[45] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_46 bl[46] br[46] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_47 bl[47] br[47] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_48 bl[48] br[48] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_49 bl[49] br[49] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_50 bl[50] br[50] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_51 bl[51] br[51] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_52 bl[52] br[52] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_53 bl[53] br[53] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_54 bl[54] br[54] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_55 bl[55] br[55] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_56 bl[56] br[56] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_57 bl[57] br[57] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_58 bl[58] br[58] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_59 bl[59] br[59] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_60 bl[60] br[60] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_61 bl[61] br[61] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_62 bl[62] br[62] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_173_63 bl[63] br[63] vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xcell_174_0 bl[0] br[0] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_1 bl[1] br[1] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_2 bl[2] br[2] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_3 bl[3] br[3] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_4 bl[4] br[4] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_5 bl[5] br[5] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_6 bl[6] br[6] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_7 bl[7] br[7] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_8 bl[8] br[8] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_9 bl[9] br[9] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_10 bl[10] br[10] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_11 bl[11] br[11] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_12 bl[12] br[12] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_13 bl[13] br[13] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_14 bl[14] br[14] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_15 bl[15] br[15] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_16 bl[16] br[16] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_17 bl[17] br[17] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_18 bl[18] br[18] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_19 bl[19] br[19] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_20 bl[20] br[20] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_21 bl[21] br[21] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_22 bl[22] br[22] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_23 bl[23] br[23] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_24 bl[24] br[24] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_25 bl[25] br[25] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_26 bl[26] br[26] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_27 bl[27] br[27] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_28 bl[28] br[28] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_29 bl[29] br[29] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_30 bl[30] br[30] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_31 bl[31] br[31] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_32 bl[32] br[32] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_33 bl[33] br[33] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_34 bl[34] br[34] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_35 bl[35] br[35] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_36 bl[36] br[36] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_37 bl[37] br[37] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_38 bl[38] br[38] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_39 bl[39] br[39] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_40 bl[40] br[40] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_41 bl[41] br[41] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_42 bl[42] br[42] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_43 bl[43] br[43] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_44 bl[44] br[44] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_45 bl[45] br[45] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_46 bl[46] br[46] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_47 bl[47] br[47] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_48 bl[48] br[48] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_49 bl[49] br[49] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_50 bl[50] br[50] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_51 bl[51] br[51] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_52 bl[52] br[52] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_53 bl[53] br[53] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_54 bl[54] br[54] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_55 bl[55] br[55] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_56 bl[56] br[56] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_57 bl[57] br[57] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_58 bl[58] br[58] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_59 bl[59] br[59] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_60 bl[60] br[60] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_61 bl[61] br[61] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_62 bl[62] br[62] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_174_63 bl[63] br[63] vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xcell_175_0 bl[0] br[0] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_1 bl[1] br[1] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_2 bl[2] br[2] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_3 bl[3] br[3] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_4 bl[4] br[4] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_5 bl[5] br[5] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_6 bl[6] br[6] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_7 bl[7] br[7] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_8 bl[8] br[8] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_9 bl[9] br[9] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_10 bl[10] br[10] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_11 bl[11] br[11] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_12 bl[12] br[12] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_13 bl[13] br[13] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_14 bl[14] br[14] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_15 bl[15] br[15] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_16 bl[16] br[16] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_17 bl[17] br[17] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_18 bl[18] br[18] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_19 bl[19] br[19] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_20 bl[20] br[20] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_21 bl[21] br[21] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_22 bl[22] br[22] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_23 bl[23] br[23] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_24 bl[24] br[24] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_25 bl[25] br[25] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_26 bl[26] br[26] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_27 bl[27] br[27] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_28 bl[28] br[28] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_29 bl[29] br[29] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_30 bl[30] br[30] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_31 bl[31] br[31] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_32 bl[32] br[32] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_33 bl[33] br[33] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_34 bl[34] br[34] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_35 bl[35] br[35] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_36 bl[36] br[36] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_37 bl[37] br[37] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_38 bl[38] br[38] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_39 bl[39] br[39] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_40 bl[40] br[40] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_41 bl[41] br[41] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_42 bl[42] br[42] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_43 bl[43] br[43] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_44 bl[44] br[44] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_45 bl[45] br[45] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_46 bl[46] br[46] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_47 bl[47] br[47] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_48 bl[48] br[48] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_49 bl[49] br[49] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_50 bl[50] br[50] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_51 bl[51] br[51] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_52 bl[52] br[52] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_53 bl[53] br[53] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_54 bl[54] br[54] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_55 bl[55] br[55] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_56 bl[56] br[56] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_57 bl[57] br[57] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_58 bl[58] br[58] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_59 bl[59] br[59] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_60 bl[60] br[60] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_61 bl[61] br[61] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_62 bl[62] br[62] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_175_63 bl[63] br[63] vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xcell_176_0 bl[0] br[0] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_1 bl[1] br[1] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_2 bl[2] br[2] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_3 bl[3] br[3] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_4 bl[4] br[4] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_5 bl[5] br[5] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_6 bl[6] br[6] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_7 bl[7] br[7] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_8 bl[8] br[8] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_9 bl[9] br[9] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_10 bl[10] br[10] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_11 bl[11] br[11] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_12 bl[12] br[12] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_13 bl[13] br[13] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_14 bl[14] br[14] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_15 bl[15] br[15] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_16 bl[16] br[16] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_17 bl[17] br[17] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_18 bl[18] br[18] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_19 bl[19] br[19] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_20 bl[20] br[20] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_21 bl[21] br[21] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_22 bl[22] br[22] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_23 bl[23] br[23] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_24 bl[24] br[24] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_25 bl[25] br[25] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_26 bl[26] br[26] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_27 bl[27] br[27] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_28 bl[28] br[28] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_29 bl[29] br[29] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_30 bl[30] br[30] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_31 bl[31] br[31] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_32 bl[32] br[32] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_33 bl[33] br[33] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_34 bl[34] br[34] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_35 bl[35] br[35] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_36 bl[36] br[36] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_37 bl[37] br[37] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_38 bl[38] br[38] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_39 bl[39] br[39] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_40 bl[40] br[40] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_41 bl[41] br[41] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_42 bl[42] br[42] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_43 bl[43] br[43] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_44 bl[44] br[44] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_45 bl[45] br[45] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_46 bl[46] br[46] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_47 bl[47] br[47] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_48 bl[48] br[48] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_49 bl[49] br[49] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_50 bl[50] br[50] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_51 bl[51] br[51] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_52 bl[52] br[52] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_53 bl[53] br[53] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_54 bl[54] br[54] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_55 bl[55] br[55] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_56 bl[56] br[56] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_57 bl[57] br[57] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_58 bl[58] br[58] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_59 bl[59] br[59] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_60 bl[60] br[60] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_61 bl[61] br[61] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_62 bl[62] br[62] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_176_63 bl[63] br[63] vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xcell_177_0 bl[0] br[0] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_1 bl[1] br[1] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_2 bl[2] br[2] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_3 bl[3] br[3] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_4 bl[4] br[4] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_5 bl[5] br[5] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_6 bl[6] br[6] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_7 bl[7] br[7] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_8 bl[8] br[8] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_9 bl[9] br[9] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_10 bl[10] br[10] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_11 bl[11] br[11] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_12 bl[12] br[12] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_13 bl[13] br[13] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_14 bl[14] br[14] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_15 bl[15] br[15] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_16 bl[16] br[16] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_17 bl[17] br[17] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_18 bl[18] br[18] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_19 bl[19] br[19] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_20 bl[20] br[20] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_21 bl[21] br[21] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_22 bl[22] br[22] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_23 bl[23] br[23] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_24 bl[24] br[24] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_25 bl[25] br[25] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_26 bl[26] br[26] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_27 bl[27] br[27] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_28 bl[28] br[28] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_29 bl[29] br[29] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_30 bl[30] br[30] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_31 bl[31] br[31] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_32 bl[32] br[32] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_33 bl[33] br[33] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_34 bl[34] br[34] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_35 bl[35] br[35] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_36 bl[36] br[36] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_37 bl[37] br[37] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_38 bl[38] br[38] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_39 bl[39] br[39] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_40 bl[40] br[40] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_41 bl[41] br[41] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_42 bl[42] br[42] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_43 bl[43] br[43] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_44 bl[44] br[44] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_45 bl[45] br[45] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_46 bl[46] br[46] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_47 bl[47] br[47] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_48 bl[48] br[48] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_49 bl[49] br[49] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_50 bl[50] br[50] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_51 bl[51] br[51] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_52 bl[52] br[52] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_53 bl[53] br[53] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_54 bl[54] br[54] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_55 bl[55] br[55] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_56 bl[56] br[56] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_57 bl[57] br[57] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_58 bl[58] br[58] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_59 bl[59] br[59] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_60 bl[60] br[60] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_61 bl[61] br[61] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_62 bl[62] br[62] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_177_63 bl[63] br[63] vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xcell_178_0 bl[0] br[0] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_1 bl[1] br[1] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_2 bl[2] br[2] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_3 bl[3] br[3] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_4 bl[4] br[4] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_5 bl[5] br[5] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_6 bl[6] br[6] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_7 bl[7] br[7] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_8 bl[8] br[8] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_9 bl[9] br[9] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_10 bl[10] br[10] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_11 bl[11] br[11] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_12 bl[12] br[12] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_13 bl[13] br[13] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_14 bl[14] br[14] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_15 bl[15] br[15] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_16 bl[16] br[16] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_17 bl[17] br[17] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_18 bl[18] br[18] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_19 bl[19] br[19] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_20 bl[20] br[20] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_21 bl[21] br[21] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_22 bl[22] br[22] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_23 bl[23] br[23] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_24 bl[24] br[24] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_25 bl[25] br[25] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_26 bl[26] br[26] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_27 bl[27] br[27] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_28 bl[28] br[28] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_29 bl[29] br[29] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_30 bl[30] br[30] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_31 bl[31] br[31] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_32 bl[32] br[32] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_33 bl[33] br[33] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_34 bl[34] br[34] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_35 bl[35] br[35] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_36 bl[36] br[36] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_37 bl[37] br[37] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_38 bl[38] br[38] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_39 bl[39] br[39] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_40 bl[40] br[40] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_41 bl[41] br[41] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_42 bl[42] br[42] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_43 bl[43] br[43] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_44 bl[44] br[44] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_45 bl[45] br[45] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_46 bl[46] br[46] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_47 bl[47] br[47] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_48 bl[48] br[48] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_49 bl[49] br[49] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_50 bl[50] br[50] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_51 bl[51] br[51] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_52 bl[52] br[52] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_53 bl[53] br[53] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_54 bl[54] br[54] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_55 bl[55] br[55] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_56 bl[56] br[56] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_57 bl[57] br[57] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_58 bl[58] br[58] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_59 bl[59] br[59] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_60 bl[60] br[60] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_61 bl[61] br[61] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_62 bl[62] br[62] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_178_63 bl[63] br[63] vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xcell_179_0 bl[0] br[0] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_1 bl[1] br[1] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_2 bl[2] br[2] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_3 bl[3] br[3] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_4 bl[4] br[4] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_5 bl[5] br[5] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_6 bl[6] br[6] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_7 bl[7] br[7] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_8 bl[8] br[8] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_9 bl[9] br[9] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_10 bl[10] br[10] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_11 bl[11] br[11] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_12 bl[12] br[12] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_13 bl[13] br[13] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_14 bl[14] br[14] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_15 bl[15] br[15] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_16 bl[16] br[16] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_17 bl[17] br[17] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_18 bl[18] br[18] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_19 bl[19] br[19] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_20 bl[20] br[20] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_21 bl[21] br[21] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_22 bl[22] br[22] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_23 bl[23] br[23] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_24 bl[24] br[24] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_25 bl[25] br[25] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_26 bl[26] br[26] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_27 bl[27] br[27] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_28 bl[28] br[28] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_29 bl[29] br[29] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_30 bl[30] br[30] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_31 bl[31] br[31] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_32 bl[32] br[32] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_33 bl[33] br[33] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_34 bl[34] br[34] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_35 bl[35] br[35] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_36 bl[36] br[36] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_37 bl[37] br[37] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_38 bl[38] br[38] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_39 bl[39] br[39] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_40 bl[40] br[40] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_41 bl[41] br[41] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_42 bl[42] br[42] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_43 bl[43] br[43] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_44 bl[44] br[44] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_45 bl[45] br[45] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_46 bl[46] br[46] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_47 bl[47] br[47] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_48 bl[48] br[48] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_49 bl[49] br[49] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_50 bl[50] br[50] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_51 bl[51] br[51] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_52 bl[52] br[52] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_53 bl[53] br[53] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_54 bl[54] br[54] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_55 bl[55] br[55] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_56 bl[56] br[56] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_57 bl[57] br[57] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_58 bl[58] br[58] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_59 bl[59] br[59] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_60 bl[60] br[60] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_61 bl[61] br[61] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_62 bl[62] br[62] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_179_63 bl[63] br[63] vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xcell_180_0 bl[0] br[0] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_1 bl[1] br[1] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_2 bl[2] br[2] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_3 bl[3] br[3] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_4 bl[4] br[4] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_5 bl[5] br[5] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_6 bl[6] br[6] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_7 bl[7] br[7] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_8 bl[8] br[8] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_9 bl[9] br[9] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_10 bl[10] br[10] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_11 bl[11] br[11] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_12 bl[12] br[12] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_13 bl[13] br[13] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_14 bl[14] br[14] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_15 bl[15] br[15] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_16 bl[16] br[16] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_17 bl[17] br[17] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_18 bl[18] br[18] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_19 bl[19] br[19] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_20 bl[20] br[20] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_21 bl[21] br[21] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_22 bl[22] br[22] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_23 bl[23] br[23] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_24 bl[24] br[24] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_25 bl[25] br[25] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_26 bl[26] br[26] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_27 bl[27] br[27] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_28 bl[28] br[28] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_29 bl[29] br[29] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_30 bl[30] br[30] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_31 bl[31] br[31] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_32 bl[32] br[32] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_33 bl[33] br[33] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_34 bl[34] br[34] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_35 bl[35] br[35] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_36 bl[36] br[36] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_37 bl[37] br[37] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_38 bl[38] br[38] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_39 bl[39] br[39] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_40 bl[40] br[40] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_41 bl[41] br[41] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_42 bl[42] br[42] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_43 bl[43] br[43] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_44 bl[44] br[44] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_45 bl[45] br[45] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_46 bl[46] br[46] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_47 bl[47] br[47] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_48 bl[48] br[48] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_49 bl[49] br[49] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_50 bl[50] br[50] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_51 bl[51] br[51] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_52 bl[52] br[52] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_53 bl[53] br[53] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_54 bl[54] br[54] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_55 bl[55] br[55] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_56 bl[56] br[56] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_57 bl[57] br[57] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_58 bl[58] br[58] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_59 bl[59] br[59] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_60 bl[60] br[60] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_61 bl[61] br[61] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_62 bl[62] br[62] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_180_63 bl[63] br[63] vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xcell_181_0 bl[0] br[0] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_1 bl[1] br[1] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_2 bl[2] br[2] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_3 bl[3] br[3] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_4 bl[4] br[4] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_5 bl[5] br[5] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_6 bl[6] br[6] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_7 bl[7] br[7] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_8 bl[8] br[8] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_9 bl[9] br[9] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_10 bl[10] br[10] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_11 bl[11] br[11] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_12 bl[12] br[12] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_13 bl[13] br[13] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_14 bl[14] br[14] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_15 bl[15] br[15] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_16 bl[16] br[16] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_17 bl[17] br[17] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_18 bl[18] br[18] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_19 bl[19] br[19] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_20 bl[20] br[20] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_21 bl[21] br[21] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_22 bl[22] br[22] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_23 bl[23] br[23] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_24 bl[24] br[24] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_25 bl[25] br[25] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_26 bl[26] br[26] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_27 bl[27] br[27] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_28 bl[28] br[28] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_29 bl[29] br[29] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_30 bl[30] br[30] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_31 bl[31] br[31] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_32 bl[32] br[32] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_33 bl[33] br[33] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_34 bl[34] br[34] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_35 bl[35] br[35] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_36 bl[36] br[36] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_37 bl[37] br[37] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_38 bl[38] br[38] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_39 bl[39] br[39] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_40 bl[40] br[40] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_41 bl[41] br[41] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_42 bl[42] br[42] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_43 bl[43] br[43] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_44 bl[44] br[44] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_45 bl[45] br[45] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_46 bl[46] br[46] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_47 bl[47] br[47] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_48 bl[48] br[48] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_49 bl[49] br[49] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_50 bl[50] br[50] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_51 bl[51] br[51] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_52 bl[52] br[52] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_53 bl[53] br[53] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_54 bl[54] br[54] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_55 bl[55] br[55] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_56 bl[56] br[56] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_57 bl[57] br[57] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_58 bl[58] br[58] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_59 bl[59] br[59] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_60 bl[60] br[60] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_61 bl[61] br[61] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_62 bl[62] br[62] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_181_63 bl[63] br[63] vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xcell_182_0 bl[0] br[0] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_1 bl[1] br[1] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_2 bl[2] br[2] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_3 bl[3] br[3] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_4 bl[4] br[4] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_5 bl[5] br[5] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_6 bl[6] br[6] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_7 bl[7] br[7] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_8 bl[8] br[8] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_9 bl[9] br[9] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_10 bl[10] br[10] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_11 bl[11] br[11] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_12 bl[12] br[12] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_13 bl[13] br[13] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_14 bl[14] br[14] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_15 bl[15] br[15] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_16 bl[16] br[16] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_17 bl[17] br[17] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_18 bl[18] br[18] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_19 bl[19] br[19] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_20 bl[20] br[20] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_21 bl[21] br[21] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_22 bl[22] br[22] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_23 bl[23] br[23] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_24 bl[24] br[24] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_25 bl[25] br[25] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_26 bl[26] br[26] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_27 bl[27] br[27] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_28 bl[28] br[28] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_29 bl[29] br[29] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_30 bl[30] br[30] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_31 bl[31] br[31] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_32 bl[32] br[32] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_33 bl[33] br[33] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_34 bl[34] br[34] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_35 bl[35] br[35] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_36 bl[36] br[36] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_37 bl[37] br[37] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_38 bl[38] br[38] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_39 bl[39] br[39] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_40 bl[40] br[40] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_41 bl[41] br[41] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_42 bl[42] br[42] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_43 bl[43] br[43] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_44 bl[44] br[44] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_45 bl[45] br[45] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_46 bl[46] br[46] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_47 bl[47] br[47] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_48 bl[48] br[48] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_49 bl[49] br[49] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_50 bl[50] br[50] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_51 bl[51] br[51] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_52 bl[52] br[52] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_53 bl[53] br[53] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_54 bl[54] br[54] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_55 bl[55] br[55] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_56 bl[56] br[56] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_57 bl[57] br[57] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_58 bl[58] br[58] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_59 bl[59] br[59] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_60 bl[60] br[60] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_61 bl[61] br[61] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_62 bl[62] br[62] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_182_63 bl[63] br[63] vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xcell_183_0 bl[0] br[0] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_1 bl[1] br[1] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_2 bl[2] br[2] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_3 bl[3] br[3] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_4 bl[4] br[4] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_5 bl[5] br[5] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_6 bl[6] br[6] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_7 bl[7] br[7] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_8 bl[8] br[8] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_9 bl[9] br[9] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_10 bl[10] br[10] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_11 bl[11] br[11] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_12 bl[12] br[12] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_13 bl[13] br[13] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_14 bl[14] br[14] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_15 bl[15] br[15] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_16 bl[16] br[16] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_17 bl[17] br[17] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_18 bl[18] br[18] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_19 bl[19] br[19] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_20 bl[20] br[20] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_21 bl[21] br[21] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_22 bl[22] br[22] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_23 bl[23] br[23] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_24 bl[24] br[24] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_25 bl[25] br[25] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_26 bl[26] br[26] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_27 bl[27] br[27] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_28 bl[28] br[28] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_29 bl[29] br[29] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_30 bl[30] br[30] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_31 bl[31] br[31] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_32 bl[32] br[32] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_33 bl[33] br[33] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_34 bl[34] br[34] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_35 bl[35] br[35] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_36 bl[36] br[36] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_37 bl[37] br[37] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_38 bl[38] br[38] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_39 bl[39] br[39] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_40 bl[40] br[40] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_41 bl[41] br[41] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_42 bl[42] br[42] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_43 bl[43] br[43] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_44 bl[44] br[44] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_45 bl[45] br[45] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_46 bl[46] br[46] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_47 bl[47] br[47] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_48 bl[48] br[48] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_49 bl[49] br[49] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_50 bl[50] br[50] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_51 bl[51] br[51] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_52 bl[52] br[52] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_53 bl[53] br[53] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_54 bl[54] br[54] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_55 bl[55] br[55] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_56 bl[56] br[56] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_57 bl[57] br[57] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_58 bl[58] br[58] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_59 bl[59] br[59] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_60 bl[60] br[60] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_61 bl[61] br[61] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_62 bl[62] br[62] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_183_63 bl[63] br[63] vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xcell_184_0 bl[0] br[0] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_1 bl[1] br[1] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_2 bl[2] br[2] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_3 bl[3] br[3] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_4 bl[4] br[4] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_5 bl[5] br[5] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_6 bl[6] br[6] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_7 bl[7] br[7] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_8 bl[8] br[8] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_9 bl[9] br[9] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_10 bl[10] br[10] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_11 bl[11] br[11] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_12 bl[12] br[12] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_13 bl[13] br[13] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_14 bl[14] br[14] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_15 bl[15] br[15] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_16 bl[16] br[16] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_17 bl[17] br[17] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_18 bl[18] br[18] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_19 bl[19] br[19] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_20 bl[20] br[20] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_21 bl[21] br[21] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_22 bl[22] br[22] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_23 bl[23] br[23] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_24 bl[24] br[24] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_25 bl[25] br[25] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_26 bl[26] br[26] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_27 bl[27] br[27] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_28 bl[28] br[28] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_29 bl[29] br[29] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_30 bl[30] br[30] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_31 bl[31] br[31] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_32 bl[32] br[32] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_33 bl[33] br[33] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_34 bl[34] br[34] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_35 bl[35] br[35] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_36 bl[36] br[36] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_37 bl[37] br[37] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_38 bl[38] br[38] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_39 bl[39] br[39] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_40 bl[40] br[40] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_41 bl[41] br[41] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_42 bl[42] br[42] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_43 bl[43] br[43] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_44 bl[44] br[44] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_45 bl[45] br[45] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_46 bl[46] br[46] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_47 bl[47] br[47] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_48 bl[48] br[48] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_49 bl[49] br[49] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_50 bl[50] br[50] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_51 bl[51] br[51] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_52 bl[52] br[52] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_53 bl[53] br[53] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_54 bl[54] br[54] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_55 bl[55] br[55] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_56 bl[56] br[56] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_57 bl[57] br[57] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_58 bl[58] br[58] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_59 bl[59] br[59] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_60 bl[60] br[60] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_61 bl[61] br[61] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_62 bl[62] br[62] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_184_63 bl[63] br[63] vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xcell_185_0 bl[0] br[0] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_1 bl[1] br[1] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_2 bl[2] br[2] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_3 bl[3] br[3] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_4 bl[4] br[4] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_5 bl[5] br[5] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_6 bl[6] br[6] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_7 bl[7] br[7] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_8 bl[8] br[8] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_9 bl[9] br[9] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_10 bl[10] br[10] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_11 bl[11] br[11] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_12 bl[12] br[12] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_13 bl[13] br[13] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_14 bl[14] br[14] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_15 bl[15] br[15] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_16 bl[16] br[16] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_17 bl[17] br[17] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_18 bl[18] br[18] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_19 bl[19] br[19] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_20 bl[20] br[20] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_21 bl[21] br[21] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_22 bl[22] br[22] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_23 bl[23] br[23] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_24 bl[24] br[24] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_25 bl[25] br[25] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_26 bl[26] br[26] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_27 bl[27] br[27] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_28 bl[28] br[28] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_29 bl[29] br[29] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_30 bl[30] br[30] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_31 bl[31] br[31] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_32 bl[32] br[32] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_33 bl[33] br[33] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_34 bl[34] br[34] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_35 bl[35] br[35] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_36 bl[36] br[36] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_37 bl[37] br[37] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_38 bl[38] br[38] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_39 bl[39] br[39] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_40 bl[40] br[40] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_41 bl[41] br[41] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_42 bl[42] br[42] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_43 bl[43] br[43] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_44 bl[44] br[44] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_45 bl[45] br[45] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_46 bl[46] br[46] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_47 bl[47] br[47] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_48 bl[48] br[48] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_49 bl[49] br[49] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_50 bl[50] br[50] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_51 bl[51] br[51] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_52 bl[52] br[52] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_53 bl[53] br[53] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_54 bl[54] br[54] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_55 bl[55] br[55] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_56 bl[56] br[56] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_57 bl[57] br[57] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_58 bl[58] br[58] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_59 bl[59] br[59] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_60 bl[60] br[60] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_61 bl[61] br[61] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_62 bl[62] br[62] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_185_63 bl[63] br[63] vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xcell_186_0 bl[0] br[0] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_1 bl[1] br[1] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_2 bl[2] br[2] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_3 bl[3] br[3] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_4 bl[4] br[4] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_5 bl[5] br[5] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_6 bl[6] br[6] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_7 bl[7] br[7] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_8 bl[8] br[8] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_9 bl[9] br[9] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_10 bl[10] br[10] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_11 bl[11] br[11] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_12 bl[12] br[12] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_13 bl[13] br[13] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_14 bl[14] br[14] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_15 bl[15] br[15] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_16 bl[16] br[16] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_17 bl[17] br[17] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_18 bl[18] br[18] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_19 bl[19] br[19] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_20 bl[20] br[20] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_21 bl[21] br[21] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_22 bl[22] br[22] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_23 bl[23] br[23] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_24 bl[24] br[24] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_25 bl[25] br[25] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_26 bl[26] br[26] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_27 bl[27] br[27] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_28 bl[28] br[28] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_29 bl[29] br[29] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_30 bl[30] br[30] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_31 bl[31] br[31] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_32 bl[32] br[32] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_33 bl[33] br[33] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_34 bl[34] br[34] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_35 bl[35] br[35] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_36 bl[36] br[36] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_37 bl[37] br[37] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_38 bl[38] br[38] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_39 bl[39] br[39] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_40 bl[40] br[40] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_41 bl[41] br[41] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_42 bl[42] br[42] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_43 bl[43] br[43] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_44 bl[44] br[44] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_45 bl[45] br[45] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_46 bl[46] br[46] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_47 bl[47] br[47] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_48 bl[48] br[48] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_49 bl[49] br[49] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_50 bl[50] br[50] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_51 bl[51] br[51] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_52 bl[52] br[52] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_53 bl[53] br[53] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_54 bl[54] br[54] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_55 bl[55] br[55] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_56 bl[56] br[56] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_57 bl[57] br[57] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_58 bl[58] br[58] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_59 bl[59] br[59] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_60 bl[60] br[60] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_61 bl[61] br[61] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_62 bl[62] br[62] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_186_63 bl[63] br[63] vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xcell_187_0 bl[0] br[0] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_1 bl[1] br[1] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_2 bl[2] br[2] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_3 bl[3] br[3] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_4 bl[4] br[4] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_5 bl[5] br[5] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_6 bl[6] br[6] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_7 bl[7] br[7] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_8 bl[8] br[8] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_9 bl[9] br[9] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_10 bl[10] br[10] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_11 bl[11] br[11] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_12 bl[12] br[12] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_13 bl[13] br[13] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_14 bl[14] br[14] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_15 bl[15] br[15] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_16 bl[16] br[16] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_17 bl[17] br[17] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_18 bl[18] br[18] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_19 bl[19] br[19] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_20 bl[20] br[20] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_21 bl[21] br[21] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_22 bl[22] br[22] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_23 bl[23] br[23] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_24 bl[24] br[24] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_25 bl[25] br[25] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_26 bl[26] br[26] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_27 bl[27] br[27] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_28 bl[28] br[28] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_29 bl[29] br[29] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_30 bl[30] br[30] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_31 bl[31] br[31] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_32 bl[32] br[32] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_33 bl[33] br[33] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_34 bl[34] br[34] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_35 bl[35] br[35] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_36 bl[36] br[36] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_37 bl[37] br[37] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_38 bl[38] br[38] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_39 bl[39] br[39] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_40 bl[40] br[40] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_41 bl[41] br[41] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_42 bl[42] br[42] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_43 bl[43] br[43] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_44 bl[44] br[44] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_45 bl[45] br[45] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_46 bl[46] br[46] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_47 bl[47] br[47] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_48 bl[48] br[48] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_49 bl[49] br[49] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_50 bl[50] br[50] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_51 bl[51] br[51] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_52 bl[52] br[52] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_53 bl[53] br[53] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_54 bl[54] br[54] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_55 bl[55] br[55] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_56 bl[56] br[56] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_57 bl[57] br[57] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_58 bl[58] br[58] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_59 bl[59] br[59] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_60 bl[60] br[60] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_61 bl[61] br[61] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_62 bl[62] br[62] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_187_63 bl[63] br[63] vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xcell_188_0 bl[0] br[0] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_1 bl[1] br[1] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_2 bl[2] br[2] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_3 bl[3] br[3] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_4 bl[4] br[4] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_5 bl[5] br[5] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_6 bl[6] br[6] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_7 bl[7] br[7] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_8 bl[8] br[8] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_9 bl[9] br[9] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_10 bl[10] br[10] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_11 bl[11] br[11] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_12 bl[12] br[12] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_13 bl[13] br[13] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_14 bl[14] br[14] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_15 bl[15] br[15] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_16 bl[16] br[16] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_17 bl[17] br[17] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_18 bl[18] br[18] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_19 bl[19] br[19] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_20 bl[20] br[20] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_21 bl[21] br[21] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_22 bl[22] br[22] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_23 bl[23] br[23] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_24 bl[24] br[24] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_25 bl[25] br[25] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_26 bl[26] br[26] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_27 bl[27] br[27] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_28 bl[28] br[28] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_29 bl[29] br[29] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_30 bl[30] br[30] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_31 bl[31] br[31] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_32 bl[32] br[32] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_33 bl[33] br[33] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_34 bl[34] br[34] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_35 bl[35] br[35] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_36 bl[36] br[36] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_37 bl[37] br[37] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_38 bl[38] br[38] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_39 bl[39] br[39] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_40 bl[40] br[40] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_41 bl[41] br[41] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_42 bl[42] br[42] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_43 bl[43] br[43] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_44 bl[44] br[44] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_45 bl[45] br[45] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_46 bl[46] br[46] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_47 bl[47] br[47] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_48 bl[48] br[48] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_49 bl[49] br[49] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_50 bl[50] br[50] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_51 bl[51] br[51] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_52 bl[52] br[52] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_53 bl[53] br[53] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_54 bl[54] br[54] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_55 bl[55] br[55] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_56 bl[56] br[56] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_57 bl[57] br[57] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_58 bl[58] br[58] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_59 bl[59] br[59] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_60 bl[60] br[60] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_61 bl[61] br[61] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_62 bl[62] br[62] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_188_63 bl[63] br[63] vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xcell_189_0 bl[0] br[0] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_1 bl[1] br[1] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_2 bl[2] br[2] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_3 bl[3] br[3] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_4 bl[4] br[4] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_5 bl[5] br[5] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_6 bl[6] br[6] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_7 bl[7] br[7] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_8 bl[8] br[8] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_9 bl[9] br[9] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_10 bl[10] br[10] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_11 bl[11] br[11] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_12 bl[12] br[12] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_13 bl[13] br[13] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_14 bl[14] br[14] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_15 bl[15] br[15] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_16 bl[16] br[16] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_17 bl[17] br[17] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_18 bl[18] br[18] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_19 bl[19] br[19] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_20 bl[20] br[20] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_21 bl[21] br[21] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_22 bl[22] br[22] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_23 bl[23] br[23] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_24 bl[24] br[24] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_25 bl[25] br[25] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_26 bl[26] br[26] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_27 bl[27] br[27] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_28 bl[28] br[28] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_29 bl[29] br[29] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_30 bl[30] br[30] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_31 bl[31] br[31] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_32 bl[32] br[32] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_33 bl[33] br[33] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_34 bl[34] br[34] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_35 bl[35] br[35] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_36 bl[36] br[36] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_37 bl[37] br[37] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_38 bl[38] br[38] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_39 bl[39] br[39] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_40 bl[40] br[40] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_41 bl[41] br[41] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_42 bl[42] br[42] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_43 bl[43] br[43] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_44 bl[44] br[44] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_45 bl[45] br[45] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_46 bl[46] br[46] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_47 bl[47] br[47] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_48 bl[48] br[48] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_49 bl[49] br[49] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_50 bl[50] br[50] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_51 bl[51] br[51] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_52 bl[52] br[52] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_53 bl[53] br[53] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_54 bl[54] br[54] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_55 bl[55] br[55] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_56 bl[56] br[56] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_57 bl[57] br[57] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_58 bl[58] br[58] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_59 bl[59] br[59] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_60 bl[60] br[60] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_61 bl[61] br[61] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_62 bl[62] br[62] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_189_63 bl[63] br[63] vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xcell_190_0 bl[0] br[0] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_1 bl[1] br[1] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_2 bl[2] br[2] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_3 bl[3] br[3] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_4 bl[4] br[4] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_5 bl[5] br[5] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_6 bl[6] br[6] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_7 bl[7] br[7] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_8 bl[8] br[8] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_9 bl[9] br[9] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_10 bl[10] br[10] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_11 bl[11] br[11] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_12 bl[12] br[12] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_13 bl[13] br[13] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_14 bl[14] br[14] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_15 bl[15] br[15] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_16 bl[16] br[16] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_17 bl[17] br[17] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_18 bl[18] br[18] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_19 bl[19] br[19] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_20 bl[20] br[20] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_21 bl[21] br[21] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_22 bl[22] br[22] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_23 bl[23] br[23] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_24 bl[24] br[24] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_25 bl[25] br[25] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_26 bl[26] br[26] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_27 bl[27] br[27] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_28 bl[28] br[28] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_29 bl[29] br[29] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_30 bl[30] br[30] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_31 bl[31] br[31] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_32 bl[32] br[32] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_33 bl[33] br[33] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_34 bl[34] br[34] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_35 bl[35] br[35] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_36 bl[36] br[36] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_37 bl[37] br[37] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_38 bl[38] br[38] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_39 bl[39] br[39] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_40 bl[40] br[40] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_41 bl[41] br[41] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_42 bl[42] br[42] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_43 bl[43] br[43] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_44 bl[44] br[44] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_45 bl[45] br[45] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_46 bl[46] br[46] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_47 bl[47] br[47] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_48 bl[48] br[48] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_49 bl[49] br[49] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_50 bl[50] br[50] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_51 bl[51] br[51] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_52 bl[52] br[52] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_53 bl[53] br[53] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_54 bl[54] br[54] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_55 bl[55] br[55] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_56 bl[56] br[56] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_57 bl[57] br[57] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_58 bl[58] br[58] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_59 bl[59] br[59] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_60 bl[60] br[60] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_61 bl[61] br[61] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_62 bl[62] br[62] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_190_63 bl[63] br[63] vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xcell_191_0 bl[0] br[0] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_1 bl[1] br[1] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_2 bl[2] br[2] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_3 bl[3] br[3] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_4 bl[4] br[4] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_5 bl[5] br[5] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_6 bl[6] br[6] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_7 bl[7] br[7] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_8 bl[8] br[8] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_9 bl[9] br[9] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_10 bl[10] br[10] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_11 bl[11] br[11] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_12 bl[12] br[12] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_13 bl[13] br[13] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_14 bl[14] br[14] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_15 bl[15] br[15] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_16 bl[16] br[16] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_17 bl[17] br[17] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_18 bl[18] br[18] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_19 bl[19] br[19] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_20 bl[20] br[20] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_21 bl[21] br[21] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_22 bl[22] br[22] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_23 bl[23] br[23] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_24 bl[24] br[24] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_25 bl[25] br[25] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_26 bl[26] br[26] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_27 bl[27] br[27] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_28 bl[28] br[28] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_29 bl[29] br[29] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_30 bl[30] br[30] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_31 bl[31] br[31] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_32 bl[32] br[32] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_33 bl[33] br[33] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_34 bl[34] br[34] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_35 bl[35] br[35] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_36 bl[36] br[36] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_37 bl[37] br[37] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_38 bl[38] br[38] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_39 bl[39] br[39] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_40 bl[40] br[40] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_41 bl[41] br[41] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_42 bl[42] br[42] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_43 bl[43] br[43] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_44 bl[44] br[44] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_45 bl[45] br[45] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_46 bl[46] br[46] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_47 bl[47] br[47] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_48 bl[48] br[48] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_49 bl[49] br[49] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_50 bl[50] br[50] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_51 bl[51] br[51] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_52 bl[52] br[52] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_53 bl[53] br[53] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_54 bl[54] br[54] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_55 bl[55] br[55] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_56 bl[56] br[56] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_57 bl[57] br[57] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_58 bl[58] br[58] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_59 bl[59] br[59] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_60 bl[60] br[60] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_61 bl[61] br[61] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_62 bl[62] br[62] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_191_63 bl[63] br[63] vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xcell_192_0 bl[0] br[0] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_1 bl[1] br[1] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_2 bl[2] br[2] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_3 bl[3] br[3] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_4 bl[4] br[4] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_5 bl[5] br[5] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_6 bl[6] br[6] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_7 bl[7] br[7] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_8 bl[8] br[8] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_9 bl[9] br[9] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_10 bl[10] br[10] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_11 bl[11] br[11] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_12 bl[12] br[12] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_13 bl[13] br[13] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_14 bl[14] br[14] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_15 bl[15] br[15] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_16 bl[16] br[16] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_17 bl[17] br[17] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_18 bl[18] br[18] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_19 bl[19] br[19] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_20 bl[20] br[20] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_21 bl[21] br[21] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_22 bl[22] br[22] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_23 bl[23] br[23] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_24 bl[24] br[24] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_25 bl[25] br[25] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_26 bl[26] br[26] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_27 bl[27] br[27] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_28 bl[28] br[28] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_29 bl[29] br[29] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_30 bl[30] br[30] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_31 bl[31] br[31] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_32 bl[32] br[32] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_33 bl[33] br[33] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_34 bl[34] br[34] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_35 bl[35] br[35] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_36 bl[36] br[36] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_37 bl[37] br[37] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_38 bl[38] br[38] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_39 bl[39] br[39] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_40 bl[40] br[40] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_41 bl[41] br[41] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_42 bl[42] br[42] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_43 bl[43] br[43] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_44 bl[44] br[44] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_45 bl[45] br[45] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_46 bl[46] br[46] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_47 bl[47] br[47] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_48 bl[48] br[48] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_49 bl[49] br[49] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_50 bl[50] br[50] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_51 bl[51] br[51] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_52 bl[52] br[52] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_53 bl[53] br[53] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_54 bl[54] br[54] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_55 bl[55] br[55] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_56 bl[56] br[56] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_57 bl[57] br[57] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_58 bl[58] br[58] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_59 bl[59] br[59] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_60 bl[60] br[60] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_61 bl[61] br[61] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_62 bl[62] br[62] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_192_63 bl[63] br[63] vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xcell_193_0 bl[0] br[0] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_1 bl[1] br[1] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_2 bl[2] br[2] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_3 bl[3] br[3] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_4 bl[4] br[4] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_5 bl[5] br[5] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_6 bl[6] br[6] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_7 bl[7] br[7] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_8 bl[8] br[8] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_9 bl[9] br[9] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_10 bl[10] br[10] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_11 bl[11] br[11] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_12 bl[12] br[12] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_13 bl[13] br[13] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_14 bl[14] br[14] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_15 bl[15] br[15] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_16 bl[16] br[16] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_17 bl[17] br[17] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_18 bl[18] br[18] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_19 bl[19] br[19] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_20 bl[20] br[20] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_21 bl[21] br[21] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_22 bl[22] br[22] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_23 bl[23] br[23] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_24 bl[24] br[24] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_25 bl[25] br[25] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_26 bl[26] br[26] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_27 bl[27] br[27] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_28 bl[28] br[28] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_29 bl[29] br[29] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_30 bl[30] br[30] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_31 bl[31] br[31] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_32 bl[32] br[32] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_33 bl[33] br[33] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_34 bl[34] br[34] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_35 bl[35] br[35] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_36 bl[36] br[36] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_37 bl[37] br[37] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_38 bl[38] br[38] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_39 bl[39] br[39] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_40 bl[40] br[40] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_41 bl[41] br[41] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_42 bl[42] br[42] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_43 bl[43] br[43] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_44 bl[44] br[44] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_45 bl[45] br[45] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_46 bl[46] br[46] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_47 bl[47] br[47] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_48 bl[48] br[48] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_49 bl[49] br[49] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_50 bl[50] br[50] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_51 bl[51] br[51] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_52 bl[52] br[52] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_53 bl[53] br[53] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_54 bl[54] br[54] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_55 bl[55] br[55] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_56 bl[56] br[56] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_57 bl[57] br[57] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_58 bl[58] br[58] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_59 bl[59] br[59] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_60 bl[60] br[60] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_61 bl[61] br[61] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_62 bl[62] br[62] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_193_63 bl[63] br[63] vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xcell_194_0 bl[0] br[0] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_1 bl[1] br[1] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_2 bl[2] br[2] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_3 bl[3] br[3] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_4 bl[4] br[4] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_5 bl[5] br[5] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_6 bl[6] br[6] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_7 bl[7] br[7] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_8 bl[8] br[8] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_9 bl[9] br[9] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_10 bl[10] br[10] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_11 bl[11] br[11] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_12 bl[12] br[12] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_13 bl[13] br[13] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_14 bl[14] br[14] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_15 bl[15] br[15] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_16 bl[16] br[16] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_17 bl[17] br[17] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_18 bl[18] br[18] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_19 bl[19] br[19] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_20 bl[20] br[20] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_21 bl[21] br[21] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_22 bl[22] br[22] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_23 bl[23] br[23] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_24 bl[24] br[24] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_25 bl[25] br[25] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_26 bl[26] br[26] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_27 bl[27] br[27] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_28 bl[28] br[28] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_29 bl[29] br[29] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_30 bl[30] br[30] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_31 bl[31] br[31] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_32 bl[32] br[32] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_33 bl[33] br[33] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_34 bl[34] br[34] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_35 bl[35] br[35] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_36 bl[36] br[36] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_37 bl[37] br[37] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_38 bl[38] br[38] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_39 bl[39] br[39] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_40 bl[40] br[40] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_41 bl[41] br[41] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_42 bl[42] br[42] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_43 bl[43] br[43] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_44 bl[44] br[44] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_45 bl[45] br[45] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_46 bl[46] br[46] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_47 bl[47] br[47] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_48 bl[48] br[48] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_49 bl[49] br[49] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_50 bl[50] br[50] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_51 bl[51] br[51] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_52 bl[52] br[52] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_53 bl[53] br[53] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_54 bl[54] br[54] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_55 bl[55] br[55] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_56 bl[56] br[56] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_57 bl[57] br[57] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_58 bl[58] br[58] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_59 bl[59] br[59] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_60 bl[60] br[60] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_61 bl[61] br[61] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_62 bl[62] br[62] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_194_63 bl[63] br[63] vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xcell_195_0 bl[0] br[0] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_1 bl[1] br[1] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_2 bl[2] br[2] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_3 bl[3] br[3] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_4 bl[4] br[4] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_5 bl[5] br[5] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_6 bl[6] br[6] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_7 bl[7] br[7] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_8 bl[8] br[8] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_9 bl[9] br[9] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_10 bl[10] br[10] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_11 bl[11] br[11] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_12 bl[12] br[12] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_13 bl[13] br[13] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_14 bl[14] br[14] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_15 bl[15] br[15] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_16 bl[16] br[16] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_17 bl[17] br[17] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_18 bl[18] br[18] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_19 bl[19] br[19] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_20 bl[20] br[20] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_21 bl[21] br[21] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_22 bl[22] br[22] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_23 bl[23] br[23] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_24 bl[24] br[24] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_25 bl[25] br[25] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_26 bl[26] br[26] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_27 bl[27] br[27] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_28 bl[28] br[28] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_29 bl[29] br[29] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_30 bl[30] br[30] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_31 bl[31] br[31] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_32 bl[32] br[32] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_33 bl[33] br[33] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_34 bl[34] br[34] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_35 bl[35] br[35] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_36 bl[36] br[36] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_37 bl[37] br[37] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_38 bl[38] br[38] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_39 bl[39] br[39] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_40 bl[40] br[40] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_41 bl[41] br[41] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_42 bl[42] br[42] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_43 bl[43] br[43] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_44 bl[44] br[44] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_45 bl[45] br[45] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_46 bl[46] br[46] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_47 bl[47] br[47] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_48 bl[48] br[48] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_49 bl[49] br[49] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_50 bl[50] br[50] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_51 bl[51] br[51] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_52 bl[52] br[52] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_53 bl[53] br[53] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_54 bl[54] br[54] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_55 bl[55] br[55] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_56 bl[56] br[56] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_57 bl[57] br[57] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_58 bl[58] br[58] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_59 bl[59] br[59] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_60 bl[60] br[60] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_61 bl[61] br[61] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_62 bl[62] br[62] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_195_63 bl[63] br[63] vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xcell_196_0 bl[0] br[0] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_1 bl[1] br[1] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_2 bl[2] br[2] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_3 bl[3] br[3] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_4 bl[4] br[4] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_5 bl[5] br[5] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_6 bl[6] br[6] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_7 bl[7] br[7] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_8 bl[8] br[8] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_9 bl[9] br[9] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_10 bl[10] br[10] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_11 bl[11] br[11] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_12 bl[12] br[12] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_13 bl[13] br[13] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_14 bl[14] br[14] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_15 bl[15] br[15] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_16 bl[16] br[16] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_17 bl[17] br[17] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_18 bl[18] br[18] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_19 bl[19] br[19] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_20 bl[20] br[20] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_21 bl[21] br[21] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_22 bl[22] br[22] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_23 bl[23] br[23] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_24 bl[24] br[24] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_25 bl[25] br[25] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_26 bl[26] br[26] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_27 bl[27] br[27] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_28 bl[28] br[28] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_29 bl[29] br[29] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_30 bl[30] br[30] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_31 bl[31] br[31] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_32 bl[32] br[32] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_33 bl[33] br[33] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_34 bl[34] br[34] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_35 bl[35] br[35] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_36 bl[36] br[36] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_37 bl[37] br[37] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_38 bl[38] br[38] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_39 bl[39] br[39] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_40 bl[40] br[40] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_41 bl[41] br[41] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_42 bl[42] br[42] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_43 bl[43] br[43] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_44 bl[44] br[44] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_45 bl[45] br[45] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_46 bl[46] br[46] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_47 bl[47] br[47] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_48 bl[48] br[48] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_49 bl[49] br[49] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_50 bl[50] br[50] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_51 bl[51] br[51] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_52 bl[52] br[52] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_53 bl[53] br[53] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_54 bl[54] br[54] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_55 bl[55] br[55] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_56 bl[56] br[56] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_57 bl[57] br[57] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_58 bl[58] br[58] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_59 bl[59] br[59] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_60 bl[60] br[60] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_61 bl[61] br[61] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_62 bl[62] br[62] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_196_63 bl[63] br[63] vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xcell_197_0 bl[0] br[0] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_1 bl[1] br[1] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_2 bl[2] br[2] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_3 bl[3] br[3] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_4 bl[4] br[4] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_5 bl[5] br[5] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_6 bl[6] br[6] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_7 bl[7] br[7] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_8 bl[8] br[8] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_9 bl[9] br[9] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_10 bl[10] br[10] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_11 bl[11] br[11] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_12 bl[12] br[12] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_13 bl[13] br[13] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_14 bl[14] br[14] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_15 bl[15] br[15] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_16 bl[16] br[16] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_17 bl[17] br[17] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_18 bl[18] br[18] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_19 bl[19] br[19] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_20 bl[20] br[20] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_21 bl[21] br[21] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_22 bl[22] br[22] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_23 bl[23] br[23] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_24 bl[24] br[24] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_25 bl[25] br[25] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_26 bl[26] br[26] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_27 bl[27] br[27] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_28 bl[28] br[28] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_29 bl[29] br[29] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_30 bl[30] br[30] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_31 bl[31] br[31] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_32 bl[32] br[32] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_33 bl[33] br[33] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_34 bl[34] br[34] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_35 bl[35] br[35] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_36 bl[36] br[36] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_37 bl[37] br[37] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_38 bl[38] br[38] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_39 bl[39] br[39] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_40 bl[40] br[40] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_41 bl[41] br[41] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_42 bl[42] br[42] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_43 bl[43] br[43] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_44 bl[44] br[44] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_45 bl[45] br[45] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_46 bl[46] br[46] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_47 bl[47] br[47] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_48 bl[48] br[48] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_49 bl[49] br[49] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_50 bl[50] br[50] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_51 bl[51] br[51] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_52 bl[52] br[52] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_53 bl[53] br[53] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_54 bl[54] br[54] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_55 bl[55] br[55] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_56 bl[56] br[56] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_57 bl[57] br[57] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_58 bl[58] br[58] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_59 bl[59] br[59] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_60 bl[60] br[60] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_61 bl[61] br[61] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_62 bl[62] br[62] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_197_63 bl[63] br[63] vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xcell_198_0 bl[0] br[0] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_1 bl[1] br[1] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_2 bl[2] br[2] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_3 bl[3] br[3] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_4 bl[4] br[4] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_5 bl[5] br[5] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_6 bl[6] br[6] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_7 bl[7] br[7] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_8 bl[8] br[8] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_9 bl[9] br[9] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_10 bl[10] br[10] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_11 bl[11] br[11] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_12 bl[12] br[12] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_13 bl[13] br[13] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_14 bl[14] br[14] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_15 bl[15] br[15] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_16 bl[16] br[16] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_17 bl[17] br[17] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_18 bl[18] br[18] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_19 bl[19] br[19] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_20 bl[20] br[20] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_21 bl[21] br[21] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_22 bl[22] br[22] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_23 bl[23] br[23] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_24 bl[24] br[24] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_25 bl[25] br[25] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_26 bl[26] br[26] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_27 bl[27] br[27] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_28 bl[28] br[28] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_29 bl[29] br[29] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_30 bl[30] br[30] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_31 bl[31] br[31] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_32 bl[32] br[32] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_33 bl[33] br[33] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_34 bl[34] br[34] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_35 bl[35] br[35] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_36 bl[36] br[36] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_37 bl[37] br[37] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_38 bl[38] br[38] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_39 bl[39] br[39] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_40 bl[40] br[40] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_41 bl[41] br[41] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_42 bl[42] br[42] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_43 bl[43] br[43] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_44 bl[44] br[44] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_45 bl[45] br[45] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_46 bl[46] br[46] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_47 bl[47] br[47] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_48 bl[48] br[48] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_49 bl[49] br[49] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_50 bl[50] br[50] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_51 bl[51] br[51] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_52 bl[52] br[52] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_53 bl[53] br[53] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_54 bl[54] br[54] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_55 bl[55] br[55] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_56 bl[56] br[56] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_57 bl[57] br[57] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_58 bl[58] br[58] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_59 bl[59] br[59] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_60 bl[60] br[60] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_61 bl[61] br[61] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_62 bl[62] br[62] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_198_63 bl[63] br[63] vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xcell_199_0 bl[0] br[0] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_1 bl[1] br[1] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_2 bl[2] br[2] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_3 bl[3] br[3] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_4 bl[4] br[4] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_5 bl[5] br[5] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_6 bl[6] br[6] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_7 bl[7] br[7] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_8 bl[8] br[8] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_9 bl[9] br[9] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_10 bl[10] br[10] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_11 bl[11] br[11] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_12 bl[12] br[12] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_13 bl[13] br[13] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_14 bl[14] br[14] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_15 bl[15] br[15] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_16 bl[16] br[16] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_17 bl[17] br[17] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_18 bl[18] br[18] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_19 bl[19] br[19] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_20 bl[20] br[20] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_21 bl[21] br[21] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_22 bl[22] br[22] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_23 bl[23] br[23] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_24 bl[24] br[24] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_25 bl[25] br[25] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_26 bl[26] br[26] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_27 bl[27] br[27] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_28 bl[28] br[28] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_29 bl[29] br[29] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_30 bl[30] br[30] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_31 bl[31] br[31] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_32 bl[32] br[32] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_33 bl[33] br[33] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_34 bl[34] br[34] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_35 bl[35] br[35] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_36 bl[36] br[36] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_37 bl[37] br[37] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_38 bl[38] br[38] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_39 bl[39] br[39] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_40 bl[40] br[40] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_41 bl[41] br[41] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_42 bl[42] br[42] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_43 bl[43] br[43] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_44 bl[44] br[44] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_45 bl[45] br[45] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_46 bl[46] br[46] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_47 bl[47] br[47] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_48 bl[48] br[48] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_49 bl[49] br[49] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_50 bl[50] br[50] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_51 bl[51] br[51] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_52 bl[52] br[52] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_53 bl[53] br[53] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_54 bl[54] br[54] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_55 bl[55] br[55] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_56 bl[56] br[56] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_57 bl[57] br[57] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_58 bl[58] br[58] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_59 bl[59] br[59] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_60 bl[60] br[60] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_61 bl[61] br[61] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_62 bl[62] br[62] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_199_63 bl[63] br[63] vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xcell_200_0 bl[0] br[0] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_1 bl[1] br[1] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_2 bl[2] br[2] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_3 bl[3] br[3] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_4 bl[4] br[4] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_5 bl[5] br[5] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_6 bl[6] br[6] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_7 bl[7] br[7] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_8 bl[8] br[8] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_9 bl[9] br[9] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_10 bl[10] br[10] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_11 bl[11] br[11] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_12 bl[12] br[12] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_13 bl[13] br[13] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_14 bl[14] br[14] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_15 bl[15] br[15] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_16 bl[16] br[16] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_17 bl[17] br[17] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_18 bl[18] br[18] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_19 bl[19] br[19] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_20 bl[20] br[20] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_21 bl[21] br[21] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_22 bl[22] br[22] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_23 bl[23] br[23] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_24 bl[24] br[24] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_25 bl[25] br[25] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_26 bl[26] br[26] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_27 bl[27] br[27] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_28 bl[28] br[28] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_29 bl[29] br[29] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_30 bl[30] br[30] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_31 bl[31] br[31] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_32 bl[32] br[32] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_33 bl[33] br[33] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_34 bl[34] br[34] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_35 bl[35] br[35] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_36 bl[36] br[36] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_37 bl[37] br[37] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_38 bl[38] br[38] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_39 bl[39] br[39] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_40 bl[40] br[40] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_41 bl[41] br[41] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_42 bl[42] br[42] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_43 bl[43] br[43] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_44 bl[44] br[44] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_45 bl[45] br[45] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_46 bl[46] br[46] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_47 bl[47] br[47] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_48 bl[48] br[48] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_49 bl[49] br[49] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_50 bl[50] br[50] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_51 bl[51] br[51] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_52 bl[52] br[52] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_53 bl[53] br[53] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_54 bl[54] br[54] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_55 bl[55] br[55] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_56 bl[56] br[56] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_57 bl[57] br[57] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_58 bl[58] br[58] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_59 bl[59] br[59] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_60 bl[60] br[60] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_61 bl[61] br[61] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_62 bl[62] br[62] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_200_63 bl[63] br[63] vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xcell_201_0 bl[0] br[0] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_1 bl[1] br[1] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_2 bl[2] br[2] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_3 bl[3] br[3] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_4 bl[4] br[4] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_5 bl[5] br[5] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_6 bl[6] br[6] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_7 bl[7] br[7] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_8 bl[8] br[8] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_9 bl[9] br[9] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_10 bl[10] br[10] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_11 bl[11] br[11] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_12 bl[12] br[12] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_13 bl[13] br[13] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_14 bl[14] br[14] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_15 bl[15] br[15] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_16 bl[16] br[16] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_17 bl[17] br[17] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_18 bl[18] br[18] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_19 bl[19] br[19] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_20 bl[20] br[20] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_21 bl[21] br[21] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_22 bl[22] br[22] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_23 bl[23] br[23] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_24 bl[24] br[24] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_25 bl[25] br[25] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_26 bl[26] br[26] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_27 bl[27] br[27] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_28 bl[28] br[28] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_29 bl[29] br[29] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_30 bl[30] br[30] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_31 bl[31] br[31] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_32 bl[32] br[32] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_33 bl[33] br[33] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_34 bl[34] br[34] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_35 bl[35] br[35] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_36 bl[36] br[36] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_37 bl[37] br[37] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_38 bl[38] br[38] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_39 bl[39] br[39] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_40 bl[40] br[40] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_41 bl[41] br[41] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_42 bl[42] br[42] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_43 bl[43] br[43] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_44 bl[44] br[44] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_45 bl[45] br[45] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_46 bl[46] br[46] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_47 bl[47] br[47] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_48 bl[48] br[48] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_49 bl[49] br[49] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_50 bl[50] br[50] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_51 bl[51] br[51] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_52 bl[52] br[52] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_53 bl[53] br[53] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_54 bl[54] br[54] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_55 bl[55] br[55] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_56 bl[56] br[56] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_57 bl[57] br[57] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_58 bl[58] br[58] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_59 bl[59] br[59] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_60 bl[60] br[60] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_61 bl[61] br[61] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_62 bl[62] br[62] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_201_63 bl[63] br[63] vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xcell_202_0 bl[0] br[0] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_1 bl[1] br[1] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_2 bl[2] br[2] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_3 bl[3] br[3] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_4 bl[4] br[4] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_5 bl[5] br[5] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_6 bl[6] br[6] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_7 bl[7] br[7] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_8 bl[8] br[8] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_9 bl[9] br[9] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_10 bl[10] br[10] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_11 bl[11] br[11] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_12 bl[12] br[12] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_13 bl[13] br[13] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_14 bl[14] br[14] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_15 bl[15] br[15] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_16 bl[16] br[16] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_17 bl[17] br[17] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_18 bl[18] br[18] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_19 bl[19] br[19] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_20 bl[20] br[20] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_21 bl[21] br[21] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_22 bl[22] br[22] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_23 bl[23] br[23] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_24 bl[24] br[24] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_25 bl[25] br[25] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_26 bl[26] br[26] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_27 bl[27] br[27] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_28 bl[28] br[28] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_29 bl[29] br[29] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_30 bl[30] br[30] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_31 bl[31] br[31] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_32 bl[32] br[32] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_33 bl[33] br[33] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_34 bl[34] br[34] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_35 bl[35] br[35] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_36 bl[36] br[36] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_37 bl[37] br[37] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_38 bl[38] br[38] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_39 bl[39] br[39] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_40 bl[40] br[40] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_41 bl[41] br[41] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_42 bl[42] br[42] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_43 bl[43] br[43] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_44 bl[44] br[44] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_45 bl[45] br[45] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_46 bl[46] br[46] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_47 bl[47] br[47] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_48 bl[48] br[48] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_49 bl[49] br[49] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_50 bl[50] br[50] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_51 bl[51] br[51] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_52 bl[52] br[52] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_53 bl[53] br[53] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_54 bl[54] br[54] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_55 bl[55] br[55] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_56 bl[56] br[56] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_57 bl[57] br[57] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_58 bl[58] br[58] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_59 bl[59] br[59] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_60 bl[60] br[60] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_61 bl[61] br[61] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_62 bl[62] br[62] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_202_63 bl[63] br[63] vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xcell_203_0 bl[0] br[0] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_1 bl[1] br[1] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_2 bl[2] br[2] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_3 bl[3] br[3] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_4 bl[4] br[4] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_5 bl[5] br[5] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_6 bl[6] br[6] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_7 bl[7] br[7] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_8 bl[8] br[8] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_9 bl[9] br[9] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_10 bl[10] br[10] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_11 bl[11] br[11] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_12 bl[12] br[12] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_13 bl[13] br[13] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_14 bl[14] br[14] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_15 bl[15] br[15] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_16 bl[16] br[16] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_17 bl[17] br[17] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_18 bl[18] br[18] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_19 bl[19] br[19] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_20 bl[20] br[20] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_21 bl[21] br[21] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_22 bl[22] br[22] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_23 bl[23] br[23] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_24 bl[24] br[24] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_25 bl[25] br[25] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_26 bl[26] br[26] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_27 bl[27] br[27] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_28 bl[28] br[28] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_29 bl[29] br[29] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_30 bl[30] br[30] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_31 bl[31] br[31] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_32 bl[32] br[32] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_33 bl[33] br[33] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_34 bl[34] br[34] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_35 bl[35] br[35] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_36 bl[36] br[36] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_37 bl[37] br[37] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_38 bl[38] br[38] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_39 bl[39] br[39] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_40 bl[40] br[40] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_41 bl[41] br[41] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_42 bl[42] br[42] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_43 bl[43] br[43] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_44 bl[44] br[44] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_45 bl[45] br[45] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_46 bl[46] br[46] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_47 bl[47] br[47] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_48 bl[48] br[48] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_49 bl[49] br[49] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_50 bl[50] br[50] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_51 bl[51] br[51] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_52 bl[52] br[52] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_53 bl[53] br[53] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_54 bl[54] br[54] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_55 bl[55] br[55] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_56 bl[56] br[56] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_57 bl[57] br[57] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_58 bl[58] br[58] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_59 bl[59] br[59] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_60 bl[60] br[60] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_61 bl[61] br[61] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_62 bl[62] br[62] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_203_63 bl[63] br[63] vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xcell_204_0 bl[0] br[0] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_1 bl[1] br[1] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_2 bl[2] br[2] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_3 bl[3] br[3] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_4 bl[4] br[4] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_5 bl[5] br[5] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_6 bl[6] br[6] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_7 bl[7] br[7] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_8 bl[8] br[8] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_9 bl[9] br[9] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_10 bl[10] br[10] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_11 bl[11] br[11] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_12 bl[12] br[12] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_13 bl[13] br[13] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_14 bl[14] br[14] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_15 bl[15] br[15] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_16 bl[16] br[16] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_17 bl[17] br[17] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_18 bl[18] br[18] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_19 bl[19] br[19] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_20 bl[20] br[20] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_21 bl[21] br[21] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_22 bl[22] br[22] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_23 bl[23] br[23] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_24 bl[24] br[24] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_25 bl[25] br[25] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_26 bl[26] br[26] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_27 bl[27] br[27] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_28 bl[28] br[28] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_29 bl[29] br[29] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_30 bl[30] br[30] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_31 bl[31] br[31] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_32 bl[32] br[32] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_33 bl[33] br[33] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_34 bl[34] br[34] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_35 bl[35] br[35] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_36 bl[36] br[36] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_37 bl[37] br[37] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_38 bl[38] br[38] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_39 bl[39] br[39] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_40 bl[40] br[40] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_41 bl[41] br[41] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_42 bl[42] br[42] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_43 bl[43] br[43] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_44 bl[44] br[44] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_45 bl[45] br[45] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_46 bl[46] br[46] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_47 bl[47] br[47] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_48 bl[48] br[48] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_49 bl[49] br[49] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_50 bl[50] br[50] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_51 bl[51] br[51] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_52 bl[52] br[52] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_53 bl[53] br[53] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_54 bl[54] br[54] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_55 bl[55] br[55] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_56 bl[56] br[56] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_57 bl[57] br[57] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_58 bl[58] br[58] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_59 bl[59] br[59] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_60 bl[60] br[60] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_61 bl[61] br[61] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_62 bl[62] br[62] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_204_63 bl[63] br[63] vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xcell_205_0 bl[0] br[0] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_1 bl[1] br[1] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_2 bl[2] br[2] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_3 bl[3] br[3] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_4 bl[4] br[4] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_5 bl[5] br[5] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_6 bl[6] br[6] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_7 bl[7] br[7] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_8 bl[8] br[8] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_9 bl[9] br[9] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_10 bl[10] br[10] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_11 bl[11] br[11] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_12 bl[12] br[12] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_13 bl[13] br[13] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_14 bl[14] br[14] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_15 bl[15] br[15] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_16 bl[16] br[16] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_17 bl[17] br[17] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_18 bl[18] br[18] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_19 bl[19] br[19] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_20 bl[20] br[20] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_21 bl[21] br[21] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_22 bl[22] br[22] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_23 bl[23] br[23] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_24 bl[24] br[24] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_25 bl[25] br[25] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_26 bl[26] br[26] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_27 bl[27] br[27] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_28 bl[28] br[28] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_29 bl[29] br[29] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_30 bl[30] br[30] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_31 bl[31] br[31] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_32 bl[32] br[32] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_33 bl[33] br[33] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_34 bl[34] br[34] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_35 bl[35] br[35] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_36 bl[36] br[36] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_37 bl[37] br[37] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_38 bl[38] br[38] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_39 bl[39] br[39] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_40 bl[40] br[40] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_41 bl[41] br[41] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_42 bl[42] br[42] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_43 bl[43] br[43] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_44 bl[44] br[44] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_45 bl[45] br[45] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_46 bl[46] br[46] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_47 bl[47] br[47] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_48 bl[48] br[48] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_49 bl[49] br[49] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_50 bl[50] br[50] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_51 bl[51] br[51] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_52 bl[52] br[52] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_53 bl[53] br[53] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_54 bl[54] br[54] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_55 bl[55] br[55] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_56 bl[56] br[56] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_57 bl[57] br[57] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_58 bl[58] br[58] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_59 bl[59] br[59] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_60 bl[60] br[60] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_61 bl[61] br[61] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_62 bl[62] br[62] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_205_63 bl[63] br[63] vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xcell_206_0 bl[0] br[0] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_1 bl[1] br[1] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_2 bl[2] br[2] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_3 bl[3] br[3] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_4 bl[4] br[4] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_5 bl[5] br[5] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_6 bl[6] br[6] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_7 bl[7] br[7] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_8 bl[8] br[8] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_9 bl[9] br[9] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_10 bl[10] br[10] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_11 bl[11] br[11] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_12 bl[12] br[12] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_13 bl[13] br[13] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_14 bl[14] br[14] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_15 bl[15] br[15] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_16 bl[16] br[16] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_17 bl[17] br[17] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_18 bl[18] br[18] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_19 bl[19] br[19] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_20 bl[20] br[20] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_21 bl[21] br[21] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_22 bl[22] br[22] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_23 bl[23] br[23] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_24 bl[24] br[24] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_25 bl[25] br[25] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_26 bl[26] br[26] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_27 bl[27] br[27] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_28 bl[28] br[28] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_29 bl[29] br[29] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_30 bl[30] br[30] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_31 bl[31] br[31] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_32 bl[32] br[32] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_33 bl[33] br[33] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_34 bl[34] br[34] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_35 bl[35] br[35] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_36 bl[36] br[36] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_37 bl[37] br[37] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_38 bl[38] br[38] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_39 bl[39] br[39] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_40 bl[40] br[40] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_41 bl[41] br[41] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_42 bl[42] br[42] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_43 bl[43] br[43] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_44 bl[44] br[44] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_45 bl[45] br[45] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_46 bl[46] br[46] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_47 bl[47] br[47] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_48 bl[48] br[48] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_49 bl[49] br[49] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_50 bl[50] br[50] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_51 bl[51] br[51] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_52 bl[52] br[52] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_53 bl[53] br[53] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_54 bl[54] br[54] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_55 bl[55] br[55] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_56 bl[56] br[56] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_57 bl[57] br[57] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_58 bl[58] br[58] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_59 bl[59] br[59] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_60 bl[60] br[60] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_61 bl[61] br[61] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_62 bl[62] br[62] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_206_63 bl[63] br[63] vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xcell_207_0 bl[0] br[0] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_1 bl[1] br[1] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_2 bl[2] br[2] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_3 bl[3] br[3] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_4 bl[4] br[4] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_5 bl[5] br[5] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_6 bl[6] br[6] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_7 bl[7] br[7] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_8 bl[8] br[8] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_9 bl[9] br[9] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_10 bl[10] br[10] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_11 bl[11] br[11] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_12 bl[12] br[12] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_13 bl[13] br[13] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_14 bl[14] br[14] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_15 bl[15] br[15] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_16 bl[16] br[16] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_17 bl[17] br[17] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_18 bl[18] br[18] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_19 bl[19] br[19] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_20 bl[20] br[20] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_21 bl[21] br[21] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_22 bl[22] br[22] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_23 bl[23] br[23] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_24 bl[24] br[24] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_25 bl[25] br[25] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_26 bl[26] br[26] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_27 bl[27] br[27] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_28 bl[28] br[28] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_29 bl[29] br[29] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_30 bl[30] br[30] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_31 bl[31] br[31] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_32 bl[32] br[32] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_33 bl[33] br[33] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_34 bl[34] br[34] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_35 bl[35] br[35] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_36 bl[36] br[36] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_37 bl[37] br[37] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_38 bl[38] br[38] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_39 bl[39] br[39] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_40 bl[40] br[40] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_41 bl[41] br[41] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_42 bl[42] br[42] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_43 bl[43] br[43] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_44 bl[44] br[44] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_45 bl[45] br[45] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_46 bl[46] br[46] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_47 bl[47] br[47] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_48 bl[48] br[48] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_49 bl[49] br[49] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_50 bl[50] br[50] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_51 bl[51] br[51] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_52 bl[52] br[52] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_53 bl[53] br[53] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_54 bl[54] br[54] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_55 bl[55] br[55] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_56 bl[56] br[56] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_57 bl[57] br[57] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_58 bl[58] br[58] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_59 bl[59] br[59] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_60 bl[60] br[60] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_61 bl[61] br[61] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_62 bl[62] br[62] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_207_63 bl[63] br[63] vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xcell_208_0 bl[0] br[0] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_1 bl[1] br[1] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_2 bl[2] br[2] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_3 bl[3] br[3] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_4 bl[4] br[4] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_5 bl[5] br[5] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_6 bl[6] br[6] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_7 bl[7] br[7] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_8 bl[8] br[8] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_9 bl[9] br[9] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_10 bl[10] br[10] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_11 bl[11] br[11] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_12 bl[12] br[12] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_13 bl[13] br[13] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_14 bl[14] br[14] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_15 bl[15] br[15] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_16 bl[16] br[16] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_17 bl[17] br[17] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_18 bl[18] br[18] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_19 bl[19] br[19] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_20 bl[20] br[20] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_21 bl[21] br[21] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_22 bl[22] br[22] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_23 bl[23] br[23] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_24 bl[24] br[24] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_25 bl[25] br[25] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_26 bl[26] br[26] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_27 bl[27] br[27] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_28 bl[28] br[28] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_29 bl[29] br[29] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_30 bl[30] br[30] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_31 bl[31] br[31] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_32 bl[32] br[32] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_33 bl[33] br[33] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_34 bl[34] br[34] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_35 bl[35] br[35] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_36 bl[36] br[36] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_37 bl[37] br[37] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_38 bl[38] br[38] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_39 bl[39] br[39] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_40 bl[40] br[40] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_41 bl[41] br[41] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_42 bl[42] br[42] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_43 bl[43] br[43] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_44 bl[44] br[44] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_45 bl[45] br[45] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_46 bl[46] br[46] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_47 bl[47] br[47] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_48 bl[48] br[48] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_49 bl[49] br[49] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_50 bl[50] br[50] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_51 bl[51] br[51] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_52 bl[52] br[52] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_53 bl[53] br[53] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_54 bl[54] br[54] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_55 bl[55] br[55] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_56 bl[56] br[56] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_57 bl[57] br[57] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_58 bl[58] br[58] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_59 bl[59] br[59] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_60 bl[60] br[60] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_61 bl[61] br[61] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_62 bl[62] br[62] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_208_63 bl[63] br[63] vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xcell_209_0 bl[0] br[0] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_1 bl[1] br[1] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_2 bl[2] br[2] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_3 bl[3] br[3] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_4 bl[4] br[4] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_5 bl[5] br[5] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_6 bl[6] br[6] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_7 bl[7] br[7] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_8 bl[8] br[8] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_9 bl[9] br[9] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_10 bl[10] br[10] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_11 bl[11] br[11] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_12 bl[12] br[12] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_13 bl[13] br[13] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_14 bl[14] br[14] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_15 bl[15] br[15] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_16 bl[16] br[16] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_17 bl[17] br[17] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_18 bl[18] br[18] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_19 bl[19] br[19] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_20 bl[20] br[20] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_21 bl[21] br[21] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_22 bl[22] br[22] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_23 bl[23] br[23] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_24 bl[24] br[24] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_25 bl[25] br[25] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_26 bl[26] br[26] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_27 bl[27] br[27] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_28 bl[28] br[28] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_29 bl[29] br[29] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_30 bl[30] br[30] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_31 bl[31] br[31] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_32 bl[32] br[32] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_33 bl[33] br[33] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_34 bl[34] br[34] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_35 bl[35] br[35] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_36 bl[36] br[36] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_37 bl[37] br[37] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_38 bl[38] br[38] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_39 bl[39] br[39] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_40 bl[40] br[40] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_41 bl[41] br[41] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_42 bl[42] br[42] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_43 bl[43] br[43] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_44 bl[44] br[44] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_45 bl[45] br[45] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_46 bl[46] br[46] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_47 bl[47] br[47] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_48 bl[48] br[48] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_49 bl[49] br[49] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_50 bl[50] br[50] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_51 bl[51] br[51] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_52 bl[52] br[52] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_53 bl[53] br[53] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_54 bl[54] br[54] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_55 bl[55] br[55] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_56 bl[56] br[56] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_57 bl[57] br[57] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_58 bl[58] br[58] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_59 bl[59] br[59] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_60 bl[60] br[60] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_61 bl[61] br[61] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_62 bl[62] br[62] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_209_63 bl[63] br[63] vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xcell_210_0 bl[0] br[0] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_1 bl[1] br[1] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_2 bl[2] br[2] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_3 bl[3] br[3] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_4 bl[4] br[4] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_5 bl[5] br[5] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_6 bl[6] br[6] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_7 bl[7] br[7] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_8 bl[8] br[8] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_9 bl[9] br[9] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_10 bl[10] br[10] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_11 bl[11] br[11] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_12 bl[12] br[12] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_13 bl[13] br[13] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_14 bl[14] br[14] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_15 bl[15] br[15] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_16 bl[16] br[16] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_17 bl[17] br[17] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_18 bl[18] br[18] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_19 bl[19] br[19] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_20 bl[20] br[20] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_21 bl[21] br[21] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_22 bl[22] br[22] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_23 bl[23] br[23] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_24 bl[24] br[24] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_25 bl[25] br[25] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_26 bl[26] br[26] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_27 bl[27] br[27] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_28 bl[28] br[28] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_29 bl[29] br[29] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_30 bl[30] br[30] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_31 bl[31] br[31] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_32 bl[32] br[32] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_33 bl[33] br[33] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_34 bl[34] br[34] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_35 bl[35] br[35] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_36 bl[36] br[36] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_37 bl[37] br[37] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_38 bl[38] br[38] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_39 bl[39] br[39] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_40 bl[40] br[40] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_41 bl[41] br[41] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_42 bl[42] br[42] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_43 bl[43] br[43] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_44 bl[44] br[44] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_45 bl[45] br[45] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_46 bl[46] br[46] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_47 bl[47] br[47] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_48 bl[48] br[48] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_49 bl[49] br[49] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_50 bl[50] br[50] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_51 bl[51] br[51] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_52 bl[52] br[52] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_53 bl[53] br[53] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_54 bl[54] br[54] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_55 bl[55] br[55] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_56 bl[56] br[56] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_57 bl[57] br[57] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_58 bl[58] br[58] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_59 bl[59] br[59] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_60 bl[60] br[60] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_61 bl[61] br[61] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_62 bl[62] br[62] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_210_63 bl[63] br[63] vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xcell_211_0 bl[0] br[0] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_1 bl[1] br[1] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_2 bl[2] br[2] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_3 bl[3] br[3] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_4 bl[4] br[4] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_5 bl[5] br[5] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_6 bl[6] br[6] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_7 bl[7] br[7] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_8 bl[8] br[8] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_9 bl[9] br[9] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_10 bl[10] br[10] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_11 bl[11] br[11] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_12 bl[12] br[12] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_13 bl[13] br[13] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_14 bl[14] br[14] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_15 bl[15] br[15] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_16 bl[16] br[16] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_17 bl[17] br[17] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_18 bl[18] br[18] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_19 bl[19] br[19] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_20 bl[20] br[20] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_21 bl[21] br[21] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_22 bl[22] br[22] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_23 bl[23] br[23] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_24 bl[24] br[24] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_25 bl[25] br[25] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_26 bl[26] br[26] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_27 bl[27] br[27] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_28 bl[28] br[28] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_29 bl[29] br[29] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_30 bl[30] br[30] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_31 bl[31] br[31] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_32 bl[32] br[32] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_33 bl[33] br[33] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_34 bl[34] br[34] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_35 bl[35] br[35] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_36 bl[36] br[36] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_37 bl[37] br[37] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_38 bl[38] br[38] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_39 bl[39] br[39] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_40 bl[40] br[40] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_41 bl[41] br[41] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_42 bl[42] br[42] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_43 bl[43] br[43] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_44 bl[44] br[44] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_45 bl[45] br[45] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_46 bl[46] br[46] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_47 bl[47] br[47] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_48 bl[48] br[48] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_49 bl[49] br[49] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_50 bl[50] br[50] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_51 bl[51] br[51] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_52 bl[52] br[52] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_53 bl[53] br[53] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_54 bl[54] br[54] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_55 bl[55] br[55] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_56 bl[56] br[56] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_57 bl[57] br[57] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_58 bl[58] br[58] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_59 bl[59] br[59] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_60 bl[60] br[60] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_61 bl[61] br[61] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_62 bl[62] br[62] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_211_63 bl[63] br[63] vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xcell_212_0 bl[0] br[0] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_1 bl[1] br[1] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_2 bl[2] br[2] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_3 bl[3] br[3] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_4 bl[4] br[4] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_5 bl[5] br[5] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_6 bl[6] br[6] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_7 bl[7] br[7] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_8 bl[8] br[8] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_9 bl[9] br[9] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_10 bl[10] br[10] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_11 bl[11] br[11] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_12 bl[12] br[12] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_13 bl[13] br[13] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_14 bl[14] br[14] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_15 bl[15] br[15] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_16 bl[16] br[16] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_17 bl[17] br[17] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_18 bl[18] br[18] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_19 bl[19] br[19] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_20 bl[20] br[20] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_21 bl[21] br[21] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_22 bl[22] br[22] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_23 bl[23] br[23] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_24 bl[24] br[24] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_25 bl[25] br[25] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_26 bl[26] br[26] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_27 bl[27] br[27] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_28 bl[28] br[28] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_29 bl[29] br[29] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_30 bl[30] br[30] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_31 bl[31] br[31] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_32 bl[32] br[32] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_33 bl[33] br[33] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_34 bl[34] br[34] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_35 bl[35] br[35] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_36 bl[36] br[36] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_37 bl[37] br[37] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_38 bl[38] br[38] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_39 bl[39] br[39] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_40 bl[40] br[40] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_41 bl[41] br[41] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_42 bl[42] br[42] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_43 bl[43] br[43] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_44 bl[44] br[44] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_45 bl[45] br[45] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_46 bl[46] br[46] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_47 bl[47] br[47] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_48 bl[48] br[48] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_49 bl[49] br[49] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_50 bl[50] br[50] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_51 bl[51] br[51] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_52 bl[52] br[52] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_53 bl[53] br[53] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_54 bl[54] br[54] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_55 bl[55] br[55] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_56 bl[56] br[56] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_57 bl[57] br[57] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_58 bl[58] br[58] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_59 bl[59] br[59] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_60 bl[60] br[60] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_61 bl[61] br[61] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_62 bl[62] br[62] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_212_63 bl[63] br[63] vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xcell_213_0 bl[0] br[0] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_1 bl[1] br[1] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_2 bl[2] br[2] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_3 bl[3] br[3] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_4 bl[4] br[4] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_5 bl[5] br[5] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_6 bl[6] br[6] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_7 bl[7] br[7] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_8 bl[8] br[8] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_9 bl[9] br[9] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_10 bl[10] br[10] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_11 bl[11] br[11] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_12 bl[12] br[12] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_13 bl[13] br[13] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_14 bl[14] br[14] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_15 bl[15] br[15] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_16 bl[16] br[16] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_17 bl[17] br[17] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_18 bl[18] br[18] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_19 bl[19] br[19] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_20 bl[20] br[20] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_21 bl[21] br[21] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_22 bl[22] br[22] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_23 bl[23] br[23] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_24 bl[24] br[24] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_25 bl[25] br[25] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_26 bl[26] br[26] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_27 bl[27] br[27] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_28 bl[28] br[28] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_29 bl[29] br[29] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_30 bl[30] br[30] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_31 bl[31] br[31] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_32 bl[32] br[32] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_33 bl[33] br[33] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_34 bl[34] br[34] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_35 bl[35] br[35] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_36 bl[36] br[36] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_37 bl[37] br[37] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_38 bl[38] br[38] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_39 bl[39] br[39] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_40 bl[40] br[40] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_41 bl[41] br[41] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_42 bl[42] br[42] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_43 bl[43] br[43] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_44 bl[44] br[44] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_45 bl[45] br[45] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_46 bl[46] br[46] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_47 bl[47] br[47] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_48 bl[48] br[48] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_49 bl[49] br[49] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_50 bl[50] br[50] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_51 bl[51] br[51] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_52 bl[52] br[52] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_53 bl[53] br[53] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_54 bl[54] br[54] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_55 bl[55] br[55] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_56 bl[56] br[56] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_57 bl[57] br[57] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_58 bl[58] br[58] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_59 bl[59] br[59] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_60 bl[60] br[60] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_61 bl[61] br[61] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_62 bl[62] br[62] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_213_63 bl[63] br[63] vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xcell_214_0 bl[0] br[0] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_1 bl[1] br[1] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_2 bl[2] br[2] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_3 bl[3] br[3] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_4 bl[4] br[4] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_5 bl[5] br[5] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_6 bl[6] br[6] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_7 bl[7] br[7] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_8 bl[8] br[8] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_9 bl[9] br[9] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_10 bl[10] br[10] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_11 bl[11] br[11] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_12 bl[12] br[12] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_13 bl[13] br[13] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_14 bl[14] br[14] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_15 bl[15] br[15] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_16 bl[16] br[16] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_17 bl[17] br[17] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_18 bl[18] br[18] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_19 bl[19] br[19] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_20 bl[20] br[20] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_21 bl[21] br[21] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_22 bl[22] br[22] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_23 bl[23] br[23] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_24 bl[24] br[24] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_25 bl[25] br[25] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_26 bl[26] br[26] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_27 bl[27] br[27] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_28 bl[28] br[28] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_29 bl[29] br[29] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_30 bl[30] br[30] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_31 bl[31] br[31] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_32 bl[32] br[32] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_33 bl[33] br[33] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_34 bl[34] br[34] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_35 bl[35] br[35] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_36 bl[36] br[36] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_37 bl[37] br[37] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_38 bl[38] br[38] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_39 bl[39] br[39] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_40 bl[40] br[40] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_41 bl[41] br[41] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_42 bl[42] br[42] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_43 bl[43] br[43] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_44 bl[44] br[44] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_45 bl[45] br[45] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_46 bl[46] br[46] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_47 bl[47] br[47] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_48 bl[48] br[48] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_49 bl[49] br[49] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_50 bl[50] br[50] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_51 bl[51] br[51] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_52 bl[52] br[52] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_53 bl[53] br[53] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_54 bl[54] br[54] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_55 bl[55] br[55] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_56 bl[56] br[56] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_57 bl[57] br[57] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_58 bl[58] br[58] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_59 bl[59] br[59] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_60 bl[60] br[60] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_61 bl[61] br[61] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_62 bl[62] br[62] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_214_63 bl[63] br[63] vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xcell_215_0 bl[0] br[0] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_1 bl[1] br[1] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_2 bl[2] br[2] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_3 bl[3] br[3] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_4 bl[4] br[4] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_5 bl[5] br[5] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_6 bl[6] br[6] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_7 bl[7] br[7] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_8 bl[8] br[8] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_9 bl[9] br[9] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_10 bl[10] br[10] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_11 bl[11] br[11] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_12 bl[12] br[12] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_13 bl[13] br[13] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_14 bl[14] br[14] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_15 bl[15] br[15] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_16 bl[16] br[16] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_17 bl[17] br[17] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_18 bl[18] br[18] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_19 bl[19] br[19] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_20 bl[20] br[20] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_21 bl[21] br[21] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_22 bl[22] br[22] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_23 bl[23] br[23] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_24 bl[24] br[24] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_25 bl[25] br[25] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_26 bl[26] br[26] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_27 bl[27] br[27] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_28 bl[28] br[28] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_29 bl[29] br[29] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_30 bl[30] br[30] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_31 bl[31] br[31] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_32 bl[32] br[32] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_33 bl[33] br[33] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_34 bl[34] br[34] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_35 bl[35] br[35] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_36 bl[36] br[36] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_37 bl[37] br[37] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_38 bl[38] br[38] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_39 bl[39] br[39] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_40 bl[40] br[40] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_41 bl[41] br[41] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_42 bl[42] br[42] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_43 bl[43] br[43] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_44 bl[44] br[44] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_45 bl[45] br[45] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_46 bl[46] br[46] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_47 bl[47] br[47] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_48 bl[48] br[48] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_49 bl[49] br[49] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_50 bl[50] br[50] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_51 bl[51] br[51] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_52 bl[52] br[52] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_53 bl[53] br[53] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_54 bl[54] br[54] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_55 bl[55] br[55] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_56 bl[56] br[56] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_57 bl[57] br[57] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_58 bl[58] br[58] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_59 bl[59] br[59] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_60 bl[60] br[60] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_61 bl[61] br[61] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_62 bl[62] br[62] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_215_63 bl[63] br[63] vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xcell_216_0 bl[0] br[0] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_1 bl[1] br[1] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_2 bl[2] br[2] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_3 bl[3] br[3] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_4 bl[4] br[4] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_5 bl[5] br[5] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_6 bl[6] br[6] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_7 bl[7] br[7] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_8 bl[8] br[8] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_9 bl[9] br[9] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_10 bl[10] br[10] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_11 bl[11] br[11] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_12 bl[12] br[12] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_13 bl[13] br[13] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_14 bl[14] br[14] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_15 bl[15] br[15] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_16 bl[16] br[16] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_17 bl[17] br[17] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_18 bl[18] br[18] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_19 bl[19] br[19] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_20 bl[20] br[20] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_21 bl[21] br[21] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_22 bl[22] br[22] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_23 bl[23] br[23] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_24 bl[24] br[24] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_25 bl[25] br[25] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_26 bl[26] br[26] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_27 bl[27] br[27] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_28 bl[28] br[28] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_29 bl[29] br[29] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_30 bl[30] br[30] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_31 bl[31] br[31] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_32 bl[32] br[32] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_33 bl[33] br[33] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_34 bl[34] br[34] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_35 bl[35] br[35] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_36 bl[36] br[36] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_37 bl[37] br[37] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_38 bl[38] br[38] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_39 bl[39] br[39] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_40 bl[40] br[40] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_41 bl[41] br[41] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_42 bl[42] br[42] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_43 bl[43] br[43] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_44 bl[44] br[44] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_45 bl[45] br[45] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_46 bl[46] br[46] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_47 bl[47] br[47] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_48 bl[48] br[48] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_49 bl[49] br[49] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_50 bl[50] br[50] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_51 bl[51] br[51] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_52 bl[52] br[52] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_53 bl[53] br[53] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_54 bl[54] br[54] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_55 bl[55] br[55] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_56 bl[56] br[56] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_57 bl[57] br[57] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_58 bl[58] br[58] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_59 bl[59] br[59] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_60 bl[60] br[60] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_61 bl[61] br[61] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_62 bl[62] br[62] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_216_63 bl[63] br[63] vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xcell_217_0 bl[0] br[0] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_1 bl[1] br[1] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_2 bl[2] br[2] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_3 bl[3] br[3] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_4 bl[4] br[4] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_5 bl[5] br[5] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_6 bl[6] br[6] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_7 bl[7] br[7] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_8 bl[8] br[8] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_9 bl[9] br[9] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_10 bl[10] br[10] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_11 bl[11] br[11] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_12 bl[12] br[12] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_13 bl[13] br[13] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_14 bl[14] br[14] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_15 bl[15] br[15] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_16 bl[16] br[16] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_17 bl[17] br[17] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_18 bl[18] br[18] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_19 bl[19] br[19] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_20 bl[20] br[20] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_21 bl[21] br[21] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_22 bl[22] br[22] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_23 bl[23] br[23] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_24 bl[24] br[24] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_25 bl[25] br[25] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_26 bl[26] br[26] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_27 bl[27] br[27] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_28 bl[28] br[28] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_29 bl[29] br[29] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_30 bl[30] br[30] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_31 bl[31] br[31] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_32 bl[32] br[32] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_33 bl[33] br[33] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_34 bl[34] br[34] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_35 bl[35] br[35] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_36 bl[36] br[36] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_37 bl[37] br[37] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_38 bl[38] br[38] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_39 bl[39] br[39] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_40 bl[40] br[40] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_41 bl[41] br[41] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_42 bl[42] br[42] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_43 bl[43] br[43] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_44 bl[44] br[44] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_45 bl[45] br[45] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_46 bl[46] br[46] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_47 bl[47] br[47] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_48 bl[48] br[48] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_49 bl[49] br[49] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_50 bl[50] br[50] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_51 bl[51] br[51] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_52 bl[52] br[52] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_53 bl[53] br[53] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_54 bl[54] br[54] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_55 bl[55] br[55] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_56 bl[56] br[56] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_57 bl[57] br[57] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_58 bl[58] br[58] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_59 bl[59] br[59] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_60 bl[60] br[60] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_61 bl[61] br[61] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_62 bl[62] br[62] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_217_63 bl[63] br[63] vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xcell_218_0 bl[0] br[0] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_1 bl[1] br[1] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_2 bl[2] br[2] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_3 bl[3] br[3] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_4 bl[4] br[4] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_5 bl[5] br[5] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_6 bl[6] br[6] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_7 bl[7] br[7] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_8 bl[8] br[8] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_9 bl[9] br[9] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_10 bl[10] br[10] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_11 bl[11] br[11] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_12 bl[12] br[12] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_13 bl[13] br[13] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_14 bl[14] br[14] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_15 bl[15] br[15] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_16 bl[16] br[16] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_17 bl[17] br[17] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_18 bl[18] br[18] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_19 bl[19] br[19] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_20 bl[20] br[20] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_21 bl[21] br[21] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_22 bl[22] br[22] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_23 bl[23] br[23] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_24 bl[24] br[24] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_25 bl[25] br[25] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_26 bl[26] br[26] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_27 bl[27] br[27] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_28 bl[28] br[28] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_29 bl[29] br[29] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_30 bl[30] br[30] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_31 bl[31] br[31] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_32 bl[32] br[32] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_33 bl[33] br[33] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_34 bl[34] br[34] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_35 bl[35] br[35] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_36 bl[36] br[36] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_37 bl[37] br[37] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_38 bl[38] br[38] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_39 bl[39] br[39] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_40 bl[40] br[40] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_41 bl[41] br[41] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_42 bl[42] br[42] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_43 bl[43] br[43] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_44 bl[44] br[44] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_45 bl[45] br[45] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_46 bl[46] br[46] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_47 bl[47] br[47] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_48 bl[48] br[48] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_49 bl[49] br[49] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_50 bl[50] br[50] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_51 bl[51] br[51] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_52 bl[52] br[52] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_53 bl[53] br[53] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_54 bl[54] br[54] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_55 bl[55] br[55] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_56 bl[56] br[56] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_57 bl[57] br[57] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_58 bl[58] br[58] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_59 bl[59] br[59] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_60 bl[60] br[60] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_61 bl[61] br[61] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_62 bl[62] br[62] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_218_63 bl[63] br[63] vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xcell_219_0 bl[0] br[0] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_1 bl[1] br[1] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_2 bl[2] br[2] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_3 bl[3] br[3] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_4 bl[4] br[4] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_5 bl[5] br[5] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_6 bl[6] br[6] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_7 bl[7] br[7] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_8 bl[8] br[8] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_9 bl[9] br[9] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_10 bl[10] br[10] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_11 bl[11] br[11] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_12 bl[12] br[12] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_13 bl[13] br[13] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_14 bl[14] br[14] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_15 bl[15] br[15] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_16 bl[16] br[16] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_17 bl[17] br[17] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_18 bl[18] br[18] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_19 bl[19] br[19] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_20 bl[20] br[20] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_21 bl[21] br[21] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_22 bl[22] br[22] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_23 bl[23] br[23] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_24 bl[24] br[24] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_25 bl[25] br[25] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_26 bl[26] br[26] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_27 bl[27] br[27] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_28 bl[28] br[28] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_29 bl[29] br[29] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_30 bl[30] br[30] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_31 bl[31] br[31] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_32 bl[32] br[32] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_33 bl[33] br[33] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_34 bl[34] br[34] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_35 bl[35] br[35] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_36 bl[36] br[36] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_37 bl[37] br[37] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_38 bl[38] br[38] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_39 bl[39] br[39] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_40 bl[40] br[40] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_41 bl[41] br[41] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_42 bl[42] br[42] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_43 bl[43] br[43] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_44 bl[44] br[44] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_45 bl[45] br[45] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_46 bl[46] br[46] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_47 bl[47] br[47] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_48 bl[48] br[48] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_49 bl[49] br[49] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_50 bl[50] br[50] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_51 bl[51] br[51] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_52 bl[52] br[52] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_53 bl[53] br[53] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_54 bl[54] br[54] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_55 bl[55] br[55] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_56 bl[56] br[56] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_57 bl[57] br[57] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_58 bl[58] br[58] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_59 bl[59] br[59] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_60 bl[60] br[60] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_61 bl[61] br[61] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_62 bl[62] br[62] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_219_63 bl[63] br[63] vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xcell_220_0 bl[0] br[0] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_1 bl[1] br[1] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_2 bl[2] br[2] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_3 bl[3] br[3] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_4 bl[4] br[4] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_5 bl[5] br[5] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_6 bl[6] br[6] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_7 bl[7] br[7] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_8 bl[8] br[8] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_9 bl[9] br[9] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_10 bl[10] br[10] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_11 bl[11] br[11] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_12 bl[12] br[12] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_13 bl[13] br[13] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_14 bl[14] br[14] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_15 bl[15] br[15] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_16 bl[16] br[16] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_17 bl[17] br[17] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_18 bl[18] br[18] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_19 bl[19] br[19] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_20 bl[20] br[20] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_21 bl[21] br[21] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_22 bl[22] br[22] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_23 bl[23] br[23] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_24 bl[24] br[24] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_25 bl[25] br[25] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_26 bl[26] br[26] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_27 bl[27] br[27] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_28 bl[28] br[28] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_29 bl[29] br[29] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_30 bl[30] br[30] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_31 bl[31] br[31] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_32 bl[32] br[32] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_33 bl[33] br[33] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_34 bl[34] br[34] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_35 bl[35] br[35] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_36 bl[36] br[36] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_37 bl[37] br[37] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_38 bl[38] br[38] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_39 bl[39] br[39] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_40 bl[40] br[40] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_41 bl[41] br[41] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_42 bl[42] br[42] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_43 bl[43] br[43] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_44 bl[44] br[44] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_45 bl[45] br[45] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_46 bl[46] br[46] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_47 bl[47] br[47] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_48 bl[48] br[48] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_49 bl[49] br[49] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_50 bl[50] br[50] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_51 bl[51] br[51] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_52 bl[52] br[52] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_53 bl[53] br[53] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_54 bl[54] br[54] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_55 bl[55] br[55] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_56 bl[56] br[56] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_57 bl[57] br[57] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_58 bl[58] br[58] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_59 bl[59] br[59] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_60 bl[60] br[60] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_61 bl[61] br[61] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_62 bl[62] br[62] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_220_63 bl[63] br[63] vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xcell_221_0 bl[0] br[0] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_1 bl[1] br[1] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_2 bl[2] br[2] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_3 bl[3] br[3] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_4 bl[4] br[4] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_5 bl[5] br[5] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_6 bl[6] br[6] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_7 bl[7] br[7] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_8 bl[8] br[8] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_9 bl[9] br[9] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_10 bl[10] br[10] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_11 bl[11] br[11] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_12 bl[12] br[12] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_13 bl[13] br[13] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_14 bl[14] br[14] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_15 bl[15] br[15] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_16 bl[16] br[16] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_17 bl[17] br[17] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_18 bl[18] br[18] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_19 bl[19] br[19] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_20 bl[20] br[20] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_21 bl[21] br[21] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_22 bl[22] br[22] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_23 bl[23] br[23] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_24 bl[24] br[24] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_25 bl[25] br[25] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_26 bl[26] br[26] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_27 bl[27] br[27] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_28 bl[28] br[28] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_29 bl[29] br[29] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_30 bl[30] br[30] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_31 bl[31] br[31] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_32 bl[32] br[32] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_33 bl[33] br[33] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_34 bl[34] br[34] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_35 bl[35] br[35] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_36 bl[36] br[36] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_37 bl[37] br[37] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_38 bl[38] br[38] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_39 bl[39] br[39] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_40 bl[40] br[40] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_41 bl[41] br[41] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_42 bl[42] br[42] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_43 bl[43] br[43] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_44 bl[44] br[44] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_45 bl[45] br[45] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_46 bl[46] br[46] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_47 bl[47] br[47] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_48 bl[48] br[48] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_49 bl[49] br[49] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_50 bl[50] br[50] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_51 bl[51] br[51] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_52 bl[52] br[52] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_53 bl[53] br[53] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_54 bl[54] br[54] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_55 bl[55] br[55] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_56 bl[56] br[56] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_57 bl[57] br[57] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_58 bl[58] br[58] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_59 bl[59] br[59] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_60 bl[60] br[60] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_61 bl[61] br[61] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_62 bl[62] br[62] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_221_63 bl[63] br[63] vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xcell_222_0 bl[0] br[0] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_1 bl[1] br[1] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_2 bl[2] br[2] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_3 bl[3] br[3] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_4 bl[4] br[4] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_5 bl[5] br[5] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_6 bl[6] br[6] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_7 bl[7] br[7] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_8 bl[8] br[8] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_9 bl[9] br[9] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_10 bl[10] br[10] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_11 bl[11] br[11] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_12 bl[12] br[12] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_13 bl[13] br[13] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_14 bl[14] br[14] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_15 bl[15] br[15] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_16 bl[16] br[16] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_17 bl[17] br[17] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_18 bl[18] br[18] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_19 bl[19] br[19] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_20 bl[20] br[20] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_21 bl[21] br[21] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_22 bl[22] br[22] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_23 bl[23] br[23] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_24 bl[24] br[24] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_25 bl[25] br[25] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_26 bl[26] br[26] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_27 bl[27] br[27] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_28 bl[28] br[28] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_29 bl[29] br[29] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_30 bl[30] br[30] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_31 bl[31] br[31] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_32 bl[32] br[32] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_33 bl[33] br[33] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_34 bl[34] br[34] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_35 bl[35] br[35] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_36 bl[36] br[36] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_37 bl[37] br[37] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_38 bl[38] br[38] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_39 bl[39] br[39] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_40 bl[40] br[40] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_41 bl[41] br[41] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_42 bl[42] br[42] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_43 bl[43] br[43] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_44 bl[44] br[44] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_45 bl[45] br[45] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_46 bl[46] br[46] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_47 bl[47] br[47] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_48 bl[48] br[48] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_49 bl[49] br[49] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_50 bl[50] br[50] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_51 bl[51] br[51] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_52 bl[52] br[52] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_53 bl[53] br[53] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_54 bl[54] br[54] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_55 bl[55] br[55] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_56 bl[56] br[56] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_57 bl[57] br[57] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_58 bl[58] br[58] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_59 bl[59] br[59] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_60 bl[60] br[60] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_61 bl[61] br[61] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_62 bl[62] br[62] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_222_63 bl[63] br[63] vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xcell_223_0 bl[0] br[0] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_1 bl[1] br[1] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_2 bl[2] br[2] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_3 bl[3] br[3] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_4 bl[4] br[4] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_5 bl[5] br[5] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_6 bl[6] br[6] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_7 bl[7] br[7] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_8 bl[8] br[8] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_9 bl[9] br[9] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_10 bl[10] br[10] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_11 bl[11] br[11] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_12 bl[12] br[12] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_13 bl[13] br[13] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_14 bl[14] br[14] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_15 bl[15] br[15] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_16 bl[16] br[16] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_17 bl[17] br[17] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_18 bl[18] br[18] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_19 bl[19] br[19] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_20 bl[20] br[20] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_21 bl[21] br[21] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_22 bl[22] br[22] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_23 bl[23] br[23] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_24 bl[24] br[24] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_25 bl[25] br[25] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_26 bl[26] br[26] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_27 bl[27] br[27] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_28 bl[28] br[28] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_29 bl[29] br[29] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_30 bl[30] br[30] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_31 bl[31] br[31] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_32 bl[32] br[32] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_33 bl[33] br[33] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_34 bl[34] br[34] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_35 bl[35] br[35] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_36 bl[36] br[36] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_37 bl[37] br[37] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_38 bl[38] br[38] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_39 bl[39] br[39] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_40 bl[40] br[40] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_41 bl[41] br[41] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_42 bl[42] br[42] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_43 bl[43] br[43] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_44 bl[44] br[44] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_45 bl[45] br[45] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_46 bl[46] br[46] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_47 bl[47] br[47] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_48 bl[48] br[48] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_49 bl[49] br[49] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_50 bl[50] br[50] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_51 bl[51] br[51] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_52 bl[52] br[52] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_53 bl[53] br[53] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_54 bl[54] br[54] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_55 bl[55] br[55] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_56 bl[56] br[56] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_57 bl[57] br[57] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_58 bl[58] br[58] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_59 bl[59] br[59] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_60 bl[60] br[60] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_61 bl[61] br[61] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_62 bl[62] br[62] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_223_63 bl[63] br[63] vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xcell_224_0 bl[0] br[0] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_1 bl[1] br[1] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_2 bl[2] br[2] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_3 bl[3] br[3] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_4 bl[4] br[4] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_5 bl[5] br[5] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_6 bl[6] br[6] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_7 bl[7] br[7] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_8 bl[8] br[8] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_9 bl[9] br[9] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_10 bl[10] br[10] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_11 bl[11] br[11] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_12 bl[12] br[12] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_13 bl[13] br[13] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_14 bl[14] br[14] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_15 bl[15] br[15] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_16 bl[16] br[16] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_17 bl[17] br[17] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_18 bl[18] br[18] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_19 bl[19] br[19] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_20 bl[20] br[20] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_21 bl[21] br[21] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_22 bl[22] br[22] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_23 bl[23] br[23] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_24 bl[24] br[24] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_25 bl[25] br[25] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_26 bl[26] br[26] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_27 bl[27] br[27] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_28 bl[28] br[28] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_29 bl[29] br[29] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_30 bl[30] br[30] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_31 bl[31] br[31] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_32 bl[32] br[32] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_33 bl[33] br[33] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_34 bl[34] br[34] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_35 bl[35] br[35] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_36 bl[36] br[36] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_37 bl[37] br[37] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_38 bl[38] br[38] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_39 bl[39] br[39] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_40 bl[40] br[40] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_41 bl[41] br[41] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_42 bl[42] br[42] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_43 bl[43] br[43] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_44 bl[44] br[44] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_45 bl[45] br[45] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_46 bl[46] br[46] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_47 bl[47] br[47] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_48 bl[48] br[48] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_49 bl[49] br[49] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_50 bl[50] br[50] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_51 bl[51] br[51] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_52 bl[52] br[52] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_53 bl[53] br[53] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_54 bl[54] br[54] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_55 bl[55] br[55] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_56 bl[56] br[56] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_57 bl[57] br[57] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_58 bl[58] br[58] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_59 bl[59] br[59] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_60 bl[60] br[60] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_61 bl[61] br[61] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_62 bl[62] br[62] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_224_63 bl[63] br[63] vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xcell_225_0 bl[0] br[0] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_1 bl[1] br[1] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_2 bl[2] br[2] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_3 bl[3] br[3] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_4 bl[4] br[4] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_5 bl[5] br[5] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_6 bl[6] br[6] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_7 bl[7] br[7] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_8 bl[8] br[8] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_9 bl[9] br[9] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_10 bl[10] br[10] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_11 bl[11] br[11] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_12 bl[12] br[12] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_13 bl[13] br[13] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_14 bl[14] br[14] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_15 bl[15] br[15] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_16 bl[16] br[16] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_17 bl[17] br[17] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_18 bl[18] br[18] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_19 bl[19] br[19] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_20 bl[20] br[20] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_21 bl[21] br[21] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_22 bl[22] br[22] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_23 bl[23] br[23] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_24 bl[24] br[24] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_25 bl[25] br[25] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_26 bl[26] br[26] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_27 bl[27] br[27] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_28 bl[28] br[28] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_29 bl[29] br[29] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_30 bl[30] br[30] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_31 bl[31] br[31] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_32 bl[32] br[32] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_33 bl[33] br[33] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_34 bl[34] br[34] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_35 bl[35] br[35] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_36 bl[36] br[36] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_37 bl[37] br[37] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_38 bl[38] br[38] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_39 bl[39] br[39] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_40 bl[40] br[40] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_41 bl[41] br[41] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_42 bl[42] br[42] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_43 bl[43] br[43] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_44 bl[44] br[44] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_45 bl[45] br[45] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_46 bl[46] br[46] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_47 bl[47] br[47] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_48 bl[48] br[48] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_49 bl[49] br[49] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_50 bl[50] br[50] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_51 bl[51] br[51] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_52 bl[52] br[52] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_53 bl[53] br[53] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_54 bl[54] br[54] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_55 bl[55] br[55] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_56 bl[56] br[56] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_57 bl[57] br[57] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_58 bl[58] br[58] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_59 bl[59] br[59] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_60 bl[60] br[60] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_61 bl[61] br[61] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_62 bl[62] br[62] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_225_63 bl[63] br[63] vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xcell_226_0 bl[0] br[0] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_1 bl[1] br[1] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_2 bl[2] br[2] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_3 bl[3] br[3] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_4 bl[4] br[4] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_5 bl[5] br[5] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_6 bl[6] br[6] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_7 bl[7] br[7] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_8 bl[8] br[8] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_9 bl[9] br[9] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_10 bl[10] br[10] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_11 bl[11] br[11] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_12 bl[12] br[12] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_13 bl[13] br[13] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_14 bl[14] br[14] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_15 bl[15] br[15] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_16 bl[16] br[16] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_17 bl[17] br[17] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_18 bl[18] br[18] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_19 bl[19] br[19] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_20 bl[20] br[20] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_21 bl[21] br[21] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_22 bl[22] br[22] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_23 bl[23] br[23] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_24 bl[24] br[24] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_25 bl[25] br[25] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_26 bl[26] br[26] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_27 bl[27] br[27] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_28 bl[28] br[28] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_29 bl[29] br[29] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_30 bl[30] br[30] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_31 bl[31] br[31] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_32 bl[32] br[32] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_33 bl[33] br[33] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_34 bl[34] br[34] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_35 bl[35] br[35] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_36 bl[36] br[36] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_37 bl[37] br[37] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_38 bl[38] br[38] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_39 bl[39] br[39] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_40 bl[40] br[40] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_41 bl[41] br[41] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_42 bl[42] br[42] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_43 bl[43] br[43] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_44 bl[44] br[44] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_45 bl[45] br[45] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_46 bl[46] br[46] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_47 bl[47] br[47] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_48 bl[48] br[48] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_49 bl[49] br[49] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_50 bl[50] br[50] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_51 bl[51] br[51] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_52 bl[52] br[52] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_53 bl[53] br[53] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_54 bl[54] br[54] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_55 bl[55] br[55] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_56 bl[56] br[56] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_57 bl[57] br[57] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_58 bl[58] br[58] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_59 bl[59] br[59] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_60 bl[60] br[60] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_61 bl[61] br[61] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_62 bl[62] br[62] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_226_63 bl[63] br[63] vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xcell_227_0 bl[0] br[0] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_1 bl[1] br[1] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_2 bl[2] br[2] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_3 bl[3] br[3] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_4 bl[4] br[4] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_5 bl[5] br[5] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_6 bl[6] br[6] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_7 bl[7] br[7] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_8 bl[8] br[8] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_9 bl[9] br[9] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_10 bl[10] br[10] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_11 bl[11] br[11] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_12 bl[12] br[12] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_13 bl[13] br[13] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_14 bl[14] br[14] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_15 bl[15] br[15] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_16 bl[16] br[16] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_17 bl[17] br[17] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_18 bl[18] br[18] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_19 bl[19] br[19] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_20 bl[20] br[20] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_21 bl[21] br[21] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_22 bl[22] br[22] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_23 bl[23] br[23] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_24 bl[24] br[24] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_25 bl[25] br[25] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_26 bl[26] br[26] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_27 bl[27] br[27] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_28 bl[28] br[28] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_29 bl[29] br[29] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_30 bl[30] br[30] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_31 bl[31] br[31] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_32 bl[32] br[32] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_33 bl[33] br[33] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_34 bl[34] br[34] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_35 bl[35] br[35] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_36 bl[36] br[36] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_37 bl[37] br[37] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_38 bl[38] br[38] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_39 bl[39] br[39] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_40 bl[40] br[40] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_41 bl[41] br[41] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_42 bl[42] br[42] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_43 bl[43] br[43] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_44 bl[44] br[44] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_45 bl[45] br[45] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_46 bl[46] br[46] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_47 bl[47] br[47] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_48 bl[48] br[48] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_49 bl[49] br[49] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_50 bl[50] br[50] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_51 bl[51] br[51] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_52 bl[52] br[52] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_53 bl[53] br[53] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_54 bl[54] br[54] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_55 bl[55] br[55] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_56 bl[56] br[56] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_57 bl[57] br[57] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_58 bl[58] br[58] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_59 bl[59] br[59] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_60 bl[60] br[60] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_61 bl[61] br[61] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_62 bl[62] br[62] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_227_63 bl[63] br[63] vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xcell_228_0 bl[0] br[0] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_1 bl[1] br[1] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_2 bl[2] br[2] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_3 bl[3] br[3] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_4 bl[4] br[4] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_5 bl[5] br[5] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_6 bl[6] br[6] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_7 bl[7] br[7] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_8 bl[8] br[8] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_9 bl[9] br[9] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_10 bl[10] br[10] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_11 bl[11] br[11] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_12 bl[12] br[12] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_13 bl[13] br[13] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_14 bl[14] br[14] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_15 bl[15] br[15] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_16 bl[16] br[16] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_17 bl[17] br[17] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_18 bl[18] br[18] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_19 bl[19] br[19] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_20 bl[20] br[20] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_21 bl[21] br[21] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_22 bl[22] br[22] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_23 bl[23] br[23] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_24 bl[24] br[24] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_25 bl[25] br[25] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_26 bl[26] br[26] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_27 bl[27] br[27] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_28 bl[28] br[28] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_29 bl[29] br[29] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_30 bl[30] br[30] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_31 bl[31] br[31] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_32 bl[32] br[32] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_33 bl[33] br[33] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_34 bl[34] br[34] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_35 bl[35] br[35] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_36 bl[36] br[36] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_37 bl[37] br[37] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_38 bl[38] br[38] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_39 bl[39] br[39] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_40 bl[40] br[40] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_41 bl[41] br[41] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_42 bl[42] br[42] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_43 bl[43] br[43] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_44 bl[44] br[44] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_45 bl[45] br[45] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_46 bl[46] br[46] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_47 bl[47] br[47] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_48 bl[48] br[48] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_49 bl[49] br[49] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_50 bl[50] br[50] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_51 bl[51] br[51] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_52 bl[52] br[52] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_53 bl[53] br[53] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_54 bl[54] br[54] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_55 bl[55] br[55] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_56 bl[56] br[56] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_57 bl[57] br[57] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_58 bl[58] br[58] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_59 bl[59] br[59] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_60 bl[60] br[60] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_61 bl[61] br[61] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_62 bl[62] br[62] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_228_63 bl[63] br[63] vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xcell_229_0 bl[0] br[0] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_1 bl[1] br[1] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_2 bl[2] br[2] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_3 bl[3] br[3] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_4 bl[4] br[4] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_5 bl[5] br[5] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_6 bl[6] br[6] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_7 bl[7] br[7] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_8 bl[8] br[8] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_9 bl[9] br[9] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_10 bl[10] br[10] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_11 bl[11] br[11] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_12 bl[12] br[12] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_13 bl[13] br[13] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_14 bl[14] br[14] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_15 bl[15] br[15] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_16 bl[16] br[16] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_17 bl[17] br[17] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_18 bl[18] br[18] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_19 bl[19] br[19] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_20 bl[20] br[20] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_21 bl[21] br[21] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_22 bl[22] br[22] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_23 bl[23] br[23] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_24 bl[24] br[24] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_25 bl[25] br[25] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_26 bl[26] br[26] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_27 bl[27] br[27] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_28 bl[28] br[28] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_29 bl[29] br[29] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_30 bl[30] br[30] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_31 bl[31] br[31] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_32 bl[32] br[32] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_33 bl[33] br[33] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_34 bl[34] br[34] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_35 bl[35] br[35] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_36 bl[36] br[36] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_37 bl[37] br[37] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_38 bl[38] br[38] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_39 bl[39] br[39] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_40 bl[40] br[40] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_41 bl[41] br[41] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_42 bl[42] br[42] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_43 bl[43] br[43] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_44 bl[44] br[44] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_45 bl[45] br[45] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_46 bl[46] br[46] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_47 bl[47] br[47] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_48 bl[48] br[48] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_49 bl[49] br[49] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_50 bl[50] br[50] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_51 bl[51] br[51] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_52 bl[52] br[52] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_53 bl[53] br[53] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_54 bl[54] br[54] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_55 bl[55] br[55] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_56 bl[56] br[56] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_57 bl[57] br[57] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_58 bl[58] br[58] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_59 bl[59] br[59] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_60 bl[60] br[60] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_61 bl[61] br[61] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_62 bl[62] br[62] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_229_63 bl[63] br[63] vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xcell_230_0 bl[0] br[0] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_1 bl[1] br[1] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_2 bl[2] br[2] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_3 bl[3] br[3] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_4 bl[4] br[4] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_5 bl[5] br[5] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_6 bl[6] br[6] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_7 bl[7] br[7] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_8 bl[8] br[8] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_9 bl[9] br[9] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_10 bl[10] br[10] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_11 bl[11] br[11] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_12 bl[12] br[12] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_13 bl[13] br[13] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_14 bl[14] br[14] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_15 bl[15] br[15] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_16 bl[16] br[16] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_17 bl[17] br[17] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_18 bl[18] br[18] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_19 bl[19] br[19] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_20 bl[20] br[20] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_21 bl[21] br[21] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_22 bl[22] br[22] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_23 bl[23] br[23] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_24 bl[24] br[24] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_25 bl[25] br[25] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_26 bl[26] br[26] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_27 bl[27] br[27] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_28 bl[28] br[28] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_29 bl[29] br[29] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_30 bl[30] br[30] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_31 bl[31] br[31] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_32 bl[32] br[32] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_33 bl[33] br[33] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_34 bl[34] br[34] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_35 bl[35] br[35] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_36 bl[36] br[36] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_37 bl[37] br[37] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_38 bl[38] br[38] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_39 bl[39] br[39] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_40 bl[40] br[40] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_41 bl[41] br[41] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_42 bl[42] br[42] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_43 bl[43] br[43] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_44 bl[44] br[44] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_45 bl[45] br[45] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_46 bl[46] br[46] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_47 bl[47] br[47] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_48 bl[48] br[48] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_49 bl[49] br[49] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_50 bl[50] br[50] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_51 bl[51] br[51] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_52 bl[52] br[52] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_53 bl[53] br[53] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_54 bl[54] br[54] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_55 bl[55] br[55] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_56 bl[56] br[56] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_57 bl[57] br[57] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_58 bl[58] br[58] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_59 bl[59] br[59] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_60 bl[60] br[60] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_61 bl[61] br[61] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_62 bl[62] br[62] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_230_63 bl[63] br[63] vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xcell_231_0 bl[0] br[0] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_1 bl[1] br[1] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_2 bl[2] br[2] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_3 bl[3] br[3] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_4 bl[4] br[4] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_5 bl[5] br[5] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_6 bl[6] br[6] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_7 bl[7] br[7] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_8 bl[8] br[8] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_9 bl[9] br[9] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_10 bl[10] br[10] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_11 bl[11] br[11] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_12 bl[12] br[12] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_13 bl[13] br[13] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_14 bl[14] br[14] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_15 bl[15] br[15] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_16 bl[16] br[16] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_17 bl[17] br[17] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_18 bl[18] br[18] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_19 bl[19] br[19] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_20 bl[20] br[20] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_21 bl[21] br[21] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_22 bl[22] br[22] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_23 bl[23] br[23] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_24 bl[24] br[24] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_25 bl[25] br[25] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_26 bl[26] br[26] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_27 bl[27] br[27] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_28 bl[28] br[28] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_29 bl[29] br[29] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_30 bl[30] br[30] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_31 bl[31] br[31] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_32 bl[32] br[32] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_33 bl[33] br[33] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_34 bl[34] br[34] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_35 bl[35] br[35] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_36 bl[36] br[36] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_37 bl[37] br[37] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_38 bl[38] br[38] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_39 bl[39] br[39] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_40 bl[40] br[40] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_41 bl[41] br[41] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_42 bl[42] br[42] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_43 bl[43] br[43] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_44 bl[44] br[44] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_45 bl[45] br[45] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_46 bl[46] br[46] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_47 bl[47] br[47] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_48 bl[48] br[48] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_49 bl[49] br[49] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_50 bl[50] br[50] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_51 bl[51] br[51] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_52 bl[52] br[52] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_53 bl[53] br[53] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_54 bl[54] br[54] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_55 bl[55] br[55] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_56 bl[56] br[56] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_57 bl[57] br[57] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_58 bl[58] br[58] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_59 bl[59] br[59] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_60 bl[60] br[60] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_61 bl[61] br[61] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_62 bl[62] br[62] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_231_63 bl[63] br[63] vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xcell_232_0 bl[0] br[0] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_1 bl[1] br[1] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_2 bl[2] br[2] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_3 bl[3] br[3] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_4 bl[4] br[4] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_5 bl[5] br[5] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_6 bl[6] br[6] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_7 bl[7] br[7] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_8 bl[8] br[8] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_9 bl[9] br[9] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_10 bl[10] br[10] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_11 bl[11] br[11] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_12 bl[12] br[12] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_13 bl[13] br[13] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_14 bl[14] br[14] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_15 bl[15] br[15] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_16 bl[16] br[16] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_17 bl[17] br[17] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_18 bl[18] br[18] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_19 bl[19] br[19] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_20 bl[20] br[20] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_21 bl[21] br[21] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_22 bl[22] br[22] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_23 bl[23] br[23] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_24 bl[24] br[24] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_25 bl[25] br[25] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_26 bl[26] br[26] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_27 bl[27] br[27] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_28 bl[28] br[28] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_29 bl[29] br[29] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_30 bl[30] br[30] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_31 bl[31] br[31] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_32 bl[32] br[32] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_33 bl[33] br[33] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_34 bl[34] br[34] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_35 bl[35] br[35] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_36 bl[36] br[36] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_37 bl[37] br[37] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_38 bl[38] br[38] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_39 bl[39] br[39] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_40 bl[40] br[40] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_41 bl[41] br[41] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_42 bl[42] br[42] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_43 bl[43] br[43] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_44 bl[44] br[44] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_45 bl[45] br[45] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_46 bl[46] br[46] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_47 bl[47] br[47] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_48 bl[48] br[48] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_49 bl[49] br[49] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_50 bl[50] br[50] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_51 bl[51] br[51] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_52 bl[52] br[52] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_53 bl[53] br[53] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_54 bl[54] br[54] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_55 bl[55] br[55] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_56 bl[56] br[56] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_57 bl[57] br[57] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_58 bl[58] br[58] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_59 bl[59] br[59] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_60 bl[60] br[60] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_61 bl[61] br[61] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_62 bl[62] br[62] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_232_63 bl[63] br[63] vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xcell_233_0 bl[0] br[0] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_1 bl[1] br[1] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_2 bl[2] br[2] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_3 bl[3] br[3] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_4 bl[4] br[4] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_5 bl[5] br[5] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_6 bl[6] br[6] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_7 bl[7] br[7] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_8 bl[8] br[8] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_9 bl[9] br[9] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_10 bl[10] br[10] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_11 bl[11] br[11] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_12 bl[12] br[12] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_13 bl[13] br[13] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_14 bl[14] br[14] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_15 bl[15] br[15] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_16 bl[16] br[16] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_17 bl[17] br[17] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_18 bl[18] br[18] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_19 bl[19] br[19] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_20 bl[20] br[20] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_21 bl[21] br[21] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_22 bl[22] br[22] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_23 bl[23] br[23] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_24 bl[24] br[24] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_25 bl[25] br[25] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_26 bl[26] br[26] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_27 bl[27] br[27] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_28 bl[28] br[28] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_29 bl[29] br[29] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_30 bl[30] br[30] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_31 bl[31] br[31] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_32 bl[32] br[32] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_33 bl[33] br[33] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_34 bl[34] br[34] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_35 bl[35] br[35] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_36 bl[36] br[36] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_37 bl[37] br[37] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_38 bl[38] br[38] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_39 bl[39] br[39] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_40 bl[40] br[40] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_41 bl[41] br[41] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_42 bl[42] br[42] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_43 bl[43] br[43] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_44 bl[44] br[44] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_45 bl[45] br[45] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_46 bl[46] br[46] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_47 bl[47] br[47] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_48 bl[48] br[48] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_49 bl[49] br[49] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_50 bl[50] br[50] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_51 bl[51] br[51] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_52 bl[52] br[52] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_53 bl[53] br[53] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_54 bl[54] br[54] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_55 bl[55] br[55] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_56 bl[56] br[56] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_57 bl[57] br[57] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_58 bl[58] br[58] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_59 bl[59] br[59] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_60 bl[60] br[60] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_61 bl[61] br[61] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_62 bl[62] br[62] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_233_63 bl[63] br[63] vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xcell_234_0 bl[0] br[0] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_1 bl[1] br[1] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_2 bl[2] br[2] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_3 bl[3] br[3] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_4 bl[4] br[4] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_5 bl[5] br[5] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_6 bl[6] br[6] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_7 bl[7] br[7] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_8 bl[8] br[8] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_9 bl[9] br[9] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_10 bl[10] br[10] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_11 bl[11] br[11] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_12 bl[12] br[12] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_13 bl[13] br[13] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_14 bl[14] br[14] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_15 bl[15] br[15] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_16 bl[16] br[16] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_17 bl[17] br[17] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_18 bl[18] br[18] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_19 bl[19] br[19] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_20 bl[20] br[20] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_21 bl[21] br[21] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_22 bl[22] br[22] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_23 bl[23] br[23] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_24 bl[24] br[24] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_25 bl[25] br[25] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_26 bl[26] br[26] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_27 bl[27] br[27] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_28 bl[28] br[28] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_29 bl[29] br[29] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_30 bl[30] br[30] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_31 bl[31] br[31] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_32 bl[32] br[32] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_33 bl[33] br[33] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_34 bl[34] br[34] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_35 bl[35] br[35] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_36 bl[36] br[36] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_37 bl[37] br[37] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_38 bl[38] br[38] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_39 bl[39] br[39] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_40 bl[40] br[40] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_41 bl[41] br[41] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_42 bl[42] br[42] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_43 bl[43] br[43] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_44 bl[44] br[44] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_45 bl[45] br[45] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_46 bl[46] br[46] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_47 bl[47] br[47] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_48 bl[48] br[48] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_49 bl[49] br[49] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_50 bl[50] br[50] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_51 bl[51] br[51] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_52 bl[52] br[52] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_53 bl[53] br[53] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_54 bl[54] br[54] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_55 bl[55] br[55] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_56 bl[56] br[56] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_57 bl[57] br[57] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_58 bl[58] br[58] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_59 bl[59] br[59] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_60 bl[60] br[60] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_61 bl[61] br[61] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_62 bl[62] br[62] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_234_63 bl[63] br[63] vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xcell_235_0 bl[0] br[0] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_1 bl[1] br[1] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_2 bl[2] br[2] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_3 bl[3] br[3] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_4 bl[4] br[4] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_5 bl[5] br[5] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_6 bl[6] br[6] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_7 bl[7] br[7] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_8 bl[8] br[8] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_9 bl[9] br[9] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_10 bl[10] br[10] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_11 bl[11] br[11] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_12 bl[12] br[12] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_13 bl[13] br[13] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_14 bl[14] br[14] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_15 bl[15] br[15] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_16 bl[16] br[16] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_17 bl[17] br[17] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_18 bl[18] br[18] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_19 bl[19] br[19] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_20 bl[20] br[20] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_21 bl[21] br[21] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_22 bl[22] br[22] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_23 bl[23] br[23] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_24 bl[24] br[24] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_25 bl[25] br[25] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_26 bl[26] br[26] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_27 bl[27] br[27] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_28 bl[28] br[28] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_29 bl[29] br[29] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_30 bl[30] br[30] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_31 bl[31] br[31] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_32 bl[32] br[32] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_33 bl[33] br[33] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_34 bl[34] br[34] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_35 bl[35] br[35] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_36 bl[36] br[36] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_37 bl[37] br[37] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_38 bl[38] br[38] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_39 bl[39] br[39] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_40 bl[40] br[40] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_41 bl[41] br[41] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_42 bl[42] br[42] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_43 bl[43] br[43] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_44 bl[44] br[44] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_45 bl[45] br[45] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_46 bl[46] br[46] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_47 bl[47] br[47] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_48 bl[48] br[48] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_49 bl[49] br[49] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_50 bl[50] br[50] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_51 bl[51] br[51] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_52 bl[52] br[52] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_53 bl[53] br[53] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_54 bl[54] br[54] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_55 bl[55] br[55] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_56 bl[56] br[56] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_57 bl[57] br[57] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_58 bl[58] br[58] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_59 bl[59] br[59] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_60 bl[60] br[60] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_61 bl[61] br[61] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_62 bl[62] br[62] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_235_63 bl[63] br[63] vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xcell_236_0 bl[0] br[0] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_1 bl[1] br[1] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_2 bl[2] br[2] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_3 bl[3] br[3] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_4 bl[4] br[4] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_5 bl[5] br[5] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_6 bl[6] br[6] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_7 bl[7] br[7] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_8 bl[8] br[8] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_9 bl[9] br[9] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_10 bl[10] br[10] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_11 bl[11] br[11] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_12 bl[12] br[12] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_13 bl[13] br[13] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_14 bl[14] br[14] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_15 bl[15] br[15] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_16 bl[16] br[16] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_17 bl[17] br[17] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_18 bl[18] br[18] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_19 bl[19] br[19] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_20 bl[20] br[20] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_21 bl[21] br[21] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_22 bl[22] br[22] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_23 bl[23] br[23] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_24 bl[24] br[24] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_25 bl[25] br[25] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_26 bl[26] br[26] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_27 bl[27] br[27] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_28 bl[28] br[28] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_29 bl[29] br[29] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_30 bl[30] br[30] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_31 bl[31] br[31] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_32 bl[32] br[32] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_33 bl[33] br[33] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_34 bl[34] br[34] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_35 bl[35] br[35] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_36 bl[36] br[36] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_37 bl[37] br[37] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_38 bl[38] br[38] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_39 bl[39] br[39] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_40 bl[40] br[40] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_41 bl[41] br[41] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_42 bl[42] br[42] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_43 bl[43] br[43] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_44 bl[44] br[44] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_45 bl[45] br[45] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_46 bl[46] br[46] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_47 bl[47] br[47] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_48 bl[48] br[48] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_49 bl[49] br[49] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_50 bl[50] br[50] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_51 bl[51] br[51] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_52 bl[52] br[52] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_53 bl[53] br[53] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_54 bl[54] br[54] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_55 bl[55] br[55] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_56 bl[56] br[56] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_57 bl[57] br[57] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_58 bl[58] br[58] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_59 bl[59] br[59] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_60 bl[60] br[60] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_61 bl[61] br[61] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_62 bl[62] br[62] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_236_63 bl[63] br[63] vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xcell_237_0 bl[0] br[0] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_1 bl[1] br[1] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_2 bl[2] br[2] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_3 bl[3] br[3] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_4 bl[4] br[4] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_5 bl[5] br[5] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_6 bl[6] br[6] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_7 bl[7] br[7] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_8 bl[8] br[8] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_9 bl[9] br[9] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_10 bl[10] br[10] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_11 bl[11] br[11] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_12 bl[12] br[12] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_13 bl[13] br[13] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_14 bl[14] br[14] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_15 bl[15] br[15] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_16 bl[16] br[16] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_17 bl[17] br[17] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_18 bl[18] br[18] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_19 bl[19] br[19] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_20 bl[20] br[20] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_21 bl[21] br[21] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_22 bl[22] br[22] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_23 bl[23] br[23] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_24 bl[24] br[24] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_25 bl[25] br[25] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_26 bl[26] br[26] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_27 bl[27] br[27] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_28 bl[28] br[28] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_29 bl[29] br[29] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_30 bl[30] br[30] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_31 bl[31] br[31] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_32 bl[32] br[32] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_33 bl[33] br[33] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_34 bl[34] br[34] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_35 bl[35] br[35] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_36 bl[36] br[36] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_37 bl[37] br[37] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_38 bl[38] br[38] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_39 bl[39] br[39] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_40 bl[40] br[40] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_41 bl[41] br[41] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_42 bl[42] br[42] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_43 bl[43] br[43] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_44 bl[44] br[44] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_45 bl[45] br[45] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_46 bl[46] br[46] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_47 bl[47] br[47] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_48 bl[48] br[48] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_49 bl[49] br[49] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_50 bl[50] br[50] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_51 bl[51] br[51] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_52 bl[52] br[52] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_53 bl[53] br[53] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_54 bl[54] br[54] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_55 bl[55] br[55] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_56 bl[56] br[56] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_57 bl[57] br[57] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_58 bl[58] br[58] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_59 bl[59] br[59] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_60 bl[60] br[60] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_61 bl[61] br[61] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_62 bl[62] br[62] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_237_63 bl[63] br[63] vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xcell_238_0 bl[0] br[0] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_1 bl[1] br[1] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_2 bl[2] br[2] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_3 bl[3] br[3] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_4 bl[4] br[4] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_5 bl[5] br[5] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_6 bl[6] br[6] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_7 bl[7] br[7] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_8 bl[8] br[8] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_9 bl[9] br[9] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_10 bl[10] br[10] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_11 bl[11] br[11] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_12 bl[12] br[12] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_13 bl[13] br[13] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_14 bl[14] br[14] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_15 bl[15] br[15] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_16 bl[16] br[16] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_17 bl[17] br[17] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_18 bl[18] br[18] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_19 bl[19] br[19] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_20 bl[20] br[20] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_21 bl[21] br[21] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_22 bl[22] br[22] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_23 bl[23] br[23] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_24 bl[24] br[24] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_25 bl[25] br[25] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_26 bl[26] br[26] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_27 bl[27] br[27] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_28 bl[28] br[28] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_29 bl[29] br[29] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_30 bl[30] br[30] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_31 bl[31] br[31] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_32 bl[32] br[32] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_33 bl[33] br[33] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_34 bl[34] br[34] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_35 bl[35] br[35] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_36 bl[36] br[36] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_37 bl[37] br[37] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_38 bl[38] br[38] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_39 bl[39] br[39] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_40 bl[40] br[40] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_41 bl[41] br[41] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_42 bl[42] br[42] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_43 bl[43] br[43] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_44 bl[44] br[44] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_45 bl[45] br[45] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_46 bl[46] br[46] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_47 bl[47] br[47] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_48 bl[48] br[48] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_49 bl[49] br[49] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_50 bl[50] br[50] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_51 bl[51] br[51] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_52 bl[52] br[52] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_53 bl[53] br[53] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_54 bl[54] br[54] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_55 bl[55] br[55] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_56 bl[56] br[56] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_57 bl[57] br[57] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_58 bl[58] br[58] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_59 bl[59] br[59] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_60 bl[60] br[60] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_61 bl[61] br[61] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_62 bl[62] br[62] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_238_63 bl[63] br[63] vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xcell_239_0 bl[0] br[0] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_1 bl[1] br[1] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_2 bl[2] br[2] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_3 bl[3] br[3] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_4 bl[4] br[4] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_5 bl[5] br[5] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_6 bl[6] br[6] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_7 bl[7] br[7] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_8 bl[8] br[8] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_9 bl[9] br[9] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_10 bl[10] br[10] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_11 bl[11] br[11] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_12 bl[12] br[12] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_13 bl[13] br[13] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_14 bl[14] br[14] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_15 bl[15] br[15] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_16 bl[16] br[16] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_17 bl[17] br[17] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_18 bl[18] br[18] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_19 bl[19] br[19] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_20 bl[20] br[20] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_21 bl[21] br[21] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_22 bl[22] br[22] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_23 bl[23] br[23] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_24 bl[24] br[24] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_25 bl[25] br[25] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_26 bl[26] br[26] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_27 bl[27] br[27] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_28 bl[28] br[28] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_29 bl[29] br[29] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_30 bl[30] br[30] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_31 bl[31] br[31] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_32 bl[32] br[32] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_33 bl[33] br[33] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_34 bl[34] br[34] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_35 bl[35] br[35] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_36 bl[36] br[36] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_37 bl[37] br[37] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_38 bl[38] br[38] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_39 bl[39] br[39] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_40 bl[40] br[40] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_41 bl[41] br[41] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_42 bl[42] br[42] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_43 bl[43] br[43] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_44 bl[44] br[44] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_45 bl[45] br[45] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_46 bl[46] br[46] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_47 bl[47] br[47] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_48 bl[48] br[48] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_49 bl[49] br[49] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_50 bl[50] br[50] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_51 bl[51] br[51] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_52 bl[52] br[52] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_53 bl[53] br[53] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_54 bl[54] br[54] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_55 bl[55] br[55] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_56 bl[56] br[56] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_57 bl[57] br[57] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_58 bl[58] br[58] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_59 bl[59] br[59] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_60 bl[60] br[60] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_61 bl[61] br[61] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_62 bl[62] br[62] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_239_63 bl[63] br[63] vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xcell_240_0 bl[0] br[0] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_1 bl[1] br[1] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_2 bl[2] br[2] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_3 bl[3] br[3] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_4 bl[4] br[4] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_5 bl[5] br[5] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_6 bl[6] br[6] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_7 bl[7] br[7] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_8 bl[8] br[8] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_9 bl[9] br[9] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_10 bl[10] br[10] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_11 bl[11] br[11] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_12 bl[12] br[12] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_13 bl[13] br[13] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_14 bl[14] br[14] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_15 bl[15] br[15] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_16 bl[16] br[16] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_17 bl[17] br[17] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_18 bl[18] br[18] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_19 bl[19] br[19] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_20 bl[20] br[20] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_21 bl[21] br[21] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_22 bl[22] br[22] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_23 bl[23] br[23] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_24 bl[24] br[24] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_25 bl[25] br[25] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_26 bl[26] br[26] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_27 bl[27] br[27] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_28 bl[28] br[28] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_29 bl[29] br[29] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_30 bl[30] br[30] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_31 bl[31] br[31] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_32 bl[32] br[32] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_33 bl[33] br[33] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_34 bl[34] br[34] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_35 bl[35] br[35] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_36 bl[36] br[36] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_37 bl[37] br[37] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_38 bl[38] br[38] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_39 bl[39] br[39] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_40 bl[40] br[40] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_41 bl[41] br[41] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_42 bl[42] br[42] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_43 bl[43] br[43] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_44 bl[44] br[44] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_45 bl[45] br[45] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_46 bl[46] br[46] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_47 bl[47] br[47] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_48 bl[48] br[48] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_49 bl[49] br[49] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_50 bl[50] br[50] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_51 bl[51] br[51] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_52 bl[52] br[52] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_53 bl[53] br[53] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_54 bl[54] br[54] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_55 bl[55] br[55] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_56 bl[56] br[56] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_57 bl[57] br[57] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_58 bl[58] br[58] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_59 bl[59] br[59] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_60 bl[60] br[60] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_61 bl[61] br[61] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_62 bl[62] br[62] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_240_63 bl[63] br[63] vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xcell_241_0 bl[0] br[0] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_1 bl[1] br[1] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_2 bl[2] br[2] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_3 bl[3] br[3] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_4 bl[4] br[4] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_5 bl[5] br[5] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_6 bl[6] br[6] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_7 bl[7] br[7] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_8 bl[8] br[8] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_9 bl[9] br[9] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_10 bl[10] br[10] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_11 bl[11] br[11] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_12 bl[12] br[12] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_13 bl[13] br[13] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_14 bl[14] br[14] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_15 bl[15] br[15] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_16 bl[16] br[16] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_17 bl[17] br[17] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_18 bl[18] br[18] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_19 bl[19] br[19] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_20 bl[20] br[20] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_21 bl[21] br[21] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_22 bl[22] br[22] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_23 bl[23] br[23] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_24 bl[24] br[24] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_25 bl[25] br[25] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_26 bl[26] br[26] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_27 bl[27] br[27] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_28 bl[28] br[28] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_29 bl[29] br[29] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_30 bl[30] br[30] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_31 bl[31] br[31] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_32 bl[32] br[32] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_33 bl[33] br[33] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_34 bl[34] br[34] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_35 bl[35] br[35] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_36 bl[36] br[36] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_37 bl[37] br[37] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_38 bl[38] br[38] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_39 bl[39] br[39] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_40 bl[40] br[40] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_41 bl[41] br[41] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_42 bl[42] br[42] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_43 bl[43] br[43] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_44 bl[44] br[44] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_45 bl[45] br[45] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_46 bl[46] br[46] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_47 bl[47] br[47] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_48 bl[48] br[48] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_49 bl[49] br[49] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_50 bl[50] br[50] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_51 bl[51] br[51] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_52 bl[52] br[52] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_53 bl[53] br[53] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_54 bl[54] br[54] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_55 bl[55] br[55] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_56 bl[56] br[56] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_57 bl[57] br[57] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_58 bl[58] br[58] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_59 bl[59] br[59] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_60 bl[60] br[60] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_61 bl[61] br[61] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_62 bl[62] br[62] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_241_63 bl[63] br[63] vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xcell_242_0 bl[0] br[0] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_1 bl[1] br[1] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_2 bl[2] br[2] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_3 bl[3] br[3] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_4 bl[4] br[4] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_5 bl[5] br[5] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_6 bl[6] br[6] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_7 bl[7] br[7] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_8 bl[8] br[8] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_9 bl[9] br[9] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_10 bl[10] br[10] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_11 bl[11] br[11] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_12 bl[12] br[12] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_13 bl[13] br[13] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_14 bl[14] br[14] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_15 bl[15] br[15] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_16 bl[16] br[16] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_17 bl[17] br[17] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_18 bl[18] br[18] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_19 bl[19] br[19] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_20 bl[20] br[20] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_21 bl[21] br[21] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_22 bl[22] br[22] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_23 bl[23] br[23] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_24 bl[24] br[24] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_25 bl[25] br[25] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_26 bl[26] br[26] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_27 bl[27] br[27] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_28 bl[28] br[28] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_29 bl[29] br[29] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_30 bl[30] br[30] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_31 bl[31] br[31] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_32 bl[32] br[32] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_33 bl[33] br[33] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_34 bl[34] br[34] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_35 bl[35] br[35] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_36 bl[36] br[36] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_37 bl[37] br[37] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_38 bl[38] br[38] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_39 bl[39] br[39] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_40 bl[40] br[40] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_41 bl[41] br[41] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_42 bl[42] br[42] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_43 bl[43] br[43] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_44 bl[44] br[44] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_45 bl[45] br[45] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_46 bl[46] br[46] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_47 bl[47] br[47] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_48 bl[48] br[48] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_49 bl[49] br[49] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_50 bl[50] br[50] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_51 bl[51] br[51] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_52 bl[52] br[52] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_53 bl[53] br[53] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_54 bl[54] br[54] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_55 bl[55] br[55] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_56 bl[56] br[56] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_57 bl[57] br[57] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_58 bl[58] br[58] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_59 bl[59] br[59] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_60 bl[60] br[60] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_61 bl[61] br[61] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_62 bl[62] br[62] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_242_63 bl[63] br[63] vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xcell_243_0 bl[0] br[0] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_1 bl[1] br[1] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_2 bl[2] br[2] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_3 bl[3] br[3] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_4 bl[4] br[4] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_5 bl[5] br[5] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_6 bl[6] br[6] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_7 bl[7] br[7] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_8 bl[8] br[8] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_9 bl[9] br[9] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_10 bl[10] br[10] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_11 bl[11] br[11] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_12 bl[12] br[12] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_13 bl[13] br[13] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_14 bl[14] br[14] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_15 bl[15] br[15] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_16 bl[16] br[16] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_17 bl[17] br[17] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_18 bl[18] br[18] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_19 bl[19] br[19] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_20 bl[20] br[20] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_21 bl[21] br[21] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_22 bl[22] br[22] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_23 bl[23] br[23] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_24 bl[24] br[24] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_25 bl[25] br[25] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_26 bl[26] br[26] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_27 bl[27] br[27] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_28 bl[28] br[28] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_29 bl[29] br[29] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_30 bl[30] br[30] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_31 bl[31] br[31] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_32 bl[32] br[32] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_33 bl[33] br[33] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_34 bl[34] br[34] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_35 bl[35] br[35] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_36 bl[36] br[36] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_37 bl[37] br[37] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_38 bl[38] br[38] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_39 bl[39] br[39] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_40 bl[40] br[40] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_41 bl[41] br[41] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_42 bl[42] br[42] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_43 bl[43] br[43] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_44 bl[44] br[44] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_45 bl[45] br[45] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_46 bl[46] br[46] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_47 bl[47] br[47] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_48 bl[48] br[48] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_49 bl[49] br[49] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_50 bl[50] br[50] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_51 bl[51] br[51] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_52 bl[52] br[52] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_53 bl[53] br[53] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_54 bl[54] br[54] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_55 bl[55] br[55] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_56 bl[56] br[56] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_57 bl[57] br[57] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_58 bl[58] br[58] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_59 bl[59] br[59] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_60 bl[60] br[60] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_61 bl[61] br[61] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_62 bl[62] br[62] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_243_63 bl[63] br[63] vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xcell_244_0 bl[0] br[0] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_1 bl[1] br[1] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_2 bl[2] br[2] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_3 bl[3] br[3] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_4 bl[4] br[4] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_5 bl[5] br[5] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_6 bl[6] br[6] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_7 bl[7] br[7] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_8 bl[8] br[8] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_9 bl[9] br[9] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_10 bl[10] br[10] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_11 bl[11] br[11] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_12 bl[12] br[12] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_13 bl[13] br[13] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_14 bl[14] br[14] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_15 bl[15] br[15] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_16 bl[16] br[16] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_17 bl[17] br[17] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_18 bl[18] br[18] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_19 bl[19] br[19] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_20 bl[20] br[20] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_21 bl[21] br[21] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_22 bl[22] br[22] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_23 bl[23] br[23] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_24 bl[24] br[24] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_25 bl[25] br[25] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_26 bl[26] br[26] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_27 bl[27] br[27] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_28 bl[28] br[28] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_29 bl[29] br[29] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_30 bl[30] br[30] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_31 bl[31] br[31] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_32 bl[32] br[32] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_33 bl[33] br[33] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_34 bl[34] br[34] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_35 bl[35] br[35] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_36 bl[36] br[36] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_37 bl[37] br[37] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_38 bl[38] br[38] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_39 bl[39] br[39] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_40 bl[40] br[40] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_41 bl[41] br[41] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_42 bl[42] br[42] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_43 bl[43] br[43] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_44 bl[44] br[44] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_45 bl[45] br[45] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_46 bl[46] br[46] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_47 bl[47] br[47] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_48 bl[48] br[48] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_49 bl[49] br[49] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_50 bl[50] br[50] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_51 bl[51] br[51] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_52 bl[52] br[52] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_53 bl[53] br[53] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_54 bl[54] br[54] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_55 bl[55] br[55] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_56 bl[56] br[56] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_57 bl[57] br[57] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_58 bl[58] br[58] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_59 bl[59] br[59] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_60 bl[60] br[60] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_61 bl[61] br[61] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_62 bl[62] br[62] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_244_63 bl[63] br[63] vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xcell_245_0 bl[0] br[0] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_1 bl[1] br[1] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_2 bl[2] br[2] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_3 bl[3] br[3] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_4 bl[4] br[4] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_5 bl[5] br[5] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_6 bl[6] br[6] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_7 bl[7] br[7] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_8 bl[8] br[8] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_9 bl[9] br[9] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_10 bl[10] br[10] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_11 bl[11] br[11] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_12 bl[12] br[12] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_13 bl[13] br[13] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_14 bl[14] br[14] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_15 bl[15] br[15] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_16 bl[16] br[16] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_17 bl[17] br[17] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_18 bl[18] br[18] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_19 bl[19] br[19] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_20 bl[20] br[20] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_21 bl[21] br[21] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_22 bl[22] br[22] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_23 bl[23] br[23] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_24 bl[24] br[24] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_25 bl[25] br[25] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_26 bl[26] br[26] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_27 bl[27] br[27] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_28 bl[28] br[28] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_29 bl[29] br[29] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_30 bl[30] br[30] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_31 bl[31] br[31] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_32 bl[32] br[32] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_33 bl[33] br[33] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_34 bl[34] br[34] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_35 bl[35] br[35] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_36 bl[36] br[36] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_37 bl[37] br[37] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_38 bl[38] br[38] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_39 bl[39] br[39] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_40 bl[40] br[40] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_41 bl[41] br[41] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_42 bl[42] br[42] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_43 bl[43] br[43] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_44 bl[44] br[44] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_45 bl[45] br[45] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_46 bl[46] br[46] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_47 bl[47] br[47] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_48 bl[48] br[48] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_49 bl[49] br[49] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_50 bl[50] br[50] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_51 bl[51] br[51] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_52 bl[52] br[52] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_53 bl[53] br[53] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_54 bl[54] br[54] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_55 bl[55] br[55] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_56 bl[56] br[56] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_57 bl[57] br[57] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_58 bl[58] br[58] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_59 bl[59] br[59] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_60 bl[60] br[60] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_61 bl[61] br[61] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_62 bl[62] br[62] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_245_63 bl[63] br[63] vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xcell_246_0 bl[0] br[0] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_1 bl[1] br[1] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_2 bl[2] br[2] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_3 bl[3] br[3] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_4 bl[4] br[4] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_5 bl[5] br[5] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_6 bl[6] br[6] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_7 bl[7] br[7] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_8 bl[8] br[8] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_9 bl[9] br[9] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_10 bl[10] br[10] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_11 bl[11] br[11] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_12 bl[12] br[12] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_13 bl[13] br[13] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_14 bl[14] br[14] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_15 bl[15] br[15] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_16 bl[16] br[16] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_17 bl[17] br[17] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_18 bl[18] br[18] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_19 bl[19] br[19] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_20 bl[20] br[20] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_21 bl[21] br[21] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_22 bl[22] br[22] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_23 bl[23] br[23] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_24 bl[24] br[24] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_25 bl[25] br[25] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_26 bl[26] br[26] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_27 bl[27] br[27] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_28 bl[28] br[28] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_29 bl[29] br[29] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_30 bl[30] br[30] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_31 bl[31] br[31] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_32 bl[32] br[32] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_33 bl[33] br[33] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_34 bl[34] br[34] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_35 bl[35] br[35] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_36 bl[36] br[36] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_37 bl[37] br[37] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_38 bl[38] br[38] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_39 bl[39] br[39] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_40 bl[40] br[40] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_41 bl[41] br[41] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_42 bl[42] br[42] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_43 bl[43] br[43] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_44 bl[44] br[44] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_45 bl[45] br[45] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_46 bl[46] br[46] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_47 bl[47] br[47] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_48 bl[48] br[48] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_49 bl[49] br[49] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_50 bl[50] br[50] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_51 bl[51] br[51] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_52 bl[52] br[52] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_53 bl[53] br[53] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_54 bl[54] br[54] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_55 bl[55] br[55] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_56 bl[56] br[56] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_57 bl[57] br[57] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_58 bl[58] br[58] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_59 bl[59] br[59] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_60 bl[60] br[60] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_61 bl[61] br[61] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_62 bl[62] br[62] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_246_63 bl[63] br[63] vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xcell_247_0 bl[0] br[0] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_1 bl[1] br[1] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_2 bl[2] br[2] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_3 bl[3] br[3] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_4 bl[4] br[4] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_5 bl[5] br[5] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_6 bl[6] br[6] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_7 bl[7] br[7] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_8 bl[8] br[8] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_9 bl[9] br[9] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_10 bl[10] br[10] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_11 bl[11] br[11] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_12 bl[12] br[12] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_13 bl[13] br[13] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_14 bl[14] br[14] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_15 bl[15] br[15] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_16 bl[16] br[16] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_17 bl[17] br[17] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_18 bl[18] br[18] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_19 bl[19] br[19] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_20 bl[20] br[20] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_21 bl[21] br[21] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_22 bl[22] br[22] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_23 bl[23] br[23] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_24 bl[24] br[24] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_25 bl[25] br[25] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_26 bl[26] br[26] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_27 bl[27] br[27] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_28 bl[28] br[28] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_29 bl[29] br[29] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_30 bl[30] br[30] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_31 bl[31] br[31] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_32 bl[32] br[32] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_33 bl[33] br[33] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_34 bl[34] br[34] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_35 bl[35] br[35] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_36 bl[36] br[36] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_37 bl[37] br[37] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_38 bl[38] br[38] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_39 bl[39] br[39] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_40 bl[40] br[40] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_41 bl[41] br[41] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_42 bl[42] br[42] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_43 bl[43] br[43] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_44 bl[44] br[44] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_45 bl[45] br[45] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_46 bl[46] br[46] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_47 bl[47] br[47] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_48 bl[48] br[48] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_49 bl[49] br[49] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_50 bl[50] br[50] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_51 bl[51] br[51] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_52 bl[52] br[52] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_53 bl[53] br[53] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_54 bl[54] br[54] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_55 bl[55] br[55] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_56 bl[56] br[56] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_57 bl[57] br[57] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_58 bl[58] br[58] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_59 bl[59] br[59] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_60 bl[60] br[60] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_61 bl[61] br[61] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_62 bl[62] br[62] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_247_63 bl[63] br[63] vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xcell_248_0 bl[0] br[0] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_1 bl[1] br[1] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_2 bl[2] br[2] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_3 bl[3] br[3] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_4 bl[4] br[4] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_5 bl[5] br[5] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_6 bl[6] br[6] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_7 bl[7] br[7] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_8 bl[8] br[8] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_9 bl[9] br[9] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_10 bl[10] br[10] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_11 bl[11] br[11] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_12 bl[12] br[12] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_13 bl[13] br[13] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_14 bl[14] br[14] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_15 bl[15] br[15] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_16 bl[16] br[16] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_17 bl[17] br[17] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_18 bl[18] br[18] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_19 bl[19] br[19] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_20 bl[20] br[20] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_21 bl[21] br[21] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_22 bl[22] br[22] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_23 bl[23] br[23] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_24 bl[24] br[24] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_25 bl[25] br[25] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_26 bl[26] br[26] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_27 bl[27] br[27] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_28 bl[28] br[28] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_29 bl[29] br[29] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_30 bl[30] br[30] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_31 bl[31] br[31] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_32 bl[32] br[32] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_33 bl[33] br[33] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_34 bl[34] br[34] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_35 bl[35] br[35] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_36 bl[36] br[36] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_37 bl[37] br[37] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_38 bl[38] br[38] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_39 bl[39] br[39] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_40 bl[40] br[40] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_41 bl[41] br[41] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_42 bl[42] br[42] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_43 bl[43] br[43] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_44 bl[44] br[44] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_45 bl[45] br[45] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_46 bl[46] br[46] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_47 bl[47] br[47] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_48 bl[48] br[48] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_49 bl[49] br[49] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_50 bl[50] br[50] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_51 bl[51] br[51] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_52 bl[52] br[52] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_53 bl[53] br[53] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_54 bl[54] br[54] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_55 bl[55] br[55] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_56 bl[56] br[56] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_57 bl[57] br[57] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_58 bl[58] br[58] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_59 bl[59] br[59] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_60 bl[60] br[60] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_61 bl[61] br[61] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_62 bl[62] br[62] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_248_63 bl[63] br[63] vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xcell_249_0 bl[0] br[0] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_1 bl[1] br[1] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_2 bl[2] br[2] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_3 bl[3] br[3] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_4 bl[4] br[4] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_5 bl[5] br[5] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_6 bl[6] br[6] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_7 bl[7] br[7] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_8 bl[8] br[8] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_9 bl[9] br[9] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_10 bl[10] br[10] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_11 bl[11] br[11] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_12 bl[12] br[12] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_13 bl[13] br[13] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_14 bl[14] br[14] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_15 bl[15] br[15] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_16 bl[16] br[16] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_17 bl[17] br[17] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_18 bl[18] br[18] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_19 bl[19] br[19] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_20 bl[20] br[20] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_21 bl[21] br[21] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_22 bl[22] br[22] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_23 bl[23] br[23] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_24 bl[24] br[24] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_25 bl[25] br[25] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_26 bl[26] br[26] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_27 bl[27] br[27] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_28 bl[28] br[28] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_29 bl[29] br[29] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_30 bl[30] br[30] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_31 bl[31] br[31] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_32 bl[32] br[32] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_33 bl[33] br[33] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_34 bl[34] br[34] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_35 bl[35] br[35] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_36 bl[36] br[36] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_37 bl[37] br[37] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_38 bl[38] br[38] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_39 bl[39] br[39] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_40 bl[40] br[40] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_41 bl[41] br[41] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_42 bl[42] br[42] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_43 bl[43] br[43] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_44 bl[44] br[44] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_45 bl[45] br[45] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_46 bl[46] br[46] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_47 bl[47] br[47] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_48 bl[48] br[48] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_49 bl[49] br[49] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_50 bl[50] br[50] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_51 bl[51] br[51] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_52 bl[52] br[52] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_53 bl[53] br[53] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_54 bl[54] br[54] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_55 bl[55] br[55] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_56 bl[56] br[56] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_57 bl[57] br[57] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_58 bl[58] br[58] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_59 bl[59] br[59] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_60 bl[60] br[60] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_61 bl[61] br[61] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_62 bl[62] br[62] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_249_63 bl[63] br[63] vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xcell_250_0 bl[0] br[0] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_1 bl[1] br[1] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_2 bl[2] br[2] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_3 bl[3] br[3] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_4 bl[4] br[4] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_5 bl[5] br[5] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_6 bl[6] br[6] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_7 bl[7] br[7] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_8 bl[8] br[8] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_9 bl[9] br[9] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_10 bl[10] br[10] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_11 bl[11] br[11] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_12 bl[12] br[12] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_13 bl[13] br[13] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_14 bl[14] br[14] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_15 bl[15] br[15] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_16 bl[16] br[16] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_17 bl[17] br[17] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_18 bl[18] br[18] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_19 bl[19] br[19] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_20 bl[20] br[20] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_21 bl[21] br[21] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_22 bl[22] br[22] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_23 bl[23] br[23] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_24 bl[24] br[24] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_25 bl[25] br[25] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_26 bl[26] br[26] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_27 bl[27] br[27] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_28 bl[28] br[28] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_29 bl[29] br[29] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_30 bl[30] br[30] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_31 bl[31] br[31] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_32 bl[32] br[32] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_33 bl[33] br[33] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_34 bl[34] br[34] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_35 bl[35] br[35] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_36 bl[36] br[36] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_37 bl[37] br[37] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_38 bl[38] br[38] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_39 bl[39] br[39] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_40 bl[40] br[40] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_41 bl[41] br[41] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_42 bl[42] br[42] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_43 bl[43] br[43] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_44 bl[44] br[44] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_45 bl[45] br[45] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_46 bl[46] br[46] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_47 bl[47] br[47] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_48 bl[48] br[48] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_49 bl[49] br[49] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_50 bl[50] br[50] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_51 bl[51] br[51] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_52 bl[52] br[52] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_53 bl[53] br[53] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_54 bl[54] br[54] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_55 bl[55] br[55] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_56 bl[56] br[56] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_57 bl[57] br[57] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_58 bl[58] br[58] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_59 bl[59] br[59] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_60 bl[60] br[60] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_61 bl[61] br[61] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_62 bl[62] br[62] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_250_63 bl[63] br[63] vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xcell_251_0 bl[0] br[0] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_1 bl[1] br[1] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_2 bl[2] br[2] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_3 bl[3] br[3] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_4 bl[4] br[4] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_5 bl[5] br[5] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_6 bl[6] br[6] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_7 bl[7] br[7] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_8 bl[8] br[8] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_9 bl[9] br[9] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_10 bl[10] br[10] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_11 bl[11] br[11] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_12 bl[12] br[12] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_13 bl[13] br[13] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_14 bl[14] br[14] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_15 bl[15] br[15] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_16 bl[16] br[16] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_17 bl[17] br[17] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_18 bl[18] br[18] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_19 bl[19] br[19] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_20 bl[20] br[20] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_21 bl[21] br[21] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_22 bl[22] br[22] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_23 bl[23] br[23] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_24 bl[24] br[24] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_25 bl[25] br[25] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_26 bl[26] br[26] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_27 bl[27] br[27] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_28 bl[28] br[28] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_29 bl[29] br[29] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_30 bl[30] br[30] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_31 bl[31] br[31] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_32 bl[32] br[32] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_33 bl[33] br[33] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_34 bl[34] br[34] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_35 bl[35] br[35] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_36 bl[36] br[36] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_37 bl[37] br[37] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_38 bl[38] br[38] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_39 bl[39] br[39] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_40 bl[40] br[40] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_41 bl[41] br[41] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_42 bl[42] br[42] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_43 bl[43] br[43] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_44 bl[44] br[44] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_45 bl[45] br[45] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_46 bl[46] br[46] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_47 bl[47] br[47] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_48 bl[48] br[48] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_49 bl[49] br[49] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_50 bl[50] br[50] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_51 bl[51] br[51] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_52 bl[52] br[52] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_53 bl[53] br[53] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_54 bl[54] br[54] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_55 bl[55] br[55] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_56 bl[56] br[56] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_57 bl[57] br[57] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_58 bl[58] br[58] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_59 bl[59] br[59] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_60 bl[60] br[60] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_61 bl[61] br[61] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_62 bl[62] br[62] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_251_63 bl[63] br[63] vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xcell_252_0 bl[0] br[0] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_1 bl[1] br[1] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_2 bl[2] br[2] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_3 bl[3] br[3] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_4 bl[4] br[4] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_5 bl[5] br[5] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_6 bl[6] br[6] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_7 bl[7] br[7] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_8 bl[8] br[8] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_9 bl[9] br[9] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_10 bl[10] br[10] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_11 bl[11] br[11] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_12 bl[12] br[12] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_13 bl[13] br[13] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_14 bl[14] br[14] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_15 bl[15] br[15] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_16 bl[16] br[16] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_17 bl[17] br[17] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_18 bl[18] br[18] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_19 bl[19] br[19] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_20 bl[20] br[20] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_21 bl[21] br[21] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_22 bl[22] br[22] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_23 bl[23] br[23] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_24 bl[24] br[24] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_25 bl[25] br[25] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_26 bl[26] br[26] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_27 bl[27] br[27] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_28 bl[28] br[28] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_29 bl[29] br[29] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_30 bl[30] br[30] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_31 bl[31] br[31] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_32 bl[32] br[32] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_33 bl[33] br[33] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_34 bl[34] br[34] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_35 bl[35] br[35] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_36 bl[36] br[36] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_37 bl[37] br[37] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_38 bl[38] br[38] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_39 bl[39] br[39] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_40 bl[40] br[40] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_41 bl[41] br[41] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_42 bl[42] br[42] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_43 bl[43] br[43] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_44 bl[44] br[44] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_45 bl[45] br[45] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_46 bl[46] br[46] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_47 bl[47] br[47] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_48 bl[48] br[48] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_49 bl[49] br[49] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_50 bl[50] br[50] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_51 bl[51] br[51] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_52 bl[52] br[52] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_53 bl[53] br[53] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_54 bl[54] br[54] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_55 bl[55] br[55] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_56 bl[56] br[56] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_57 bl[57] br[57] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_58 bl[58] br[58] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_59 bl[59] br[59] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_60 bl[60] br[60] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_61 bl[61] br[61] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_62 bl[62] br[62] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_252_63 bl[63] br[63] vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xcell_253_0 bl[0] br[0] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_1 bl[1] br[1] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_2 bl[2] br[2] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_3 bl[3] br[3] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_4 bl[4] br[4] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_5 bl[5] br[5] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_6 bl[6] br[6] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_7 bl[7] br[7] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_8 bl[8] br[8] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_9 bl[9] br[9] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_10 bl[10] br[10] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_11 bl[11] br[11] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_12 bl[12] br[12] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_13 bl[13] br[13] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_14 bl[14] br[14] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_15 bl[15] br[15] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_16 bl[16] br[16] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_17 bl[17] br[17] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_18 bl[18] br[18] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_19 bl[19] br[19] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_20 bl[20] br[20] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_21 bl[21] br[21] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_22 bl[22] br[22] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_23 bl[23] br[23] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_24 bl[24] br[24] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_25 bl[25] br[25] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_26 bl[26] br[26] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_27 bl[27] br[27] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_28 bl[28] br[28] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_29 bl[29] br[29] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_30 bl[30] br[30] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_31 bl[31] br[31] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_32 bl[32] br[32] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_33 bl[33] br[33] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_34 bl[34] br[34] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_35 bl[35] br[35] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_36 bl[36] br[36] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_37 bl[37] br[37] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_38 bl[38] br[38] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_39 bl[39] br[39] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_40 bl[40] br[40] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_41 bl[41] br[41] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_42 bl[42] br[42] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_43 bl[43] br[43] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_44 bl[44] br[44] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_45 bl[45] br[45] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_46 bl[46] br[46] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_47 bl[47] br[47] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_48 bl[48] br[48] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_49 bl[49] br[49] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_50 bl[50] br[50] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_51 bl[51] br[51] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_52 bl[52] br[52] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_53 bl[53] br[53] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_54 bl[54] br[54] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_55 bl[55] br[55] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_56 bl[56] br[56] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_57 bl[57] br[57] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_58 bl[58] br[58] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_59 bl[59] br[59] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_60 bl[60] br[60] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_61 bl[61] br[61] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_62 bl[62] br[62] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_253_63 bl[63] br[63] vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xcell_254_0 bl[0] br[0] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_1 bl[1] br[1] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_2 bl[2] br[2] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_3 bl[3] br[3] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_4 bl[4] br[4] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_5 bl[5] br[5] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_6 bl[6] br[6] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_7 bl[7] br[7] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_8 bl[8] br[8] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_9 bl[9] br[9] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_10 bl[10] br[10] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_11 bl[11] br[11] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_12 bl[12] br[12] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_13 bl[13] br[13] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_14 bl[14] br[14] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_15 bl[15] br[15] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_16 bl[16] br[16] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_17 bl[17] br[17] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_18 bl[18] br[18] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_19 bl[19] br[19] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_20 bl[20] br[20] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_21 bl[21] br[21] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_22 bl[22] br[22] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_23 bl[23] br[23] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_24 bl[24] br[24] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_25 bl[25] br[25] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_26 bl[26] br[26] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_27 bl[27] br[27] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_28 bl[28] br[28] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_29 bl[29] br[29] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_30 bl[30] br[30] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_31 bl[31] br[31] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_32 bl[32] br[32] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_33 bl[33] br[33] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_34 bl[34] br[34] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_35 bl[35] br[35] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_36 bl[36] br[36] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_37 bl[37] br[37] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_38 bl[38] br[38] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_39 bl[39] br[39] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_40 bl[40] br[40] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_41 bl[41] br[41] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_42 bl[42] br[42] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_43 bl[43] br[43] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_44 bl[44] br[44] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_45 bl[45] br[45] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_46 bl[46] br[46] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_47 bl[47] br[47] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_48 bl[48] br[48] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_49 bl[49] br[49] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_50 bl[50] br[50] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_51 bl[51] br[51] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_52 bl[52] br[52] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_53 bl[53] br[53] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_54 bl[54] br[54] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_55 bl[55] br[55] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_56 bl[56] br[56] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_57 bl[57] br[57] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_58 bl[58] br[58] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_59 bl[59] br[59] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_60 bl[60] br[60] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_61 bl[61] br[61] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_62 bl[62] br[62] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_254_63 bl[63] br[63] vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xcell_255_0 bl[0] br[0] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_1 bl[1] br[1] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_2 bl[2] br[2] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_3 bl[3] br[3] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_4 bl[4] br[4] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_5 bl[5] br[5] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_6 bl[6] br[6] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_7 bl[7] br[7] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_8 bl[8] br[8] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_9 bl[9] br[9] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_10 bl[10] br[10] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_11 bl[11] br[11] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_12 bl[12] br[12] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_13 bl[13] br[13] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_14 bl[14] br[14] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_15 bl[15] br[15] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_16 bl[16] br[16] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_17 bl[17] br[17] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_18 bl[18] br[18] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_19 bl[19] br[19] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_20 bl[20] br[20] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_21 bl[21] br[21] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_22 bl[22] br[22] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_23 bl[23] br[23] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_24 bl[24] br[24] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_25 bl[25] br[25] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_26 bl[26] br[26] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_27 bl[27] br[27] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_28 bl[28] br[28] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_29 bl[29] br[29] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_30 bl[30] br[30] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_31 bl[31] br[31] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_32 bl[32] br[32] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_33 bl[33] br[33] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_34 bl[34] br[34] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_35 bl[35] br[35] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_36 bl[36] br[36] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_37 bl[37] br[37] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_38 bl[38] br[38] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_39 bl[39] br[39] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_40 bl[40] br[40] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_41 bl[41] br[41] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_42 bl[42] br[42] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_43 bl[43] br[43] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_44 bl[44] br[44] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_45 bl[45] br[45] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_46 bl[46] br[46] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_47 bl[47] br[47] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_48 bl[48] br[48] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_49 bl[49] br[49] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_50 bl[50] br[50] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_51 bl[51] br[51] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_52 bl[52] br[52] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_53 bl[53] br[53] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_54 bl[54] br[54] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_55 bl[55] br[55] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_56 bl[56] br[56] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_57 bl[57] br[57] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_58 bl[58] br[58] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_59 bl[59] br[59] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_60 bl[60] br[60] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_61 bl[61] br[61] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_62 bl[62] br[62] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xcell_255_63 bl[63] br[63] vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_0 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_0 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_1 dummy_bl dummy_br vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_1 vdd vdd vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_2 dummy_bl dummy_br vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_2 vdd vdd vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_3 dummy_bl dummy_br vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_3 vdd vdd vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_4 dummy_bl dummy_br vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_4 vdd vdd vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_5 dummy_bl dummy_br vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_5 vdd vdd vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_6 dummy_bl dummy_br vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_6 vdd vdd vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_7 dummy_bl dummy_br vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_7 vdd vdd vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_8 dummy_bl dummy_br vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_8 vdd vdd vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_9 dummy_bl dummy_br vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_9 vdd vdd vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_10 dummy_bl dummy_br vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_10 vdd vdd vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_11 dummy_bl dummy_br vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_11 vdd vdd vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_12 dummy_bl dummy_br vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_12 vdd vdd vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_13 dummy_bl dummy_br vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_13 vdd vdd vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_14 dummy_bl dummy_br vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_14 vdd vdd vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_15 dummy_bl dummy_br vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_15 vdd vdd vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_16 dummy_bl dummy_br vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_16 vdd vdd vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_17 dummy_bl dummy_br vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_17 vdd vdd vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_18 dummy_bl dummy_br vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_18 vdd vdd vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_19 dummy_bl dummy_br vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_19 vdd vdd vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_20 dummy_bl dummy_br vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_20 vdd vdd vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_21 dummy_bl dummy_br vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_21 vdd vdd vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_22 dummy_bl dummy_br vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_22 vdd vdd vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_23 dummy_bl dummy_br vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_23 vdd vdd vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_24 dummy_bl dummy_br vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_24 vdd vdd vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_25 dummy_bl dummy_br vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_25 vdd vdd vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_26 dummy_bl dummy_br vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_26 vdd vdd vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_27 dummy_bl dummy_br vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_27 vdd vdd vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_28 dummy_bl dummy_br vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_28 vdd vdd vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_29 dummy_bl dummy_br vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_29 vdd vdd vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_30 dummy_bl dummy_br vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_30 vdd vdd vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_31 dummy_bl dummy_br vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_31 vdd vdd vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_32 dummy_bl dummy_br vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_32 vdd vdd vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_33 dummy_bl dummy_br vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_33 vdd vdd vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_34 dummy_bl dummy_br vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_34 vdd vdd vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_35 dummy_bl dummy_br vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_35 vdd vdd vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_36 dummy_bl dummy_br vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_36 vdd vdd vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_37 dummy_bl dummy_br vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_37 vdd vdd vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_38 dummy_bl dummy_br vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_38 vdd vdd vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_39 dummy_bl dummy_br vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_39 vdd vdd vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_40 dummy_bl dummy_br vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_40 vdd vdd vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_41 dummy_bl dummy_br vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_41 vdd vdd vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_42 dummy_bl dummy_br vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_42 vdd vdd vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_43 dummy_bl dummy_br vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_43 vdd vdd vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_44 dummy_bl dummy_br vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_44 vdd vdd vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_45 dummy_bl dummy_br vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_45 vdd vdd vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_46 dummy_bl dummy_br vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_46 vdd vdd vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_47 dummy_bl dummy_br vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_47 vdd vdd vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_48 dummy_bl dummy_br vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_48 vdd vdd vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_49 dummy_bl dummy_br vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_49 vdd vdd vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_50 dummy_bl dummy_br vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_50 vdd vdd vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_51 dummy_bl dummy_br vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_51 vdd vdd vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_52 dummy_bl dummy_br vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_52 vdd vdd vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_53 dummy_bl dummy_br vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_53 vdd vdd vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_54 dummy_bl dummy_br vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_54 vdd vdd vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_55 dummy_bl dummy_br vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_55 vdd vdd vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_56 dummy_bl dummy_br vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_56 vdd vdd vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_57 dummy_bl dummy_br vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_57 vdd vdd vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_58 dummy_bl dummy_br vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_58 vdd vdd vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_59 dummy_bl dummy_br vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_59 vdd vdd vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_60 dummy_bl dummy_br vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_60 vdd vdd vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_61 dummy_bl dummy_br vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_61 vdd vdd vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_62 dummy_bl dummy_br vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_62 vdd vdd vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_63 dummy_bl dummy_br vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_63 vdd vdd vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_64 dummy_bl dummy_br vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_64 vdd vdd vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_65 dummy_bl dummy_br vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_65 vdd vdd vdd vss wl[64] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_66 dummy_bl dummy_br vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_66 vdd vdd vdd vss wl[65] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_67 dummy_bl dummy_br vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_67 vdd vdd vdd vss wl[66] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_68 dummy_bl dummy_br vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_68 vdd vdd vdd vss wl[67] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_69 dummy_bl dummy_br vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_69 vdd vdd vdd vss wl[68] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_70 dummy_bl dummy_br vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_70 vdd vdd vdd vss wl[69] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_71 dummy_bl dummy_br vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_71 vdd vdd vdd vss wl[70] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_72 dummy_bl dummy_br vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_72 vdd vdd vdd vss wl[71] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_73 dummy_bl dummy_br vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_73 vdd vdd vdd vss wl[72] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_74 dummy_bl dummy_br vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_74 vdd vdd vdd vss wl[73] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_75 dummy_bl dummy_br vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_75 vdd vdd vdd vss wl[74] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_76 dummy_bl dummy_br vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_76 vdd vdd vdd vss wl[75] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_77 dummy_bl dummy_br vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_77 vdd vdd vdd vss wl[76] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_78 dummy_bl dummy_br vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_78 vdd vdd vdd vss wl[77] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_79 dummy_bl dummy_br vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_79 vdd vdd vdd vss wl[78] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_80 dummy_bl dummy_br vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_80 vdd vdd vdd vss wl[79] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_81 dummy_bl dummy_br vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_81 vdd vdd vdd vss wl[80] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_82 dummy_bl dummy_br vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_82 vdd vdd vdd vss wl[81] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_83 dummy_bl dummy_br vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_83 vdd vdd vdd vss wl[82] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_84 dummy_bl dummy_br vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_84 vdd vdd vdd vss wl[83] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_85 dummy_bl dummy_br vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_85 vdd vdd vdd vss wl[84] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_86 dummy_bl dummy_br vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_86 vdd vdd vdd vss wl[85] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_87 dummy_bl dummy_br vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_87 vdd vdd vdd vss wl[86] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_88 dummy_bl dummy_br vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_88 vdd vdd vdd vss wl[87] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_89 dummy_bl dummy_br vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_89 vdd vdd vdd vss wl[88] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_90 dummy_bl dummy_br vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_90 vdd vdd vdd vss wl[89] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_91 dummy_bl dummy_br vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_91 vdd vdd vdd vss wl[90] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_92 dummy_bl dummy_br vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_92 vdd vdd vdd vss wl[91] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_93 dummy_bl dummy_br vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_93 vdd vdd vdd vss wl[92] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_94 dummy_bl dummy_br vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_94 vdd vdd vdd vss wl[93] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_95 dummy_bl dummy_br vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_95 vdd vdd vdd vss wl[94] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_96 dummy_bl dummy_br vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_96 vdd vdd vdd vss wl[95] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_97 dummy_bl dummy_br vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_97 vdd vdd vdd vss wl[96] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_98 dummy_bl dummy_br vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_98 vdd vdd vdd vss wl[97] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_99 dummy_bl dummy_br vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_99 vdd vdd vdd vss wl[98] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_100 dummy_bl dummy_br vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_100 vdd vdd vdd vss wl[99] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_101 dummy_bl dummy_br vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_101 vdd vdd vdd vss wl[100] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_102 dummy_bl dummy_br vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_102 vdd vdd vdd vss wl[101] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_103 dummy_bl dummy_br vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_103 vdd vdd vdd vss wl[102] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_104 dummy_bl dummy_br vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_104 vdd vdd vdd vss wl[103] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_105 dummy_bl dummy_br vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_105 vdd vdd vdd vss wl[104] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_106 dummy_bl dummy_br vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_106 vdd vdd vdd vss wl[105] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_107 dummy_bl dummy_br vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_107 vdd vdd vdd vss wl[106] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_108 dummy_bl dummy_br vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_108 vdd vdd vdd vss wl[107] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_109 dummy_bl dummy_br vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_109 vdd vdd vdd vss wl[108] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_110 dummy_bl dummy_br vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_110 vdd vdd vdd vss wl[109] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_111 dummy_bl dummy_br vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_111 vdd vdd vdd vss wl[110] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_112 dummy_bl dummy_br vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_112 vdd vdd vdd vss wl[111] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_113 dummy_bl dummy_br vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_113 vdd vdd vdd vss wl[112] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_114 dummy_bl dummy_br vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_114 vdd vdd vdd vss wl[113] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_115 dummy_bl dummy_br vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_115 vdd vdd vdd vss wl[114] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_116 dummy_bl dummy_br vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_116 vdd vdd vdd vss wl[115] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_117 dummy_bl dummy_br vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_117 vdd vdd vdd vss wl[116] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_118 dummy_bl dummy_br vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_118 vdd vdd vdd vss wl[117] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_119 dummy_bl dummy_br vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_119 vdd vdd vdd vss wl[118] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_120 dummy_bl dummy_br vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_120 vdd vdd vdd vss wl[119] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_121 dummy_bl dummy_br vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_121 vdd vdd vdd vss wl[120] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_122 dummy_bl dummy_br vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_122 vdd vdd vdd vss wl[121] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_123 dummy_bl dummy_br vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_123 vdd vdd vdd vss wl[122] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_124 dummy_bl dummy_br vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_124 vdd vdd vdd vss wl[123] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_125 dummy_bl dummy_br vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_125 vdd vdd vdd vss wl[124] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_126 dummy_bl dummy_br vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_126 vdd vdd vdd vss wl[125] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_127 dummy_bl dummy_br vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_127 vdd vdd vdd vss wl[126] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_128 dummy_bl dummy_br vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_128 vdd vdd vdd vss wl[127] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_129 dummy_bl dummy_br vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_129 vdd vdd vdd vss wl[128] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_130 dummy_bl dummy_br vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_130 vdd vdd vdd vss wl[129] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_131 dummy_bl dummy_br vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_131 vdd vdd vdd vss wl[130] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_132 dummy_bl dummy_br vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_132 vdd vdd vdd vss wl[131] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_133 dummy_bl dummy_br vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_133 vdd vdd vdd vss wl[132] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_134 dummy_bl dummy_br vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_134 vdd vdd vdd vss wl[133] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_135 dummy_bl dummy_br vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_135 vdd vdd vdd vss wl[134] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_136 dummy_bl dummy_br vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_136 vdd vdd vdd vss wl[135] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_137 dummy_bl dummy_br vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_137 vdd vdd vdd vss wl[136] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_138 dummy_bl dummy_br vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_138 vdd vdd vdd vss wl[137] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_139 dummy_bl dummy_br vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_139 vdd vdd vdd vss wl[138] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_140 dummy_bl dummy_br vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_140 vdd vdd vdd vss wl[139] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_141 dummy_bl dummy_br vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_141 vdd vdd vdd vss wl[140] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_142 dummy_bl dummy_br vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_142 vdd vdd vdd vss wl[141] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_143 dummy_bl dummy_br vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_143 vdd vdd vdd vss wl[142] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_144 dummy_bl dummy_br vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_144 vdd vdd vdd vss wl[143] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_145 dummy_bl dummy_br vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_145 vdd vdd vdd vss wl[144] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_146 dummy_bl dummy_br vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_146 vdd vdd vdd vss wl[145] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_147 dummy_bl dummy_br vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_147 vdd vdd vdd vss wl[146] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_148 dummy_bl dummy_br vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_148 vdd vdd vdd vss wl[147] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_149 dummy_bl dummy_br vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_149 vdd vdd vdd vss wl[148] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_150 dummy_bl dummy_br vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_150 vdd vdd vdd vss wl[149] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_151 dummy_bl dummy_br vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_151 vdd vdd vdd vss wl[150] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_152 dummy_bl dummy_br vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_152 vdd vdd vdd vss wl[151] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_153 dummy_bl dummy_br vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_153 vdd vdd vdd vss wl[152] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_154 dummy_bl dummy_br vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_154 vdd vdd vdd vss wl[153] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_155 dummy_bl dummy_br vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_155 vdd vdd vdd vss wl[154] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_156 dummy_bl dummy_br vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_156 vdd vdd vdd vss wl[155] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_157 dummy_bl dummy_br vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_157 vdd vdd vdd vss wl[156] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_158 dummy_bl dummy_br vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_158 vdd vdd vdd vss wl[157] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_159 dummy_bl dummy_br vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_159 vdd vdd vdd vss wl[158] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_160 dummy_bl dummy_br vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_160 vdd vdd vdd vss wl[159] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_161 dummy_bl dummy_br vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_161 vdd vdd vdd vss wl[160] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_162 dummy_bl dummy_br vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_162 vdd vdd vdd vss wl[161] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_163 dummy_bl dummy_br vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_163 vdd vdd vdd vss wl[162] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_164 dummy_bl dummy_br vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_164 vdd vdd vdd vss wl[163] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_165 dummy_bl dummy_br vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_165 vdd vdd vdd vss wl[164] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_166 dummy_bl dummy_br vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_166 vdd vdd vdd vss wl[165] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_167 dummy_bl dummy_br vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_167 vdd vdd vdd vss wl[166] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_168 dummy_bl dummy_br vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_168 vdd vdd vdd vss wl[167] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_169 dummy_bl dummy_br vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_169 vdd vdd vdd vss wl[168] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_170 dummy_bl dummy_br vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_170 vdd vdd vdd vss wl[169] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_171 dummy_bl dummy_br vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_171 vdd vdd vdd vss wl[170] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_172 dummy_bl dummy_br vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_172 vdd vdd vdd vss wl[171] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_173 dummy_bl dummy_br vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_173 vdd vdd vdd vss wl[172] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_174 dummy_bl dummy_br vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_174 vdd vdd vdd vss wl[173] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_175 dummy_bl dummy_br vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_175 vdd vdd vdd vss wl[174] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_176 dummy_bl dummy_br vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_176 vdd vdd vdd vss wl[175] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_177 dummy_bl dummy_br vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_177 vdd vdd vdd vss wl[176] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_178 dummy_bl dummy_br vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_178 vdd vdd vdd vss wl[177] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_179 dummy_bl dummy_br vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_179 vdd vdd vdd vss wl[178] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_180 dummy_bl dummy_br vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_180 vdd vdd vdd vss wl[179] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_181 dummy_bl dummy_br vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_181 vdd vdd vdd vss wl[180] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_182 dummy_bl dummy_br vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_182 vdd vdd vdd vss wl[181] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_183 dummy_bl dummy_br vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_183 vdd vdd vdd vss wl[182] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_184 dummy_bl dummy_br vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_184 vdd vdd vdd vss wl[183] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_185 dummy_bl dummy_br vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_185 vdd vdd vdd vss wl[184] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_186 dummy_bl dummy_br vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_186 vdd vdd vdd vss wl[185] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_187 dummy_bl dummy_br vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_187 vdd vdd vdd vss wl[186] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_188 dummy_bl dummy_br vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_188 vdd vdd vdd vss wl[187] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_189 dummy_bl dummy_br vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_189 vdd vdd vdd vss wl[188] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_190 dummy_bl dummy_br vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_190 vdd vdd vdd vss wl[189] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_191 dummy_bl dummy_br vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_191 vdd vdd vdd vss wl[190] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_192 dummy_bl dummy_br vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_192 vdd vdd vdd vss wl[191] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_193 dummy_bl dummy_br vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_193 vdd vdd vdd vss wl[192] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_194 dummy_bl dummy_br vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_194 vdd vdd vdd vss wl[193] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_195 dummy_bl dummy_br vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_195 vdd vdd vdd vss wl[194] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_196 dummy_bl dummy_br vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_196 vdd vdd vdd vss wl[195] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_197 dummy_bl dummy_br vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_197 vdd vdd vdd vss wl[196] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_198 dummy_bl dummy_br vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_198 vdd vdd vdd vss wl[197] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_199 dummy_bl dummy_br vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_199 vdd vdd vdd vss wl[198] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_200 dummy_bl dummy_br vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_200 vdd vdd vdd vss wl[199] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_201 dummy_bl dummy_br vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_201 vdd vdd vdd vss wl[200] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_202 dummy_bl dummy_br vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_202 vdd vdd vdd vss wl[201] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_203 dummy_bl dummy_br vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_203 vdd vdd vdd vss wl[202] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_204 dummy_bl dummy_br vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_204 vdd vdd vdd vss wl[203] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_205 dummy_bl dummy_br vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_205 vdd vdd vdd vss wl[204] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_206 dummy_bl dummy_br vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_206 vdd vdd vdd vss wl[205] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_207 dummy_bl dummy_br vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_207 vdd vdd vdd vss wl[206] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_208 dummy_bl dummy_br vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_208 vdd vdd vdd vss wl[207] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_209 dummy_bl dummy_br vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_209 vdd vdd vdd vss wl[208] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_210 dummy_bl dummy_br vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_210 vdd vdd vdd vss wl[209] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_211 dummy_bl dummy_br vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_211 vdd vdd vdd vss wl[210] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_212 dummy_bl dummy_br vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_212 vdd vdd vdd vss wl[211] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_213 dummy_bl dummy_br vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_213 vdd vdd vdd vss wl[212] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_214 dummy_bl dummy_br vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_214 vdd vdd vdd vss wl[213] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_215 dummy_bl dummy_br vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_215 vdd vdd vdd vss wl[214] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_216 dummy_bl dummy_br vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_216 vdd vdd vdd vss wl[215] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_217 dummy_bl dummy_br vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_217 vdd vdd vdd vss wl[216] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_218 dummy_bl dummy_br vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_218 vdd vdd vdd vss wl[217] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_219 dummy_bl dummy_br vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_219 vdd vdd vdd vss wl[218] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_220 dummy_bl dummy_br vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_220 vdd vdd vdd vss wl[219] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_221 dummy_bl dummy_br vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_221 vdd vdd vdd vss wl[220] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_222 dummy_bl dummy_br vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_222 vdd vdd vdd vss wl[221] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_223 dummy_bl dummy_br vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_223 vdd vdd vdd vss wl[222] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_224 dummy_bl dummy_br vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_224 vdd vdd vdd vss wl[223] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_225 dummy_bl dummy_br vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_225 vdd vdd vdd vss wl[224] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_226 dummy_bl dummy_br vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_226 vdd vdd vdd vss wl[225] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_227 dummy_bl dummy_br vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_227 vdd vdd vdd vss wl[226] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_228 dummy_bl dummy_br vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_228 vdd vdd vdd vss wl[227] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_229 dummy_bl dummy_br vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_229 vdd vdd vdd vss wl[228] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_230 dummy_bl dummy_br vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_230 vdd vdd vdd vss wl[229] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_231 dummy_bl dummy_br vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_231 vdd vdd vdd vss wl[230] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_232 dummy_bl dummy_br vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_232 vdd vdd vdd vss wl[231] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_233 dummy_bl dummy_br vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_233 vdd vdd vdd vss wl[232] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_234 dummy_bl dummy_br vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_234 vdd vdd vdd vss wl[233] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_235 dummy_bl dummy_br vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_235 vdd vdd vdd vss wl[234] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_236 dummy_bl dummy_br vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_236 vdd vdd vdd vss wl[235] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_237 dummy_bl dummy_br vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_237 vdd vdd vdd vss wl[236] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_238 dummy_bl dummy_br vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_238 vdd vdd vdd vss wl[237] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_239 dummy_bl dummy_br vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_239 vdd vdd vdd vss wl[238] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_240 dummy_bl dummy_br vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_240 vdd vdd vdd vss wl[239] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_241 dummy_bl dummy_br vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_241 vdd vdd vdd vss wl[240] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_242 dummy_bl dummy_br vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_242 vdd vdd vdd vss wl[241] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_243 dummy_bl dummy_br vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_243 vdd vdd vdd vss wl[242] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_244 dummy_bl dummy_br vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_244 vdd vdd vdd vss wl[243] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_245 dummy_bl dummy_br vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_245 vdd vdd vdd vss wl[244] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_246 dummy_bl dummy_br vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_246 vdd vdd vdd vss wl[245] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_247 dummy_bl dummy_br vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_247 vdd vdd vdd vss wl[246] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_248 dummy_bl dummy_br vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_248 vdd vdd vdd vss wl[247] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_249 dummy_bl dummy_br vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_249 vdd vdd vdd vss wl[248] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_250 dummy_bl dummy_br vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_250 vdd vdd vdd vss wl[249] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_251 dummy_bl dummy_br vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_251 vdd vdd vdd vss wl[250] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_252 dummy_bl dummy_br vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_252 vdd vdd vdd vss wl[251] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_253 dummy_bl dummy_br vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_253 vdd vdd vdd vss wl[252] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_254 dummy_bl dummy_br vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_254 vdd vdd vdd vss wl[253] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_255 dummy_bl dummy_br vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_255 vdd vdd vdd vss wl[254] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_256 dummy_bl dummy_br vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_256 vdd vdd vdd vss wl[255] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_257 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_257 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xcolend_top_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xcolend_bot_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xhstrap_0_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_65 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xcolend_bot_65 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xhstrap_0_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_17_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_18_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_19_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_20_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_21_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_22_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_23_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_24_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_25_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_26_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_27_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_28_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_29_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_30_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_31_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_32_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_33_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_34_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_35_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_36_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_37_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_38_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_39_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_40_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_41_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_42_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_43_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_44_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_45_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_46_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_47_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_48_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_49_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_50_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_51_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_52_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_53_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_54_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_55_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_56_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_57_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_58_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_59_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_60_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_61_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_62_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_63_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_64_65 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhoriz_wlstrap_0_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_17_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_18_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_19_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_20_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_21_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_22_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_23_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_24_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_25_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_26_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_27_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_28_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_29_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_30_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_31_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_32_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_33_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_34_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_35_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_36_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_37_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_38_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_39_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_40_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_41_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_42_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_43_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_44_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_45_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_46_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_47_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_48_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_49_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_50_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_51_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_52_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_53_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_54_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_55_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_56_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_57_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_58_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_59_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_60_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_61_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_62_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_63_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_64_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper

.ENDS sp_cell_array

.SUBCKT dff_array_13 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] d[8] d[9] d[10] d[11] d[12] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] q[8] q[9] q[10] q[11] q[12] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7] qn[8] qn[9] qn[10] qn[11] qn[12]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_8 clk d[8] rb vss vss vdd vdd q[8] qn[8] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_9 clk d[9] rb vss vss vdd vdd q[9] qn[9] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_10 clk d[10] rb vss vss vdd vdd q[10] qn[10] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_11 clk d[11] rb vss vss vdd vdd q[11] qn[11] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_12 clk d[12] rb vss vss vdd vdd q[12] qn[12] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_13

.SUBCKT sram_sp_cell_replica BL BR VSS VDD VPB VNB WL

  X0 VDD WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q VDD VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 VDD WL VDD VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q VDD VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q VDD VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell_replica

.SUBCKT sram_sp_cell_replica_wrapper BL BR VSS VDD VPB VNB WL

  X0 BL BR VSS VDD VPB VNB WL sram_sp_cell_replica

.ENDS sram_sp_cell_replica_wrapper

.SUBCKT replica_cell_array vdd vss rbl rbr rwl

  Xcell_0_0 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_0_1 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_1_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_1_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_6_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_6_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_7_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_7_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_8_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_8_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_9_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_9_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_10_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_10_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_11_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_11_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_12_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_12_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_13_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_13_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_14_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_14_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_15_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_15_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_16_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_16_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_17_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_17_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_18_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_18_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_19_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_19_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_20_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_20_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_21_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_21_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_22_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_22_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_23_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_23_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_24_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_24_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_25_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_25_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_26_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_26_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_27_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_27_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_28_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_28_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_29_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_29_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_30_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_30_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_31_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_31_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_32_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_32_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_33_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_33_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_34_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_34_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_35_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_35_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_36_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_36_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_37_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_37_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_38_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_38_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_39_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_39_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_40_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_40_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_41_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_41_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_42_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_42_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_43_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_43_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_44_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_44_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_45_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_45_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcolend_0_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_0_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xrowtapend_0_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_0_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_0_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_0_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_1_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_1_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_1_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_2_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_2_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_2_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_3_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_3_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_3_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_4_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_4_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_4_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_5_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_5_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_5_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_6_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_6_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_6_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_7_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_7_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_7_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_8_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_8_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_8_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_9_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_9_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_9_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_10_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_10_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_10_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_11_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_11_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_11_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper

.ENDS replica_cell_array

.SUBCKT decoder_stage vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] wl_en in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15]

  Xgate_0_0_0 vdd wl_en in[0] y[0] y_b[0] vss and2
  Xgate_0_1_0 vdd wl_en in[1] y[1] y_b[1] vss and2
  Xgate_0_2_0 vdd wl_en in[2] y[2] y_b[2] vss and2
  Xgate_0_3_0 vdd wl_en in[3] y[3] y_b[3] vss and2
  Xgate_0_4_0 vdd wl_en in[4] y[4] y_b[4] vss and2
  Xgate_0_5_0 vdd wl_en in[5] y[5] y_b[5] vss and2
  Xgate_0_6_0 vdd wl_en in[6] y[6] y_b[6] vss and2
  Xgate_0_7_0 vdd wl_en in[7] y[7] y_b[7] vss and2
  Xgate_0_8_0 vdd wl_en in[8] y[8] y_b[8] vss and2
  Xgate_0_9_0 vdd wl_en in[9] y[9] y_b[9] vss and2
  Xgate_0_10_0 vdd wl_en in[10] y[10] y_b[10] vss and2
  Xgate_0_11_0 vdd wl_en in[11] y[11] y_b[11] vss and2
  Xgate_0_12_0 vdd wl_en in[12] y[12] y_b[12] vss and2
  Xgate_0_13_0 vdd wl_en in[13] y[13] y_b[13] vss and2
  Xgate_0_14_0 vdd wl_en in[14] y[14] y_b[14] vss and2
  Xgate_0_15_0 vdd wl_en in[15] y[15] y_b[15] vss and2

.ENDS decoder_stage

.SUBCKT multi_finger_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_7

.SUBCKT decoder_stage_4 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_7
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_7

.ENDS decoder_stage_4

.SUBCKT mos_w1650_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.650


.ENDS mos_w1650_l150_m1_nf1_id1

.SUBCKT precharge vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w1650_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w1650_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w1000_l150_m1_nf1_id1

.ENDS precharge

.SUBCKT sram22_inner vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] addr[10] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7]

  Xaddr_gate vdd vss addr_gated[0] addr_gated[1] addr_gated[2] addr_gated[3] addr_gated[4] addr_gated[5] addr_gated[6] addr_gated[7] addr_b_gated[0] addr_b_gated[1] addr_b_gated[2] addr_b_gated[3] addr_b_gated[4] addr_b_gated[5] addr_b_gated[6] addr_b_gated[7] addr_gate_y_b_noconn[0] addr_gate_y_b_noconn[1] addr_gate_y_b_noconn[2] addr_gate_y_b_noconn[3] addr_gate_y_b_noconn[4] addr_gate_y_b_noconn[5] addr_gate_y_b_noconn[6] addr_gate_y_b_noconn[7] addr_gate_y_b_noconn[8] addr_gate_y_b_noconn[9] addr_gate_y_b_noconn[10] addr_gate_y_b_noconn[11] addr_gate_y_b_noconn[12] addr_gate_y_b_noconn[13] addr_gate_y_b_noconn[14] addr_gate_y_b_noconn[15] wl_en addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in[9] addr_in[10] addr_in_b[3] addr_in_b[4] addr_in_b[5] addr_in_b[6] addr_in_b[7] addr_in_b[8] addr_in_b[9] addr_in_b[10] decoder_stage
  Xdecoder vdd vss wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] wl_b[0] wl_b[1] wl_b[2] wl_b[3] wl_b[4] wl_b[5] wl_b[6] wl_b[7] wl_b[8] wl_b[9] wl_b[10] wl_b[11] wl_b[12] wl_b[13] wl_b[14] wl_b[15] wl_b[16] wl_b[17] wl_b[18] wl_b[19] wl_b[20] wl_b[21] wl_b[22] wl_b[23] wl_b[24] wl_b[25] wl_b[26] wl_b[27] wl_b[28] wl_b[29] wl_b[30] wl_b[31] wl_b[32] wl_b[33] wl_b[34] wl_b[35] wl_b[36] wl_b[37] wl_b[38] wl_b[39] wl_b[40] wl_b[41] wl_b[42] wl_b[43] wl_b[44] wl_b[45] wl_b[46] wl_b[47] wl_b[48] wl_b[49] wl_b[50] wl_b[51] wl_b[52] wl_b[53] wl_b[54] wl_b[55] wl_b[56] wl_b[57] wl_b[58] wl_b[59] wl_b[60] wl_b[61] wl_b[62] wl_b[63] wl_b[64] wl_b[65] wl_b[66] wl_b[67] wl_b[68] wl_b[69] wl_b[70] wl_b[71] wl_b[72] wl_b[73] wl_b[74] wl_b[75] wl_b[76] wl_b[77] wl_b[78] wl_b[79] wl_b[80] wl_b[81] wl_b[82] wl_b[83] wl_b[84] wl_b[85] wl_b[86] wl_b[87] wl_b[88] wl_b[89] wl_b[90] wl_b[91] wl_b[92] wl_b[93] wl_b[94] wl_b[95] wl_b[96] wl_b[97] wl_b[98] wl_b[99] wl_b[100] wl_b[101] wl_b[102] wl_b[103] wl_b[104] wl_b[105] wl_b[106] wl_b[107] wl_b[108] wl_b[109] wl_b[110] wl_b[111] wl_b[112] wl_b[113] wl_b[114] wl_b[115] wl_b[116] wl_b[117] wl_b[118] wl_b[119] wl_b[120] wl_b[121] wl_b[122] wl_b[123] wl_b[124] wl_b[125] wl_b[126] wl_b[127] wl_b[128] wl_b[129] wl_b[130] wl_b[131] wl_b[132] wl_b[133] wl_b[134] wl_b[135] wl_b[136] wl_b[137] wl_b[138] wl_b[139] wl_b[140] wl_b[141] wl_b[142] wl_b[143] wl_b[144] wl_b[145] wl_b[146] wl_b[147] wl_b[148] wl_b[149] wl_b[150] wl_b[151] wl_b[152] wl_b[153] wl_b[154] wl_b[155] wl_b[156] wl_b[157] wl_b[158] wl_b[159] wl_b[160] wl_b[161] wl_b[162] wl_b[163] wl_b[164] wl_b[165] wl_b[166] wl_b[167] wl_b[168] wl_b[169] wl_b[170] wl_b[171] wl_b[172] wl_b[173] wl_b[174] wl_b[175] wl_b[176] wl_b[177] wl_b[178] wl_b[179] wl_b[180] wl_b[181] wl_b[182] wl_b[183] wl_b[184] wl_b[185] wl_b[186] wl_b[187] wl_b[188] wl_b[189] wl_b[190] wl_b[191] wl_b[192] wl_b[193] wl_b[194] wl_b[195] wl_b[196] wl_b[197] wl_b[198] wl_b[199] wl_b[200] wl_b[201] wl_b[202] wl_b[203] wl_b[204] wl_b[205] wl_b[206] wl_b[207] wl_b[208] wl_b[209] wl_b[210] wl_b[211] wl_b[212] wl_b[213] wl_b[214] wl_b[215] wl_b[216] wl_b[217] wl_b[218] wl_b[219] wl_b[220] wl_b[221] wl_b[222] wl_b[223] wl_b[224] wl_b[225] wl_b[226] wl_b[227] wl_b[228] wl_b[229] wl_b[230] wl_b[231] wl_b[232] wl_b[233] wl_b[234] wl_b[235] wl_b[236] wl_b[237] wl_b[238] wl_b[239] wl_b[240] wl_b[241] wl_b[242] wl_b[243] wl_b[244] wl_b[245] wl_b[246] wl_b[247] wl_b[248] wl_b[249] wl_b[250] wl_b[251] wl_b[252] wl_b[253] wl_b[254] wl_b[255] addr_b_gated[0] addr_gated[0] addr_b_gated[1] addr_gated[1] addr_b_gated[2] addr_gated[2] addr_b_gated[3] addr_gated[3] addr_b_gated[4] addr_gated[4] addr_b_gated[5] addr_gated[5] addr_b_gated[6] addr_gated[6] addr_b_gated[7] addr_gated[7] decoder
  Xcolumn_decoder vdd vss col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel[4] col_sel[5] col_sel[6] col_sel[7] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] col_sel_b[4] col_sel_b[5] col_sel_b[6] col_sel_b[7] addr_in_b[0] addr_in[0] addr_in_b[1] addr_in[1] addr_in_b[2] addr_in[2] decoder_1
  Xcontrol_logic clk ce_in we_in rstb rbl sense_en0 pc_b0 rwl wl_en0 write_driver_en0 vdd vss control_logic_replica_v2
  Xpc_b_buffer vdd vss pc_b pc pc_b0 decoder_stage_1
  Xwlen_buffer vdd vss wl_en wl_en_b wl_en0 decoder_stage_2
  Xwrite_driver_en_buffer vdd vss write_driver_en write_driver_en_b write_driver_en0 decoder_stage_3
  Xsense_en_buffer vdd vss sense_en sense_en_b sense_en0 decoder_stage_4
  Xaddr_we_ce_dffs vdd vss clk rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] addr[10] we ce addr_in[0] addr_in[1] addr_in[2] addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in[9] addr_in[10] we_in ce_in addr_in_b[0] addr_in_b[1] addr_in_b[2] addr_in_b[3] addr_in_b[4] addr_in_b[5] addr_in_b[6] addr_in_b[7] addr_in_b[8] addr_in_b[9] addr_in_b[10] we_in_b ce_in_b dff_array_13
  Xbitcell_array vdd vss vdd vdd bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] sp_cell_array
  Xreplica_bitcell_array vdd vss rbl rbr rwl replica_cell_array
  Xcol_circuitry clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] pc_b col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel[4] col_sel[5] col_sel[6] col_sel[7] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] col_sel_b[4] col_sel_b[5] col_sel_b[6] col_sel_b[7] write_driver_en wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] col_peripherals
  Xreplica_precharge_0 vdd rbl rbr pc_b0 precharge
  Xreplica_precharge_1 vdd rbl rbr pc_b0 precharge
  Xreplica_mos vdd vss rbl replica_column_mos

.ENDS sram22_inner

.SUBCKT sram22_2048x8m8w1 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] addr[10] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7]

  X0 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] addr[10] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] sram22_inner

.ENDS sram22_2048x8m8w1

