VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sramgen_sram_4096x8m8w8_replica_v1
  CLASS BLOCK ;
  ORIGIN 93.555 1025.97 ;
  FOREIGN sramgen_sram_4096x8m8w8_replica_v1 -93.555 -1025.97 ;
  SIZE 276.015 BY 1037.685 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -88.2 -1025.57 -87.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -86.6 -1025.57 -86.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -85 -1025.57 -84.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -83.4 -1025.57 -83 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -81.8 -993.54 -81.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -80.2 -1012.62 -79.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -78.6 -1025.57 -78.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -77 -1007.32 -76.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -77 -1025.57 -76.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -75.4 -1008.38 -75 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.8 -1012.62 -73.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.8 -1025.57 -73.4 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.2 -1025.57 -71.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.6 -1006.26 -70.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.6 -1025.57 -70.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -69 -1012.62 -68.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -1012.62 -67 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -1025.57 -67 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.8 -1025.57 -65.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -1006.26 -63.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -1025.57 -63.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.6 -1012.62 -62.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -61 -1025.57 -60.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -1004.14 -59 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -1025.57 -59 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.8 -1012.62 -57.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -1012.62 -55.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -1025.57 -55.8 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.6 -1025.57 -54.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -1003.08 -52.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -1025.57 -52.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.4 -1012.62 -51 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -1012.62 -49.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -1025.57 -49.4 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.2 -1025.57 -47.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -1003.08 -46.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -1025.57 -46.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -1012.62 -44.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -1025.57 -44.6 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.4 -1025.57 -43 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -1002.02 -41.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -1025.57 -41.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.2 -1012.62 -39.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -1012.62 -38.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -1025.57 -38.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -37 -1025.57 -36.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -1000.96 -35 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -1025.57 -35 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.8 -1012.62 -33.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.2 -1025.57 -31.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -999.9 -30.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -1025.57 -30.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -999.9 -28.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -1025.57 -28.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -1012.62 -27 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -1025.57 -27 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.8 -1025.57 -25.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -998.84 -23.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -1025.57 -23.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.6 -1012.62 -22.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -1012.62 -20.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -1025.57 -20.6 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.4 -1025.57 -19 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -997.78 -17.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -1025.57 -17.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.2 -1012.62 -15.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.6 -1025.57 -14.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -996.72 -12.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -1025.57 -12.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -996.72 -11 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -1025.57 -11 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -818.64 -9.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -1012.62 -9.4 -975.94 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -1025.57 -9.4 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.2 -1025.57 -7.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -992.48 -6.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -1025.57 -6.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -5 -1025.57 -4.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.4 -1025.57 -3 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 2.86 -1.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 -1025.57 -1.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 2.86 0.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 -1025.57 0.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 2.86 1.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 -1025.57 1.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 2.86 3.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 -1025.57 3.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 2.86 5 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 -1025.57 5 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 2.86 6.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -1025.57 6.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 2.86 8.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -1025.57 8.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 2.86 9.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -1025.57 9.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 2.86 11.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -862.1 11.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -1025.57 11.4 -973.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 2.86 13 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -828.18 13 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -898.14 13 -889.02 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 2.86 14.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -839.84 14.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -1025.57 14.6 -904.92 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 2.86 16.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 -1025.57 16.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 2.86 17.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 -1025.57 17.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 2.86 19.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -1025.57 19.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 2.86 21 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -1025.57 21 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 2.86 22.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 -904.5 22.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 2.86 24.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 -903.44 24.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 -1025.57 24.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 2.86 25.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 -1025.57 25.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 2.86 27.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 -1025.57 27.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 2.86 29 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -1025.57 29 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 2.86 30.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -1025.57 30.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 2.86 32.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 -1025.57 32.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 2.86 33.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -828.18 33.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -898.14 33.8 -889.02 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 2.86 35.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -828.18 35.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -1025.57 35.4 -913.4 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 2.86 37 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -1025.57 37 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 2.86 38.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -1025.57 38.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 2.86 40.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -1025.57 40.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 2.86 41.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 -1025.57 41.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 2.86 43.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 -1025.57 43.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 2.86 45 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 -1025.57 45 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 2.86 46.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 -1025.57 46.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 2.86 48.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -1025.57 48.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 2.86 49.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -1025.57 49.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 2.86 51.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 -1025.57 51.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 2.86 53 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -828.18 53 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -898.14 53 -889.02 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 2.86 54.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -839.84 54.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -1025.57 54.6 -904.92 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 2.86 56.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 -1025.57 56.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 2.86 57.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 -1025.57 57.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 2.86 59.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -1025.57 59.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 2.86 61 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -1025.57 61 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 2.86 62.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 -904.5 62.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 2.86 64.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -903.44 64.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -1025.57 64.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 2.86 65.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 -1025.57 65.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 2.86 67.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 -1025.57 67.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 2.86 69 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -1025.57 69 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 2.86 70.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -1025.57 70.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 2.86 72.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 -1025.57 72.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 2.86 73.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -828.18 73.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -898.14 73.8 -889.02 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 2.86 75.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -828.18 75.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -1025.57 75.4 -913.4 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 2.86 77 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 -1025.57 77 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 2.86 78.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -1025.57 78.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 2.86 80.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -1025.57 80.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 2.86 81.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 -1025.57 81.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 2.86 83.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 -1025.57 83.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 2.86 85 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 -1025.57 85 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 2.86 86.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 -1025.57 86.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 2.86 88.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -1025.57 88.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 2.86 89.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -1025.57 89.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 2.86 91.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 -1025.57 91.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 2.86 93 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -828.18 93 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -898.14 93 -889.02 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 2.86 94.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -839.84 94.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -1025.57 94.6 -904.92 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 2.86 96.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 -1025.57 96.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 2.86 97.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 -1025.57 97.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 2.86 99.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -1025.57 99.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 2.86 101 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -1025.57 101 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 2.86 102.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 -904.5 102.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 2.86 104.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -903.44 104.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -1025.57 104.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 2.86 105.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 -1025.57 105.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 2.86 107.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 -1025.57 107.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 2.86 109 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -1025.57 109 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 2.86 110.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -1025.57 110.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 2.86 112.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 -1025.57 112.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 2.86 113.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -828.18 113.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -898.14 113.8 -889.02 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 2.86 115.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -828.18 115.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -1025.57 115.4 -913.4 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 2.86 117 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 -1025.57 117 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 2.86 118.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -1025.57 118.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 2.86 120.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -1025.57 120.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 2.86 121.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 -1025.57 121.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 2.86 123.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 -1025.57 123.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 2.86 125 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 -1025.57 125 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 2.86 126.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 -1025.57 126.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 2.86 128.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -1025.57 128.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 2.86 129.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -1025.57 129.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 2.86 131.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 -1025.57 131.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 2.86 133 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -828.18 133 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -898.14 133 -889.02 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 2.86 134.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -839.84 134.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -1025.57 134.6 -904.92 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 2.86 136.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 -1025.57 136.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 2.86 137.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 -1025.57 137.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 2.86 139.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -1025.57 139.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 2.86 141 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -1025.57 141 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 2.86 142.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 -904.5 142.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 2.86 144.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -903.44 144.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -1025.57 144.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 2.86 145.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 -1025.57 145.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 2.86 147.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 -1025.57 147.4 -818 ;
        RECT 146.95 -901.37 147.4 -901.04 ;
        RECT 146.95 -915.51 147.4 -915.18 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 2.86 149 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -1025.57 149 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 2.86 150.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -1025.57 150.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 2.86 152.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 -1025.57 152.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 2.86 153.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -828.18 153.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -898.14 153.8 -889.02 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 2.86 155.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -828.18 155.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -1025.57 155.4 -913.4 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 2.86 157 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 -1025.57 157 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 2.86 158.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -1025.57 158.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 2.86 160.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -1025.57 160.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 2.86 161.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 -1025.57 161.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 2.86 163.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 -1025.57 163.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 2.86 165 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 -1025.57 165 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 2.86 166.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 -1025.57 166.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 2.86 168.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -1025.57 168.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 2.86 169.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -1025.57 169.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 -1025.57 171.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -1025.57 173 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -1025.57 174.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 -1025.57 176.2 11.315 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -87.4 -1024.03 -87 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -85.8 -1024.03 -85.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -84.2 -1024.03 -83.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -82.6 -1024.03 -82.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -81 -993.54 -80.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.4 -1012.62 -79 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.4 -1024.03 -79 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -77.8 -1024.03 -77.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -76.2 -1007.32 -75.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -76.2 -1024.03 -75.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.6 -1012.62 -74.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -73 -1024.03 -72.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.4 -1006.26 -71 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.4 -1024.03 -71 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.8 -1007.32 -69.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.8 -1024.03 -69.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -1012.62 -67.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -1024.03 -67.8 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.6 -1024.03 -66.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -1005.2 -64.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -1024.03 -64.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.4 -1012.62 -63 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -1012.62 -61.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -1024.03 -61.4 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.2 -1024.03 -59.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -1004.14 -58.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -1024.03 -58.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -57 -1012.62 -56.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.4 -1024.03 -55 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -1003.08 -53.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -1024.03 -53.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.2 -1004.14 -51.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -1012.62 -50.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -1024.03 -50.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -49 -1024.03 -48.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -1002.02 -47 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -1024.03 -47 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.8 -1012.62 -45.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -1012.62 -43.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -1024.03 -43.8 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.6 -1024.03 -42.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -1002.02 -40.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -1024.03 -40.6 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.4 -1012.62 -39 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.8 -1024.03 -37.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -1000.96 -35.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -1024.03 -35.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.6 -1000.96 -34.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -1012.62 -32.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -1024.03 -32.6 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.4 -1024.03 -31 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -999.9 -29.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -1024.03 -29.4 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.2 -1012.62 -27.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -1012.62 -26.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -1024.03 -26.2 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -25 -1024.03 -24.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -998.84 -23 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -1024.03 -23 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.8 -1012.62 -21.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.2 -1024.03 -19.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -997.78 -18.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -1024.03 -18.2 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -17 -997.78 -16.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -1012.62 -15 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -1024.03 -15 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.8 -1024.03 -13.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -996.72 -11.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -1024.03 -11.8 -1015.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -818.64 -10.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -1012.62 -10.2 -975.94 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -1012.62 -8.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -1024.03 -8.6 -1018.34 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.4 -1024.03 -7 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -992.48 -5.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -1024.03 -5.4 -1015.16 ;
        RECT -5.825 -1017.025 -5.4 -1016.695 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.2 -1024.03 -3.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.6 -1024.03 -2.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 2.86 -0.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 -1024.03 -0.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 2.86 1 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 -1024.03 1 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 2.86 2.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 -1024.03 2.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 2.86 4.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 -1024.03 4.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 2.86 5.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -1024.03 5.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 2.86 7.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 -1024.03 7.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 2.86 9 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -1024.03 9 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 2.86 10.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -1024.03 10.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 2.86 12.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 -1024.03 12.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 2.86 13.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -828.18 13.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -898.14 13.8 -889.02 ;
        RECT 13.435 -898.14 13.765 -888.98 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 2.86 15.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -828.18 15.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -1024.03 15.4 -904.92 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 2.86 17 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 -1024.03 17 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 2.86 18.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -1024.03 18.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 2.86 20.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -1024.03 20.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 2.86 21.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -904.5 21.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 2.86 23.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 -903.44 23.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 2.86 25 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 -1024.03 25 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 2.86 26.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 -1024.03 26.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 2.86 28.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -1024.03 28.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 2.86 29.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -1024.03 29.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 2.86 31.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 -1024.03 31.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 2.86 33 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -828.18 33 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -898.14 33 -889.02 ;
        RECT 32.635 -898.14 32.965 -888.98 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 2.86 34.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -839.84 34.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -1024.03 34.6 -913.4 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 2.86 36.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -1024.03 36.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 2.86 37.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 -1024.03 37.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 2.86 39.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -1024.03 39.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 2.86 41 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -1024.03 41 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 2.86 42.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 -1024.03 42.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 2.86 44.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 -1024.03 44.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 2.86 45.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 -1024.03 45.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 2.86 47.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 -1024.03 47.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 2.86 49 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -1024.03 49 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 2.86 50.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -1024.03 50.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 2.86 52.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 -1024.03 52.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 2.86 53.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -828.18 53.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -898.14 53.8 -889.02 ;
        RECT 53.435 -898.14 53.765 -888.98 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 2.86 55.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -828.18 55.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -1024.03 55.4 -904.92 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 2.86 57 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 -1024.03 57 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 2.86 58.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -1024.03 58.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 2.86 60.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -1024.03 60.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 2.86 61.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 -904.5 61.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 2.86 63.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 -903.44 63.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 2.86 65 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 -1024.03 65 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 2.86 66.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 -1024.03 66.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 2.86 68.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -1024.03 68.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 2.86 69.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -1024.03 69.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 2.86 71.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 -1024.03 71.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 2.86 73 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -828.18 73 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -898.14 73 -889.02 ;
        RECT 72.635 -898.14 72.965 -888.98 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 2.86 74.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -839.84 74.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -1024.03 74.6 -913.4 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 2.86 76.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 -1024.03 76.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 2.86 77.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 -1024.03 77.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 2.86 79.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -1024.03 79.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 2.86 81 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -1024.03 81 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 2.86 82.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 -1024.03 82.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 2.86 84.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 -1024.03 84.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 2.86 85.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 -1024.03 85.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 2.86 87.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 -1024.03 87.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 2.86 89 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -1024.03 89 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 2.86 90.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -1024.03 90.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 2.86 92.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 -1024.03 92.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 2.86 93.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -828.18 93.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -898.14 93.8 -889.02 ;
        RECT 93.435 -898.14 93.765 -888.98 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 2.86 95.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -828.18 95.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -1024.03 95.4 -904.92 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 2.86 97 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 -1024.03 97 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 2.86 98.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -1024.03 98.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 2.86 100.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -1024.03 100.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 2.86 101.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -904.5 101.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 2.86 103.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 -903.44 103.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 2.86 105 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 -1024.03 105 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 2.86 106.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 -1024.03 106.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 2.86 108.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -1024.03 108.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 2.86 109.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -1024.03 109.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 2.86 111.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 -1024.03 111.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 2.86 113 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -828.18 113 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -898.14 113 -889.02 ;
        RECT 112.635 -898.14 112.965 -888.98 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 2.86 114.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -839.84 114.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -1024.03 114.6 -913.4 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 2.86 116.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 -1024.03 116.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 2.86 117.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 -1024.03 117.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 2.86 119.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -1024.03 119.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 2.86 121 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -1024.03 121 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 2.86 122.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 -1024.03 122.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 2.86 124.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 -1024.03 124.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 2.86 125.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 -1024.03 125.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 2.86 127.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 -1024.03 127.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 2.86 129 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -1024.03 129 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 2.86 130.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -1024.03 130.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 2.86 132.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 -1024.03 132.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 2.86 133.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -828.18 133.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -898.14 133.8 -889.02 ;
        RECT 133.435 -898.14 133.765 -888.98 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 2.86 135.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -828.18 135.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -1024.03 135.4 -904.92 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 2.86 137 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 -1024.03 137 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 2.86 138.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -1024.03 138.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 2.86 140.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -1024.03 140.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 2.86 141.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 -904.5 141.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 2.86 143.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 -903.44 143.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 2.86 145 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 -1024.03 145 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 2.86 146.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 -1024.03 146.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 2.86 148.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -1024.03 148.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 2.86 149.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -1024.03 149.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 2.86 151.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 -1024.03 151.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 2.86 153 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -828.18 153 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -898.14 153 -889.02 ;
        RECT 152.635 -898.14 152.965 -888.98 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 2.86 154.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -839.84 154.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -1024.03 154.6 -913.4 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 2.86 156.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 -1024.03 156.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 2.86 157.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 -1024.03 157.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 2.86 159.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -1024.03 159.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 2.86 161 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -1024.03 161 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 2.86 162.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 -1024.03 162.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 2.86 164.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 -1024.03 164.2 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 2.86 165.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 -1024.03 165.8 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 2.86 167.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 -1024.03 167.4 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 2.86 169 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -1024.03 169 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 2.86 170.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -1024.03 170.6 -818 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 -1024.03 172.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -1024.03 173.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -1024.03 175.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 -1024.03 177 9.775 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -16.46 -1025.97 -16.16 -1025.67 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -74.86 -1025.97 -74.56 -1025.67 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -80.7 -1025.97 -80.4 -1025.67 ;
    END
  END addr[11]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -22.3 -1025.97 -22 -1025.67 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.14 -1025.97 -27.84 -1025.67 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -33.98 -1025.97 -33.68 -1025.67 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -39.82 -1025.97 -39.52 -1025.67 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -45.66 -1025.97 -45.36 -1025.67 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -51.5 -1025.97 -51.2 -1025.67 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -57.34 -1025.97 -57.04 -1025.67 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -63.18 -1025.97 -62.88 -1025.67 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -69.02 -1025.97 -68.72 -1025.67 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -81.72 -1025.97 -81.3 -1025.55 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.015 -1025.97 22.315 -1025.67 ;
    END
  END din[0]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.63 -1025.97 22.93 -1025.67 ;
    END
  END din[1]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.015 -1025.97 62.315 -1025.67 ;
    END
  END din[2]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.63 -1025.97 62.93 -1025.67 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.015 -1025.97 102.315 -1025.67 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.63 -1025.97 102.93 -1025.67 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.015 -1025.97 142.315 -1025.67 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.63 -1025.97 142.93 -1025.67 ;
    END
  END din[7]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 13.285 -1025.97 13.585 -1025.67 ;
    END
  END dout[0]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 33.285 -1025.97 33.585 -1025.67 ;
    END
  END dout[1]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.285 -1025.97 53.585 -1025.67 ;
    END
  END dout[2]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 73.285 -1025.97 73.585 -1025.67 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 93.285 -1025.97 93.585 -1025.67 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.285 -1025.97 113.585 -1025.67 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.285 -1025.97 133.585 -1025.67 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 153.285 -1025.97 153.585 -1025.67 ;
    END
  END dout[7]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -10.62 -1025.97 -10.32 -1025.67 ;
    END
  END we
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -93.555 -1025.97 182.46 11.715 ;
    LAYER met2 SPACING 0.14 ;
      RECT -93.555 -1025.97 182.46 11.715 ;
    LAYER met3 SPACING 0.3 ;
      RECT 155.115 -873.025 155.445 -872.695 ;
      RECT 155.13 -888.455 155.43 -872.695 ;
      RECT 155.115 -888.455 155.445 -888.125 ;
      RECT 155.13 -869.24 155.43 -829.2 ;
      RECT 155.115 -831.175 155.445 -830.845 ;
      RECT 155.115 -868.83 155.445 -868.5 ;
      RECT 154.515 -912.345 154.815 -840.535 ;
      RECT 154.5 -840.91 154.83 -840.58 ;
      RECT 154.5 -856.61 154.83 -856.28 ;
      RECT 154.5 -912.345 154.83 -912.015 ;
      RECT 153.9 -851.95 154.2 -841.165 ;
      RECT 153.885 -841.54 154.215 -841.21 ;
      RECT 153.885 -851.95 154.215 -851.62 ;
      RECT 153.27 -899.43 153.6 -899.1 ;
      RECT 153.285 -1025.18 153.585 -899.1 ;
      RECT 153.27 -873.485 153.6 -873.155 ;
      RECT 153.285 -888.455 153.585 -873.155 ;
      RECT 153.27 -888.455 153.6 -888.125 ;
      RECT 153.285 -869.26 153.585 -829.2 ;
      RECT 153.27 -829.575 153.6 -829.245 ;
      RECT 153.27 -869.26 153.6 -868.93 ;
      RECT 143.245 -904.82 143.575 -904.49 ;
      RECT 143.26 -1017.91 143.56 -904.49 ;
      RECT 143.245 -912.06 143.575 -911.73 ;
      RECT 143.245 -1017.865 143.575 -1017.535 ;
      RECT 142.615 -911.26 142.945 -910.93 ;
      RECT 142.63 -1025.18 142.93 -910.93 ;
      RECT 142 -905.62 142.33 -905.29 ;
      RECT 142.015 -1025.18 142.315 -905.29 ;
      RECT 135.115 -873.025 135.445 -872.695 ;
      RECT 135.13 -888.455 135.43 -872.695 ;
      RECT 135.115 -888.455 135.445 -888.125 ;
      RECT 135.13 -869.24 135.43 -829.2 ;
      RECT 135.115 -831.175 135.445 -830.845 ;
      RECT 135.115 -868.83 135.445 -868.5 ;
      RECT 134.515 -904.335 134.815 -840.535 ;
      RECT 134.5 -840.91 134.83 -840.58 ;
      RECT 134.5 -856.61 134.83 -856.28 ;
      RECT 134.5 -904.335 134.83 -904.005 ;
      RECT 133.9 -851.95 134.2 -841.165 ;
      RECT 133.885 -841.54 134.215 -841.21 ;
      RECT 133.885 -851.95 134.215 -851.62 ;
      RECT 133.27 -899.43 133.6 -899.1 ;
      RECT 133.285 -1025.18 133.585 -899.1 ;
      RECT 133.27 -873.485 133.6 -873.155 ;
      RECT 133.285 -888.455 133.585 -873.155 ;
      RECT 133.27 -888.455 133.6 -888.125 ;
      RECT 133.285 -869.26 133.585 -829.2 ;
      RECT 133.27 -829.575 133.6 -829.245 ;
      RECT 133.27 -869.26 133.6 -868.93 ;
      RECT 115.115 -873.025 115.445 -872.695 ;
      RECT 115.13 -888.455 115.43 -872.695 ;
      RECT 115.115 -888.455 115.445 -888.125 ;
      RECT 115.13 -869.24 115.43 -829.2 ;
      RECT 115.115 -831.175 115.445 -830.845 ;
      RECT 115.115 -868.83 115.445 -868.5 ;
      RECT 114.515 -912.345 114.815 -840.535 ;
      RECT 114.5 -840.91 114.83 -840.58 ;
      RECT 114.5 -856.61 114.83 -856.28 ;
      RECT 114.5 -912.345 114.83 -912.015 ;
      RECT 113.9 -851.95 114.2 -841.165 ;
      RECT 113.885 -841.54 114.215 -841.21 ;
      RECT 113.885 -851.95 114.215 -851.62 ;
      RECT 113.27 -899.43 113.6 -899.1 ;
      RECT 113.285 -1025.18 113.585 -899.1 ;
      RECT 113.27 -873.485 113.6 -873.155 ;
      RECT 113.285 -888.455 113.585 -873.155 ;
      RECT 113.27 -888.455 113.6 -888.125 ;
      RECT 113.285 -869.26 113.585 -829.2 ;
      RECT 113.27 -829.575 113.6 -829.245 ;
      RECT 113.27 -869.26 113.6 -868.93 ;
      RECT 103.245 -904.82 103.575 -904.49 ;
      RECT 103.26 -1017.91 103.56 -904.49 ;
      RECT 103.245 -912.06 103.575 -911.73 ;
      RECT 103.245 -1017.865 103.575 -1017.535 ;
      RECT 102.615 -911.26 102.945 -910.93 ;
      RECT 102.63 -1025.18 102.93 -910.93 ;
      RECT 102 -905.62 102.33 -905.29 ;
      RECT 102.015 -1025.18 102.315 -905.29 ;
      RECT 95.115 -873.025 95.445 -872.695 ;
      RECT 95.13 -888.455 95.43 -872.695 ;
      RECT 95.115 -888.455 95.445 -888.125 ;
      RECT 95.13 -869.24 95.43 -829.2 ;
      RECT 95.115 -831.175 95.445 -830.845 ;
      RECT 95.115 -868.83 95.445 -868.5 ;
      RECT 94.515 -904.335 94.815 -840.535 ;
      RECT 94.5 -840.91 94.83 -840.58 ;
      RECT 94.5 -856.61 94.83 -856.28 ;
      RECT 94.5 -904.335 94.83 -904.005 ;
      RECT 93.9 -851.95 94.2 -841.165 ;
      RECT 93.885 -841.54 94.215 -841.21 ;
      RECT 93.885 -851.95 94.215 -851.62 ;
      RECT 93.27 -899.43 93.6 -899.1 ;
      RECT 93.285 -1025.18 93.585 -899.1 ;
      RECT 93.27 -873.485 93.6 -873.155 ;
      RECT 93.285 -888.455 93.585 -873.155 ;
      RECT 93.27 -888.455 93.6 -888.125 ;
      RECT 93.285 -869.26 93.585 -829.2 ;
      RECT 93.27 -829.575 93.6 -829.245 ;
      RECT 93.27 -869.26 93.6 -868.93 ;
      RECT 75.115 -873.025 75.445 -872.695 ;
      RECT 75.13 -888.455 75.43 -872.695 ;
      RECT 75.115 -888.455 75.445 -888.125 ;
      RECT 75.13 -869.24 75.43 -829.2 ;
      RECT 75.115 -831.175 75.445 -830.845 ;
      RECT 75.115 -868.83 75.445 -868.5 ;
      RECT 74.515 -912.345 74.815 -840.535 ;
      RECT 74.5 -840.91 74.83 -840.58 ;
      RECT 74.5 -856.61 74.83 -856.28 ;
      RECT 74.5 -912.345 74.83 -912.015 ;
      RECT 73.9 -851.95 74.2 -841.165 ;
      RECT 73.885 -841.54 74.215 -841.21 ;
      RECT 73.885 -851.95 74.215 -851.62 ;
      RECT 73.27 -899.43 73.6 -899.1 ;
      RECT 73.285 -1025.18 73.585 -899.1 ;
      RECT 73.27 -873.485 73.6 -873.155 ;
      RECT 73.285 -888.455 73.585 -873.155 ;
      RECT 73.27 -888.455 73.6 -888.125 ;
      RECT 73.285 -869.26 73.585 -829.2 ;
      RECT 73.27 -829.575 73.6 -829.245 ;
      RECT 73.27 -869.26 73.6 -868.93 ;
      RECT 63.245 -904.82 63.575 -904.49 ;
      RECT 63.26 -1017.91 63.56 -904.49 ;
      RECT 63.245 -912.06 63.575 -911.73 ;
      RECT 63.245 -1017.865 63.575 -1017.535 ;
      RECT 62.615 -911.26 62.945 -910.93 ;
      RECT 62.63 -1025.18 62.93 -910.93 ;
      RECT 62 -905.62 62.33 -905.29 ;
      RECT 62.015 -1025.18 62.315 -905.29 ;
      RECT 55.115 -873.025 55.445 -872.695 ;
      RECT 55.13 -888.455 55.43 -872.695 ;
      RECT 55.115 -888.455 55.445 -888.125 ;
      RECT 55.13 -869.24 55.43 -829.2 ;
      RECT 55.115 -831.175 55.445 -830.845 ;
      RECT 55.115 -868.83 55.445 -868.5 ;
      RECT 54.515 -904.335 54.815 -840.535 ;
      RECT 54.5 -840.91 54.83 -840.58 ;
      RECT 54.5 -856.61 54.83 -856.28 ;
      RECT 54.5 -904.335 54.83 -904.005 ;
      RECT 53.9 -851.95 54.2 -841.165 ;
      RECT 53.885 -841.54 54.215 -841.21 ;
      RECT 53.885 -851.95 54.215 -851.62 ;
      RECT 53.27 -899.43 53.6 -899.1 ;
      RECT 53.285 -1025.18 53.585 -899.1 ;
      RECT 53.27 -873.485 53.6 -873.155 ;
      RECT 53.285 -888.455 53.585 -873.155 ;
      RECT 53.27 -888.455 53.6 -888.125 ;
      RECT 53.285 -869.26 53.585 -829.2 ;
      RECT 53.27 -829.575 53.6 -829.245 ;
      RECT 53.27 -869.26 53.6 -868.93 ;
      RECT 35.115 -873.025 35.445 -872.695 ;
      RECT 35.13 -888.455 35.43 -872.695 ;
      RECT 35.115 -888.455 35.445 -888.125 ;
      RECT 35.13 -869.24 35.43 -829.2 ;
      RECT 35.115 -831.175 35.445 -830.845 ;
      RECT 35.115 -868.83 35.445 -868.5 ;
      RECT 34.515 -912.345 34.815 -840.535 ;
      RECT 34.5 -840.91 34.83 -840.58 ;
      RECT 34.5 -856.61 34.83 -856.28 ;
      RECT 34.5 -912.345 34.83 -912.015 ;
      RECT 33.9 -851.95 34.2 -841.165 ;
      RECT 33.885 -841.54 34.215 -841.21 ;
      RECT 33.885 -851.95 34.215 -851.62 ;
      RECT 33.27 -899.43 33.6 -899.1 ;
      RECT 33.285 -1025.18 33.585 -899.1 ;
      RECT 33.27 -873.485 33.6 -873.155 ;
      RECT 33.285 -888.455 33.585 -873.155 ;
      RECT 33.27 -888.455 33.6 -888.125 ;
      RECT 33.285 -869.26 33.585 -829.2 ;
      RECT 33.27 -829.575 33.6 -829.245 ;
      RECT 33.27 -869.26 33.6 -868.93 ;
      RECT 23.245 -904.82 23.575 -904.49 ;
      RECT 23.26 -1017.91 23.56 -904.49 ;
      RECT 23.245 -912.06 23.575 -911.73 ;
      RECT 23.245 -1017.865 23.575 -1017.535 ;
      RECT 22.615 -911.26 22.945 -910.93 ;
      RECT 22.63 -1025.18 22.93 -910.93 ;
      RECT 22 -905.62 22.33 -905.29 ;
      RECT 22.015 -1025.18 22.315 -905.29 ;
      RECT 15.115 -873.025 15.445 -872.695 ;
      RECT 15.13 -888.455 15.43 -872.695 ;
      RECT 15.115 -888.455 15.445 -888.125 ;
      RECT 15.13 -869.24 15.43 -829.2 ;
      RECT 15.115 -831.175 15.445 -830.845 ;
      RECT 15.115 -868.83 15.445 -868.5 ;
      RECT 14.515 -904.335 14.815 -840.535 ;
      RECT 14.5 -840.91 14.83 -840.58 ;
      RECT 14.5 -856.61 14.83 -856.28 ;
      RECT 14.5 -904.335 14.83 -904.005 ;
      RECT 13.9 -851.95 14.2 -841.165 ;
      RECT 13.885 -841.54 14.215 -841.21 ;
      RECT 13.885 -851.95 14.215 -851.62 ;
      RECT 13.27 -899.43 13.6 -899.1 ;
      RECT 13.285 -1025.18 13.585 -899.1 ;
      RECT 13.27 -873.485 13.6 -873.155 ;
      RECT 13.285 -888.455 13.585 -873.155 ;
      RECT 13.27 -888.455 13.6 -888.125 ;
      RECT 13.285 -869.26 13.585 -829.2 ;
      RECT 13.27 -829.575 13.6 -829.245 ;
      RECT 13.27 -869.26 13.6 -868.93 ;
      RECT 11.005 -863.245 11.335 -862.915 ;
      RECT 11.02 -972.98 11.32 -862.915 ;
      RECT 11.005 -972.98 11.335 -972.65 ;
      RECT -5.91 -993.415 -5.58 -993.085 ;
      RECT -5.895 -1013.85 -5.595 -993.085 ;
      RECT -5.91 -1013.85 -5.58 -1013.52 ;
      RECT -9.505 -1013.405 -9.175 -1013.075 ;
      RECT -9.49 -1017.91 -9.19 -1013.075 ;
      RECT -9.505 -1017.865 -9.175 -1017.535 ;
      RECT -10.34 -819.74 -10.01 -819.41 ;
      RECT -10.325 -974.77 -10.025 -819.41 ;
      RECT -10.34 -974.77 -10.01 -974.44 ;
      RECT -10.635 -1014.205 -10.305 -1013.875 ;
      RECT -10.62 -1025.18 -10.32 -1013.875 ;
      RECT -11.75 -998.18 -11.42 -997.85 ;
      RECT -11.735 -1013.85 -11.435 -997.85 ;
      RECT -11.75 -1013.85 -11.42 -1013.52 ;
      RECT -12.385 -997.68 -12.055 -997.35 ;
      RECT -12.37 -1014.605 -12.07 -997.35 ;
      RECT -12.385 -1014.605 -12.055 -1014.275 ;
      RECT -15.345 -1013.405 -15.015 -1013.075 ;
      RECT -15.33 -1017.91 -15.03 -1013.075 ;
      RECT -15.345 -1017.865 -15.015 -1017.535 ;
      RECT -16.475 -1014.205 -16.145 -1013.875 ;
      RECT -16.46 -1025.18 -16.16 -1013.875 ;
      RECT -17.59 -999.18 -17.26 -998.85 ;
      RECT -17.575 -1013.85 -17.275 -998.85 ;
      RECT -17.59 -1013.85 -17.26 -1013.52 ;
      RECT -18.225 -998.68 -17.895 -998.35 ;
      RECT -18.21 -1014.605 -17.91 -998.35 ;
      RECT -18.225 -1014.605 -17.895 -1014.275 ;
      RECT -21.185 -1013.405 -20.855 -1013.075 ;
      RECT -21.17 -1017.91 -20.87 -1013.075 ;
      RECT -21.185 -1017.865 -20.855 -1017.535 ;
      RECT -22.315 -1014.205 -21.985 -1013.875 ;
      RECT -22.3 -1025.18 -22 -1013.875 ;
      RECT -23.43 -1000.18 -23.1 -999.85 ;
      RECT -23.415 -1013.85 -23.115 -999.85 ;
      RECT -23.43 -1013.85 -23.1 -1013.52 ;
      RECT -24.065 -999.68 -23.735 -999.35 ;
      RECT -24.05 -1014.605 -23.75 -999.35 ;
      RECT -24.065 -1014.605 -23.735 -1014.275 ;
      RECT -27.025 -1013.405 -26.695 -1013.075 ;
      RECT -27.01 -1017.91 -26.71 -1013.075 ;
      RECT -27.025 -1017.865 -26.695 -1017.535 ;
      RECT -28.155 -1014.205 -27.825 -1013.875 ;
      RECT -28.14 -1025.18 -27.84 -1013.875 ;
      RECT -29.27 -1001.18 -28.94 -1000.85 ;
      RECT -29.255 -1013.85 -28.955 -1000.85 ;
      RECT -29.27 -1013.85 -28.94 -1013.52 ;
      RECT -29.905 -1000.68 -29.575 -1000.35 ;
      RECT -29.89 -1014.605 -29.59 -1000.35 ;
      RECT -29.905 -1014.605 -29.575 -1014.275 ;
      RECT -32.865 -1013.405 -32.535 -1013.075 ;
      RECT -32.85 -1017.91 -32.55 -1013.075 ;
      RECT -32.865 -1017.865 -32.535 -1017.535 ;
      RECT -33.995 -1014.205 -33.665 -1013.875 ;
      RECT -33.98 -1025.18 -33.68 -1013.875 ;
      RECT -35.11 -1002.18 -34.78 -1001.85 ;
      RECT -35.095 -1013.85 -34.795 -1001.85 ;
      RECT -35.11 -1013.85 -34.78 -1013.52 ;
      RECT -35.745 -1001.68 -35.415 -1001.35 ;
      RECT -35.73 -1014.605 -35.43 -1001.35 ;
      RECT -35.745 -1014.605 -35.415 -1014.275 ;
      RECT -38.705 -1013.405 -38.375 -1013.075 ;
      RECT -38.69 -1017.91 -38.39 -1013.075 ;
      RECT -38.705 -1017.865 -38.375 -1017.535 ;
      RECT -39.835 -1014.205 -39.505 -1013.875 ;
      RECT -39.82 -1025.18 -39.52 -1013.875 ;
      RECT -40.95 -1003.18 -40.62 -1002.85 ;
      RECT -40.935 -1013.85 -40.635 -1002.85 ;
      RECT -40.95 -1013.85 -40.62 -1013.52 ;
      RECT -41.585 -1002.68 -41.255 -1002.35 ;
      RECT -41.57 -1014.605 -41.27 -1002.35 ;
      RECT -41.585 -1014.605 -41.255 -1014.275 ;
      RECT -44.545 -1013.405 -44.215 -1013.075 ;
      RECT -44.53 -1017.91 -44.23 -1013.075 ;
      RECT -44.545 -1017.865 -44.215 -1017.535 ;
      RECT -45.675 -1014.205 -45.345 -1013.875 ;
      RECT -45.66 -1025.18 -45.36 -1013.875 ;
      RECT -46.79 -1004.18 -46.46 -1003.85 ;
      RECT -46.775 -1013.85 -46.475 -1003.85 ;
      RECT -46.79 -1013.85 -46.46 -1013.52 ;
      RECT -47.425 -1003.68 -47.095 -1003.35 ;
      RECT -47.41 -1014.605 -47.11 -1003.35 ;
      RECT -47.425 -1014.605 -47.095 -1014.275 ;
      RECT -50.385 -1013.405 -50.055 -1013.075 ;
      RECT -50.37 -1017.91 -50.07 -1013.075 ;
      RECT -50.385 -1017.865 -50.055 -1017.535 ;
      RECT -51.515 -1014.205 -51.185 -1013.875 ;
      RECT -51.5 -1025.18 -51.2 -1013.875 ;
      RECT -52.63 -1005.18 -52.3 -1004.85 ;
      RECT -52.615 -1013.85 -52.315 -1004.85 ;
      RECT -52.63 -1013.85 -52.3 -1013.52 ;
      RECT -53.265 -1004.68 -52.935 -1004.35 ;
      RECT -53.25 -1014.605 -52.95 -1004.35 ;
      RECT -53.265 -1014.605 -52.935 -1014.275 ;
      RECT -56.225 -1013.405 -55.895 -1013.075 ;
      RECT -56.21 -1017.91 -55.91 -1013.075 ;
      RECT -56.225 -1017.865 -55.895 -1017.535 ;
      RECT -57.355 -1014.205 -57.025 -1013.875 ;
      RECT -57.34 -1025.18 -57.04 -1013.875 ;
      RECT -58.47 -1006.18 -58.14 -1005.85 ;
      RECT -58.455 -1013.85 -58.155 -1005.85 ;
      RECT -58.47 -1013.85 -58.14 -1013.52 ;
      RECT -59.105 -1005.68 -58.775 -1005.35 ;
      RECT -59.09 -1014.605 -58.79 -1005.35 ;
      RECT -59.105 -1014.605 -58.775 -1014.275 ;
      RECT -62.065 -1013.405 -61.735 -1013.075 ;
      RECT -62.05 -1017.91 -61.75 -1013.075 ;
      RECT -62.065 -1017.865 -61.735 -1017.535 ;
      RECT -63.195 -1014.205 -62.865 -1013.875 ;
      RECT -63.18 -1025.18 -62.88 -1013.875 ;
      RECT -64.31 -1007.18 -63.98 -1006.85 ;
      RECT -64.295 -1013.85 -63.995 -1006.85 ;
      RECT -64.31 -1013.85 -63.98 -1013.52 ;
      RECT -64.945 -1006.68 -64.615 -1006.35 ;
      RECT -64.93 -1014.605 -64.63 -1006.35 ;
      RECT -64.945 -1014.605 -64.615 -1014.275 ;
      RECT -67.905 -1013.405 -67.575 -1013.075 ;
      RECT -67.89 -1017.91 -67.59 -1013.075 ;
      RECT -67.905 -1017.865 -67.575 -1017.535 ;
      RECT -69.035 -1014.205 -68.705 -1013.875 ;
      RECT -69.02 -1025.18 -68.72 -1013.875 ;
      RECT -70.15 -1008.18 -69.82 -1007.85 ;
      RECT -70.135 -1013.85 -69.835 -1007.85 ;
      RECT -70.15 -1013.85 -69.82 -1013.52 ;
      RECT -70.785 -1007.68 -70.455 -1007.35 ;
      RECT -70.77 -1014.605 -70.47 -1007.35 ;
      RECT -70.785 -1014.605 -70.455 -1014.275 ;
      RECT -73.745 -1013.405 -73.415 -1013.075 ;
      RECT -73.73 -1017.91 -73.43 -1013.075 ;
      RECT -73.745 -1017.865 -73.415 -1017.535 ;
      RECT -74.875 -1014.205 -74.545 -1013.875 ;
      RECT -74.86 -1025.18 -74.56 -1013.875 ;
      RECT -75.99 -1009.18 -75.66 -1008.85 ;
      RECT -75.975 -1013.85 -75.675 -1008.85 ;
      RECT -75.99 -1013.85 -75.66 -1013.52 ;
      RECT -76.625 -1008.68 -76.295 -1008.35 ;
      RECT -76.61 -1014.605 -76.31 -1008.35 ;
      RECT -76.625 -1014.605 -76.295 -1014.275 ;
      RECT -79.585 -1013.405 -79.255 -1013.075 ;
      RECT -79.57 -1017.91 -79.27 -1013.075 ;
      RECT -79.585 -1017.865 -79.255 -1017.535 ;
      RECT -80.715 -1014.205 -80.385 -1013.875 ;
      RECT -80.7 -1025.18 -80.4 -1013.875 ;
      RECT -81.58 -1017.91 -81.18 -994.725 ;
      RECT -81.72 -1025.06 -81.3 -1017.49 ;
  END
END sramgen_sram_4096x8m8w8_replica_v1

END LIBRARY
