VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_64x22m4w22
    CLASS BLOCK  ;
    FOREIGN sram22_64x22m4w22   ;
    SIZE 286.880 BY 193.720 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 139.150 0.000 139.290 0.140 ;
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 145.250 0.000 145.390 0.140 ;
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 151.350 0.000 151.490 0.140 ;
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 157.450 0.000 157.590 0.140 ;
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.550 0.000 163.690 0.140 ;
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 169.650 0.000 169.790 0.140 ;
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 175.750 0.000 175.890 0.140 ;
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 181.850 0.000 181.990 0.140 ;
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 187.950 0.000 188.090 0.140 ;
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.050 0.000 194.190 0.140 ;
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 200.150 0.000 200.290 0.140 ;
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 206.250 0.000 206.390 0.140 ;
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 212.350 0.000 212.490 0.140 ;
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 218.450 0.000 218.590 0.140 ;
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 224.550 0.000 224.690 0.140 ;
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 230.650 0.000 230.790 0.140 ;
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 236.750 0.000 236.890 0.140 ;
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 242.850 0.000 242.990 0.140 ;
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 248.950 0.000 249.090 0.140 ;
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 255.050 0.000 255.190 0.140 ;
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 261.150 0.000 261.290 0.140 ;
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.471200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 267.250 0.000 267.390 0.140 ;
        END 
    END dout[21] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 138.730 0.000 138.870 0.140 ;
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 144.830 0.000 144.970 0.140 ;
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 150.930 0.000 151.070 0.140 ;
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 157.030 0.000 157.170 0.140 ;
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.130 0.000 163.270 0.140 ;
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 169.230 0.000 169.370 0.140 ;
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 175.330 0.000 175.470 0.140 ;
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 181.430 0.000 181.570 0.140 ;
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 187.530 0.000 187.670 0.140 ;
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 193.630 0.000 193.770 0.140 ;
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 199.730 0.000 199.870 0.140 ;
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 205.830 0.000 205.970 0.140 ;
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 211.930 0.000 212.070 0.140 ;
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 218.030 0.000 218.170 0.140 ;
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 224.130 0.000 224.270 0.140 ;
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 230.230 0.000 230.370 0.140 ;
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 236.330 0.000 236.470 0.140 ;
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 242.430 0.000 242.570 0.140 ;
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 248.530 0.000 248.670 0.140 ;
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 254.630 0.000 254.770 0.140 ;
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 260.730 0.000 260.870 0.140 ;
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.437300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.192800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 266.830 0.000 266.970 0.140 ;
        END 
    END din[21] 
    PIN wmask 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.247700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 138.380 0.000 138.520 0.140 ;
        END 
    END wmask 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 97.040 0.000 97.360 0.320 ;
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 90.920 0.000 91.240 0.320 ;
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 84.800 0.000 85.120 0.320 ;
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 78.680 0.000 79.000 0.320 ;
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 72.560 0.000 72.880 0.320 ;
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 66.440 0.000 66.760 0.320 ;
        END 
    END addr[5] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 109.280 0.000 109.600 0.320 ;
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 103.160 0.000 103.480 0.320 ;
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 15.345000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 112.000 0.000 112.320 0.320 ;
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 19.251000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 112.680 0.000 113.000 0.320 ;
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 138.160 6.240 ;
                RECT 139.880 5.920 144.280 6.240 ;
                RECT 146.000 5.920 150.400 6.240 ;
                RECT 152.120 5.920 156.520 6.240 ;
                RECT 158.240 5.920 162.640 6.240 ;
                RECT 164.360 5.920 168.760 6.240 ;
                RECT 170.480 5.920 174.880 6.240 ;
                RECT 176.600 5.920 181.000 6.240 ;
                RECT 182.720 5.920 187.120 6.240 ;
                RECT 188.840 5.920 193.240 6.240 ;
                RECT 194.960 5.920 199.360 6.240 ;
                RECT 201.080 5.920 205.480 6.240 ;
                RECT 207.200 5.920 211.600 6.240 ;
                RECT 213.320 5.920 217.720 6.240 ;
                RECT 219.440 5.920 223.840 6.240 ;
                RECT 225.560 5.920 229.960 6.240 ;
                RECT 231.680 5.920 236.080 6.240 ;
                RECT 237.800 5.920 242.200 6.240 ;
                RECT 243.920 5.920 248.320 6.240 ;
                RECT 250.040 5.920 254.440 6.240 ;
                RECT 256.160 5.920 260.560 6.240 ;
                RECT 262.280 5.920 266.680 6.240 ;
                RECT 268.400 5.920 286.720 6.240 ;
                RECT 0.160 7.280 286.720 7.600 ;
                RECT 0.160 8.640 286.720 8.960 ;
                RECT 0.160 10.000 111.640 10.320 ;
                RECT 134.440 10.000 286.720 10.320 ;
                RECT 0.160 11.360 286.720 11.680 ;
                RECT 0.160 12.720 286.720 13.040 ;
                RECT 0.160 14.080 62.680 14.400 ;
                RECT 113.360 14.080 286.720 14.400 ;
                RECT 0.160 15.440 286.720 15.760 ;
                RECT 0.160 16.800 286.720 17.120 ;
                RECT 0.160 18.160 62.680 18.480 ;
                RECT 112.680 18.160 286.720 18.480 ;
                RECT 0.160 19.520 286.720 19.840 ;
                RECT 0.160 20.880 286.720 21.200 ;
                RECT 0.160 22.240 127.960 22.560 ;
                RECT 276.560 22.240 286.720 22.560 ;
                RECT 0.160 23.600 127.960 23.920 ;
                RECT 276.560 23.600 286.720 23.920 ;
                RECT 0.160 24.960 127.960 25.280 ;
                RECT 276.560 24.960 286.720 25.280 ;
                RECT 0.160 26.320 127.960 26.640 ;
                RECT 276.560 26.320 286.720 26.640 ;
                RECT 0.160 27.680 127.960 28.000 ;
                RECT 276.560 27.680 286.720 28.000 ;
                RECT 0.160 29.040 127.960 29.360 ;
                RECT 276.560 29.040 286.720 29.360 ;
                RECT 0.160 30.400 127.960 30.720 ;
                RECT 276.560 30.400 286.720 30.720 ;
                RECT 0.160 31.760 79.000 32.080 ;
                RECT 90.240 31.760 127.960 32.080 ;
                RECT 276.560 31.760 286.720 32.080 ;
                RECT 0.160 33.120 77.640 33.440 ;
                RECT 96.360 33.120 127.960 33.440 ;
                RECT 276.560 33.120 286.720 33.440 ;
                RECT 0.160 34.480 57.920 34.800 ;
                RECT 113.360 34.480 127.960 34.800 ;
                RECT 276.560 34.480 286.720 34.800 ;
                RECT 0.160 35.840 57.240 36.160 ;
                RECT 109.280 35.840 127.960 36.160 ;
                RECT 276.560 35.840 286.720 36.160 ;
                RECT 0.160 37.200 127.960 37.520 ;
                RECT 276.560 37.200 286.720 37.520 ;
                RECT 0.160 38.560 127.960 38.880 ;
                RECT 276.560 38.560 286.720 38.880 ;
                RECT 0.160 39.920 127.280 40.240 ;
                RECT 276.560 39.920 286.720 40.240 ;
                RECT 0.160 41.280 127.960 41.600 ;
                RECT 276.560 41.280 286.720 41.600 ;
                RECT 0.160 42.640 53.160 42.960 ;
                RECT 64.400 42.640 127.960 42.960 ;
                RECT 276.560 42.640 286.720 42.960 ;
                RECT 0.160 44.000 54.520 44.320 ;
                RECT 60.320 44.000 68.120 44.320 ;
                RECT 70.520 44.000 127.960 44.320 ;
                RECT 276.560 44.000 286.720 44.320 ;
                RECT 0.160 45.360 55.880 45.680 ;
                RECT 59.640 45.360 127.960 45.680 ;
                RECT 276.560 45.360 286.720 45.680 ;
                RECT 0.160 46.720 62.680 47.040 ;
                RECT 69.840 46.720 127.960 47.040 ;
                RECT 276.560 46.720 286.720 47.040 ;
                RECT 0.160 48.080 65.400 48.400 ;
                RECT 71.200 48.080 106.880 48.400 ;
                RECT 111.320 48.080 127.960 48.400 ;
                RECT 276.560 48.080 286.720 48.400 ;
                RECT 0.160 49.440 55.200 49.760 ;
                RECT 64.400 49.440 106.880 49.760 ;
                RECT 276.560 49.440 286.720 49.760 ;
                RECT 0.160 50.800 58.600 51.120 ;
                RECT 63.720 50.800 106.880 51.120 ;
                RECT 111.320 50.800 127.960 51.120 ;
                RECT 276.560 50.800 286.720 51.120 ;
                RECT 0.160 52.160 106.880 52.480 ;
                RECT 111.320 52.160 127.960 52.480 ;
                RECT 276.560 52.160 286.720 52.480 ;
                RECT 0.160 53.520 54.520 53.840 ;
                RECT 64.400 53.520 127.960 53.840 ;
                RECT 276.560 53.520 286.720 53.840 ;
                RECT 0.160 54.880 62.000 55.200 ;
                RECT 70.520 54.880 127.960 55.200 ;
                RECT 276.560 54.880 286.720 55.200 ;
                RECT 0.160 56.240 127.960 56.560 ;
                RECT 276.560 56.240 286.720 56.560 ;
                RECT 0.160 57.600 62.680 57.920 ;
                RECT 68.480 57.600 88.520 57.920 ;
                RECT 110.640 57.600 127.960 57.920 ;
                RECT 276.560 57.600 286.720 57.920 ;
                RECT 0.160 58.960 65.400 59.280 ;
                RECT 70.520 58.960 78.320 59.280 ;
                RECT 82.760 58.960 88.520 59.280 ;
                RECT 110.640 58.960 127.960 59.280 ;
                RECT 276.560 58.960 286.720 59.280 ;
                RECT 0.160 60.320 59.280 60.640 ;
                RECT 64.400 60.320 79.680 60.640 ;
                RECT 82.080 60.320 88.520 60.640 ;
                RECT 118.800 60.320 127.960 60.640 ;
                RECT 276.560 60.320 286.720 60.640 ;
                RECT 0.160 61.680 88.520 62.000 ;
                RECT 120.160 61.680 127.960 62.000 ;
                RECT 276.560 61.680 286.720 62.000 ;
                RECT 0.160 63.040 53.160 63.360 ;
                RECT 75.960 63.040 88.520 63.360 ;
                RECT 120.160 63.040 127.960 63.360 ;
                RECT 276.560 63.040 286.720 63.360 ;
                RECT 0.160 64.400 62.680 64.720 ;
                RECT 70.520 64.400 88.520 64.720 ;
                RECT 118.800 64.400 127.960 64.720 ;
                RECT 276.560 64.400 286.720 64.720 ;
                RECT 0.160 65.760 62.000 66.080 ;
                RECT 64.400 65.760 71.520 66.080 ;
                RECT 78.000 65.760 88.520 66.080 ;
                RECT 120.160 65.760 127.960 66.080 ;
                RECT 276.560 65.760 286.720 66.080 ;
                RECT 0.160 67.120 53.160 67.440 ;
                RECT 67.120 67.120 88.520 67.440 ;
                RECT 110.640 67.120 127.960 67.440 ;
                RECT 276.560 67.120 286.720 67.440 ;
                RECT 0.160 68.480 62.000 68.800 ;
                RECT 70.520 68.480 88.520 68.800 ;
                RECT 122.880 68.480 127.960 68.800 ;
                RECT 276.560 68.480 286.720 68.800 ;
                RECT 0.160 69.840 59.960 70.160 ;
                RECT 63.720 69.840 88.520 70.160 ;
                RECT 122.880 69.840 127.960 70.160 ;
                RECT 276.560 69.840 286.720 70.160 ;
                RECT 0.160 71.200 55.200 71.520 ;
                RECT 59.640 71.200 62.680 71.520 ;
                RECT 71.200 71.200 88.520 71.520 ;
                RECT 121.520 71.200 127.960 71.520 ;
                RECT 276.560 71.200 286.720 71.520 ;
                RECT 0.160 72.560 57.920 72.880 ;
                RECT 61.680 72.560 88.520 72.880 ;
                RECT 122.880 72.560 127.960 72.880 ;
                RECT 276.560 72.560 286.720 72.880 ;
                RECT 0.160 73.920 54.520 74.240 ;
                RECT 58.280 73.920 88.520 74.240 ;
                RECT 122.880 73.920 127.960 74.240 ;
                RECT 276.560 73.920 286.720 74.240 ;
                RECT 0.160 75.280 58.600 75.600 ;
                RECT 64.400 75.280 88.520 75.600 ;
                RECT 110.640 75.280 127.960 75.600 ;
                RECT 276.560 75.280 286.720 75.600 ;
                RECT 0.160 76.640 54.520 76.960 ;
                RECT 70.520 76.640 88.520 76.960 ;
                RECT 125.600 76.640 127.960 76.960 ;
                RECT 276.560 76.640 286.720 76.960 ;
                RECT 0.160 78.000 62.000 78.320 ;
                RECT 66.440 78.000 88.520 78.320 ;
                RECT 124.240 78.000 127.960 78.320 ;
                RECT 276.560 78.000 286.720 78.320 ;
                RECT 0.160 79.360 88.520 79.680 ;
                RECT 125.600 79.360 127.960 79.680 ;
                RECT 276.560 79.360 286.720 79.680 ;
                RECT 0.160 80.720 62.680 81.040 ;
                RECT 66.440 80.720 88.520 81.040 ;
                RECT 125.600 80.720 127.960 81.040 ;
                RECT 276.560 80.720 286.720 81.040 ;
                RECT 0.160 82.080 53.160 82.400 ;
                RECT 60.320 82.080 88.520 82.400 ;
                RECT 125.600 82.080 127.960 82.400 ;
                RECT 276.560 82.080 286.720 82.400 ;
                RECT 0.160 83.440 59.280 83.760 ;
                RECT 64.400 83.440 88.520 83.760 ;
                RECT 124.240 83.440 127.960 83.760 ;
                RECT 276.560 83.440 286.720 83.760 ;
                RECT 0.160 84.800 56.560 85.120 ;
                RECT 63.720 84.800 88.520 85.120 ;
                RECT 110.640 84.800 127.960 85.120 ;
                RECT 276.560 84.800 286.720 85.120 ;
                RECT 0.160 86.160 62.000 86.480 ;
                RECT 65.080 86.160 88.520 86.480 ;
                RECT 276.560 86.160 286.720 86.480 ;
                RECT 0.160 87.520 58.600 87.840 ;
                RECT 70.520 87.520 88.520 87.840 ;
                RECT 276.560 87.520 286.720 87.840 ;
                RECT 0.160 88.880 88.520 89.200 ;
                RECT 276.560 88.880 286.720 89.200 ;
                RECT 0.160 90.240 49.760 90.560 ;
                RECT 67.120 90.240 88.520 90.560 ;
                RECT 276.560 90.240 286.720 90.560 ;
                RECT 0.160 91.600 88.520 91.920 ;
                RECT 276.560 91.600 286.720 91.920 ;
                RECT 0.160 92.960 88.520 93.280 ;
                RECT 110.640 92.960 127.960 93.280 ;
                RECT 276.560 92.960 286.720 93.280 ;
                RECT 0.160 94.320 127.960 94.640 ;
                RECT 276.560 94.320 286.720 94.640 ;
                RECT 0.160 95.680 65.400 96.000 ;
                RECT 73.240 95.680 127.960 96.000 ;
                RECT 276.560 95.680 286.720 96.000 ;
                RECT 0.160 97.040 68.800 97.360 ;
                RECT 71.200 97.040 127.960 97.360 ;
                RECT 276.560 97.040 286.720 97.360 ;
                RECT 0.160 98.400 127.960 98.720 ;
                RECT 276.560 98.400 286.720 98.720 ;
                RECT 0.160 99.760 53.160 100.080 ;
                RECT 58.280 99.760 76.960 100.080 ;
                RECT 88.200 99.760 91.240 100.080 ;
                RECT 111.320 99.760 127.960 100.080 ;
                RECT 276.560 99.760 286.720 100.080 ;
                RECT 0.160 101.120 91.240 101.440 ;
                RECT 111.320 101.120 127.960 101.440 ;
                RECT 276.560 101.120 286.720 101.440 ;
                RECT 0.160 102.480 91.240 102.800 ;
                RECT 111.320 102.480 127.960 102.800 ;
                RECT 276.560 102.480 286.720 102.800 ;
                RECT 0.160 103.840 91.240 104.160 ;
                RECT 111.320 103.840 127.960 104.160 ;
                RECT 276.560 103.840 286.720 104.160 ;
                RECT 0.160 105.200 62.000 105.520 ;
                RECT 70.520 105.200 91.240 105.520 ;
                RECT 111.320 105.200 127.960 105.520 ;
                RECT 276.560 105.200 286.720 105.520 ;
                RECT 0.160 106.560 91.240 106.880 ;
                RECT 111.320 106.560 127.960 106.880 ;
                RECT 276.560 106.560 286.720 106.880 ;
                RECT 0.160 107.920 91.240 108.240 ;
                RECT 111.320 107.920 127.960 108.240 ;
                RECT 276.560 107.920 286.720 108.240 ;
                RECT 0.160 109.280 55.200 109.600 ;
                RECT 60.320 109.280 91.240 109.600 ;
                RECT 111.320 109.280 127.960 109.600 ;
                RECT 276.560 109.280 286.720 109.600 ;
                RECT 0.160 110.640 91.240 110.960 ;
                RECT 111.320 110.640 127.960 110.960 ;
                RECT 276.560 110.640 286.720 110.960 ;
                RECT 0.160 112.000 31.400 112.320 ;
                RECT 50.120 112.000 58.600 112.320 ;
                RECT 61.000 112.000 91.240 112.320 ;
                RECT 276.560 112.000 286.720 112.320 ;
                RECT 0.160 113.360 31.400 113.680 ;
                RECT 50.120 113.360 91.240 113.680 ;
                RECT 111.320 113.360 125.240 113.680 ;
                RECT 276.560 113.360 286.720 113.680 ;
                RECT 0.160 114.720 31.400 115.040 ;
                RECT 50.120 114.720 91.240 115.040 ;
                RECT 111.320 114.720 122.520 115.040 ;
                RECT 276.560 114.720 286.720 115.040 ;
                RECT 0.160 116.080 31.400 116.400 ;
                RECT 50.120 116.080 54.520 116.400 ;
                RECT 57.600 116.080 91.240 116.400 ;
                RECT 111.320 116.080 119.800 116.400 ;
                RECT 276.560 116.080 286.720 116.400 ;
                RECT 0.160 117.440 31.400 117.760 ;
                RECT 50.120 117.440 55.200 117.760 ;
                RECT 60.320 117.440 91.240 117.760 ;
                RECT 111.320 117.440 117.080 117.760 ;
                RECT 276.560 117.440 286.720 117.760 ;
                RECT 0.160 118.800 31.400 119.120 ;
                RECT 50.800 118.800 91.240 119.120 ;
                RECT 111.320 118.800 127.960 119.120 ;
                RECT 276.560 118.800 286.720 119.120 ;
                RECT 0.160 120.160 31.400 120.480 ;
                RECT 50.120 120.160 127.960 120.480 ;
                RECT 276.560 120.160 286.720 120.480 ;
                RECT 0.160 121.520 31.400 121.840 ;
                RECT 50.120 121.520 127.960 121.840 ;
                RECT 276.560 121.520 286.720 121.840 ;
                RECT 0.160 122.880 31.400 123.200 ;
                RECT 50.120 122.880 127.960 123.200 ;
                RECT 276.560 122.880 286.720 123.200 ;
                RECT 0.160 124.240 31.400 124.560 ;
                RECT 50.120 124.240 127.960 124.560 ;
                RECT 276.560 124.240 286.720 124.560 ;
                RECT 0.160 125.600 31.400 125.920 ;
                RECT 50.120 125.600 91.240 125.920 ;
                RECT 111.320 125.600 127.960 125.920 ;
                RECT 276.560 125.600 286.720 125.920 ;
                RECT 0.160 126.960 31.400 127.280 ;
                RECT 50.120 126.960 91.240 127.280 ;
                RECT 111.320 126.960 118.440 127.280 ;
                RECT 276.560 126.960 286.720 127.280 ;
                RECT 0.160 128.320 31.400 128.640 ;
                RECT 50.120 128.320 56.560 128.640 ;
                RECT 60.320 128.320 91.240 128.640 ;
                RECT 111.320 128.320 121.160 128.640 ;
                RECT 276.560 128.320 286.720 128.640 ;
                RECT 0.160 129.680 91.240 130.000 ;
                RECT 111.320 129.680 123.880 130.000 ;
                RECT 276.560 129.680 286.720 130.000 ;
                RECT 0.160 131.040 91.240 131.360 ;
                RECT 111.320 131.040 126.600 131.360 ;
                RECT 276.560 131.040 286.720 131.360 ;
                RECT 0.160 132.400 58.600 132.720 ;
                RECT 65.080 132.400 91.240 132.720 ;
                RECT 276.560 132.400 286.720 132.720 ;
                RECT 0.160 133.760 15.080 134.080 ;
                RECT 31.760 133.760 37.520 134.080 ;
                RECT 45.360 133.760 91.240 134.080 ;
                RECT 111.320 133.760 127.960 134.080 ;
                RECT 276.560 133.760 286.720 134.080 ;
                RECT 0.160 135.120 15.080 135.440 ;
                RECT 49.440 135.120 91.240 135.440 ;
                RECT 111.320 135.120 127.960 135.440 ;
                RECT 276.560 135.120 286.720 135.440 ;
                RECT 0.160 136.480 15.080 136.800 ;
                RECT 49.440 136.480 91.240 136.800 ;
                RECT 276.560 136.480 286.720 136.800 ;
                RECT 0.160 137.840 15.080 138.160 ;
                RECT 31.760 137.840 37.520 138.160 ;
                RECT 45.360 137.840 57.240 138.160 ;
                RECT 63.720 137.840 91.240 138.160 ;
                RECT 276.560 137.840 286.720 138.160 ;
                RECT 0.160 139.200 15.760 139.520 ;
                RECT 44.680 139.200 91.240 139.520 ;
                RECT 111.320 139.200 286.720 139.520 ;
                RECT 0.160 140.560 44.320 140.880 ;
                RECT 88.880 140.560 286.720 140.880 ;
                RECT 0.160 141.920 125.240 142.240 ;
                RECT 279.280 141.920 286.720 142.240 ;
                RECT 0.160 143.280 125.240 143.600 ;
                RECT 279.280 143.280 286.720 143.600 ;
                RECT 0.160 144.640 125.240 144.960 ;
                RECT 279.280 144.640 286.720 144.960 ;
                RECT 0.160 146.000 28.680 146.320 ;
                RECT 35.160 146.000 36.840 146.320 ;
                RECT 46.040 146.000 74.240 146.320 ;
                RECT 279.280 146.000 286.720 146.320 ;
                RECT 0.160 147.360 26.640 147.680 ;
                RECT 44.680 147.360 55.880 147.680 ;
                RECT 57.600 147.360 74.240 147.680 ;
                RECT 279.280 147.360 286.720 147.680 ;
                RECT 0.160 148.720 26.640 149.040 ;
                RECT 37.200 148.720 55.880 149.040 ;
                RECT 59.640 148.720 74.240 149.040 ;
                RECT 279.280 148.720 286.720 149.040 ;
                RECT 0.160 150.080 26.640 150.400 ;
                RECT 37.200 150.080 55.880 150.400 ;
                RECT 60.320 150.080 74.240 150.400 ;
                RECT 279.280 150.080 286.720 150.400 ;
                RECT 0.160 151.440 55.880 151.760 ;
                RECT 61.000 151.440 74.240 151.760 ;
                RECT 279.280 151.440 286.720 151.760 ;
                RECT 0.160 152.800 26.640 153.120 ;
                RECT 37.200 152.800 55.880 153.120 ;
                RECT 57.600 152.800 74.240 153.120 ;
                RECT 279.280 152.800 286.720 153.120 ;
                RECT 0.160 154.160 26.640 154.480 ;
                RECT 37.200 154.160 74.240 154.480 ;
                RECT 279.280 154.160 286.720 154.480 ;
                RECT 0.160 155.520 74.240 155.840 ;
                RECT 279.280 155.520 286.720 155.840 ;
                RECT 0.160 156.880 74.240 157.200 ;
                RECT 279.280 156.880 286.720 157.200 ;
                RECT 0.160 158.240 14.400 158.560 ;
                RECT 22.240 158.240 74.240 158.560 ;
                RECT 279.280 158.240 286.720 158.560 ;
                RECT 0.160 159.600 74.240 159.920 ;
                RECT 279.280 159.600 286.720 159.920 ;
                RECT 0.160 160.960 13.720 161.280 ;
                RECT 22.240 160.960 35.480 161.280 ;
                RECT 38.560 160.960 74.240 161.280 ;
                RECT 279.280 160.960 286.720 161.280 ;
                RECT 0.160 162.320 13.040 162.640 ;
                RECT 22.240 162.320 35.480 162.640 ;
                RECT 45.360 162.320 74.240 162.640 ;
                RECT 279.280 162.320 286.720 162.640 ;
                RECT 0.160 163.680 12.360 164.000 ;
                RECT 22.240 163.680 35.480 164.000 ;
                RECT 44.680 163.680 55.880 164.000 ;
                RECT 57.600 163.680 74.240 164.000 ;
                RECT 279.280 163.680 286.720 164.000 ;
                RECT 0.160 165.040 55.880 165.360 ;
                RECT 58.280 165.040 74.240 165.360 ;
                RECT 279.280 165.040 286.720 165.360 ;
                RECT 0.160 166.400 11.680 166.720 ;
                RECT 22.240 166.400 35.480 166.720 ;
                RECT 40.600 166.400 55.880 166.720 ;
                RECT 58.280 166.400 74.240 166.720 ;
                RECT 279.280 166.400 286.720 166.720 ;
                RECT 0.160 167.760 11.000 168.080 ;
                RECT 22.240 167.760 55.880 168.080 ;
                RECT 58.960 167.760 74.240 168.080 ;
                RECT 279.280 167.760 286.720 168.080 ;
                RECT 0.160 169.120 10.320 169.440 ;
                RECT 22.240 169.120 55.880 169.440 ;
                RECT 59.640 169.120 74.240 169.440 ;
                RECT 279.280 169.120 286.720 169.440 ;
                RECT 0.160 170.480 9.640 170.800 ;
                RECT 22.240 170.480 74.240 170.800 ;
                RECT 279.280 170.480 286.720 170.800 ;
                RECT 0.160 171.840 74.240 172.160 ;
                RECT 279.280 171.840 286.720 172.160 ;
                RECT 0.160 173.200 74.240 173.520 ;
                RECT 279.280 173.200 286.720 173.520 ;
                RECT 0.160 174.560 74.240 174.880 ;
                RECT 279.280 174.560 286.720 174.880 ;
                RECT 0.160 175.920 74.240 176.240 ;
                RECT 279.280 175.920 286.720 176.240 ;
                RECT 0.160 177.280 74.240 177.600 ;
                RECT 279.280 177.280 286.720 177.600 ;
                RECT 0.160 178.640 74.240 178.960 ;
                RECT 279.280 178.640 286.720 178.960 ;
                RECT 0.160 180.000 125.240 180.320 ;
                RECT 279.280 180.000 286.720 180.320 ;
                RECT 0.160 181.360 125.240 181.680 ;
                RECT 279.280 181.360 286.720 181.680 ;
                RECT 0.160 182.720 125.240 183.040 ;
                RECT 279.280 182.720 286.720 183.040 ;
                RECT 0.160 184.080 286.720 184.400 ;
                RECT 0.160 185.440 286.720 185.760 ;
                RECT 0.160 186.800 286.720 187.120 ;
                RECT 0.160 188.160 286.720 188.480 ;
                RECT 0.160 0.160 286.720 1.520 ;
                RECT 0.160 192.200 286.720 193.560 ;
                RECT 129.380 43.695 135.180 45.065 ;
                RECT 269.080 43.695 274.880 45.065 ;
                RECT 129.380 49.385 135.180 51.255 ;
                RECT 269.080 49.385 274.880 51.255 ;
                RECT 129.380 55.205 135.180 56.605 ;
                RECT 269.080 55.205 274.880 56.605 ;
                RECT 129.380 60.315 135.180 61.715 ;
                RECT 269.080 60.315 274.880 61.715 ;
                RECT 129.380 68.490 274.880 70.290 ;
                RECT 129.380 134.745 274.880 135.545 ;
                RECT 129.380 120.420 274.880 121.290 ;
                RECT 129.380 87.860 274.880 88.660 ;
                RECT 129.380 98.165 274.880 98.455 ;
                RECT 129.380 79.960 274.880 80.760 ;
                RECT 129.380 94.085 274.880 94.885 ;
                RECT 129.380 82.970 274.880 83.770 ;
                RECT 129.380 27.940 274.880 29.740 ;
                RECT 80.980 145.715 82.900 178.895 ;
                RECT 84.820 145.715 86.740 178.895 ;
                RECT 101.775 145.715 103.695 178.895 ;
                RECT 105.615 145.715 107.535 178.895 ;
                RECT 109.455 145.715 111.375 178.895 ;
                RECT 113.295 145.715 115.215 178.895 ;
                RECT 117.135 145.715 119.055 178.895 ;
                RECT 120.975 145.715 122.895 178.895 ;
                RECT 92.165 57.820 94.085 93.220 ;
                RECT 99.785 57.820 101.705 93.220 ;
                RECT 108.050 57.820 109.970 93.220 ;
                RECT 95.370 125.020 97.290 139.080 ;
                RECT 102.215 125.020 103.965 139.080 ;
                RECT 108.675 125.020 110.595 139.080 ;
                RECT 95.155 99.220 97.075 119.020 ;
                RECT 102.215 99.220 103.965 119.020 ;
                RECT 108.675 99.220 110.595 119.020 ;
                RECT 109.640 48.240 110.960 51.820 ;
                RECT 27.260 147.985 36.420 148.735 ;
                RECT 27.260 152.610 36.420 154.360 ;
                RECT 32.910 135.770 48.950 136.570 ;
                RECT 16.110 136.480 30.950 138.170 ;
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 138.160 5.560 ;
                RECT 139.880 5.240 144.280 5.560 ;
                RECT 146.000 5.240 150.400 5.560 ;
                RECT 152.120 5.240 156.520 5.560 ;
                RECT 158.240 5.240 162.640 5.560 ;
                RECT 164.360 5.240 168.760 5.560 ;
                RECT 170.480 5.240 174.880 5.560 ;
                RECT 176.600 5.240 181.000 5.560 ;
                RECT 182.720 5.240 187.120 5.560 ;
                RECT 188.840 5.240 193.240 5.560 ;
                RECT 194.960 5.240 199.360 5.560 ;
                RECT 201.080 5.240 205.480 5.560 ;
                RECT 207.200 5.240 211.600 5.560 ;
                RECT 213.320 5.240 217.720 5.560 ;
                RECT 219.440 5.240 223.840 5.560 ;
                RECT 225.560 5.240 229.960 5.560 ;
                RECT 231.680 5.240 236.080 5.560 ;
                RECT 237.800 5.240 242.200 5.560 ;
                RECT 243.920 5.240 248.320 5.560 ;
                RECT 250.040 5.240 254.440 5.560 ;
                RECT 256.160 5.240 260.560 5.560 ;
                RECT 262.280 5.240 266.680 5.560 ;
                RECT 268.400 5.240 284.000 5.560 ;
                RECT 2.880 6.600 284.000 6.920 ;
                RECT 2.880 7.960 284.000 8.280 ;
                RECT 2.880 9.320 112.320 9.640 ;
                RECT 133.760 9.320 284.000 9.640 ;
                RECT 2.880 10.680 284.000 11.000 ;
                RECT 2.880 12.040 284.000 12.360 ;
                RECT 2.880 13.400 62.680 13.720 ;
                RECT 113.360 13.400 284.000 13.720 ;
                RECT 2.880 14.760 284.000 15.080 ;
                RECT 2.880 16.120 284.000 16.440 ;
                RECT 2.880 17.480 62.680 17.800 ;
                RECT 112.680 17.480 284.000 17.800 ;
                RECT 2.880 18.840 284.000 19.160 ;
                RECT 2.880 20.200 284.000 20.520 ;
                RECT 2.880 21.560 127.960 21.880 ;
                RECT 276.560 21.560 284.000 21.880 ;
                RECT 2.880 22.920 127.960 23.240 ;
                RECT 276.560 22.920 284.000 23.240 ;
                RECT 2.880 24.280 127.960 24.600 ;
                RECT 276.560 24.280 284.000 24.600 ;
                RECT 2.880 25.640 127.960 25.960 ;
                RECT 276.560 25.640 284.000 25.960 ;
                RECT 2.880 27.000 127.960 27.320 ;
                RECT 276.560 27.000 284.000 27.320 ;
                RECT 2.880 28.360 127.960 28.680 ;
                RECT 276.560 28.360 284.000 28.680 ;
                RECT 2.880 29.720 127.960 30.040 ;
                RECT 276.560 29.720 284.000 30.040 ;
                RECT 2.880 31.080 79.680 31.400 ;
                RECT 91.600 31.080 127.960 31.400 ;
                RECT 276.560 31.080 284.000 31.400 ;
                RECT 2.880 32.440 78.320 32.760 ;
                RECT 97.720 32.440 127.960 32.760 ;
                RECT 276.560 32.440 284.000 32.760 ;
                RECT 2.880 33.800 55.200 34.120 ;
                RECT 112.680 33.800 127.960 34.120 ;
                RECT 276.560 33.800 284.000 34.120 ;
                RECT 2.880 35.160 55.880 35.480 ;
                RECT 103.160 35.160 127.960 35.480 ;
                RECT 276.560 35.160 284.000 35.480 ;
                RECT 2.880 36.520 127.960 36.840 ;
                RECT 276.560 36.520 284.000 36.840 ;
                RECT 2.880 37.880 127.960 38.200 ;
                RECT 276.560 37.880 284.000 38.200 ;
                RECT 2.880 39.240 127.280 39.560 ;
                RECT 276.560 39.240 284.000 39.560 ;
                RECT 2.880 40.600 127.960 40.920 ;
                RECT 276.560 40.600 284.000 40.920 ;
                RECT 2.880 41.960 53.160 42.280 ;
                RECT 64.400 41.960 127.960 42.280 ;
                RECT 276.560 41.960 284.000 42.280 ;
                RECT 2.880 43.320 54.520 43.640 ;
                RECT 56.920 43.320 127.960 43.640 ;
                RECT 276.560 43.320 284.000 43.640 ;
                RECT 2.880 44.680 55.880 45.000 ;
                RECT 60.320 44.680 68.120 45.000 ;
                RECT 70.520 44.680 127.960 45.000 ;
                RECT 276.560 44.680 284.000 45.000 ;
                RECT 2.880 46.040 55.880 46.360 ;
                RECT 59.640 46.040 127.960 46.360 ;
                RECT 276.560 46.040 284.000 46.360 ;
                RECT 2.880 47.400 62.680 47.720 ;
                RECT 71.200 47.400 127.960 47.720 ;
                RECT 276.560 47.400 284.000 47.720 ;
                RECT 2.880 48.760 57.920 49.080 ;
                RECT 64.400 48.760 106.880 49.080 ;
                RECT 111.320 48.760 127.960 49.080 ;
                RECT 276.560 48.760 284.000 49.080 ;
                RECT 2.880 50.120 55.200 50.440 ;
                RECT 64.400 50.120 106.880 50.440 ;
                RECT 276.560 50.120 284.000 50.440 ;
                RECT 2.880 51.480 76.280 51.800 ;
                RECT 111.320 51.480 127.960 51.800 ;
                RECT 276.560 51.480 284.000 51.800 ;
                RECT 2.880 52.840 54.520 53.160 ;
                RECT 64.400 52.840 127.960 53.160 ;
                RECT 276.560 52.840 284.000 53.160 ;
                RECT 2.880 54.200 62.680 54.520 ;
                RECT 70.520 54.200 127.960 54.520 ;
                RECT 276.560 54.200 284.000 54.520 ;
                RECT 2.880 55.560 62.000 55.880 ;
                RECT 64.400 55.560 127.960 55.880 ;
                RECT 276.560 55.560 284.000 55.880 ;
                RECT 2.880 56.920 127.960 57.240 ;
                RECT 276.560 56.920 284.000 57.240 ;
                RECT 2.880 58.280 62.680 58.600 ;
                RECT 70.520 58.280 77.640 58.600 ;
                RECT 83.440 58.280 88.520 58.600 ;
                RECT 110.640 58.280 127.960 58.600 ;
                RECT 276.560 58.280 284.000 58.600 ;
                RECT 2.880 59.640 59.280 59.960 ;
                RECT 64.400 59.640 79.000 59.960 ;
                RECT 82.760 59.640 88.520 59.960 ;
                RECT 120.160 59.640 127.960 59.960 ;
                RECT 276.560 59.640 284.000 59.960 ;
                RECT 2.880 61.000 62.000 61.320 ;
                RECT 64.400 61.000 88.520 61.320 ;
                RECT 120.160 61.000 127.960 61.320 ;
                RECT 276.560 61.000 284.000 61.320 ;
                RECT 2.880 62.360 65.400 62.680 ;
                RECT 75.960 62.360 88.520 62.680 ;
                RECT 118.800 62.360 127.960 62.680 ;
                RECT 276.560 62.360 284.000 62.680 ;
                RECT 2.880 63.720 53.160 64.040 ;
                RECT 70.520 63.720 88.520 64.040 ;
                RECT 120.160 63.720 127.960 64.040 ;
                RECT 276.560 63.720 284.000 64.040 ;
                RECT 2.880 65.080 71.520 65.400 ;
                RECT 77.320 65.080 88.520 65.400 ;
                RECT 120.160 65.080 127.960 65.400 ;
                RECT 276.560 65.080 284.000 65.400 ;
                RECT 2.880 66.440 62.000 66.760 ;
                RECT 64.400 66.440 74.240 66.760 ;
                RECT 78.000 66.440 88.520 66.760 ;
                RECT 118.800 66.440 127.960 66.760 ;
                RECT 276.560 66.440 284.000 66.760 ;
                RECT 2.880 67.800 53.160 68.120 ;
                RECT 67.120 67.800 88.520 68.120 ;
                RECT 122.880 67.800 127.960 68.120 ;
                RECT 276.560 67.800 284.000 68.120 ;
                RECT 2.880 69.160 62.000 69.480 ;
                RECT 70.520 69.160 88.520 69.480 ;
                RECT 121.520 69.160 127.960 69.480 ;
                RECT 276.560 69.160 284.000 69.480 ;
                RECT 2.880 70.520 59.960 70.840 ;
                RECT 71.200 70.520 88.520 70.840 ;
                RECT 122.880 70.520 127.960 70.840 ;
                RECT 276.560 70.520 284.000 70.840 ;
                RECT 2.880 71.880 55.200 72.200 ;
                RECT 61.680 71.880 88.520 72.200 ;
                RECT 122.880 71.880 127.960 72.200 ;
                RECT 276.560 71.880 284.000 72.200 ;
                RECT 2.880 73.240 88.520 73.560 ;
                RECT 110.640 73.240 127.960 73.560 ;
                RECT 276.560 73.240 284.000 73.560 ;
                RECT 2.880 74.600 54.520 74.920 ;
                RECT 58.280 74.600 88.520 74.920 ;
                RECT 121.520 74.600 127.960 74.920 ;
                RECT 276.560 74.600 284.000 74.920 ;
                RECT 2.880 75.960 54.520 76.280 ;
                RECT 64.400 75.960 88.520 76.280 ;
                RECT 110.640 75.960 127.960 76.280 ;
                RECT 276.560 75.960 284.000 76.280 ;
                RECT 2.880 77.320 58.600 77.640 ;
                RECT 70.520 77.320 88.520 77.640 ;
                RECT 125.600 77.320 127.960 77.640 ;
                RECT 276.560 77.320 284.000 77.640 ;
                RECT 2.880 78.680 62.000 79.000 ;
                RECT 66.440 78.680 88.520 79.000 ;
                RECT 125.600 78.680 127.960 79.000 ;
                RECT 276.560 78.680 284.000 79.000 ;
                RECT 2.880 80.040 62.680 80.360 ;
                RECT 66.440 80.040 88.520 80.360 ;
                RECT 125.600 80.040 127.960 80.360 ;
                RECT 276.560 80.040 284.000 80.360 ;
                RECT 2.880 81.400 88.520 81.720 ;
                RECT 124.240 81.400 127.960 81.720 ;
                RECT 276.560 81.400 284.000 81.720 ;
                RECT 2.880 82.760 53.160 83.080 ;
                RECT 60.320 82.760 88.520 83.080 ;
                RECT 125.600 82.760 127.960 83.080 ;
                RECT 276.560 82.760 284.000 83.080 ;
                RECT 2.880 84.120 56.560 84.440 ;
                RECT 64.400 84.120 88.520 84.440 ;
                RECT 110.640 84.120 127.960 84.440 ;
                RECT 276.560 84.120 284.000 84.440 ;
                RECT 2.880 85.480 62.000 85.800 ;
                RECT 65.080 85.480 88.520 85.800 ;
                RECT 276.560 85.480 284.000 85.800 ;
                RECT 2.880 86.840 88.520 87.160 ;
                RECT 276.560 86.840 284.000 87.160 ;
                RECT 2.880 88.200 58.600 88.520 ;
                RECT 70.520 88.200 88.520 88.520 ;
                RECT 276.560 88.200 284.000 88.520 ;
                RECT 2.880 89.560 49.760 89.880 ;
                RECT 63.720 89.560 88.520 89.880 ;
                RECT 276.560 89.560 284.000 89.880 ;
                RECT 2.880 90.920 59.960 91.240 ;
                RECT 67.120 90.920 88.520 91.240 ;
                RECT 276.560 90.920 284.000 91.240 ;
                RECT 2.880 92.280 88.520 92.600 ;
                RECT 276.560 92.280 284.000 92.600 ;
                RECT 2.880 93.640 127.960 93.960 ;
                RECT 276.560 93.640 284.000 93.960 ;
                RECT 2.880 95.000 65.400 95.320 ;
                RECT 73.240 95.000 127.960 95.320 ;
                RECT 276.560 95.000 284.000 95.320 ;
                RECT 2.880 96.360 127.960 96.680 ;
                RECT 276.560 96.360 284.000 96.680 ;
                RECT 2.880 97.720 68.800 98.040 ;
                RECT 71.200 97.720 127.960 98.040 ;
                RECT 276.560 97.720 284.000 98.040 ;
                RECT 2.880 99.080 55.200 99.400 ;
                RECT 58.280 99.080 91.240 99.400 ;
                RECT 111.320 99.080 127.960 99.400 ;
                RECT 276.560 99.080 284.000 99.400 ;
                RECT 2.880 100.440 53.160 100.760 ;
                RECT 56.920 100.440 91.240 100.760 ;
                RECT 111.320 100.440 127.960 100.760 ;
                RECT 276.560 100.440 284.000 100.760 ;
                RECT 2.880 101.800 91.240 102.120 ;
                RECT 111.320 101.800 127.960 102.120 ;
                RECT 276.560 101.800 284.000 102.120 ;
                RECT 2.880 103.160 91.240 103.480 ;
                RECT 111.320 103.160 127.960 103.480 ;
                RECT 276.560 103.160 284.000 103.480 ;
                RECT 2.880 104.520 91.240 104.840 ;
                RECT 111.320 104.520 127.960 104.840 ;
                RECT 276.560 104.520 284.000 104.840 ;
                RECT 2.880 105.880 62.000 106.200 ;
                RECT 70.520 105.880 91.240 106.200 ;
                RECT 111.320 105.880 127.960 106.200 ;
                RECT 276.560 105.880 284.000 106.200 ;
                RECT 2.880 107.240 91.240 107.560 ;
                RECT 111.320 107.240 127.960 107.560 ;
                RECT 276.560 107.240 284.000 107.560 ;
                RECT 2.880 108.600 55.200 108.920 ;
                RECT 60.320 108.600 91.240 108.920 ;
                RECT 111.320 108.600 127.960 108.920 ;
                RECT 276.560 108.600 284.000 108.920 ;
                RECT 2.880 109.960 91.240 110.280 ;
                RECT 111.320 109.960 127.960 110.280 ;
                RECT 276.560 109.960 284.000 110.280 ;
                RECT 2.880 111.320 31.400 111.640 ;
                RECT 50.120 111.320 58.600 111.640 ;
                RECT 61.000 111.320 91.240 111.640 ;
                RECT 111.320 111.320 127.960 111.640 ;
                RECT 276.560 111.320 284.000 111.640 ;
                RECT 2.880 112.680 31.400 113.000 ;
                RECT 50.120 112.680 91.240 113.000 ;
                RECT 276.560 112.680 284.000 113.000 ;
                RECT 2.880 114.040 31.400 114.360 ;
                RECT 50.120 114.040 91.240 114.360 ;
                RECT 111.320 114.040 125.240 114.360 ;
                RECT 276.560 114.040 284.000 114.360 ;
                RECT 2.880 115.400 31.400 115.720 ;
                RECT 50.120 115.400 54.520 115.720 ;
                RECT 57.600 115.400 91.240 115.720 ;
                RECT 111.320 115.400 122.520 115.720 ;
                RECT 276.560 115.400 284.000 115.720 ;
                RECT 2.880 116.760 31.400 117.080 ;
                RECT 50.120 116.760 55.200 117.080 ;
                RECT 60.320 116.760 91.240 117.080 ;
                RECT 111.320 116.760 117.080 117.080 ;
                RECT 276.560 116.760 284.000 117.080 ;
                RECT 2.880 118.120 31.400 118.440 ;
                RECT 50.120 118.120 91.240 118.440 ;
                RECT 111.320 118.120 117.080 118.440 ;
                RECT 276.560 118.120 284.000 118.440 ;
                RECT 2.880 119.480 31.400 119.800 ;
                RECT 50.120 119.480 127.960 119.800 ;
                RECT 276.560 119.480 284.000 119.800 ;
                RECT 2.880 120.840 31.400 121.160 ;
                RECT 50.120 120.840 127.960 121.160 ;
                RECT 276.560 120.840 284.000 121.160 ;
                RECT 2.880 122.200 31.400 122.520 ;
                RECT 50.120 122.200 127.960 122.520 ;
                RECT 276.560 122.200 284.000 122.520 ;
                RECT 2.880 123.560 31.400 123.880 ;
                RECT 50.120 123.560 127.960 123.880 ;
                RECT 276.560 123.560 284.000 123.880 ;
                RECT 2.880 124.920 31.400 125.240 ;
                RECT 50.120 124.920 91.240 125.240 ;
                RECT 111.320 124.920 127.960 125.240 ;
                RECT 276.560 124.920 284.000 125.240 ;
                RECT 2.880 126.280 31.400 126.600 ;
                RECT 50.120 126.280 91.240 126.600 ;
                RECT 111.320 126.280 118.440 126.600 ;
                RECT 276.560 126.280 284.000 126.600 ;
                RECT 2.880 127.640 31.400 127.960 ;
                RECT 50.120 127.640 56.560 127.960 ;
                RECT 60.320 127.640 91.240 127.960 ;
                RECT 111.320 127.640 118.440 127.960 ;
                RECT 276.560 127.640 284.000 127.960 ;
                RECT 2.880 129.000 31.400 129.320 ;
                RECT 50.120 129.000 91.240 129.320 ;
                RECT 111.320 129.000 121.160 129.320 ;
                RECT 276.560 129.000 284.000 129.320 ;
                RECT 2.880 130.360 91.240 130.680 ;
                RECT 111.320 130.360 123.880 130.680 ;
                RECT 276.560 130.360 284.000 130.680 ;
                RECT 2.880 131.720 91.240 132.040 ;
                RECT 276.560 131.720 284.000 132.040 ;
                RECT 2.880 133.080 15.080 133.400 ;
                RECT 31.760 133.080 58.600 133.400 ;
                RECT 65.080 133.080 91.240 133.400 ;
                RECT 276.560 133.080 284.000 133.400 ;
                RECT 2.880 134.440 15.080 134.760 ;
                RECT 31.760 134.440 37.520 134.760 ;
                RECT 45.360 134.440 91.240 134.760 ;
                RECT 111.320 134.440 127.960 134.760 ;
                RECT 276.560 134.440 284.000 134.760 ;
                RECT 2.880 135.800 15.080 136.120 ;
                RECT 49.440 135.800 91.240 136.120 ;
                RECT 111.320 135.800 127.960 136.120 ;
                RECT 276.560 135.800 284.000 136.120 ;
                RECT 2.880 137.160 15.080 137.480 ;
                RECT 31.760 137.160 91.240 137.480 ;
                RECT 276.560 137.160 284.000 137.480 ;
                RECT 2.880 138.520 15.080 138.840 ;
                RECT 45.360 138.520 57.240 138.840 ;
                RECT 63.720 138.520 91.240 138.840 ;
                RECT 111.320 138.520 127.960 138.840 ;
                RECT 276.560 138.520 284.000 138.840 ;
                RECT 2.880 139.880 37.520 140.200 ;
                RECT 57.600 139.880 284.000 140.200 ;
                RECT 2.880 141.240 33.440 141.560 ;
                RECT 56.920 141.240 284.000 141.560 ;
                RECT 2.880 142.600 125.240 142.920 ;
                RECT 279.280 142.600 284.000 142.920 ;
                RECT 2.880 143.960 125.240 144.280 ;
                RECT 279.280 143.960 284.000 144.280 ;
                RECT 2.880 145.320 28.680 145.640 ;
                RECT 35.160 145.320 74.240 145.640 ;
                RECT 279.280 145.320 284.000 145.640 ;
                RECT 2.880 146.680 26.640 147.000 ;
                RECT 45.360 146.680 74.240 147.000 ;
                RECT 279.280 146.680 284.000 147.000 ;
                RECT 2.880 148.040 26.640 148.360 ;
                RECT 44.680 148.040 55.880 148.360 ;
                RECT 57.600 148.040 74.240 148.360 ;
                RECT 279.280 148.040 284.000 148.360 ;
                RECT 2.880 149.400 55.880 149.720 ;
                RECT 57.600 149.400 74.240 149.720 ;
                RECT 279.280 149.400 284.000 149.720 ;
                RECT 2.880 150.760 26.640 151.080 ;
                RECT 37.200 150.760 55.880 151.080 ;
                RECT 60.320 150.760 74.240 151.080 ;
                RECT 279.280 150.760 284.000 151.080 ;
                RECT 2.880 152.120 26.640 152.440 ;
                RECT 37.200 152.120 55.880 152.440 ;
                RECT 61.000 152.120 74.240 152.440 ;
                RECT 279.280 152.120 284.000 152.440 ;
                RECT 2.880 153.480 26.640 153.800 ;
                RECT 37.200 153.480 55.880 153.800 ;
                RECT 61.680 153.480 74.240 153.800 ;
                RECT 279.280 153.480 284.000 153.800 ;
                RECT 2.880 154.840 74.240 155.160 ;
                RECT 279.280 154.840 284.000 155.160 ;
                RECT 2.880 156.200 74.240 156.520 ;
                RECT 279.280 156.200 284.000 156.520 ;
                RECT 2.880 157.560 74.240 157.880 ;
                RECT 279.280 157.560 284.000 157.880 ;
                RECT 2.880 158.920 14.400 159.240 ;
                RECT 22.240 158.920 35.480 159.240 ;
                RECT 37.880 158.920 74.240 159.240 ;
                RECT 279.280 158.920 284.000 159.240 ;
                RECT 2.880 160.280 13.720 160.600 ;
                RECT 22.240 160.280 74.240 160.600 ;
                RECT 279.280 160.280 284.000 160.600 ;
                RECT 2.880 161.640 13.040 161.960 ;
                RECT 22.240 161.640 39.560 161.960 ;
                RECT 46.040 161.640 74.240 161.960 ;
                RECT 279.280 161.640 284.000 161.960 ;
                RECT 2.880 163.000 12.360 163.320 ;
                RECT 22.240 163.000 40.920 163.320 ;
                RECT 44.680 163.000 74.240 163.320 ;
                RECT 279.280 163.000 284.000 163.320 ;
                RECT 2.880 164.360 55.880 164.680 ;
                RECT 58.280 164.360 74.240 164.680 ;
                RECT 279.280 164.360 284.000 164.680 ;
                RECT 2.880 165.720 11.680 166.040 ;
                RECT 22.240 165.720 55.880 166.040 ;
                RECT 58.280 165.720 74.240 166.040 ;
                RECT 279.280 165.720 284.000 166.040 ;
                RECT 2.880 167.080 55.880 167.400 ;
                RECT 58.960 167.080 74.240 167.400 ;
                RECT 279.280 167.080 284.000 167.400 ;
                RECT 2.880 168.440 11.000 168.760 ;
                RECT 22.240 168.440 35.480 168.760 ;
                RECT 41.280 168.440 55.880 168.760 ;
                RECT 57.600 168.440 74.240 168.760 ;
                RECT 279.280 168.440 284.000 168.760 ;
                RECT 2.880 169.800 10.320 170.120 ;
                RECT 22.240 169.800 35.480 170.120 ;
                RECT 41.960 169.800 55.880 170.120 ;
                RECT 59.640 169.800 74.240 170.120 ;
                RECT 279.280 169.800 284.000 170.120 ;
                RECT 2.880 171.160 9.640 171.480 ;
                RECT 22.240 171.160 35.480 171.480 ;
                RECT 42.640 171.160 74.240 171.480 ;
                RECT 279.280 171.160 284.000 171.480 ;
                RECT 2.880 172.520 74.240 172.840 ;
                RECT 279.280 172.520 284.000 172.840 ;
                RECT 2.880 173.880 74.240 174.200 ;
                RECT 279.280 173.880 284.000 174.200 ;
                RECT 2.880 175.240 74.240 175.560 ;
                RECT 279.280 175.240 284.000 175.560 ;
                RECT 2.880 176.600 74.240 176.920 ;
                RECT 279.280 176.600 284.000 176.920 ;
                RECT 2.880 177.960 74.240 178.280 ;
                RECT 279.280 177.960 284.000 178.280 ;
                RECT 2.880 179.320 125.240 179.640 ;
                RECT 279.280 179.320 284.000 179.640 ;
                RECT 2.880 180.680 125.240 181.000 ;
                RECT 279.280 180.680 284.000 181.000 ;
                RECT 2.880 182.040 125.240 182.360 ;
                RECT 279.280 182.040 284.000 182.360 ;
                RECT 2.880 183.400 284.000 183.720 ;
                RECT 2.880 184.760 284.000 185.080 ;
                RECT 2.880 186.120 284.000 186.440 ;
                RECT 2.880 187.480 284.000 187.800 ;
                RECT 2.880 2.880 284.000 4.240 ;
                RECT 2.880 189.480 284.000 190.840 ;
                RECT 129.380 41.050 135.180 42.170 ;
                RECT 269.080 41.050 274.880 42.170 ;
                RECT 129.380 46.940 135.180 47.760 ;
                RECT 269.080 46.940 274.880 47.760 ;
                RECT 129.380 53.285 135.180 53.915 ;
                RECT 269.080 53.285 274.880 53.915 ;
                RECT 129.380 58.395 135.180 59.025 ;
                RECT 269.080 58.395 274.880 59.025 ;
                RECT 129.380 72.230 274.880 74.030 ;
                RECT 129.380 89.180 274.880 89.980 ;
                RECT 129.380 124.700 274.880 124.945 ;
                RECT 129.380 92.365 274.880 93.165 ;
                RECT 129.380 84.290 274.880 85.090 ;
                RECT 129.380 85.970 274.880 86.770 ;
                RECT 129.380 81.280 274.880 82.080 ;
                RECT 129.380 110.725 274.880 111.015 ;
                RECT 129.380 31.680 274.880 33.480 ;
                RECT 75.245 145.715 77.165 178.895 ;
                RECT 91.910 145.715 93.830 178.895 ;
                RECT 95.750 145.715 97.670 178.895 ;
                RECT 89.540 57.820 90.430 93.220 ;
                RECT 96.405 57.820 97.515 93.220 ;
                RECT 104.455 57.820 105.565 93.220 ;
                RECT 92.205 125.020 93.315 139.080 ;
                RECT 99.720 125.020 100.610 139.080 ;
                RECT 106.050 125.020 106.940 139.080 ;
                RECT 91.775 99.220 92.885 119.020 ;
                RECT 99.720 99.220 100.610 119.020 ;
                RECT 106.050 99.220 106.940 119.020 ;
                RECT 107.680 48.240 108.360 51.820 ;
                RECT 27.260 146.780 36.420 147.150 ;
                RECT 27.260 150.115 36.420 151.005 ;
                RECT 16.110 133.140 30.950 133.810 ;
                RECT 16.110 134.440 30.950 135.450 ;
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 286.880 193.720 ;
        LAYER met2 ;
            RECT 0.000 0.000 286.880 193.720 ;
    END 
END sram22_64x22m4w22 
END LIBRARY 

