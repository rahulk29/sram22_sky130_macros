VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_64x32m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_64x32m4w8   ;
    SIZE 360.320 BY 191.000 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 152.070 0.000 152.210 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 158.170 0.000 158.310 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 164.270 0.000 164.410 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 170.370 0.000 170.510 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 176.470 0.000 176.610 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 182.570 0.000 182.710 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 188.670 0.000 188.810 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.770 0.000 194.910 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 200.870 0.000 201.010 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 206.970 0.000 207.110 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 213.070 0.000 213.210 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 219.170 0.000 219.310 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 225.270 0.000 225.410 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 231.370 0.000 231.510 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 237.470 0.000 237.610 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 243.570 0.000 243.710 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 249.670 0.000 249.810 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 255.770 0.000 255.910 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 261.870 0.000 262.010 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 267.970 0.000 268.110 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 274.070 0.000 274.210 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 280.170 0.000 280.310 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 286.270 0.000 286.410 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 292.370 0.000 292.510 0.140 ; 
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 298.470 0.000 298.610 0.140 ; 
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 304.570 0.000 304.710 0.140 ; 
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 310.670 0.000 310.810 0.140 ; 
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 316.770 0.000 316.910 0.140 ; 
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 322.870 0.000 323.010 0.140 ; 
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 328.970 0.000 329.110 0.140 ; 
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 335.070 0.000 335.210 0.140 ; 
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 341.170 0.000 341.310 0.140 ; 
        END 
    END dout[31] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 151.650 0.000 151.790 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 157.750 0.000 157.890 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.850 0.000 163.990 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 169.950 0.000 170.090 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 176.050 0.000 176.190 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 182.150 0.000 182.290 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 188.250 0.000 188.390 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.350 0.000 194.490 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 200.450 0.000 200.590 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 206.550 0.000 206.690 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 212.650 0.000 212.790 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 218.750 0.000 218.890 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 224.850 0.000 224.990 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 230.950 0.000 231.090 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 237.050 0.000 237.190 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 243.150 0.000 243.290 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 249.250 0.000 249.390 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 255.350 0.000 255.490 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 261.450 0.000 261.590 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 267.550 0.000 267.690 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 273.650 0.000 273.790 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 279.750 0.000 279.890 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 285.850 0.000 285.990 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 291.950 0.000 292.090 0.140 ; 
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 298.050 0.000 298.190 0.140 ; 
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 304.150 0.000 304.290 0.140 ; 
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 310.250 0.000 310.390 0.140 ; 
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 316.350 0.000 316.490 0.140 ; 
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 322.450 0.000 322.590 0.140 ; 
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 328.550 0.000 328.690 0.140 ; 
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 334.650 0.000 334.790 0.140 ; 
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 340.750 0.000 340.890 0.140 ; 
        END 
    END din[31] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.048900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 151.300 0.000 151.440 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.048900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 200.100 0.000 200.240 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.048900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 248.900 0.000 249.040 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.048900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 297.700 0.000 297.840 0.140 ; 
        END 
    END wmask[3] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 109.960 0.000 110.280 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 103.840 0.000 104.160 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 97.720 0.000 98.040 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 91.600 0.000 91.920 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 85.480 0.000 85.800 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 79.360 0.000 79.680 0.320 ; 
        END 
    END addr[5] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 122.200 0.000 122.520 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 116.080 0.000 116.400 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 21.762000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 124.920 0.000 125.240 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 25.668000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 125.600 0.000 125.920 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 151.080 6.240 ; 
                RECT 152.800 5.920 157.200 6.240 ; 
                RECT 158.920 5.920 163.320 6.240 ; 
                RECT 165.040 5.920 169.440 6.240 ; 
                RECT 171.160 5.920 175.560 6.240 ; 
                RECT 177.280 5.920 181.680 6.240 ; 
                RECT 183.400 5.920 187.800 6.240 ; 
                RECT 189.520 5.920 193.920 6.240 ; 
                RECT 195.640 5.920 200.040 6.240 ; 
                RECT 201.760 5.920 206.160 6.240 ; 
                RECT 207.880 5.920 212.280 6.240 ; 
                RECT 214.000 5.920 218.400 6.240 ; 
                RECT 220.120 5.920 224.520 6.240 ; 
                RECT 226.240 5.920 230.640 6.240 ; 
                RECT 232.360 5.920 236.760 6.240 ; 
                RECT 238.480 5.920 242.880 6.240 ; 
                RECT 244.600 5.920 249.000 6.240 ; 
                RECT 250.720 5.920 255.120 6.240 ; 
                RECT 256.840 5.920 261.240 6.240 ; 
                RECT 262.960 5.920 267.360 6.240 ; 
                RECT 269.080 5.920 273.480 6.240 ; 
                RECT 275.200 5.920 279.600 6.240 ; 
                RECT 281.320 5.920 285.720 6.240 ; 
                RECT 287.440 5.920 291.840 6.240 ; 
                RECT 292.880 5.920 297.960 6.240 ; 
                RECT 299.000 5.920 304.080 6.240 ; 
                RECT 305.120 5.920 310.200 6.240 ; 
                RECT 311.240 5.920 316.320 6.240 ; 
                RECT 317.360 5.920 322.440 6.240 ; 
                RECT 323.480 5.920 328.560 6.240 ; 
                RECT 329.600 5.920 334.680 6.240 ; 
                RECT 335.720 5.920 340.800 6.240 ; 
                RECT 341.840 5.920 360.160 6.240 ; 
                RECT 0.160 7.280 360.160 7.600 ; 
                RECT 0.160 8.640 360.160 8.960 ; 
                RECT 0.160 10.000 124.560 10.320 ; 
                RECT 147.360 10.000 360.160 10.320 ; 
                RECT 0.160 11.360 360.160 11.680 ; 
                RECT 0.160 12.720 360.160 13.040 ; 
                RECT 0.160 14.080 75.600 14.400 ; 
                RECT 126.280 14.080 360.160 14.400 ; 
                RECT 0.160 15.440 360.160 15.760 ; 
                RECT 0.160 16.800 360.160 17.120 ; 
                RECT 0.160 18.160 75.600 18.480 ; 
                RECT 125.600 18.160 360.160 18.480 ; 
                RECT 0.160 19.520 360.160 19.840 ; 
                RECT 0.160 20.880 140.880 21.200 ; 
                RECT 350.680 20.880 360.160 21.200 ; 
                RECT 0.160 22.240 140.880 22.560 ; 
                RECT 350.680 22.240 360.160 22.560 ; 
                RECT 0.160 23.600 140.880 23.920 ; 
                RECT 350.680 23.600 360.160 23.920 ; 
                RECT 0.160 24.960 140.880 25.280 ; 
                RECT 350.680 24.960 360.160 25.280 ; 
                RECT 0.160 26.320 140.880 26.640 ; 
                RECT 350.680 26.320 360.160 26.640 ; 
                RECT 0.160 27.680 140.880 28.000 ; 
                RECT 350.680 27.680 360.160 28.000 ; 
                RECT 0.160 29.040 140.880 29.360 ; 
                RECT 350.680 29.040 360.160 29.360 ; 
                RECT 0.160 30.400 140.880 30.720 ; 
                RECT 350.680 30.400 360.160 30.720 ; 
                RECT 0.160 31.760 89.880 32.080 ; 
                RECT 103.160 31.760 140.880 32.080 ; 
                RECT 350.680 31.760 360.160 32.080 ; 
                RECT 0.160 33.120 88.520 33.440 ; 
                RECT 109.280 33.120 140.880 33.440 ; 
                RECT 350.680 33.120 360.160 33.440 ; 
                RECT 0.160 34.480 68.800 34.800 ; 
                RECT 126.280 34.480 140.880 34.800 ; 
                RECT 350.680 34.480 360.160 34.800 ; 
                RECT 0.160 35.840 68.120 36.160 ; 
                RECT 122.200 35.840 140.880 36.160 ; 
                RECT 350.680 35.840 360.160 36.160 ; 
                RECT 0.160 37.200 140.880 37.520 ; 
                RECT 350.680 37.200 360.160 37.520 ; 
                RECT 0.160 38.560 140.200 38.880 ; 
                RECT 350.680 38.560 360.160 38.880 ; 
                RECT 0.160 39.920 140.880 40.240 ; 
                RECT 350.680 39.920 360.160 40.240 ; 
                RECT 0.160 41.280 140.880 41.600 ; 
                RECT 350.680 41.280 360.160 41.600 ; 
                RECT 0.160 42.640 64.040 42.960 ; 
                RECT 75.280 42.640 140.880 42.960 ; 
                RECT 350.680 42.640 360.160 42.960 ; 
                RECT 0.160 44.000 65.400 44.320 ; 
                RECT 71.200 44.000 79.000 44.320 ; 
                RECT 81.400 44.000 140.880 44.320 ; 
                RECT 350.680 44.000 360.160 44.320 ; 
                RECT 0.160 45.360 66.760 45.680 ; 
                RECT 70.520 45.360 140.880 45.680 ; 
                RECT 350.680 45.360 360.160 45.680 ; 
                RECT 0.160 46.720 117.080 47.040 ; 
                RECT 123.560 46.720 140.880 47.040 ; 
                RECT 350.680 46.720 360.160 47.040 ; 
                RECT 0.160 48.080 73.560 48.400 ; 
                RECT 82.080 48.080 117.080 48.400 ; 
                RECT 350.680 48.080 360.160 48.400 ; 
                RECT 0.160 49.440 66.080 49.760 ; 
                RECT 75.280 49.440 117.080 49.760 ; 
                RECT 123.560 49.440 140.880 49.760 ; 
                RECT 350.680 49.440 360.160 49.760 ; 
                RECT 0.160 50.800 69.480 51.120 ; 
                RECT 74.600 50.800 117.080 51.120 ; 
                RECT 123.560 50.800 140.880 51.120 ; 
                RECT 350.680 50.800 360.160 51.120 ; 
                RECT 0.160 52.160 140.880 52.480 ; 
                RECT 350.680 52.160 360.160 52.480 ; 
                RECT 0.160 53.520 65.400 53.840 ; 
                RECT 75.280 53.520 140.880 53.840 ; 
                RECT 350.680 53.520 360.160 53.840 ; 
                RECT 0.160 54.880 72.200 55.200 ; 
                RECT 81.400 54.880 140.880 55.200 ; 
                RECT 350.680 54.880 360.160 55.200 ; 
                RECT 0.160 56.240 99.400 56.560 ; 
                RECT 122.880 56.240 140.880 56.560 ; 
                RECT 350.680 56.240 360.160 56.560 ; 
                RECT 0.160 57.600 73.560 57.920 ; 
                RECT 79.360 57.600 89.200 57.920 ; 
                RECT 93.640 57.600 99.400 57.920 ; 
                RECT 122.880 57.600 140.880 57.920 ; 
                RECT 350.680 57.600 360.160 57.920 ; 
                RECT 0.160 58.960 76.280 59.280 ; 
                RECT 81.400 58.960 90.560 59.280 ; 
                RECT 92.960 58.960 99.400 59.280 ; 
                RECT 133.080 58.960 140.880 59.280 ; 
                RECT 350.680 58.960 360.160 59.280 ; 
                RECT 0.160 60.320 70.160 60.640 ; 
                RECT 75.280 60.320 99.400 60.640 ; 
                RECT 133.080 60.320 140.880 60.640 ; 
                RECT 350.680 60.320 360.160 60.640 ; 
                RECT 0.160 61.680 99.400 62.000 ; 
                RECT 133.080 61.680 140.880 62.000 ; 
                RECT 350.680 61.680 360.160 62.000 ; 
                RECT 0.160 63.040 64.040 63.360 ; 
                RECT 86.840 63.040 99.400 63.360 ; 
                RECT 131.720 63.040 140.880 63.360 ; 
                RECT 350.680 63.040 360.160 63.360 ; 
                RECT 0.160 64.400 73.560 64.720 ; 
                RECT 81.400 64.400 99.400 64.720 ; 
                RECT 133.080 64.400 140.880 64.720 ; 
                RECT 350.680 64.400 360.160 64.720 ; 
                RECT 0.160 65.760 72.200 66.080 ; 
                RECT 75.280 65.760 82.400 66.080 ; 
                RECT 88.880 65.760 99.400 66.080 ; 
                RECT 122.880 65.760 140.880 66.080 ; 
                RECT 350.680 65.760 360.160 66.080 ; 
                RECT 0.160 67.120 64.040 67.440 ; 
                RECT 78.000 67.120 99.400 67.440 ; 
                RECT 135.800 67.120 140.880 67.440 ; 
                RECT 350.680 67.120 360.160 67.440 ; 
                RECT 0.160 68.480 72.200 68.800 ; 
                RECT 81.400 68.480 99.400 68.800 ; 
                RECT 135.800 68.480 140.880 68.800 ; 
                RECT 350.680 68.480 360.160 68.800 ; 
                RECT 0.160 69.840 70.840 70.160 ; 
                RECT 74.600 69.840 99.400 70.160 ; 
                RECT 134.440 69.840 140.880 70.160 ; 
                RECT 350.680 69.840 360.160 70.160 ; 
                RECT 0.160 71.200 66.080 71.520 ; 
                RECT 70.520 71.200 73.560 71.520 ; 
                RECT 82.080 71.200 99.400 71.520 ; 
                RECT 135.800 71.200 140.880 71.520 ; 
                RECT 350.680 71.200 360.160 71.520 ; 
                RECT 0.160 72.560 68.800 72.880 ; 
                RECT 72.560 72.560 99.400 72.880 ; 
                RECT 135.800 72.560 140.880 72.880 ; 
                RECT 350.680 72.560 360.160 72.880 ; 
                RECT 0.160 73.920 65.400 74.240 ; 
                RECT 69.160 73.920 99.400 74.240 ; 
                RECT 134.440 73.920 140.880 74.240 ; 
                RECT 350.680 73.920 360.160 74.240 ; 
                RECT 0.160 75.280 69.480 75.600 ; 
                RECT 75.280 75.280 99.400 75.600 ; 
                RECT 138.520 75.280 140.880 75.600 ; 
                RECT 350.680 75.280 360.160 75.600 ; 
                RECT 0.160 76.640 65.400 76.960 ; 
                RECT 81.400 76.640 99.400 76.960 ; 
                RECT 137.160 76.640 140.880 76.960 ; 
                RECT 350.680 76.640 360.160 76.960 ; 
                RECT 0.160 78.000 73.560 78.320 ; 
                RECT 77.320 78.000 99.400 78.320 ; 
                RECT 138.520 78.000 140.880 78.320 ; 
                RECT 350.680 78.000 360.160 78.320 ; 
                RECT 0.160 79.360 72.880 79.680 ; 
                RECT 75.280 79.360 99.400 79.680 ; 
                RECT 138.520 79.360 140.880 79.680 ; 
                RECT 350.680 79.360 360.160 79.680 ; 
                RECT 0.160 80.720 73.560 81.040 ; 
                RECT 77.320 80.720 99.400 81.040 ; 
                RECT 122.880 80.720 140.880 81.040 ; 
                RECT 350.680 80.720 360.160 81.040 ; 
                RECT 0.160 82.080 64.040 82.400 ; 
                RECT 71.200 82.080 99.400 82.400 ; 
                RECT 137.160 82.080 140.880 82.400 ; 
                RECT 350.680 82.080 360.160 82.400 ; 
                RECT 0.160 83.440 64.040 83.760 ; 
                RECT 75.280 83.440 99.400 83.760 ; 
                RECT 122.880 83.440 140.880 83.760 ; 
                RECT 350.680 83.440 360.160 83.760 ; 
                RECT 0.160 84.800 67.440 85.120 ; 
                RECT 73.920 84.800 99.400 85.120 ; 
                RECT 350.680 84.800 360.160 85.120 ; 
                RECT 0.160 86.160 72.880 86.480 ; 
                RECT 75.280 86.160 99.400 86.480 ; 
                RECT 350.680 86.160 360.160 86.480 ; 
                RECT 0.160 87.520 69.480 87.840 ; 
                RECT 81.400 87.520 99.400 87.840 ; 
                RECT 350.680 87.520 360.160 87.840 ; 
                RECT 0.160 88.880 99.400 89.200 ; 
                RECT 350.680 88.880 360.160 89.200 ; 
                RECT 0.160 90.240 60.640 90.560 ; 
                RECT 78.000 90.240 99.400 90.560 ; 
                RECT 350.680 90.240 360.160 90.560 ; 
                RECT 0.160 91.600 99.400 91.920 ; 
                RECT 122.880 91.600 140.880 91.920 ; 
                RECT 350.680 91.600 360.160 91.920 ; 
                RECT 0.160 92.960 140.880 93.280 ; 
                RECT 350.680 92.960 360.160 93.280 ; 
                RECT 0.160 94.320 140.880 94.640 ; 
                RECT 350.680 94.320 360.160 94.640 ; 
                RECT 0.160 95.680 76.280 96.000 ; 
                RECT 84.120 95.680 140.880 96.000 ; 
                RECT 350.680 95.680 360.160 96.000 ; 
                RECT 0.160 97.040 79.680 97.360 ; 
                RECT 82.080 97.040 140.880 97.360 ; 
                RECT 350.680 97.040 360.160 97.360 ; 
                RECT 0.160 98.400 87.840 98.720 ; 
                RECT 99.760 98.400 102.120 98.720 ; 
                RECT 123.560 98.400 140.880 98.720 ; 
                RECT 350.680 98.400 360.160 98.720 ; 
                RECT 0.160 99.760 64.040 100.080 ; 
                RECT 69.160 99.760 102.120 100.080 ; 
                RECT 123.560 99.760 140.880 100.080 ; 
                RECT 350.680 99.760 360.160 100.080 ; 
                RECT 0.160 101.120 102.120 101.440 ; 
                RECT 123.560 101.120 140.880 101.440 ; 
                RECT 350.680 101.120 360.160 101.440 ; 
                RECT 0.160 102.480 102.120 102.800 ; 
                RECT 123.560 102.480 140.880 102.800 ; 
                RECT 350.680 102.480 360.160 102.800 ; 
                RECT 0.160 103.840 102.120 104.160 ; 
                RECT 123.560 103.840 140.880 104.160 ; 
                RECT 350.680 103.840 360.160 104.160 ; 
                RECT 0.160 105.200 72.200 105.520 ; 
                RECT 81.400 105.200 102.120 105.520 ; 
                RECT 123.560 105.200 140.880 105.520 ; 
                RECT 350.680 105.200 360.160 105.520 ; 
                RECT 0.160 106.560 102.120 106.880 ; 
                RECT 123.560 106.560 140.880 106.880 ; 
                RECT 350.680 106.560 360.160 106.880 ; 
                RECT 0.160 107.920 102.120 108.240 ; 
                RECT 123.560 107.920 140.880 108.240 ; 
                RECT 350.680 107.920 360.160 108.240 ; 
                RECT 0.160 109.280 66.080 109.600 ; 
                RECT 71.200 109.280 102.120 109.600 ; 
                RECT 350.680 109.280 360.160 109.600 ; 
                RECT 0.160 110.640 102.120 110.960 ; 
                RECT 123.560 110.640 138.160 110.960 ; 
                RECT 350.680 110.640 360.160 110.960 ; 
                RECT 0.160 112.000 102.120 112.320 ; 
                RECT 123.560 112.000 135.440 112.320 ; 
                RECT 350.680 112.000 360.160 112.320 ; 
                RECT 0.160 113.360 102.120 113.680 ; 
                RECT 123.560 113.360 132.720 113.680 ; 
                RECT 350.680 113.360 360.160 113.680 ; 
                RECT 0.160 114.720 42.280 115.040 ; 
                RECT 61.000 114.720 68.800 115.040 ; 
                RECT 71.200 114.720 102.120 115.040 ; 
                RECT 123.560 114.720 130.000 115.040 ; 
                RECT 350.680 114.720 360.160 115.040 ; 
                RECT 0.160 116.080 42.280 116.400 ; 
                RECT 61.000 116.080 65.400 116.400 ; 
                RECT 68.480 116.080 102.120 116.400 ; 
                RECT 123.560 116.080 140.880 116.400 ; 
                RECT 350.680 116.080 360.160 116.400 ; 
                RECT 0.160 117.440 42.280 117.760 ; 
                RECT 61.000 117.440 102.120 117.760 ; 
                RECT 123.560 117.440 140.880 117.760 ; 
                RECT 350.680 117.440 360.160 117.760 ; 
                RECT 0.160 118.800 42.280 119.120 ; 
                RECT 61.000 118.800 140.880 119.120 ; 
                RECT 350.680 118.800 360.160 119.120 ; 
                RECT 0.160 120.160 42.280 120.480 ; 
                RECT 61.680 120.160 140.880 120.480 ; 
                RECT 350.680 120.160 360.160 120.480 ; 
                RECT 0.160 121.520 42.280 121.840 ; 
                RECT 61.000 121.520 140.880 121.840 ; 
                RECT 350.680 121.520 360.160 121.840 ; 
                RECT 0.160 122.880 42.280 123.200 ; 
                RECT 61.000 122.880 140.880 123.200 ; 
                RECT 350.680 122.880 360.160 123.200 ; 
                RECT 0.160 124.240 42.280 124.560 ; 
                RECT 61.000 124.240 101.440 124.560 ; 
                RECT 123.560 124.240 131.360 124.560 ; 
                RECT 350.680 124.240 360.160 124.560 ; 
                RECT 0.160 125.600 42.280 125.920 ; 
                RECT 61.000 125.600 67.440 125.920 ; 
                RECT 71.200 125.600 101.440 125.920 ; 
                RECT 123.560 125.600 134.080 125.920 ; 
                RECT 350.680 125.600 360.160 125.920 ; 
                RECT 0.160 126.960 101.440 127.280 ; 
                RECT 123.560 126.960 136.800 127.280 ; 
                RECT 350.680 126.960 360.160 127.280 ; 
                RECT 0.160 128.320 101.440 128.640 ; 
                RECT 123.560 128.320 139.520 128.640 ; 
                RECT 350.680 128.320 360.160 128.640 ; 
                RECT 0.160 129.680 69.480 130.000 ; 
                RECT 75.280 129.680 101.440 130.000 ; 
                RECT 350.680 129.680 360.160 130.000 ; 
                RECT 0.160 131.040 25.960 131.360 ; 
                RECT 42.640 131.040 48.400 131.360 ; 
                RECT 55.560 131.040 101.440 131.360 ; 
                RECT 123.560 131.040 140.880 131.360 ; 
                RECT 350.680 131.040 360.160 131.360 ; 
                RECT 0.160 132.400 25.960 132.720 ; 
                RECT 60.320 132.400 101.440 132.720 ; 
                RECT 123.560 132.400 140.880 132.720 ; 
                RECT 350.680 132.400 360.160 132.720 ; 
                RECT 0.160 133.760 25.960 134.080 ; 
                RECT 60.320 133.760 101.440 134.080 ; 
                RECT 350.680 133.760 360.160 134.080 ; 
                RECT 0.160 135.120 25.960 135.440 ; 
                RECT 42.640 135.120 48.400 135.440 ; 
                RECT 55.560 135.120 64.040 135.440 ; 
                RECT 73.920 135.120 101.440 135.440 ; 
                RECT 123.560 135.120 127.280 135.440 ; 
                RECT 350.680 135.120 360.160 135.440 ; 
                RECT 0.160 136.480 26.640 136.800 ; 
                RECT 54.880 136.480 101.440 136.800 ; 
                RECT 123.560 136.480 360.160 136.800 ; 
                RECT 0.160 137.840 54.520 138.160 ; 
                RECT 98.400 137.840 360.160 138.160 ; 
                RECT 0.160 139.200 138.160 139.520 ; 
                RECT 352.720 139.200 360.160 139.520 ; 
                RECT 0.160 140.560 138.160 140.880 ; 
                RECT 352.720 140.560 360.160 140.880 ; 
                RECT 0.160 141.920 138.160 142.240 ; 
                RECT 352.720 141.920 360.160 142.240 ; 
                RECT 0.160 143.280 23.240 143.600 ; 
                RECT 29.720 143.280 32.080 143.600 ; 
                RECT 40.600 143.280 71.520 143.600 ; 
                RECT 352.720 143.280 360.160 143.600 ; 
                RECT 0.160 144.640 21.200 144.960 ; 
                RECT 31.760 144.640 33.440 144.960 ; 
                RECT 39.920 144.640 51.120 144.960 ; 
                RECT 52.160 144.640 71.520 144.960 ; 
                RECT 352.720 144.640 360.160 144.960 ; 
                RECT 0.160 146.000 21.200 146.320 ; 
                RECT 31.760 146.000 51.120 146.320 ; 
                RECT 54.880 146.000 71.520 146.320 ; 
                RECT 352.720 146.000 360.160 146.320 ; 
                RECT 0.160 147.360 21.200 147.680 ; 
                RECT 31.760 147.360 51.120 147.680 ; 
                RECT 55.560 147.360 71.520 147.680 ; 
                RECT 352.720 147.360 360.160 147.680 ; 
                RECT 0.160 148.720 51.120 149.040 ; 
                RECT 55.560 148.720 71.520 149.040 ; 
                RECT 352.720 148.720 360.160 149.040 ; 
                RECT 0.160 150.080 21.200 150.400 ; 
                RECT 31.760 150.080 51.120 150.400 ; 
                RECT 52.160 150.080 71.520 150.400 ; 
                RECT 352.720 150.080 360.160 150.400 ; 
                RECT 0.160 151.440 21.200 151.760 ; 
                RECT 31.760 151.440 71.520 151.760 ; 
                RECT 352.720 151.440 360.160 151.760 ; 
                RECT 0.160 152.800 71.520 153.120 ; 
                RECT 352.720 152.800 360.160 153.120 ; 
                RECT 0.160 154.160 71.520 154.480 ; 
                RECT 352.720 154.160 360.160 154.480 ; 
                RECT 0.160 155.520 14.400 155.840 ; 
                RECT 16.800 155.520 71.520 155.840 ; 
                RECT 352.720 155.520 360.160 155.840 ; 
                RECT 0.160 156.880 71.520 157.200 ; 
                RECT 352.720 156.880 360.160 157.200 ; 
                RECT 0.160 158.240 13.720 158.560 ; 
                RECT 16.800 158.240 30.040 158.560 ; 
                RECT 33.800 158.240 71.520 158.560 ; 
                RECT 352.720 158.240 360.160 158.560 ; 
                RECT 0.160 159.600 13.040 159.920 ; 
                RECT 16.800 159.600 30.040 159.920 ; 
                RECT 39.920 159.600 71.520 159.920 ; 
                RECT 352.720 159.600 360.160 159.920 ; 
                RECT 0.160 160.960 12.360 161.280 ; 
                RECT 16.800 160.960 30.040 161.280 ; 
                RECT 39.240 160.960 51.120 161.280 ; 
                RECT 52.160 160.960 71.520 161.280 ; 
                RECT 352.720 160.960 360.160 161.280 ; 
                RECT 0.160 162.320 51.120 162.640 ; 
                RECT 52.840 162.320 71.520 162.640 ; 
                RECT 352.720 162.320 360.160 162.640 ; 
                RECT 0.160 163.680 11.680 164.000 ; 
                RECT 16.800 163.680 30.040 164.000 ; 
                RECT 35.840 163.680 51.120 164.000 ; 
                RECT 53.520 163.680 71.520 164.000 ; 
                RECT 352.720 163.680 360.160 164.000 ; 
                RECT 0.160 165.040 11.000 165.360 ; 
                RECT 16.800 165.040 51.120 165.360 ; 
                RECT 54.200 165.040 71.520 165.360 ; 
                RECT 352.720 165.040 360.160 165.360 ; 
                RECT 0.160 166.400 10.320 166.720 ; 
                RECT 16.800 166.400 51.120 166.720 ; 
                RECT 54.200 166.400 71.520 166.720 ; 
                RECT 352.720 166.400 360.160 166.720 ; 
                RECT 0.160 167.760 9.640 168.080 ; 
                RECT 16.800 167.760 71.520 168.080 ; 
                RECT 352.720 167.760 360.160 168.080 ; 
                RECT 0.160 169.120 71.520 169.440 ; 
                RECT 352.720 169.120 360.160 169.440 ; 
                RECT 0.160 170.480 71.520 170.800 ; 
                RECT 352.720 170.480 360.160 170.800 ; 
                RECT 0.160 171.840 71.520 172.160 ; 
                RECT 352.720 171.840 360.160 172.160 ; 
                RECT 0.160 173.200 71.520 173.520 ; 
                RECT 352.720 173.200 360.160 173.520 ; 
                RECT 0.160 174.560 71.520 174.880 ; 
                RECT 352.720 174.560 360.160 174.880 ; 
                RECT 0.160 175.920 71.520 176.240 ; 
                RECT 352.720 175.920 360.160 176.240 ; 
                RECT 0.160 177.280 138.160 177.600 ; 
                RECT 352.720 177.280 360.160 177.600 ; 
                RECT 0.160 178.640 138.160 178.960 ; 
                RECT 352.720 178.640 360.160 178.960 ; 
                RECT 0.160 180.000 138.160 180.320 ; 
                RECT 352.720 180.000 360.160 180.320 ; 
                RECT 0.160 181.360 360.160 181.680 ; 
                RECT 0.160 182.720 360.160 183.040 ; 
                RECT 0.160 184.080 360.160 184.400 ; 
                RECT 0.160 185.440 360.160 185.760 ; 
                RECT 0.160 0.160 360.160 1.520 ; 
                RECT 0.160 189.480 360.160 190.840 ; 
                RECT 142.300 42.275 148.100 43.645 ; 
                RECT 343.000 42.275 348.800 43.645 ; 
                RECT 142.300 47.315 148.100 48.685 ; 
                RECT 343.000 47.315 348.800 48.685 ; 
                RECT 142.300 52.415 148.100 53.835 ; 
                RECT 343.000 52.415 348.800 53.835 ; 
                RECT 142.300 57.585 148.100 59.005 ; 
                RECT 343.000 57.585 348.800 59.005 ; 
                RECT 142.300 91.365 348.800 92.165 ; 
                RECT 142.300 95.445 348.800 95.735 ; 
                RECT 142.300 80.250 348.800 81.050 ; 
                RECT 142.300 77.240 348.800 78.040 ; 
                RECT 142.300 117.700 348.800 118.570 ; 
                RECT 142.300 85.140 348.800 85.940 ; 
                RECT 142.300 65.770 348.800 67.570 ; 
                RECT 142.300 132.025 348.800 132.825 ; 
                RECT 142.300 26.520 348.800 28.320 ; 
                RECT 78.435 142.995 80.355 176.175 ; 
                RECT 82.275 142.995 84.195 176.175 ; 
                RECT 86.115 142.995 88.035 176.175 ; 
                RECT 106.555 142.995 108.475 176.175 ; 
                RECT 110.395 142.995 112.315 176.175 ; 
                RECT 114.235 142.995 116.155 176.175 ; 
                RECT 118.075 142.995 119.995 176.175 ; 
                RECT 121.915 142.995 123.835 176.175 ; 
                RECT 125.755 142.995 127.675 176.175 ; 
                RECT 129.595 142.995 131.515 176.175 ; 
                RECT 133.435 142.995 135.355 176.175 ; 
                RECT 103.580 56.680 105.500 92.080 ; 
                RECT 110.555 56.680 112.475 92.080 ; 
                RECT 120.110 56.680 122.030 92.080 ; 
                RECT 105.495 123.880 107.415 136.360 ; 
                RECT 112.555 123.880 114.305 136.360 ; 
                RECT 120.735 123.880 122.655 136.360 ; 
                RECT 106.570 98.080 108.490 117.880 ; 
                RECT 113.845 98.080 115.595 117.880 ; 
                RECT 121.165 98.080 123.085 117.880 ; 
                RECT 121.185 47.100 123.105 50.680 ; 
                RECT 21.950 145.265 31.110 146.015 ; 
                RECT 21.950 149.890 31.110 151.640 ; 
                RECT 43.680 133.050 59.720 133.850 ; 
                RECT 26.880 133.760 41.720 135.450 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 151.080 5.560 ; 
                RECT 152.800 5.240 157.200 5.560 ; 
                RECT 158.920 5.240 163.320 5.560 ; 
                RECT 165.040 5.240 169.440 5.560 ; 
                RECT 171.160 5.240 175.560 5.560 ; 
                RECT 177.280 5.240 181.680 5.560 ; 
                RECT 183.400 5.240 187.800 5.560 ; 
                RECT 189.520 5.240 193.920 5.560 ; 
                RECT 195.640 5.240 200.040 5.560 ; 
                RECT 201.760 5.240 206.160 5.560 ; 
                RECT 207.880 5.240 212.280 5.560 ; 
                RECT 214.000 5.240 218.400 5.560 ; 
                RECT 220.120 5.240 224.520 5.560 ; 
                RECT 226.240 5.240 230.640 5.560 ; 
                RECT 232.360 5.240 236.760 5.560 ; 
                RECT 238.480 5.240 242.880 5.560 ; 
                RECT 244.600 5.240 249.000 5.560 ; 
                RECT 250.720 5.240 255.120 5.560 ; 
                RECT 256.840 5.240 261.240 5.560 ; 
                RECT 262.960 5.240 267.360 5.560 ; 
                RECT 269.080 5.240 273.480 5.560 ; 
                RECT 275.200 5.240 279.600 5.560 ; 
                RECT 281.320 5.240 285.720 5.560 ; 
                RECT 287.440 5.240 291.840 5.560 ; 
                RECT 292.880 5.240 297.960 5.560 ; 
                RECT 299.000 5.240 304.080 5.560 ; 
                RECT 305.120 5.240 310.200 5.560 ; 
                RECT 311.240 5.240 316.320 5.560 ; 
                RECT 317.360 5.240 322.440 5.560 ; 
                RECT 323.480 5.240 328.560 5.560 ; 
                RECT 329.600 5.240 334.680 5.560 ; 
                RECT 335.720 5.240 340.800 5.560 ; 
                RECT 341.840 5.240 357.440 5.560 ; 
                RECT 2.880 6.600 357.440 6.920 ; 
                RECT 2.880 7.960 357.440 8.280 ; 
                RECT 2.880 9.320 125.240 9.640 ; 
                RECT 146.680 9.320 357.440 9.640 ; 
                RECT 2.880 10.680 357.440 11.000 ; 
                RECT 2.880 12.040 357.440 12.360 ; 
                RECT 2.880 13.400 75.600 13.720 ; 
                RECT 126.280 13.400 357.440 13.720 ; 
                RECT 2.880 14.760 357.440 15.080 ; 
                RECT 2.880 16.120 357.440 16.440 ; 
                RECT 2.880 17.480 75.600 17.800 ; 
                RECT 125.600 17.480 357.440 17.800 ; 
                RECT 2.880 18.840 357.440 19.160 ; 
                RECT 2.880 20.200 140.880 20.520 ; 
                RECT 350.680 20.200 357.440 20.520 ; 
                RECT 2.880 21.560 140.880 21.880 ; 
                RECT 350.680 21.560 357.440 21.880 ; 
                RECT 2.880 22.920 140.880 23.240 ; 
                RECT 350.680 22.920 357.440 23.240 ; 
                RECT 2.880 24.280 140.880 24.600 ; 
                RECT 350.680 24.280 357.440 24.600 ; 
                RECT 2.880 25.640 140.880 25.960 ; 
                RECT 350.680 25.640 357.440 25.960 ; 
                RECT 2.880 27.000 140.880 27.320 ; 
                RECT 350.680 27.000 357.440 27.320 ; 
                RECT 2.880 28.360 140.880 28.680 ; 
                RECT 350.680 28.360 357.440 28.680 ; 
                RECT 2.880 29.720 140.880 30.040 ; 
                RECT 350.680 29.720 357.440 30.040 ; 
                RECT 2.880 31.080 90.560 31.400 ; 
                RECT 104.520 31.080 140.880 31.400 ; 
                RECT 350.680 31.080 357.440 31.400 ; 
                RECT 2.880 32.440 89.200 32.760 ; 
                RECT 110.640 32.440 140.880 32.760 ; 
                RECT 350.680 32.440 357.440 32.760 ; 
                RECT 2.880 33.800 66.080 34.120 ; 
                RECT 125.600 33.800 140.880 34.120 ; 
                RECT 350.680 33.800 357.440 34.120 ; 
                RECT 2.880 35.160 66.760 35.480 ; 
                RECT 116.080 35.160 140.880 35.480 ; 
                RECT 350.680 35.160 357.440 35.480 ; 
                RECT 2.880 36.520 140.880 36.840 ; 
                RECT 350.680 36.520 357.440 36.840 ; 
                RECT 2.880 37.880 140.200 38.200 ; 
                RECT 350.680 37.880 357.440 38.200 ; 
                RECT 2.880 39.240 140.880 39.560 ; 
                RECT 350.680 39.240 357.440 39.560 ; 
                RECT 2.880 40.600 140.880 40.920 ; 
                RECT 350.680 40.600 357.440 40.920 ; 
                RECT 2.880 41.960 64.040 42.280 ; 
                RECT 75.280 41.960 140.880 42.280 ; 
                RECT 350.680 41.960 357.440 42.280 ; 
                RECT 2.880 43.320 65.400 43.640 ; 
                RECT 67.800 43.320 140.880 43.640 ; 
                RECT 350.680 43.320 357.440 43.640 ; 
                RECT 2.880 44.680 66.760 45.000 ; 
                RECT 71.200 44.680 79.000 45.000 ; 
                RECT 81.400 44.680 140.880 45.000 ; 
                RECT 350.680 44.680 357.440 45.000 ; 
                RECT 2.880 46.040 66.760 46.360 ; 
                RECT 70.520 46.040 140.880 46.360 ; 
                RECT 350.680 46.040 357.440 46.360 ; 
                RECT 2.880 47.400 73.560 47.720 ; 
                RECT 82.080 47.400 117.080 47.720 ; 
                RECT 123.560 47.400 140.880 47.720 ; 
                RECT 350.680 47.400 357.440 47.720 ; 
                RECT 2.880 48.760 68.800 49.080 ; 
                RECT 75.280 48.760 117.080 49.080 ; 
                RECT 350.680 48.760 357.440 49.080 ; 
                RECT 2.880 50.120 66.080 50.440 ; 
                RECT 75.280 50.120 87.160 50.440 ; 
                RECT 114.040 50.120 117.080 50.440 ; 
                RECT 123.560 50.120 140.880 50.440 ; 
                RECT 350.680 50.120 357.440 50.440 ; 
                RECT 2.880 51.480 140.880 51.800 ; 
                RECT 350.680 51.480 357.440 51.800 ; 
                RECT 2.880 52.840 65.400 53.160 ; 
                RECT 75.280 52.840 140.880 53.160 ; 
                RECT 350.680 52.840 357.440 53.160 ; 
                RECT 2.880 54.200 73.560 54.520 ; 
                RECT 81.400 54.200 140.880 54.520 ; 
                RECT 350.680 54.200 357.440 54.520 ; 
                RECT 2.880 55.560 72.200 55.880 ; 
                RECT 75.280 55.560 140.880 55.880 ; 
                RECT 350.680 55.560 357.440 55.880 ; 
                RECT 2.880 56.920 88.520 57.240 ; 
                RECT 94.320 56.920 99.400 57.240 ; 
                RECT 122.880 56.920 140.880 57.240 ; 
                RECT 350.680 56.920 357.440 57.240 ; 
                RECT 2.880 58.280 73.560 58.600 ; 
                RECT 81.400 58.280 89.880 58.600 ; 
                RECT 92.960 58.280 99.400 58.600 ; 
                RECT 133.080 58.280 140.880 58.600 ; 
                RECT 350.680 58.280 357.440 58.600 ; 
                RECT 2.880 59.640 70.160 59.960 ; 
                RECT 75.280 59.640 99.400 59.960 ; 
                RECT 131.720 59.640 140.880 59.960 ; 
                RECT 350.680 59.640 357.440 59.960 ; 
                RECT 2.880 61.000 72.200 61.320 ; 
                RECT 75.280 61.000 99.400 61.320 ; 
                RECT 133.080 61.000 140.880 61.320 ; 
                RECT 350.680 61.000 357.440 61.320 ; 
                RECT 2.880 62.360 99.400 62.680 ; 
                RECT 133.080 62.360 140.880 62.680 ; 
                RECT 350.680 62.360 357.440 62.680 ; 
                RECT 2.880 63.720 64.040 64.040 ; 
                RECT 86.840 63.720 99.400 64.040 ; 
                RECT 133.080 63.720 140.880 64.040 ; 
                RECT 350.680 63.720 357.440 64.040 ; 
                RECT 2.880 65.080 82.400 65.400 ; 
                RECT 88.200 65.080 99.400 65.400 ; 
                RECT 131.720 65.080 140.880 65.400 ; 
                RECT 350.680 65.080 357.440 65.400 ; 
                RECT 2.880 66.440 72.200 66.760 ; 
                RECT 75.280 66.440 85.120 66.760 ; 
                RECT 88.880 66.440 99.400 66.760 ; 
                RECT 122.880 66.440 140.880 66.760 ; 
                RECT 350.680 66.440 357.440 66.760 ; 
                RECT 2.880 67.800 64.040 68.120 ; 
                RECT 78.000 67.800 99.400 68.120 ; 
                RECT 134.440 67.800 140.880 68.120 ; 
                RECT 350.680 67.800 357.440 68.120 ; 
                RECT 2.880 69.160 72.200 69.480 ; 
                RECT 81.400 69.160 99.400 69.480 ; 
                RECT 135.800 69.160 140.880 69.480 ; 
                RECT 350.680 69.160 357.440 69.480 ; 
                RECT 2.880 70.520 70.840 70.840 ; 
                RECT 82.080 70.520 99.400 70.840 ; 
                RECT 135.800 70.520 140.880 70.840 ; 
                RECT 350.680 70.520 357.440 70.840 ; 
                RECT 2.880 71.880 66.080 72.200 ; 
                RECT 72.560 71.880 99.400 72.200 ; 
                RECT 134.440 71.880 140.880 72.200 ; 
                RECT 350.680 71.880 357.440 72.200 ; 
                RECT 2.880 73.240 99.400 73.560 ; 
                RECT 135.800 73.240 140.880 73.560 ; 
                RECT 350.680 73.240 357.440 73.560 ; 
                RECT 2.880 74.600 65.400 74.920 ; 
                RECT 69.160 74.600 99.400 74.920 ; 
                RECT 122.880 74.600 140.880 74.920 ; 
                RECT 350.680 74.600 357.440 74.920 ; 
                RECT 2.880 75.960 65.400 76.280 ; 
                RECT 75.280 75.960 99.400 76.280 ; 
                RECT 138.520 75.960 140.880 76.280 ; 
                RECT 350.680 75.960 357.440 76.280 ; 
                RECT 2.880 77.320 69.480 77.640 ; 
                RECT 81.400 77.320 99.400 77.640 ; 
                RECT 138.520 77.320 140.880 77.640 ; 
                RECT 350.680 77.320 357.440 77.640 ; 
                RECT 2.880 78.680 72.880 79.000 ; 
                RECT 77.320 78.680 99.400 79.000 ; 
                RECT 137.160 78.680 140.880 79.000 ; 
                RECT 350.680 78.680 357.440 79.000 ; 
                RECT 2.880 80.040 73.560 80.360 ; 
                RECT 77.320 80.040 99.400 80.360 ; 
                RECT 138.520 80.040 140.880 80.360 ; 
                RECT 350.680 80.040 357.440 80.360 ; 
                RECT 2.880 81.400 99.400 81.720 ; 
                RECT 138.520 81.400 140.880 81.720 ; 
                RECT 350.680 81.400 357.440 81.720 ; 
                RECT 2.880 82.760 64.040 83.080 ; 
                RECT 71.200 82.760 99.400 83.080 ; 
                RECT 122.880 82.760 140.880 83.080 ; 
                RECT 350.680 82.760 357.440 83.080 ; 
                RECT 2.880 84.120 64.040 84.440 ; 
                RECT 75.280 84.120 99.400 84.440 ; 
                RECT 350.680 84.120 357.440 84.440 ; 
                RECT 2.880 85.480 72.880 85.800 ; 
                RECT 75.280 85.480 99.400 85.800 ; 
                RECT 122.880 85.480 140.880 85.800 ; 
                RECT 350.680 85.480 357.440 85.800 ; 
                RECT 2.880 86.840 99.400 87.160 ; 
                RECT 350.680 86.840 357.440 87.160 ; 
                RECT 2.880 88.200 69.480 88.520 ; 
                RECT 81.400 88.200 99.400 88.520 ; 
                RECT 350.680 88.200 357.440 88.520 ; 
                RECT 2.880 89.560 60.640 89.880 ; 
                RECT 73.920 89.560 99.400 89.880 ; 
                RECT 350.680 89.560 357.440 89.880 ; 
                RECT 2.880 90.920 70.840 91.240 ; 
                RECT 78.000 90.920 99.400 91.240 ; 
                RECT 350.680 90.920 357.440 91.240 ; 
                RECT 2.880 92.280 99.400 92.600 ; 
                RECT 122.880 92.280 140.880 92.600 ; 
                RECT 350.680 92.280 357.440 92.600 ; 
                RECT 2.880 93.640 140.880 93.960 ; 
                RECT 350.680 93.640 357.440 93.960 ; 
                RECT 2.880 95.000 76.280 95.320 ; 
                RECT 84.120 95.000 140.880 95.320 ; 
                RECT 350.680 95.000 357.440 95.320 ; 
                RECT 2.880 96.360 140.880 96.680 ; 
                RECT 350.680 96.360 357.440 96.680 ; 
                RECT 2.880 97.720 79.680 98.040 ; 
                RECT 82.080 97.720 102.120 98.040 ; 
                RECT 123.560 97.720 140.880 98.040 ; 
                RECT 350.680 97.720 357.440 98.040 ; 
                RECT 2.880 99.080 66.080 99.400 ; 
                RECT 69.160 99.080 102.120 99.400 ; 
                RECT 123.560 99.080 140.880 99.400 ; 
                RECT 350.680 99.080 357.440 99.400 ; 
                RECT 2.880 100.440 64.040 100.760 ; 
                RECT 67.800 100.440 102.120 100.760 ; 
                RECT 123.560 100.440 140.880 100.760 ; 
                RECT 350.680 100.440 357.440 100.760 ; 
                RECT 2.880 101.800 102.120 102.120 ; 
                RECT 123.560 101.800 140.880 102.120 ; 
                RECT 350.680 101.800 357.440 102.120 ; 
                RECT 2.880 103.160 102.120 103.480 ; 
                RECT 123.560 103.160 140.880 103.480 ; 
                RECT 350.680 103.160 357.440 103.480 ; 
                RECT 2.880 104.520 102.120 104.840 ; 
                RECT 123.560 104.520 140.880 104.840 ; 
                RECT 350.680 104.520 357.440 104.840 ; 
                RECT 2.880 105.880 72.200 106.200 ; 
                RECT 81.400 105.880 102.120 106.200 ; 
                RECT 123.560 105.880 140.880 106.200 ; 
                RECT 350.680 105.880 357.440 106.200 ; 
                RECT 2.880 107.240 102.120 107.560 ; 
                RECT 123.560 107.240 140.880 107.560 ; 
                RECT 350.680 107.240 357.440 107.560 ; 
                RECT 2.880 108.600 66.080 108.920 ; 
                RECT 71.200 108.600 102.120 108.920 ; 
                RECT 123.560 108.600 140.880 108.920 ; 
                RECT 350.680 108.600 357.440 108.920 ; 
                RECT 2.880 109.960 102.120 110.280 ; 
                RECT 350.680 109.960 357.440 110.280 ; 
                RECT 2.880 111.320 102.120 111.640 ; 
                RECT 123.560 111.320 138.160 111.640 ; 
                RECT 350.680 111.320 357.440 111.640 ; 
                RECT 2.880 112.680 102.120 113.000 ; 
                RECT 123.560 112.680 135.440 113.000 ; 
                RECT 350.680 112.680 357.440 113.000 ; 
                RECT 2.880 114.040 68.800 114.360 ; 
                RECT 71.200 114.040 102.120 114.360 ; 
                RECT 123.560 114.040 130.000 114.360 ; 
                RECT 350.680 114.040 357.440 114.360 ; 
                RECT 2.880 115.400 42.280 115.720 ; 
                RECT 61.000 115.400 65.400 115.720 ; 
                RECT 68.480 115.400 102.120 115.720 ; 
                RECT 123.560 115.400 130.000 115.720 ; 
                RECT 350.680 115.400 357.440 115.720 ; 
                RECT 2.880 116.760 42.280 117.080 ; 
                RECT 61.000 116.760 102.120 117.080 ; 
                RECT 123.560 116.760 140.880 117.080 ; 
                RECT 350.680 116.760 357.440 117.080 ; 
                RECT 2.880 118.120 42.280 118.440 ; 
                RECT 61.000 118.120 102.120 118.440 ; 
                RECT 123.560 118.120 140.880 118.440 ; 
                RECT 350.680 118.120 357.440 118.440 ; 
                RECT 2.880 119.480 42.280 119.800 ; 
                RECT 61.680 119.480 140.880 119.800 ; 
                RECT 350.680 119.480 357.440 119.800 ; 
                RECT 2.880 120.840 42.280 121.160 ; 
                RECT 61.000 120.840 140.880 121.160 ; 
                RECT 350.680 120.840 357.440 121.160 ; 
                RECT 2.880 122.200 42.280 122.520 ; 
                RECT 61.000 122.200 140.880 122.520 ; 
                RECT 350.680 122.200 357.440 122.520 ; 
                RECT 2.880 123.560 42.280 123.880 ; 
                RECT 61.000 123.560 101.440 123.880 ; 
                RECT 123.560 123.560 131.360 123.880 ; 
                RECT 350.680 123.560 357.440 123.880 ; 
                RECT 2.880 124.920 42.280 125.240 ; 
                RECT 61.000 124.920 67.440 125.240 ; 
                RECT 71.200 124.920 101.440 125.240 ; 
                RECT 123.560 124.920 131.360 125.240 ; 
                RECT 350.680 124.920 357.440 125.240 ; 
                RECT 2.880 126.280 42.280 126.600 ; 
                RECT 61.000 126.280 101.440 126.600 ; 
                RECT 123.560 126.280 134.080 126.600 ; 
                RECT 350.680 126.280 357.440 126.600 ; 
                RECT 2.880 127.640 101.440 127.960 ; 
                RECT 123.560 127.640 136.800 127.960 ; 
                RECT 350.680 127.640 357.440 127.960 ; 
                RECT 2.880 129.000 101.440 129.320 ; 
                RECT 350.680 129.000 357.440 129.320 ; 
                RECT 2.880 130.360 25.960 130.680 ; 
                RECT 42.640 130.360 69.480 130.680 ; 
                RECT 75.280 130.360 101.440 130.680 ; 
                RECT 350.680 130.360 357.440 130.680 ; 
                RECT 2.880 131.720 25.960 132.040 ; 
                RECT 42.640 131.720 48.400 132.040 ; 
                RECT 55.560 131.720 101.440 132.040 ; 
                RECT 123.560 131.720 140.880 132.040 ; 
                RECT 350.680 131.720 357.440 132.040 ; 
                RECT 2.880 133.080 25.960 133.400 ; 
                RECT 60.320 133.080 101.440 133.400 ; 
                RECT 123.560 133.080 140.880 133.400 ; 
                RECT 350.680 133.080 357.440 133.400 ; 
                RECT 2.880 134.440 25.960 134.760 ; 
                RECT 42.640 134.440 101.440 134.760 ; 
                RECT 350.680 134.440 357.440 134.760 ; 
                RECT 2.880 135.800 25.960 136.120 ; 
                RECT 55.560 135.800 64.040 136.120 ; 
                RECT 73.920 135.800 101.440 136.120 ; 
                RECT 123.560 135.800 140.880 136.120 ; 
                RECT 350.680 135.800 357.440 136.120 ; 
                RECT 2.880 137.160 48.400 137.480 ; 
                RECT 68.480 137.160 357.440 137.480 ; 
                RECT 2.880 138.520 28.000 138.840 ; 
                RECT 67.800 138.520 357.440 138.840 ; 
                RECT 2.880 139.880 138.160 140.200 ; 
                RECT 352.720 139.880 357.440 140.200 ; 
                RECT 2.880 141.240 138.160 141.560 ; 
                RECT 352.720 141.240 357.440 141.560 ; 
                RECT 2.880 142.600 23.240 142.920 ; 
                RECT 29.720 142.600 71.520 142.920 ; 
                RECT 352.720 142.600 357.440 142.920 ; 
                RECT 2.880 143.960 21.200 144.280 ; 
                RECT 39.920 143.960 71.520 144.280 ; 
                RECT 352.720 143.960 357.440 144.280 ; 
                RECT 2.880 145.320 21.200 145.640 ; 
                RECT 39.240 145.320 51.120 145.640 ; 
                RECT 52.160 145.320 71.520 145.640 ; 
                RECT 352.720 145.320 357.440 145.640 ; 
                RECT 2.880 146.680 51.120 147.000 ; 
                RECT 52.160 146.680 71.520 147.000 ; 
                RECT 352.720 146.680 357.440 147.000 ; 
                RECT 2.880 148.040 21.200 148.360 ; 
                RECT 31.760 148.040 51.120 148.360 ; 
                RECT 55.560 148.040 71.520 148.360 ; 
                RECT 352.720 148.040 357.440 148.360 ; 
                RECT 2.880 149.400 21.200 149.720 ; 
                RECT 31.760 149.400 51.120 149.720 ; 
                RECT 55.560 149.400 71.520 149.720 ; 
                RECT 352.720 149.400 357.440 149.720 ; 
                RECT 2.880 150.760 21.200 151.080 ; 
                RECT 31.760 150.760 51.120 151.080 ; 
                RECT 56.240 150.760 71.520 151.080 ; 
                RECT 352.720 150.760 357.440 151.080 ; 
                RECT 2.880 152.120 71.520 152.440 ; 
                RECT 352.720 152.120 357.440 152.440 ; 
                RECT 2.880 153.480 71.520 153.800 ; 
                RECT 352.720 153.480 357.440 153.800 ; 
                RECT 2.880 154.840 71.520 155.160 ; 
                RECT 352.720 154.840 357.440 155.160 ; 
                RECT 2.880 156.200 14.400 156.520 ; 
                RECT 16.800 156.200 30.040 156.520 ; 
                RECT 33.120 156.200 71.520 156.520 ; 
                RECT 352.720 156.200 357.440 156.520 ; 
                RECT 2.880 157.560 13.720 157.880 ; 
                RECT 16.800 157.560 71.520 157.880 ; 
                RECT 352.720 157.560 357.440 157.880 ; 
                RECT 2.880 158.920 13.040 159.240 ; 
                RECT 16.800 158.920 34.800 159.240 ; 
                RECT 40.600 158.920 71.520 159.240 ; 
                RECT 352.720 158.920 357.440 159.240 ; 
                RECT 2.880 160.280 12.360 160.600 ; 
                RECT 16.800 160.280 36.160 160.600 ; 
                RECT 39.920 160.280 71.520 160.600 ; 
                RECT 352.720 160.280 357.440 160.600 ; 
                RECT 2.880 161.640 51.120 161.960 ; 
                RECT 52.840 161.640 71.520 161.960 ; 
                RECT 352.720 161.640 357.440 161.960 ; 
                RECT 2.880 163.000 11.680 163.320 ; 
                RECT 16.800 163.000 51.120 163.320 ; 
                RECT 53.520 163.000 71.520 163.320 ; 
                RECT 352.720 163.000 357.440 163.320 ; 
                RECT 2.880 164.360 51.120 164.680 ; 
                RECT 54.200 164.360 71.520 164.680 ; 
                RECT 352.720 164.360 357.440 164.680 ; 
                RECT 2.880 165.720 11.000 166.040 ; 
                RECT 16.800 165.720 30.040 166.040 ; 
                RECT 36.520 165.720 51.120 166.040 ; 
                RECT 52.160 165.720 71.520 166.040 ; 
                RECT 352.720 165.720 357.440 166.040 ; 
                RECT 2.880 167.080 10.320 167.400 ; 
                RECT 16.800 167.080 30.040 167.400 ; 
                RECT 37.200 167.080 51.120 167.400 ; 
                RECT 54.200 167.080 71.520 167.400 ; 
                RECT 352.720 167.080 357.440 167.400 ; 
                RECT 2.880 168.440 9.640 168.760 ; 
                RECT 16.800 168.440 30.040 168.760 ; 
                RECT 37.880 168.440 71.520 168.760 ; 
                RECT 352.720 168.440 357.440 168.760 ; 
                RECT 2.880 169.800 71.520 170.120 ; 
                RECT 352.720 169.800 357.440 170.120 ; 
                RECT 2.880 171.160 71.520 171.480 ; 
                RECT 352.720 171.160 357.440 171.480 ; 
                RECT 2.880 172.520 71.520 172.840 ; 
                RECT 352.720 172.520 357.440 172.840 ; 
                RECT 2.880 173.880 71.520 174.200 ; 
                RECT 352.720 173.880 357.440 174.200 ; 
                RECT 2.880 175.240 71.520 175.560 ; 
                RECT 352.720 175.240 357.440 175.560 ; 
                RECT 2.880 176.600 138.160 176.920 ; 
                RECT 352.720 176.600 357.440 176.920 ; 
                RECT 2.880 177.960 138.160 178.280 ; 
                RECT 352.720 177.960 357.440 178.280 ; 
                RECT 2.880 179.320 138.160 179.640 ; 
                RECT 352.720 179.320 357.440 179.640 ; 
                RECT 2.880 180.680 357.440 181.000 ; 
                RECT 2.880 182.040 357.440 182.360 ; 
                RECT 2.880 183.400 357.440 183.720 ; 
                RECT 2.880 184.760 357.440 185.080 ; 
                RECT 2.880 2.880 357.440 4.240 ; 
                RECT 2.880 186.760 357.440 188.120 ; 
                RECT 142.300 39.630 148.100 40.750 ; 
                RECT 343.000 39.630 348.800 40.750 ; 
                RECT 142.300 45.420 148.100 46.040 ; 
                RECT 343.000 45.420 348.800 46.040 ; 
                RECT 142.300 50.470 148.100 51.110 ; 
                RECT 343.000 50.470 348.800 51.110 ; 
                RECT 142.300 55.640 148.100 56.280 ; 
                RECT 343.000 55.640 348.800 56.280 ; 
                RECT 142.300 89.645 348.800 90.445 ; 
                RECT 142.300 81.570 348.800 82.370 ; 
                RECT 142.300 69.510 348.800 71.310 ; 
                RECT 142.300 86.460 348.800 87.260 ; 
                RECT 142.300 83.250 348.800 84.050 ; 
                RECT 142.300 78.560 348.800 79.360 ; 
                RECT 142.300 121.980 348.800 122.225 ; 
                RECT 142.300 108.005 348.800 108.295 ; 
                RECT 142.300 30.260 348.800 32.060 ; 
                RECT 72.470 142.995 74.390 176.175 ; 
                RECT 92.590 142.995 94.510 176.175 ; 
                RECT 96.430 142.995 98.350 176.175 ; 
                RECT 100.270 142.995 102.190 176.175 ; 
                RECT 100.415 56.680 101.525 92.080 ; 
                RECT 107.930 56.680 108.820 92.080 ; 
                RECT 115.010 56.680 116.550 92.080 ; 
                RECT 102.115 123.880 103.225 136.360 ; 
                RECT 110.060 123.880 110.950 136.360 ; 
                RECT 116.605 123.880 117.925 136.360 ; 
                RECT 102.975 98.080 104.085 117.880 ; 
                RECT 111.350 98.080 112.240 117.880 ; 
                RECT 117.785 98.080 118.895 117.880 ; 
                RECT 117.805 47.100 118.915 50.680 ; 
                RECT 21.950 144.060 31.110 144.430 ; 
                RECT 21.950 147.395 31.110 148.285 ; 
                RECT 26.880 130.420 41.720 131.090 ; 
                RECT 26.880 131.720 41.720 132.730 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 360.320 191.000 ; 
        LAYER met2 ;
            RECT 0.000 0.000 360.320 191.000 ; 
    END 
END sram22_64x32m4w8 
END LIBRARY 

