VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sramgen_sram_64x32m4w32_replica_v1
  CLASS BLOCK ;
  ORIGIN 72.135 136.07 ;
  FOREIGN sramgen_sram_64x32m4w32_replica_v1 -72.135 -136.07 ;
  SIZE 414.595 BY 147.785 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -65.8 -135.67 -65.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -135.67 -63.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.6 -135.67 -62.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -61 -135.67 -60.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -135.67 -59 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.8 -135.67 -57.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -135.67 -55.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.6 -135.67 -54.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -135.67 -52.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.4 -135.67 -51 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -135.67 -49.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.2 -135.67 -47.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -101.02 -46.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -112.68 -44.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -135.67 -44.6 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.4 -135.67 -43 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -108.44 -41.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -135.67 -41.4 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.2 -113.74 -39.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -112.68 -38.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -135.67 -38.2 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -37 -135.67 -36.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -107.38 -35 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -135.67 -35 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.8 -113.74 -33.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.2 -135.67 -31.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -106.32 -30.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -135.67 -30.2 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -106.32 -28.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -135.67 -28.6 -115.22 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -112.68 -27 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -135.67 -27 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.8 -135.67 -25.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -105.26 -23.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -135.67 -23.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.6 -113.74 -22.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -112.68 -20.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -135.67 -20.6 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.4 -135.67 -19 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -104.2 -17.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -135.67 -17.4 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.2 -113.74 -15.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.6 -135.67 -14.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -103.14 -12.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -135.67 -12.6 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -104.2 -11 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -135.67 -11 -115.22 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -35.3 -9.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -112.68 -9.4 -82.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -135.67 -9.4 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.2 -135.67 -7.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -98.9 -6.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -135.67 -6.2 -115.22 ;
    END
    PORT
      LAYER met3 ;
        RECT -5 -135.67 -4.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.4 -135.67 -3 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 2.86 -1.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 -135.67 -1.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 2.86 0.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 -135.67 0.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 2.86 1.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 -135.67 1.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 2.86 3.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 -135.67 3.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 2.86 5 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 -135.67 5 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 2.86 6.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -73.46 6.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -135.67 6.6 -80.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 2.86 8.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -44.84 8.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -109.5 8.2 -100.38 ;
        RECT 7.84 -109.535 8.17 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 2.86 9.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -53.32 9.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -135.67 9.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 2.86 11.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -135.67 11.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 2.86 13 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -114.8 13 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 2.86 14.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -135.67 14.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 2.86 16.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 -135.67 16.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 2.86 17.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 -135.67 17.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 2.86 19.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -53.32 19.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -135.67 19.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 2.86 21 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -44.84 21 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -135.67 21 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 2.86 22.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 -135.67 22.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 2.86 24.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 -135.67 24.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 2.86 25.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 -135.67 25.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 2.86 27.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 -135.67 27.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 2.86 29 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -44.84 29 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -109.5 29 -100.38 ;
        RECT 28.635 -109.535 28.965 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 2.86 30.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -44.84 30.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -135.67 30.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 2.86 32.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 -115.86 32.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 2.86 33.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -114.8 33.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -135.67 33.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 2.86 35.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -135.67 35.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 2.86 37 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -135.67 37 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 2.86 38.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -44.84 38.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -109.5 38.6 -100.38 ;
        RECT 38.235 -109.535 38.565 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 2.86 40.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -44.84 40.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -135.67 40.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 2.86 41.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 -135.67 41.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 2.86 43.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 -135.67 43.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 2.86 45 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 -135.67 45 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 2.86 46.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 -135.67 46.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 2.86 48.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -44.84 48.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -109.5 48.2 -100.38 ;
        RECT 47.835 -109.535 48.165 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 2.86 49.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -53.32 49.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -135.67 49.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 2.86 51.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 -135.67 51.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 2.86 53 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -114.8 53 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 2.86 54.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -135.67 54.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 2.86 56.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 -135.67 56.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 2.86 57.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 -135.67 57.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 2.86 59.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -53.32 59.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -135.67 59.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 2.86 61 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -44.84 61 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -135.67 61 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 2.86 62.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 -135.67 62.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 2.86 64.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -135.67 64.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 2.86 65.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 -135.67 65.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 2.86 67.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 -135.67 67.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 2.86 69 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -44.84 69 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -109.5 69 -100.38 ;
        RECT 68.635 -109.535 68.965 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 2.86 70.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -44.84 70.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -135.67 70.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 2.86 72.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 -115.86 72.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 2.86 73.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -114.8 73.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -135.67 73.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 2.86 75.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -135.67 75.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 2.86 77 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 -135.67 77 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 2.86 78.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -44.84 78.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -109.5 78.6 -100.38 ;
        RECT 78.235 -109.535 78.565 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 2.86 80.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -44.84 80.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -135.67 80.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 2.86 81.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 -135.67 81.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 2.86 83.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 -135.67 83.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 2.86 85 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 -135.67 85 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 2.86 86.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 -135.67 86.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 2.86 88.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -44.84 88.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -109.5 88.2 -100.38 ;
        RECT 87.835 -109.535 88.165 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 2.86 89.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -53.32 89.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -135.67 89.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 2.86 91.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 -135.67 91.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 2.86 93 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -114.8 93 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 2.86 94.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -135.67 94.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 2.86 96.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 -135.67 96.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 2.86 97.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 -135.67 97.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 2.86 99.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -53.32 99.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -135.67 99.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 2.86 101 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -44.84 101 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -135.67 101 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 2.86 102.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 -135.67 102.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 2.86 104.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -135.67 104.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 2.86 105.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 -135.67 105.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 2.86 107.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 -135.67 107.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 2.86 109 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -44.84 109 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -109.5 109 -100.38 ;
        RECT 108.635 -109.535 108.965 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 2.86 110.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -44.84 110.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -135.67 110.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 2.86 112.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 -115.86 112.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 2.86 113.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -114.8 113.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -135.67 113.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 2.86 115.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -135.67 115.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 2.86 117 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 -135.67 117 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 2.86 118.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -44.84 118.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -109.5 118.6 -100.38 ;
        RECT 118.235 -109.535 118.565 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 2.86 120.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -44.84 120.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -135.67 120.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 2.86 121.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 -135.67 121.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 2.86 123.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 -135.67 123.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 2.86 125 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 -135.67 125 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 2.86 126.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 -135.67 126.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 2.86 128.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -44.84 128.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -109.5 128.2 -100.38 ;
        RECT 127.835 -109.535 128.165 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 2.86 129.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -53.32 129.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -135.67 129.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 2.86 131.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 -135.67 131.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 2.86 133 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -114.8 133 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 2.86 134.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -135.67 134.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 2.86 136.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 -135.67 136.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 2.86 137.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 -135.67 137.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 2.86 139.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -53.32 139.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -135.67 139.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 2.86 141 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -44.84 141 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -135.67 141 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 2.86 142.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 -135.67 142.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 2.86 144.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -135.67 144.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 2.86 145.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 -135.67 145.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 2.86 147.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 -135.67 147.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 2.86 149 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -44.84 149 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -109.5 149 -100.38 ;
        RECT 148.635 -109.535 148.965 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 2.86 150.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -44.84 150.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -135.67 150.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 2.86 152.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 -115.86 152.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 2.86 153.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -114.8 153.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -135.67 153.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 2.86 155.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -135.67 155.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 2.86 157 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 -135.67 157 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 2.86 158.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -44.84 158.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -109.5 158.6 -100.38 ;
        RECT 158.235 -109.535 158.565 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 2.86 160.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -44.84 160.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -135.67 160.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 2.86 161.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 -135.67 161.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 2.86 163.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 -135.67 163.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 2.86 165 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 -135.67 165 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 2.86 166.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 -135.67 166.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 2.86 168.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -44.84 168.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -109.5 168.2 -100.38 ;
        RECT 167.835 -109.535 168.165 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 2.86 169.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -53.32 169.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -135.67 169.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 2.86 171.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 -135.67 171.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 2.86 173 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -114.8 173 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 2.86 174.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -135.67 174.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 2.86 176.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 -135.67 176.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 2.86 177.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 -135.67 177.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 2.86 179.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 -53.32 179.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 -135.67 179.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 2.86 181 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 -44.84 181 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 -135.67 181 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 2.86 182.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 -135.67 182.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 2.86 184.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 -135.67 184.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 2.86 185.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 -135.67 185.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 2.86 187.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 -135.67 187.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 2.86 189 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 -44.84 189 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 -109.5 189 -100.38 ;
        RECT 188.635 -109.535 188.965 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 2.86 190.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 -44.84 190.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 -135.67 190.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 2.86 192.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 -115.86 192.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 2.86 193.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -114.8 193.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -135.67 193.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 2.86 195.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -135.67 195.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 2.86 197 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 -135.67 197 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 2.86 198.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 -44.84 198.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 -109.5 198.6 -100.38 ;
        RECT 198.235 -109.535 198.565 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 2.86 200.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 -44.84 200.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 -135.67 200.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 2.86 201.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 -135.67 201.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 2.86 203.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 -135.67 203.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 2.86 205 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 -135.67 205 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 2.86 206.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 -135.67 206.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 2.86 208.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 -44.84 208.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 -109.5 208.2 -100.38 ;
        RECT 207.835 -109.535 208.165 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 2.86 209.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 -53.32 209.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 -135.67 209.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 2.86 211.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 -135.67 211.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 2.86 213 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 -114.8 213 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 2.86 214.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 -135.67 214.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 2.86 216.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 -135.67 216.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 2.86 217.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 -135.67 217.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 2.86 219.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 -53.32 219.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 -135.67 219.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 2.86 221 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 -44.84 221 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 -135.67 221 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 2.86 222.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 -135.67 222.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 2.86 224.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 -135.67 224.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 2.86 225.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 -135.67 225.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 2.86 227.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 -135.67 227.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 2.86 229 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 -44.84 229 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 -109.5 229 -100.38 ;
        RECT 228.635 -109.535 228.965 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 2.86 230.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 -44.84 230.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 -135.67 230.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 2.86 232.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 -115.86 232.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 2.86 233.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -114.8 233.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -135.67 233.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 2.86 235.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 -135.67 235.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 2.86 237 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 -135.67 237 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 2.86 238.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 -44.84 238.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 -109.5 238.6 -100.38 ;
        RECT 238.235 -109.535 238.565 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 2.86 240.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 -44.84 240.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 -135.67 240.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 2.86 241.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 -135.67 241.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 2.86 243.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 -135.67 243.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 2.86 245 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 -135.67 245 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 2.86 246.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 -135.67 246.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 2.86 248.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 -44.84 248.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 -109.5 248.2 -100.38 ;
        RECT 247.835 -109.535 248.165 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 2.86 249.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -53.32 249.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -135.67 249.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 2.86 251.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 -135.67 251.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 2.86 253 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 -114.8 253 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 2.86 254.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 -135.67 254.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 2.86 256.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 -135.67 256.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 2.86 257.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 -135.67 257.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 2.86 259.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 -53.32 259.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 -135.67 259.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 2.86 261 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 -44.84 261 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 -135.67 261 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 2.86 262.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 -135.67 262.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 2.86 264.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 -135.67 264.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 2.86 265.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 -135.67 265.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 2.86 267.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 -135.67 267.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 2.86 269 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 -44.84 269 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 -109.5 269 -100.38 ;
        RECT 268.635 -109.535 268.965 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 2.86 270.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 -44.84 270.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 -135.67 270.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 2.86 272.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 -115.86 272.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 2.86 273.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -114.8 273.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -135.67 273.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 2.86 275.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 -135.67 275.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 2.86 277 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 -135.67 277 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 2.86 278.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 -44.84 278.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 -109.5 278.6 -100.38 ;
        RECT 278.235 -109.535 278.565 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 2.86 280.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 -44.84 280.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 -135.67 280.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 2.86 281.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 -135.67 281.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 2.86 283.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 -135.67 283.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 2.86 285 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 -135.67 285 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 2.86 286.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 -135.67 286.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 2.86 288.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 -44.84 288.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 -109.5 288.2 -100.38 ;
        RECT 287.835 -109.535 288.165 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 2.86 289.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 -53.32 289.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 -135.67 289.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 2.86 291.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 -135.67 291.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 2.86 293 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 -114.8 293 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 2.86 294.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 -135.67 294.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 2.86 296.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 -135.67 296.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 2.86 297.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 -135.67 297.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 2.86 299.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 -53.32 299.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 -135.67 299.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 2.86 301 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 -44.84 301 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 -135.67 301 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 2.86 302.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 -135.67 302.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 2.86 304.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 -135.67 304.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 2.86 305.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 -135.67 305.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 2.86 307.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 -135.67 307.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 2.86 309 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 -44.84 309 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 -109.5 309 -100.38 ;
        RECT 308.635 -109.535 308.965 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 2.86 310.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 -44.84 310.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 -135.67 310.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 2.86 312.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 -115.86 312.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 2.86 313.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -114.8 313.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -135.67 313.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 2.86 315.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 -135.67 315.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 2.86 317 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 -135.67 317 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 2.86 318.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 -44.84 318.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 -109.5 318.6 -100.38 ;
        RECT 318.235 -109.535 318.565 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 2.86 320.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 -44.84 320.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 -135.67 320.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 2.86 321.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 -135.67 321.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 2.86 323.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 -135.67 323.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 2.86 325 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 -135.67 325 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 2.86 326.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 -135.67 326.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 2.86 328.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 -135.67 328.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 2.86 329.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 -135.67 329.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 331 -135.67 331.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 -135.67 333 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 -135.67 334.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.8 -135.67 336.2 11.315 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -66.6 -134.13 -66.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -134.13 -64.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.4 -134.13 -63 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -134.13 -61.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.2 -134.13 -59.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -134.13 -58.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -57 -134.13 -56.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.4 -134.13 -55 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -134.13 -53.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.2 -134.13 -51.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -134.13 -50.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -49 -134.13 -48.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -134.13 -47 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.8 -113.74 -45.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -112.68 -43.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -134.13 -43.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.6 -134.13 -42.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -108.44 -40.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -134.13 -40.6 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.4 -112.68 -39 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.8 -134.13 -37.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -107.38 -35.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -134.13 -35.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.6 -107.38 -34.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -112.68 -32.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -134.13 -32.6 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.4 -134.13 -31 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -106.32 -29.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -134.13 -29.4 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.2 -113.74 -27.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -112.68 -26.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -134.13 -26.2 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -25 -134.13 -24.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -105.26 -23 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -134.13 -23 -115.22 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.8 -112.68 -21.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.2 -134.13 -19.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -104.2 -18.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -134.13 -18.2 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -17 -105.26 -16.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -112.68 -15 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -134.13 -15 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.8 -134.13 -13.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -103.14 -11.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -134.13 -11.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -35.3 -10.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -113.74 -10.2 -82.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -112.68 -8.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -134.13 -8.6 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.4 -134.13 -7 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -98.9 -5.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -134.13 -5.4 -115.22 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.2 -134.13 -3.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.6 -134.13 -2.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 2.86 -0.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 -134.13 -0.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 2.86 1 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 -134.13 1 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 2.86 2.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 -134.13 2.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 2.86 4.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 -134.13 4.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 2.86 5.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -73.46 5.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -134.13 5.8 -80.24 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 2.86 7.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 -134.13 7.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 2.86 9 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -44.84 9 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -109.5 9 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 2.86 10.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -44.84 10.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -134.13 10.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 2.86 12.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 -115.86 12.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 2.86 13.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -114.8 13.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -134.13 13.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 2.86 15.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -134.13 15.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 2.86 17 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 -134.13 17 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 2.86 18.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -44.84 18.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -109.5 18.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 2.86 20.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -44.84 20.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -134.13 20.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 2.86 21.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -134.13 21.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 2.86 23.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 -134.13 23.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 2.86 25 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 -134.13 25 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 2.86 26.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 -134.13 26.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 2.86 28.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -44.84 28.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -109.5 28.2 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 2.86 29.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -53.32 29.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -134.13 29.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 2.86 31.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 -134.13 31.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 2.86 33 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -114.8 33 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 2.86 34.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -134.13 34.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 2.86 36.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -134.13 36.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 2.86 37.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 -134.13 37.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 2.86 39.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -53.32 39.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -134.13 39.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 2.86 41 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -44.84 41 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -134.13 41 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 2.86 42.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 -134.13 42.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 2.86 44.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 -134.13 44.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 2.86 45.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 -134.13 45.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 2.86 47.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 -134.13 47.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 2.86 49 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -44.84 49 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -109.5 49 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 2.86 50.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -44.84 50.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -134.13 50.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 2.86 52.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 -115.86 52.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 2.86 53.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -114.8 53.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -134.13 53.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 2.86 55.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -134.13 55.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 2.86 57 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 -134.13 57 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 2.86 58.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -44.84 58.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -109.5 58.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 2.86 60.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -44.84 60.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -134.13 60.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 2.86 61.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 -134.13 61.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 2.86 63.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 -134.13 63.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 2.86 65 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 -134.13 65 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 2.86 66.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 -134.13 66.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 2.86 68.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -44.84 68.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -109.5 68.2 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 2.86 69.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -53.32 69.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -134.13 69.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 2.86 71.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 -134.13 71.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 2.86 73 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -114.8 73 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 2.86 74.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -134.13 74.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 2.86 76.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 -134.13 76.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 2.86 77.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 -134.13 77.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 2.86 79.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -53.32 79.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -134.13 79.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 2.86 81 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -44.84 81 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -134.13 81 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 2.86 82.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 -134.13 82.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 2.86 84.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 -134.13 84.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 2.86 85.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 -134.13 85.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 2.86 87.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 -134.13 87.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 2.86 89 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -44.84 89 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -109.5 89 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 2.86 90.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -44.84 90.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -134.13 90.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 2.86 92.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 -115.86 92.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 2.86 93.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -114.8 93.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -134.13 93.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 2.86 95.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -134.13 95.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 2.86 97 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 -134.13 97 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 2.86 98.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -44.84 98.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -109.5 98.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 2.86 100.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -44.84 100.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -134.13 100.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 2.86 101.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -134.13 101.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 2.86 103.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 -134.13 103.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 2.86 105 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 -134.13 105 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 2.86 106.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 -134.13 106.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 2.86 108.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -44.84 108.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -109.5 108.2 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 2.86 109.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -53.32 109.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -134.13 109.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 2.86 111.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 -134.13 111.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 2.86 113 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -114.8 113 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 2.86 114.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -134.13 114.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 2.86 116.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 -134.13 116.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 2.86 117.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 -134.13 117.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 2.86 119.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -53.32 119.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -134.13 119.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 2.86 121 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -44.84 121 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -134.13 121 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 2.86 122.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 -134.13 122.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 2.86 124.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 -134.13 124.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 2.86 125.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 -134.13 125.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 2.86 127.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 -134.13 127.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 2.86 129 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -44.84 129 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -109.5 129 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 2.86 130.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -44.84 130.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -134.13 130.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 2.86 132.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 -115.86 132.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 2.86 133.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -114.8 133.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -134.13 133.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 2.86 135.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -134.13 135.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 2.86 137 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 -134.13 137 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 2.86 138.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -44.84 138.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -109.5 138.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 2.86 140.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -44.84 140.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -134.13 140.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 2.86 141.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 -134.13 141.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 2.86 143.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 -134.13 143.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 2.86 145 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 -134.13 145 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 2.86 146.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 -134.13 146.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 2.86 148.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -44.84 148.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -109.5 148.2 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 2.86 149.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -53.32 149.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -134.13 149.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 2.86 151.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 -134.13 151.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 2.86 153 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -114.8 153 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 2.86 154.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -134.13 154.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 2.86 156.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 -134.13 156.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 2.86 157.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 -134.13 157.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 2.86 159.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -53.32 159.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -134.13 159.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 2.86 161 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -44.84 161 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -134.13 161 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 2.86 162.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 -134.13 162.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 2.86 164.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 -134.13 164.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 2.86 165.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 -134.13 165.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 2.86 167.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 -134.13 167.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 2.86 169 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -44.84 169 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -109.5 169 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 2.86 170.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -44.84 170.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -134.13 170.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 2.86 172.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 -115.86 172.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 2.86 173.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -114.8 173.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -134.13 173.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 2.86 175.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -134.13 175.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 2.86 177 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 -134.13 177 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 2.86 178.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 -44.84 178.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 -109.5 178.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 2.86 180.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 -44.84 180.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 -134.13 180.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 2.86 181.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 -134.13 181.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 2.86 183.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 -134.13 183.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 2.86 185 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 -134.13 185 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 2.86 186.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 -134.13 186.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 2.86 188.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 -44.84 188.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 -109.5 188.2 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 2.86 189.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 -53.32 189.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 -134.13 189.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 2.86 191.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 -134.13 191.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 2.86 193 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 -114.8 193 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 2.86 194.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 -134.13 194.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 2.86 196.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 -134.13 196.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 2.86 197.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 -134.13 197.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 2.86 199.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 -53.32 199.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 -134.13 199.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 2.86 201 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 -44.84 201 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 -134.13 201 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 2.86 202.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 -134.13 202.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 2.86 204.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 -134.13 204.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 2.86 205.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 -134.13 205.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 2.86 207.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 -134.13 207.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 2.86 209 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 -44.84 209 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 -109.5 209 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 2.86 210.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 -44.84 210.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 -134.13 210.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 2.86 212.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 -115.86 212.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 2.86 213.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -114.8 213.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -134.13 213.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 2.86 215.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 -134.13 215.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 2.86 217 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 -134.13 217 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 2.86 218.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 -44.84 218.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 -109.5 218.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 2.86 220.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 -44.84 220.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 -134.13 220.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 2.86 221.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 -134.13 221.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 2.86 223.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 -134.13 223.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 2.86 225 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 -134.13 225 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 2.86 226.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 -134.13 226.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 2.86 228.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 -44.84 228.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 -109.5 228.2 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 2.86 229.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 -53.32 229.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 -134.13 229.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 2.86 231.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 -134.13 231.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 2.86 233 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 -114.8 233 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 2.86 234.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 -134.13 234.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 2.86 236.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 -134.13 236.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 2.86 237.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 -134.13 237.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 2.86 239.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 -53.32 239.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 -134.13 239.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 2.86 241 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 -44.84 241 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 -134.13 241 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 2.86 242.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 -134.13 242.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 2.86 244.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 -134.13 244.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 2.86 245.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 -134.13 245.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 2.86 247.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 -134.13 247.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 2.86 249 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 -44.84 249 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 -109.5 249 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 2.86 250.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 -44.84 250.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 -134.13 250.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 2.86 252.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 -115.86 252.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 2.86 253.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -114.8 253.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -134.13 253.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 2.86 255.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 -134.13 255.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 2.86 257 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 -134.13 257 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 2.86 258.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 -44.84 258.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 -109.5 258.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 2.86 260.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 -44.84 260.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 -134.13 260.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 2.86 261.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 -134.13 261.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 2.86 263.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 -134.13 263.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 2.86 265 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 -134.13 265 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 2.86 266.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 -134.13 266.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 2.86 268.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 -44.84 268.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 -109.5 268.2 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 2.86 269.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 -53.32 269.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 -134.13 269.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 2.86 271.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 -134.13 271.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 2.86 273 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 -114.8 273 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 2.86 274.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 -134.13 274.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 2.86 276.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 -134.13 276.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 2.86 277.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 -134.13 277.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 2.86 279.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 -53.32 279.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 -134.13 279.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 2.86 281 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 -44.84 281 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 -134.13 281 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 2.86 282.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 -134.13 282.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 2.86 284.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 -134.13 284.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 2.86 285.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 -134.13 285.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 2.86 287.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 -134.13 287.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 2.86 289 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 -44.84 289 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 -109.5 289 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 2.86 290.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -44.84 290.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -134.13 290.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 2.86 292.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 -115.86 292.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 2.86 293.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -114.8 293.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -134.13 293.8 -129 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 2.86 295.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 -134.13 295.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 2.86 297 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 -134.13 297 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 2.86 298.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 -44.84 298.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 -109.5 298.6 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 2.86 300.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 -44.84 300.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 -134.13 300.2 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 2.86 301.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 -134.13 301.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 2.86 303.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 -134.13 303.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 2.86 305 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 -134.13 305 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 2.86 306.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 -134.13 306.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 2.86 308.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 -44.84 308.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 -109.5 308.2 -100.38 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 2.86 309.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 -53.32 309.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 -134.13 309.8 -116.28 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 2.86 311.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 -134.13 311.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 2.86 313 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 -114.8 313 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 2.86 314.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 -134.13 314.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 2.86 316.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 -134.13 316.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 2.86 317.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 -134.13 317.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 2.86 319.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 -53.32 319.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 -134.13 319.4 -124.76 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 2.86 321 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 -44.84 321 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 -134.13 321 -100.38 ;
        RECT 320.58 -100.785 321 -100.455 ;
        RECT 320.58 -106.395 321 -106.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 2.86 322.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 -134.13 322.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 2.86 324.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 -134.13 324.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 2.86 325.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 -134.13 325.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 2.86 327.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 -134.13 327.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 2.86 329 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 -134.13 329 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 2.86 330.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 -134.13 330.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.8 -134.13 332.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 -134.13 333.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 -134.13 335.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.6 -134.13 337 9.775 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -16.46 -136.07 -16.16 -135.77 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -22.3 -136.07 -22 -135.77 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.14 -136.07 -27.84 -135.77 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -33.98 -136.07 -33.68 -135.77 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -39.82 -136.07 -39.52 -135.77 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -45.66 -136.07 -45.36 -135.77 ;
    END
  END addr[5]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -46.68 -136.07 -46.26 -135.65 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.015 -136.07 12.315 -135.77 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.015 -136.07 112.315 -135.77 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.63 -136.07 112.93 -135.77 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.015 -136.07 132.315 -135.77 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.63 -136.07 132.93 -135.77 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.015 -136.07 152.315 -135.77 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.63 -136.07 152.93 -135.77 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 172.015 -136.07 172.315 -135.77 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 172.63 -136.07 172.93 -135.77 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 192.015 -136.07 192.315 -135.77 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 192.63 -136.07 192.93 -135.77 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.63 -136.07 12.93 -135.77 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.015 -136.07 212.315 -135.77 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.63 -136.07 212.93 -135.77 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.015 -136.07 232.315 -135.77 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.63 -136.07 232.93 -135.77 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 252.015 -136.07 252.315 -135.77 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 252.63 -136.07 252.93 -135.77 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 272.015 -136.07 272.315 -135.77 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 272.63 -136.07 272.93 -135.77 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 292.015 -136.07 292.315 -135.77 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 292.63 -136.07 292.93 -135.77 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 32.015 -136.07 32.315 -135.77 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 312.015 -136.07 312.315 -135.77 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 312.63 -136.07 312.93 -135.77 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 32.63 -136.07 32.93 -135.77 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.015 -136.07 52.315 -135.77 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.63 -136.07 52.93 -135.77 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.015 -136.07 72.315 -135.77 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.63 -136.07 72.93 -135.77 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 92.015 -136.07 92.315 -135.77 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 92.63 -136.07 92.93 -135.77 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.285 -136.07 8.585 -135.77 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.285 -136.07 108.585 -135.77 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.285 -136.07 118.585 -135.77 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.285 -136.07 128.585 -135.77 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.285 -136.07 138.585 -135.77 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.285 -136.07 148.585 -135.77 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.285 -136.07 158.585 -135.77 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 168.285 -136.07 168.585 -135.77 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.285 -136.07 178.585 -135.77 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 188.285 -136.07 188.585 -135.77 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 198.285 -136.07 198.585 -135.77 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.285 -136.07 18.585 -135.77 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 208.285 -136.07 208.585 -135.77 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.285 -136.07 218.585 -135.77 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 228.285 -136.07 228.585 -135.77 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 238.285 -136.07 238.585 -135.77 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 248.285 -136.07 248.585 -135.77 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 258.285 -136.07 258.585 -135.77 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.285 -136.07 268.585 -135.77 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 278.285 -136.07 278.585 -135.77 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 288.285 -136.07 288.585 -135.77 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 298.285 -136.07 298.585 -135.77 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.285 -136.07 28.585 -135.77 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.285 -136.07 308.585 -135.77 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 318.285 -136.07 318.585 -135.77 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 38.285 -136.07 38.585 -135.77 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.285 -136.07 48.585 -135.77 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.285 -136.07 58.585 -135.77 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.285 -136.07 68.585 -135.77 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.285 -136.07 78.585 -135.77 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 88.285 -136.07 88.585 -135.77 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 98.285 -136.07 98.585 -135.77 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -10.62 -136.07 -10.32 -135.77 ;
    END
  END we
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -72.135 -136.07 342.46 11.715 ;
    LAYER met2 SPACING 0.14 ;
      RECT -72.135 -136.07 342.46 11.715 ;
    LAYER met3 SPACING 0.3 ;
      RECT 320.115 -84.585 320.445 -84.255 ;
      RECT 320.13 -100.015 320.43 -84.255 ;
      RECT 320.115 -100.015 320.445 -99.685 ;
      RECT 320.13 -80.8 320.43 -45.52 ;
      RECT 320.115 -47.495 320.445 -47.165 ;
      RECT 320.115 -80.39 320.445 -80.06 ;
      RECT 319.515 -123.905 319.815 -54.615 ;
      RECT 319.5 -54.99 319.83 -54.66 ;
      RECT 319.5 -68.17 319.83 -67.84 ;
      RECT 319.5 -123.905 319.83 -123.575 ;
      RECT 318.9 -63.51 319.2 -55.245 ;
      RECT 318.885 -55.62 319.215 -55.29 ;
      RECT 318.885 -63.51 319.215 -63.18 ;
      RECT 318.27 -110.99 318.6 -110.66 ;
      RECT 318.285 -135.28 318.585 -110.66 ;
      RECT 318.27 -85.045 318.6 -84.715 ;
      RECT 318.285 -100.015 318.585 -84.715 ;
      RECT 318.27 -100.015 318.6 -99.685 ;
      RECT 318.285 -80.82 318.585 -45.52 ;
      RECT 318.27 -45.895 318.6 -45.565 ;
      RECT 318.27 -80.82 318.6 -80.49 ;
      RECT 313.245 -116.38 313.575 -116.05 ;
      RECT 313.26 -128.01 313.56 -116.05 ;
      RECT 313.245 -123.62 313.575 -123.29 ;
      RECT 313.245 -127.965 313.575 -127.635 ;
      RECT 312.615 -122.82 312.945 -122.49 ;
      RECT 312.63 -135.28 312.93 -122.49 ;
      RECT 312 -117.18 312.33 -116.85 ;
      RECT 312.015 -135.28 312.315 -116.85 ;
      RECT 310.115 -84.585 310.445 -84.255 ;
      RECT 310.13 -100.015 310.43 -84.255 ;
      RECT 310.115 -100.015 310.445 -99.685 ;
      RECT 310.13 -80.8 310.43 -45.52 ;
      RECT 310.115 -47.495 310.445 -47.165 ;
      RECT 310.115 -80.39 310.445 -80.06 ;
      RECT 309.515 -115.895 309.815 -54.615 ;
      RECT 309.5 -54.99 309.83 -54.66 ;
      RECT 309.5 -68.17 309.83 -67.84 ;
      RECT 309.5 -115.895 309.83 -115.565 ;
      RECT 308.9 -63.51 309.2 -55.245 ;
      RECT 308.885 -55.62 309.215 -55.29 ;
      RECT 308.885 -63.51 309.215 -63.18 ;
      RECT 308.27 -110.99 308.6 -110.66 ;
      RECT 308.285 -135.28 308.585 -110.66 ;
      RECT 308.27 -85.045 308.6 -84.715 ;
      RECT 308.285 -100.015 308.585 -84.715 ;
      RECT 308.27 -100.015 308.6 -99.685 ;
      RECT 308.285 -80.82 308.585 -45.52 ;
      RECT 308.27 -45.895 308.6 -45.565 ;
      RECT 308.27 -80.82 308.6 -80.49 ;
      RECT 300.115 -84.585 300.445 -84.255 ;
      RECT 300.13 -100.015 300.43 -84.255 ;
      RECT 300.115 -100.015 300.445 -99.685 ;
      RECT 300.13 -80.8 300.43 -45.52 ;
      RECT 300.115 -47.495 300.445 -47.165 ;
      RECT 300.115 -80.39 300.445 -80.06 ;
      RECT 299.515 -123.905 299.815 -54.615 ;
      RECT 299.5 -54.99 299.83 -54.66 ;
      RECT 299.5 -68.17 299.83 -67.84 ;
      RECT 299.5 -123.905 299.83 -123.575 ;
      RECT 298.9 -63.51 299.2 -55.245 ;
      RECT 298.885 -55.62 299.215 -55.29 ;
      RECT 298.885 -63.51 299.215 -63.18 ;
      RECT 298.27 -110.99 298.6 -110.66 ;
      RECT 298.285 -135.28 298.585 -110.66 ;
      RECT 298.27 -85.045 298.6 -84.715 ;
      RECT 298.285 -100.015 298.585 -84.715 ;
      RECT 298.27 -100.015 298.6 -99.685 ;
      RECT 298.285 -80.82 298.585 -45.52 ;
      RECT 298.27 -45.895 298.6 -45.565 ;
      RECT 298.27 -80.82 298.6 -80.49 ;
      RECT 293.245 -116.38 293.575 -116.05 ;
      RECT 293.26 -128.01 293.56 -116.05 ;
      RECT 293.245 -123.62 293.575 -123.29 ;
      RECT 293.245 -127.965 293.575 -127.635 ;
      RECT 292.615 -122.82 292.945 -122.49 ;
      RECT 292.63 -135.28 292.93 -122.49 ;
      RECT 292 -117.18 292.33 -116.85 ;
      RECT 292.015 -135.28 292.315 -116.85 ;
      RECT 290.115 -84.585 290.445 -84.255 ;
      RECT 290.13 -100.015 290.43 -84.255 ;
      RECT 290.115 -100.015 290.445 -99.685 ;
      RECT 290.13 -80.8 290.43 -45.52 ;
      RECT 290.115 -47.495 290.445 -47.165 ;
      RECT 290.115 -80.39 290.445 -80.06 ;
      RECT 289.515 -115.895 289.815 -54.615 ;
      RECT 289.5 -54.99 289.83 -54.66 ;
      RECT 289.5 -68.17 289.83 -67.84 ;
      RECT 289.5 -115.895 289.83 -115.565 ;
      RECT 288.9 -63.51 289.2 -55.245 ;
      RECT 288.885 -55.62 289.215 -55.29 ;
      RECT 288.885 -63.51 289.215 -63.18 ;
      RECT 288.27 -110.99 288.6 -110.66 ;
      RECT 288.285 -135.28 288.585 -110.66 ;
      RECT 288.27 -85.045 288.6 -84.715 ;
      RECT 288.285 -100.015 288.585 -84.715 ;
      RECT 288.27 -100.015 288.6 -99.685 ;
      RECT 288.285 -80.82 288.585 -45.52 ;
      RECT 288.27 -45.895 288.6 -45.565 ;
      RECT 288.27 -80.82 288.6 -80.49 ;
      RECT 280.115 -84.585 280.445 -84.255 ;
      RECT 280.13 -100.015 280.43 -84.255 ;
      RECT 280.115 -100.015 280.445 -99.685 ;
      RECT 280.13 -80.8 280.43 -45.52 ;
      RECT 280.115 -47.495 280.445 -47.165 ;
      RECT 280.115 -80.39 280.445 -80.06 ;
      RECT 279.515 -123.905 279.815 -54.615 ;
      RECT 279.5 -54.99 279.83 -54.66 ;
      RECT 279.5 -68.17 279.83 -67.84 ;
      RECT 279.5 -123.905 279.83 -123.575 ;
      RECT 278.9 -63.51 279.2 -55.245 ;
      RECT 278.885 -55.62 279.215 -55.29 ;
      RECT 278.885 -63.51 279.215 -63.18 ;
      RECT 278.27 -110.99 278.6 -110.66 ;
      RECT 278.285 -135.28 278.585 -110.66 ;
      RECT 278.27 -85.045 278.6 -84.715 ;
      RECT 278.285 -100.015 278.585 -84.715 ;
      RECT 278.27 -100.015 278.6 -99.685 ;
      RECT 278.285 -80.82 278.585 -45.52 ;
      RECT 278.27 -45.895 278.6 -45.565 ;
      RECT 278.27 -80.82 278.6 -80.49 ;
      RECT 273.245 -116.38 273.575 -116.05 ;
      RECT 273.26 -128.01 273.56 -116.05 ;
      RECT 273.245 -123.62 273.575 -123.29 ;
      RECT 273.245 -127.965 273.575 -127.635 ;
      RECT 272.615 -122.82 272.945 -122.49 ;
      RECT 272.63 -135.28 272.93 -122.49 ;
      RECT 272 -117.18 272.33 -116.85 ;
      RECT 272.015 -135.28 272.315 -116.85 ;
      RECT 270.115 -84.585 270.445 -84.255 ;
      RECT 270.13 -100.015 270.43 -84.255 ;
      RECT 270.115 -100.015 270.445 -99.685 ;
      RECT 270.13 -80.8 270.43 -45.52 ;
      RECT 270.115 -47.495 270.445 -47.165 ;
      RECT 270.115 -80.39 270.445 -80.06 ;
      RECT 269.515 -115.895 269.815 -54.615 ;
      RECT 269.5 -54.99 269.83 -54.66 ;
      RECT 269.5 -68.17 269.83 -67.84 ;
      RECT 269.5 -115.895 269.83 -115.565 ;
      RECT 268.9 -63.51 269.2 -55.245 ;
      RECT 268.885 -55.62 269.215 -55.29 ;
      RECT 268.885 -63.51 269.215 -63.18 ;
      RECT 268.27 -110.99 268.6 -110.66 ;
      RECT 268.285 -135.28 268.585 -110.66 ;
      RECT 268.27 -85.045 268.6 -84.715 ;
      RECT 268.285 -100.015 268.585 -84.715 ;
      RECT 268.27 -100.015 268.6 -99.685 ;
      RECT 268.285 -80.82 268.585 -45.52 ;
      RECT 268.27 -45.895 268.6 -45.565 ;
      RECT 268.27 -80.82 268.6 -80.49 ;
      RECT 260.115 -84.585 260.445 -84.255 ;
      RECT 260.13 -100.015 260.43 -84.255 ;
      RECT 260.115 -100.015 260.445 -99.685 ;
      RECT 260.13 -80.8 260.43 -45.52 ;
      RECT 260.115 -47.495 260.445 -47.165 ;
      RECT 260.115 -80.39 260.445 -80.06 ;
      RECT 259.515 -123.905 259.815 -54.615 ;
      RECT 259.5 -54.99 259.83 -54.66 ;
      RECT 259.5 -68.17 259.83 -67.84 ;
      RECT 259.5 -123.905 259.83 -123.575 ;
      RECT 258.9 -63.51 259.2 -55.245 ;
      RECT 258.885 -55.62 259.215 -55.29 ;
      RECT 258.885 -63.51 259.215 -63.18 ;
      RECT 258.27 -110.99 258.6 -110.66 ;
      RECT 258.285 -135.28 258.585 -110.66 ;
      RECT 258.27 -85.045 258.6 -84.715 ;
      RECT 258.285 -100.015 258.585 -84.715 ;
      RECT 258.27 -100.015 258.6 -99.685 ;
      RECT 258.285 -80.82 258.585 -45.52 ;
      RECT 258.27 -45.895 258.6 -45.565 ;
      RECT 258.27 -80.82 258.6 -80.49 ;
      RECT 253.245 -116.38 253.575 -116.05 ;
      RECT 253.26 -128.01 253.56 -116.05 ;
      RECT 253.245 -123.62 253.575 -123.29 ;
      RECT 253.245 -127.965 253.575 -127.635 ;
      RECT 252.615 -122.82 252.945 -122.49 ;
      RECT 252.63 -135.28 252.93 -122.49 ;
      RECT 252 -117.18 252.33 -116.85 ;
      RECT 252.015 -135.28 252.315 -116.85 ;
      RECT 250.115 -84.585 250.445 -84.255 ;
      RECT 250.13 -100.015 250.43 -84.255 ;
      RECT 250.115 -100.015 250.445 -99.685 ;
      RECT 250.13 -80.8 250.43 -45.52 ;
      RECT 250.115 -47.495 250.445 -47.165 ;
      RECT 250.115 -80.39 250.445 -80.06 ;
      RECT 249.515 -115.895 249.815 -54.615 ;
      RECT 249.5 -54.99 249.83 -54.66 ;
      RECT 249.5 -68.17 249.83 -67.84 ;
      RECT 249.5 -115.895 249.83 -115.565 ;
      RECT 248.9 -63.51 249.2 -55.245 ;
      RECT 248.885 -55.62 249.215 -55.29 ;
      RECT 248.885 -63.51 249.215 -63.18 ;
      RECT 248.27 -110.99 248.6 -110.66 ;
      RECT 248.285 -135.28 248.585 -110.66 ;
      RECT 248.27 -85.045 248.6 -84.715 ;
      RECT 248.285 -100.015 248.585 -84.715 ;
      RECT 248.27 -100.015 248.6 -99.685 ;
      RECT 248.285 -80.82 248.585 -45.52 ;
      RECT 248.27 -45.895 248.6 -45.565 ;
      RECT 248.27 -80.82 248.6 -80.49 ;
      RECT 240.115 -84.585 240.445 -84.255 ;
      RECT 240.13 -100.015 240.43 -84.255 ;
      RECT 240.115 -100.015 240.445 -99.685 ;
      RECT 240.13 -80.8 240.43 -45.52 ;
      RECT 240.115 -47.495 240.445 -47.165 ;
      RECT 240.115 -80.39 240.445 -80.06 ;
      RECT 239.515 -123.905 239.815 -54.615 ;
      RECT 239.5 -54.99 239.83 -54.66 ;
      RECT 239.5 -68.17 239.83 -67.84 ;
      RECT 239.5 -123.905 239.83 -123.575 ;
      RECT 238.9 -63.51 239.2 -55.245 ;
      RECT 238.885 -55.62 239.215 -55.29 ;
      RECT 238.885 -63.51 239.215 -63.18 ;
      RECT 238.27 -110.99 238.6 -110.66 ;
      RECT 238.285 -135.28 238.585 -110.66 ;
      RECT 238.27 -85.045 238.6 -84.715 ;
      RECT 238.285 -100.015 238.585 -84.715 ;
      RECT 238.27 -100.015 238.6 -99.685 ;
      RECT 238.285 -80.82 238.585 -45.52 ;
      RECT 238.27 -45.895 238.6 -45.565 ;
      RECT 238.27 -80.82 238.6 -80.49 ;
      RECT 233.245 -116.38 233.575 -116.05 ;
      RECT 233.26 -128.01 233.56 -116.05 ;
      RECT 233.245 -123.62 233.575 -123.29 ;
      RECT 233.245 -127.965 233.575 -127.635 ;
      RECT 232.615 -122.82 232.945 -122.49 ;
      RECT 232.63 -135.28 232.93 -122.49 ;
      RECT 232 -117.18 232.33 -116.85 ;
      RECT 232.015 -135.28 232.315 -116.85 ;
      RECT 230.115 -84.585 230.445 -84.255 ;
      RECT 230.13 -100.015 230.43 -84.255 ;
      RECT 230.115 -100.015 230.445 -99.685 ;
      RECT 230.13 -80.8 230.43 -45.52 ;
      RECT 230.115 -47.495 230.445 -47.165 ;
      RECT 230.115 -80.39 230.445 -80.06 ;
      RECT 229.515 -115.895 229.815 -54.615 ;
      RECT 229.5 -54.99 229.83 -54.66 ;
      RECT 229.5 -68.17 229.83 -67.84 ;
      RECT 229.5 -115.895 229.83 -115.565 ;
      RECT 228.9 -63.51 229.2 -55.245 ;
      RECT 228.885 -55.62 229.215 -55.29 ;
      RECT 228.885 -63.51 229.215 -63.18 ;
      RECT 228.27 -110.99 228.6 -110.66 ;
      RECT 228.285 -135.28 228.585 -110.66 ;
      RECT 228.27 -85.045 228.6 -84.715 ;
      RECT 228.285 -100.015 228.585 -84.715 ;
      RECT 228.27 -100.015 228.6 -99.685 ;
      RECT 228.285 -80.82 228.585 -45.52 ;
      RECT 228.27 -45.895 228.6 -45.565 ;
      RECT 228.27 -80.82 228.6 -80.49 ;
      RECT 220.115 -84.585 220.445 -84.255 ;
      RECT 220.13 -100.015 220.43 -84.255 ;
      RECT 220.115 -100.015 220.445 -99.685 ;
      RECT 220.13 -80.8 220.43 -45.52 ;
      RECT 220.115 -47.495 220.445 -47.165 ;
      RECT 220.115 -80.39 220.445 -80.06 ;
      RECT 219.515 -123.905 219.815 -54.615 ;
      RECT 219.5 -54.99 219.83 -54.66 ;
      RECT 219.5 -68.17 219.83 -67.84 ;
      RECT 219.5 -123.905 219.83 -123.575 ;
      RECT 218.9 -63.51 219.2 -55.245 ;
      RECT 218.885 -55.62 219.215 -55.29 ;
      RECT 218.885 -63.51 219.215 -63.18 ;
      RECT 218.27 -110.99 218.6 -110.66 ;
      RECT 218.285 -135.28 218.585 -110.66 ;
      RECT 218.27 -85.045 218.6 -84.715 ;
      RECT 218.285 -100.015 218.585 -84.715 ;
      RECT 218.27 -100.015 218.6 -99.685 ;
      RECT 218.285 -80.82 218.585 -45.52 ;
      RECT 218.27 -45.895 218.6 -45.565 ;
      RECT 218.27 -80.82 218.6 -80.49 ;
      RECT 213.245 -116.38 213.575 -116.05 ;
      RECT 213.26 -128.01 213.56 -116.05 ;
      RECT 213.245 -123.62 213.575 -123.29 ;
      RECT 213.245 -127.965 213.575 -127.635 ;
      RECT 212.615 -122.82 212.945 -122.49 ;
      RECT 212.63 -135.28 212.93 -122.49 ;
      RECT 212 -117.18 212.33 -116.85 ;
      RECT 212.015 -135.28 212.315 -116.85 ;
      RECT 210.115 -84.585 210.445 -84.255 ;
      RECT 210.13 -100.015 210.43 -84.255 ;
      RECT 210.115 -100.015 210.445 -99.685 ;
      RECT 210.13 -80.8 210.43 -45.52 ;
      RECT 210.115 -47.495 210.445 -47.165 ;
      RECT 210.115 -80.39 210.445 -80.06 ;
      RECT 209.515 -115.895 209.815 -54.615 ;
      RECT 209.5 -54.99 209.83 -54.66 ;
      RECT 209.5 -68.17 209.83 -67.84 ;
      RECT 209.5 -115.895 209.83 -115.565 ;
      RECT 208.9 -63.51 209.2 -55.245 ;
      RECT 208.885 -55.62 209.215 -55.29 ;
      RECT 208.885 -63.51 209.215 -63.18 ;
      RECT 208.27 -110.99 208.6 -110.66 ;
      RECT 208.285 -135.28 208.585 -110.66 ;
      RECT 208.27 -85.045 208.6 -84.715 ;
      RECT 208.285 -100.015 208.585 -84.715 ;
      RECT 208.27 -100.015 208.6 -99.685 ;
      RECT 208.285 -80.82 208.585 -45.52 ;
      RECT 208.27 -45.895 208.6 -45.565 ;
      RECT 208.27 -80.82 208.6 -80.49 ;
      RECT 200.115 -84.585 200.445 -84.255 ;
      RECT 200.13 -100.015 200.43 -84.255 ;
      RECT 200.115 -100.015 200.445 -99.685 ;
      RECT 200.13 -80.8 200.43 -45.52 ;
      RECT 200.115 -47.495 200.445 -47.165 ;
      RECT 200.115 -80.39 200.445 -80.06 ;
      RECT 199.515 -123.905 199.815 -54.615 ;
      RECT 199.5 -54.99 199.83 -54.66 ;
      RECT 199.5 -68.17 199.83 -67.84 ;
      RECT 199.5 -123.905 199.83 -123.575 ;
      RECT 198.9 -63.51 199.2 -55.245 ;
      RECT 198.885 -55.62 199.215 -55.29 ;
      RECT 198.885 -63.51 199.215 -63.18 ;
      RECT 198.27 -110.99 198.6 -110.66 ;
      RECT 198.285 -135.28 198.585 -110.66 ;
      RECT 198.27 -85.045 198.6 -84.715 ;
      RECT 198.285 -100.015 198.585 -84.715 ;
      RECT 198.27 -100.015 198.6 -99.685 ;
      RECT 198.285 -80.82 198.585 -45.52 ;
      RECT 198.27 -45.895 198.6 -45.565 ;
      RECT 198.27 -80.82 198.6 -80.49 ;
      RECT 193.245 -116.38 193.575 -116.05 ;
      RECT 193.26 -128.01 193.56 -116.05 ;
      RECT 193.245 -123.62 193.575 -123.29 ;
      RECT 193.245 -127.965 193.575 -127.635 ;
      RECT 192.615 -122.82 192.945 -122.49 ;
      RECT 192.63 -135.28 192.93 -122.49 ;
      RECT 192 -117.18 192.33 -116.85 ;
      RECT 192.015 -135.28 192.315 -116.85 ;
      RECT 190.115 -84.585 190.445 -84.255 ;
      RECT 190.13 -100.015 190.43 -84.255 ;
      RECT 190.115 -100.015 190.445 -99.685 ;
      RECT 190.13 -80.8 190.43 -45.52 ;
      RECT 190.115 -47.495 190.445 -47.165 ;
      RECT 190.115 -80.39 190.445 -80.06 ;
      RECT 189.515 -115.895 189.815 -54.615 ;
      RECT 189.5 -54.99 189.83 -54.66 ;
      RECT 189.5 -68.17 189.83 -67.84 ;
      RECT 189.5 -115.895 189.83 -115.565 ;
      RECT 188.9 -63.51 189.2 -55.245 ;
      RECT 188.885 -55.62 189.215 -55.29 ;
      RECT 188.885 -63.51 189.215 -63.18 ;
      RECT 188.27 -110.99 188.6 -110.66 ;
      RECT 188.285 -135.28 188.585 -110.66 ;
      RECT 188.27 -85.045 188.6 -84.715 ;
      RECT 188.285 -100.015 188.585 -84.715 ;
      RECT 188.27 -100.015 188.6 -99.685 ;
      RECT 188.285 -80.82 188.585 -45.52 ;
      RECT 188.27 -45.895 188.6 -45.565 ;
      RECT 188.27 -80.82 188.6 -80.49 ;
      RECT 180.115 -84.585 180.445 -84.255 ;
      RECT 180.13 -100.015 180.43 -84.255 ;
      RECT 180.115 -100.015 180.445 -99.685 ;
      RECT 180.13 -80.8 180.43 -45.52 ;
      RECT 180.115 -47.495 180.445 -47.165 ;
      RECT 180.115 -80.39 180.445 -80.06 ;
      RECT 179.515 -123.905 179.815 -54.615 ;
      RECT 179.5 -54.99 179.83 -54.66 ;
      RECT 179.5 -68.17 179.83 -67.84 ;
      RECT 179.5 -123.905 179.83 -123.575 ;
      RECT 178.9 -63.51 179.2 -55.245 ;
      RECT 178.885 -55.62 179.215 -55.29 ;
      RECT 178.885 -63.51 179.215 -63.18 ;
      RECT 178.27 -110.99 178.6 -110.66 ;
      RECT 178.285 -135.28 178.585 -110.66 ;
      RECT 178.27 -85.045 178.6 -84.715 ;
      RECT 178.285 -100.015 178.585 -84.715 ;
      RECT 178.27 -100.015 178.6 -99.685 ;
      RECT 178.285 -80.82 178.585 -45.52 ;
      RECT 178.27 -45.895 178.6 -45.565 ;
      RECT 178.27 -80.82 178.6 -80.49 ;
      RECT 173.245 -116.38 173.575 -116.05 ;
      RECT 173.26 -128.01 173.56 -116.05 ;
      RECT 173.245 -123.62 173.575 -123.29 ;
      RECT 173.245 -127.965 173.575 -127.635 ;
      RECT 172.615 -122.82 172.945 -122.49 ;
      RECT 172.63 -135.28 172.93 -122.49 ;
      RECT 172 -117.18 172.33 -116.85 ;
      RECT 172.015 -135.28 172.315 -116.85 ;
      RECT 170.115 -84.585 170.445 -84.255 ;
      RECT 170.13 -100.015 170.43 -84.255 ;
      RECT 170.115 -100.015 170.445 -99.685 ;
      RECT 170.13 -80.8 170.43 -45.52 ;
      RECT 170.115 -47.495 170.445 -47.165 ;
      RECT 170.115 -80.39 170.445 -80.06 ;
      RECT 169.515 -115.895 169.815 -54.615 ;
      RECT 169.5 -54.99 169.83 -54.66 ;
      RECT 169.5 -68.17 169.83 -67.84 ;
      RECT 169.5 -115.895 169.83 -115.565 ;
      RECT 168.9 -63.51 169.2 -55.245 ;
      RECT 168.885 -55.62 169.215 -55.29 ;
      RECT 168.885 -63.51 169.215 -63.18 ;
      RECT 168.27 -110.99 168.6 -110.66 ;
      RECT 168.285 -135.28 168.585 -110.66 ;
      RECT 168.27 -85.045 168.6 -84.715 ;
      RECT 168.285 -100.015 168.585 -84.715 ;
      RECT 168.27 -100.015 168.6 -99.685 ;
      RECT 168.285 -80.82 168.585 -45.52 ;
      RECT 168.27 -45.895 168.6 -45.565 ;
      RECT 168.27 -80.82 168.6 -80.49 ;
      RECT 160.115 -84.585 160.445 -84.255 ;
      RECT 160.13 -100.015 160.43 -84.255 ;
      RECT 160.115 -100.015 160.445 -99.685 ;
      RECT 160.13 -80.8 160.43 -45.52 ;
      RECT 160.115 -47.495 160.445 -47.165 ;
      RECT 160.115 -80.39 160.445 -80.06 ;
      RECT 159.515 -123.905 159.815 -54.615 ;
      RECT 159.5 -54.99 159.83 -54.66 ;
      RECT 159.5 -68.17 159.83 -67.84 ;
      RECT 159.5 -123.905 159.83 -123.575 ;
      RECT 158.9 -63.51 159.2 -55.245 ;
      RECT 158.885 -55.62 159.215 -55.29 ;
      RECT 158.885 -63.51 159.215 -63.18 ;
      RECT 158.27 -110.99 158.6 -110.66 ;
      RECT 158.285 -135.28 158.585 -110.66 ;
      RECT 158.27 -85.045 158.6 -84.715 ;
      RECT 158.285 -100.015 158.585 -84.715 ;
      RECT 158.27 -100.015 158.6 -99.685 ;
      RECT 158.285 -80.82 158.585 -45.52 ;
      RECT 158.27 -45.895 158.6 -45.565 ;
      RECT 158.27 -80.82 158.6 -80.49 ;
      RECT 153.245 -116.38 153.575 -116.05 ;
      RECT 153.26 -128.01 153.56 -116.05 ;
      RECT 153.245 -123.62 153.575 -123.29 ;
      RECT 153.245 -127.965 153.575 -127.635 ;
      RECT 152.615 -122.82 152.945 -122.49 ;
      RECT 152.63 -135.28 152.93 -122.49 ;
      RECT 152 -117.18 152.33 -116.85 ;
      RECT 152.015 -135.28 152.315 -116.85 ;
      RECT 150.115 -84.585 150.445 -84.255 ;
      RECT 150.13 -100.015 150.43 -84.255 ;
      RECT 150.115 -100.015 150.445 -99.685 ;
      RECT 150.13 -80.8 150.43 -45.52 ;
      RECT 150.115 -47.495 150.445 -47.165 ;
      RECT 150.115 -80.39 150.445 -80.06 ;
      RECT 149.515 -115.895 149.815 -54.615 ;
      RECT 149.5 -54.99 149.83 -54.66 ;
      RECT 149.5 -68.17 149.83 -67.84 ;
      RECT 149.5 -115.895 149.83 -115.565 ;
      RECT 148.9 -63.51 149.2 -55.245 ;
      RECT 148.885 -55.62 149.215 -55.29 ;
      RECT 148.885 -63.51 149.215 -63.18 ;
      RECT 148.27 -110.99 148.6 -110.66 ;
      RECT 148.285 -135.28 148.585 -110.66 ;
      RECT 148.27 -85.045 148.6 -84.715 ;
      RECT 148.285 -100.015 148.585 -84.715 ;
      RECT 148.27 -100.015 148.6 -99.685 ;
      RECT 148.285 -80.82 148.585 -45.52 ;
      RECT 148.27 -45.895 148.6 -45.565 ;
      RECT 148.27 -80.82 148.6 -80.49 ;
      RECT 140.115 -84.585 140.445 -84.255 ;
      RECT 140.13 -100.015 140.43 -84.255 ;
      RECT 140.115 -100.015 140.445 -99.685 ;
      RECT 140.13 -80.8 140.43 -45.52 ;
      RECT 140.115 -47.495 140.445 -47.165 ;
      RECT 140.115 -80.39 140.445 -80.06 ;
      RECT 139.515 -123.905 139.815 -54.615 ;
      RECT 139.5 -54.99 139.83 -54.66 ;
      RECT 139.5 -68.17 139.83 -67.84 ;
      RECT 139.5 -123.905 139.83 -123.575 ;
      RECT 138.9 -63.51 139.2 -55.245 ;
      RECT 138.885 -55.62 139.215 -55.29 ;
      RECT 138.885 -63.51 139.215 -63.18 ;
      RECT 138.27 -110.99 138.6 -110.66 ;
      RECT 138.285 -135.28 138.585 -110.66 ;
      RECT 138.27 -85.045 138.6 -84.715 ;
      RECT 138.285 -100.015 138.585 -84.715 ;
      RECT 138.27 -100.015 138.6 -99.685 ;
      RECT 138.285 -80.82 138.585 -45.52 ;
      RECT 138.27 -45.895 138.6 -45.565 ;
      RECT 138.27 -80.82 138.6 -80.49 ;
      RECT 133.245 -116.38 133.575 -116.05 ;
      RECT 133.26 -128.01 133.56 -116.05 ;
      RECT 133.245 -123.62 133.575 -123.29 ;
      RECT 133.245 -127.965 133.575 -127.635 ;
      RECT 132.615 -122.82 132.945 -122.49 ;
      RECT 132.63 -135.28 132.93 -122.49 ;
      RECT 132 -117.18 132.33 -116.85 ;
      RECT 132.015 -135.28 132.315 -116.85 ;
      RECT 130.115 -84.585 130.445 -84.255 ;
      RECT 130.13 -100.015 130.43 -84.255 ;
      RECT 130.115 -100.015 130.445 -99.685 ;
      RECT 130.13 -80.8 130.43 -45.52 ;
      RECT 130.115 -47.495 130.445 -47.165 ;
      RECT 130.115 -80.39 130.445 -80.06 ;
      RECT 129.515 -115.895 129.815 -54.615 ;
      RECT 129.5 -54.99 129.83 -54.66 ;
      RECT 129.5 -68.17 129.83 -67.84 ;
      RECT 129.5 -115.895 129.83 -115.565 ;
      RECT 128.9 -63.51 129.2 -55.245 ;
      RECT 128.885 -55.62 129.215 -55.29 ;
      RECT 128.885 -63.51 129.215 -63.18 ;
      RECT 128.27 -110.99 128.6 -110.66 ;
      RECT 128.285 -135.28 128.585 -110.66 ;
      RECT 128.27 -85.045 128.6 -84.715 ;
      RECT 128.285 -100.015 128.585 -84.715 ;
      RECT 128.27 -100.015 128.6 -99.685 ;
      RECT 128.285 -80.82 128.585 -45.52 ;
      RECT 128.27 -45.895 128.6 -45.565 ;
      RECT 128.27 -80.82 128.6 -80.49 ;
      RECT 120.115 -84.585 120.445 -84.255 ;
      RECT 120.13 -100.015 120.43 -84.255 ;
      RECT 120.115 -100.015 120.445 -99.685 ;
      RECT 120.13 -80.8 120.43 -45.52 ;
      RECT 120.115 -47.495 120.445 -47.165 ;
      RECT 120.115 -80.39 120.445 -80.06 ;
      RECT 119.515 -123.905 119.815 -54.615 ;
      RECT 119.5 -54.99 119.83 -54.66 ;
      RECT 119.5 -68.17 119.83 -67.84 ;
      RECT 119.5 -123.905 119.83 -123.575 ;
      RECT 118.9 -63.51 119.2 -55.245 ;
      RECT 118.885 -55.62 119.215 -55.29 ;
      RECT 118.885 -63.51 119.215 -63.18 ;
      RECT 118.27 -110.99 118.6 -110.66 ;
      RECT 118.285 -135.28 118.585 -110.66 ;
      RECT 118.27 -85.045 118.6 -84.715 ;
      RECT 118.285 -100.015 118.585 -84.715 ;
      RECT 118.27 -100.015 118.6 -99.685 ;
      RECT 118.285 -80.82 118.585 -45.52 ;
      RECT 118.27 -45.895 118.6 -45.565 ;
      RECT 118.27 -80.82 118.6 -80.49 ;
      RECT 113.245 -116.38 113.575 -116.05 ;
      RECT 113.26 -128.01 113.56 -116.05 ;
      RECT 113.245 -123.62 113.575 -123.29 ;
      RECT 113.245 -127.965 113.575 -127.635 ;
      RECT 112.615 -122.82 112.945 -122.49 ;
      RECT 112.63 -135.28 112.93 -122.49 ;
      RECT 112 -117.18 112.33 -116.85 ;
      RECT 112.015 -135.28 112.315 -116.85 ;
      RECT 110.115 -84.585 110.445 -84.255 ;
      RECT 110.13 -100.015 110.43 -84.255 ;
      RECT 110.115 -100.015 110.445 -99.685 ;
      RECT 110.13 -80.8 110.43 -45.52 ;
      RECT 110.115 -47.495 110.445 -47.165 ;
      RECT 110.115 -80.39 110.445 -80.06 ;
      RECT 109.515 -115.895 109.815 -54.615 ;
      RECT 109.5 -54.99 109.83 -54.66 ;
      RECT 109.5 -68.17 109.83 -67.84 ;
      RECT 109.5 -115.895 109.83 -115.565 ;
      RECT 108.9 -63.51 109.2 -55.245 ;
      RECT 108.885 -55.62 109.215 -55.29 ;
      RECT 108.885 -63.51 109.215 -63.18 ;
      RECT 108.27 -110.99 108.6 -110.66 ;
      RECT 108.285 -135.28 108.585 -110.66 ;
      RECT 108.27 -85.045 108.6 -84.715 ;
      RECT 108.285 -100.015 108.585 -84.715 ;
      RECT 108.27 -100.015 108.6 -99.685 ;
      RECT 108.285 -80.82 108.585 -45.52 ;
      RECT 108.27 -45.895 108.6 -45.565 ;
      RECT 108.27 -80.82 108.6 -80.49 ;
      RECT 100.115 -84.585 100.445 -84.255 ;
      RECT 100.13 -100.015 100.43 -84.255 ;
      RECT 100.115 -100.015 100.445 -99.685 ;
      RECT 100.13 -80.8 100.43 -45.52 ;
      RECT 100.115 -47.495 100.445 -47.165 ;
      RECT 100.115 -80.39 100.445 -80.06 ;
      RECT 99.515 -123.905 99.815 -54.615 ;
      RECT 99.5 -54.99 99.83 -54.66 ;
      RECT 99.5 -68.17 99.83 -67.84 ;
      RECT 99.5 -123.905 99.83 -123.575 ;
      RECT 98.9 -63.51 99.2 -55.245 ;
      RECT 98.885 -55.62 99.215 -55.29 ;
      RECT 98.885 -63.51 99.215 -63.18 ;
      RECT 98.27 -110.99 98.6 -110.66 ;
      RECT 98.285 -135.28 98.585 -110.66 ;
      RECT 98.27 -85.045 98.6 -84.715 ;
      RECT 98.285 -100.015 98.585 -84.715 ;
      RECT 98.27 -100.015 98.6 -99.685 ;
      RECT 98.285 -80.82 98.585 -45.52 ;
      RECT 98.27 -45.895 98.6 -45.565 ;
      RECT 98.27 -80.82 98.6 -80.49 ;
      RECT 93.245 -116.38 93.575 -116.05 ;
      RECT 93.26 -128.01 93.56 -116.05 ;
      RECT 93.245 -123.62 93.575 -123.29 ;
      RECT 93.245 -127.965 93.575 -127.635 ;
      RECT 92.615 -122.82 92.945 -122.49 ;
      RECT 92.63 -135.28 92.93 -122.49 ;
      RECT 92 -117.18 92.33 -116.85 ;
      RECT 92.015 -135.28 92.315 -116.85 ;
      RECT 90.115 -84.585 90.445 -84.255 ;
      RECT 90.13 -100.015 90.43 -84.255 ;
      RECT 90.115 -100.015 90.445 -99.685 ;
      RECT 90.13 -80.8 90.43 -45.52 ;
      RECT 90.115 -47.495 90.445 -47.165 ;
      RECT 90.115 -80.39 90.445 -80.06 ;
      RECT 89.515 -115.895 89.815 -54.615 ;
      RECT 89.5 -54.99 89.83 -54.66 ;
      RECT 89.5 -68.17 89.83 -67.84 ;
      RECT 89.5 -115.895 89.83 -115.565 ;
      RECT 88.9 -63.51 89.2 -55.245 ;
      RECT 88.885 -55.62 89.215 -55.29 ;
      RECT 88.885 -63.51 89.215 -63.18 ;
      RECT 88.27 -110.99 88.6 -110.66 ;
      RECT 88.285 -135.28 88.585 -110.66 ;
      RECT 88.27 -85.045 88.6 -84.715 ;
      RECT 88.285 -100.015 88.585 -84.715 ;
      RECT 88.27 -100.015 88.6 -99.685 ;
      RECT 88.285 -80.82 88.585 -45.52 ;
      RECT 88.27 -45.895 88.6 -45.565 ;
      RECT 88.27 -80.82 88.6 -80.49 ;
      RECT 80.115 -84.585 80.445 -84.255 ;
      RECT 80.13 -100.015 80.43 -84.255 ;
      RECT 80.115 -100.015 80.445 -99.685 ;
      RECT 80.13 -80.8 80.43 -45.52 ;
      RECT 80.115 -47.495 80.445 -47.165 ;
      RECT 80.115 -80.39 80.445 -80.06 ;
      RECT 79.515 -123.905 79.815 -54.615 ;
      RECT 79.5 -54.99 79.83 -54.66 ;
      RECT 79.5 -68.17 79.83 -67.84 ;
      RECT 79.5 -123.905 79.83 -123.575 ;
      RECT 78.9 -63.51 79.2 -55.245 ;
      RECT 78.885 -55.62 79.215 -55.29 ;
      RECT 78.885 -63.51 79.215 -63.18 ;
      RECT 78.27 -110.99 78.6 -110.66 ;
      RECT 78.285 -135.28 78.585 -110.66 ;
      RECT 78.27 -85.045 78.6 -84.715 ;
      RECT 78.285 -100.015 78.585 -84.715 ;
      RECT 78.27 -100.015 78.6 -99.685 ;
      RECT 78.285 -80.82 78.585 -45.52 ;
      RECT 78.27 -45.895 78.6 -45.565 ;
      RECT 78.27 -80.82 78.6 -80.49 ;
      RECT 73.245 -116.38 73.575 -116.05 ;
      RECT 73.26 -128.01 73.56 -116.05 ;
      RECT 73.245 -123.62 73.575 -123.29 ;
      RECT 73.245 -127.965 73.575 -127.635 ;
      RECT 72.615 -122.82 72.945 -122.49 ;
      RECT 72.63 -135.28 72.93 -122.49 ;
      RECT 72 -117.18 72.33 -116.85 ;
      RECT 72.015 -135.28 72.315 -116.85 ;
      RECT 70.115 -84.585 70.445 -84.255 ;
      RECT 70.13 -100.015 70.43 -84.255 ;
      RECT 70.115 -100.015 70.445 -99.685 ;
      RECT 70.13 -80.8 70.43 -45.52 ;
      RECT 70.115 -47.495 70.445 -47.165 ;
      RECT 70.115 -80.39 70.445 -80.06 ;
      RECT 69.515 -115.895 69.815 -54.615 ;
      RECT 69.5 -54.99 69.83 -54.66 ;
      RECT 69.5 -68.17 69.83 -67.84 ;
      RECT 69.5 -115.895 69.83 -115.565 ;
      RECT 68.9 -63.51 69.2 -55.245 ;
      RECT 68.885 -55.62 69.215 -55.29 ;
      RECT 68.885 -63.51 69.215 -63.18 ;
      RECT 68.27 -110.99 68.6 -110.66 ;
      RECT 68.285 -135.28 68.585 -110.66 ;
      RECT 68.27 -85.045 68.6 -84.715 ;
      RECT 68.285 -100.015 68.585 -84.715 ;
      RECT 68.27 -100.015 68.6 -99.685 ;
      RECT 68.285 -80.82 68.585 -45.52 ;
      RECT 68.27 -45.895 68.6 -45.565 ;
      RECT 68.27 -80.82 68.6 -80.49 ;
      RECT 60.115 -84.585 60.445 -84.255 ;
      RECT 60.13 -100.015 60.43 -84.255 ;
      RECT 60.115 -100.015 60.445 -99.685 ;
      RECT 60.13 -80.8 60.43 -45.52 ;
      RECT 60.115 -47.495 60.445 -47.165 ;
      RECT 60.115 -80.39 60.445 -80.06 ;
      RECT 59.515 -123.905 59.815 -54.615 ;
      RECT 59.5 -54.99 59.83 -54.66 ;
      RECT 59.5 -68.17 59.83 -67.84 ;
      RECT 59.5 -123.905 59.83 -123.575 ;
      RECT 58.9 -63.51 59.2 -55.245 ;
      RECT 58.885 -55.62 59.215 -55.29 ;
      RECT 58.885 -63.51 59.215 -63.18 ;
      RECT 58.27 -110.99 58.6 -110.66 ;
      RECT 58.285 -135.28 58.585 -110.66 ;
      RECT 58.27 -85.045 58.6 -84.715 ;
      RECT 58.285 -100.015 58.585 -84.715 ;
      RECT 58.27 -100.015 58.6 -99.685 ;
      RECT 58.285 -80.82 58.585 -45.52 ;
      RECT 58.27 -45.895 58.6 -45.565 ;
      RECT 58.27 -80.82 58.6 -80.49 ;
      RECT 53.245 -116.38 53.575 -116.05 ;
      RECT 53.26 -128.01 53.56 -116.05 ;
      RECT 53.245 -123.62 53.575 -123.29 ;
      RECT 53.245 -127.965 53.575 -127.635 ;
      RECT 52.615 -122.82 52.945 -122.49 ;
      RECT 52.63 -135.28 52.93 -122.49 ;
      RECT 52 -117.18 52.33 -116.85 ;
      RECT 52.015 -135.28 52.315 -116.85 ;
      RECT 50.115 -84.585 50.445 -84.255 ;
      RECT 50.13 -100.015 50.43 -84.255 ;
      RECT 50.115 -100.015 50.445 -99.685 ;
      RECT 50.13 -80.8 50.43 -45.52 ;
      RECT 50.115 -47.495 50.445 -47.165 ;
      RECT 50.115 -80.39 50.445 -80.06 ;
      RECT 49.515 -115.895 49.815 -54.615 ;
      RECT 49.5 -54.99 49.83 -54.66 ;
      RECT 49.5 -68.17 49.83 -67.84 ;
      RECT 49.5 -115.895 49.83 -115.565 ;
      RECT 48.9 -63.51 49.2 -55.245 ;
      RECT 48.885 -55.62 49.215 -55.29 ;
      RECT 48.885 -63.51 49.215 -63.18 ;
      RECT 48.27 -110.99 48.6 -110.66 ;
      RECT 48.285 -135.28 48.585 -110.66 ;
      RECT 48.27 -85.045 48.6 -84.715 ;
      RECT 48.285 -100.015 48.585 -84.715 ;
      RECT 48.27 -100.015 48.6 -99.685 ;
      RECT 48.285 -80.82 48.585 -45.52 ;
      RECT 48.27 -45.895 48.6 -45.565 ;
      RECT 48.27 -80.82 48.6 -80.49 ;
      RECT 40.115 -84.585 40.445 -84.255 ;
      RECT 40.13 -100.015 40.43 -84.255 ;
      RECT 40.115 -100.015 40.445 -99.685 ;
      RECT 40.13 -80.8 40.43 -45.52 ;
      RECT 40.115 -47.495 40.445 -47.165 ;
      RECT 40.115 -80.39 40.445 -80.06 ;
      RECT 39.515 -123.905 39.815 -54.615 ;
      RECT 39.5 -54.99 39.83 -54.66 ;
      RECT 39.5 -68.17 39.83 -67.84 ;
      RECT 39.5 -123.905 39.83 -123.575 ;
      RECT 38.9 -63.51 39.2 -55.245 ;
      RECT 38.885 -55.62 39.215 -55.29 ;
      RECT 38.885 -63.51 39.215 -63.18 ;
      RECT 38.27 -110.99 38.6 -110.66 ;
      RECT 38.285 -135.28 38.585 -110.66 ;
      RECT 38.27 -85.045 38.6 -84.715 ;
      RECT 38.285 -100.015 38.585 -84.715 ;
      RECT 38.27 -100.015 38.6 -99.685 ;
      RECT 38.285 -80.82 38.585 -45.52 ;
      RECT 38.27 -45.895 38.6 -45.565 ;
      RECT 38.27 -80.82 38.6 -80.49 ;
      RECT 33.245 -116.38 33.575 -116.05 ;
      RECT 33.26 -128.01 33.56 -116.05 ;
      RECT 33.245 -123.62 33.575 -123.29 ;
      RECT 33.245 -127.965 33.575 -127.635 ;
      RECT 32.615 -122.82 32.945 -122.49 ;
      RECT 32.63 -135.28 32.93 -122.49 ;
      RECT 32 -117.18 32.33 -116.85 ;
      RECT 32.015 -135.28 32.315 -116.85 ;
      RECT 30.115 -84.585 30.445 -84.255 ;
      RECT 30.13 -100.015 30.43 -84.255 ;
      RECT 30.115 -100.015 30.445 -99.685 ;
      RECT 30.13 -80.8 30.43 -45.52 ;
      RECT 30.115 -47.495 30.445 -47.165 ;
      RECT 30.115 -80.39 30.445 -80.06 ;
      RECT 29.515 -115.895 29.815 -54.615 ;
      RECT 29.5 -54.99 29.83 -54.66 ;
      RECT 29.5 -68.17 29.83 -67.84 ;
      RECT 29.5 -115.895 29.83 -115.565 ;
      RECT 28.9 -63.51 29.2 -55.245 ;
      RECT 28.885 -55.62 29.215 -55.29 ;
      RECT 28.885 -63.51 29.215 -63.18 ;
      RECT 28.27 -110.99 28.6 -110.66 ;
      RECT 28.285 -135.28 28.585 -110.66 ;
      RECT 28.27 -85.045 28.6 -84.715 ;
      RECT 28.285 -100.015 28.585 -84.715 ;
      RECT 28.27 -100.015 28.6 -99.685 ;
      RECT 28.285 -80.82 28.585 -45.52 ;
      RECT 28.27 -45.895 28.6 -45.565 ;
      RECT 28.27 -80.82 28.6 -80.49 ;
      RECT 20.115 -84.585 20.445 -84.255 ;
      RECT 20.13 -100.015 20.43 -84.255 ;
      RECT 20.115 -100.015 20.445 -99.685 ;
      RECT 20.13 -80.8 20.43 -45.52 ;
      RECT 20.115 -47.495 20.445 -47.165 ;
      RECT 20.115 -80.39 20.445 -80.06 ;
      RECT 19.515 -123.905 19.815 -54.615 ;
      RECT 19.5 -54.99 19.83 -54.66 ;
      RECT 19.5 -68.17 19.83 -67.84 ;
      RECT 19.5 -123.905 19.83 -123.575 ;
      RECT 18.9 -63.51 19.2 -55.245 ;
      RECT 18.885 -55.62 19.215 -55.29 ;
      RECT 18.885 -63.51 19.215 -63.18 ;
      RECT 18.27 -110.99 18.6 -110.66 ;
      RECT 18.285 -135.28 18.585 -110.66 ;
      RECT 18.27 -85.045 18.6 -84.715 ;
      RECT 18.285 -100.015 18.585 -84.715 ;
      RECT 18.27 -100.015 18.6 -99.685 ;
      RECT 18.285 -80.82 18.585 -45.52 ;
      RECT 18.27 -45.895 18.6 -45.565 ;
      RECT 18.27 -80.82 18.6 -80.49 ;
      RECT 13.245 -116.38 13.575 -116.05 ;
      RECT 13.26 -128.01 13.56 -116.05 ;
      RECT 13.245 -123.62 13.575 -123.29 ;
      RECT 13.245 -127.965 13.575 -127.635 ;
      RECT 12.615 -122.82 12.945 -122.49 ;
      RECT 12.63 -135.28 12.93 -122.49 ;
      RECT 12 -117.18 12.33 -116.85 ;
      RECT 12.015 -135.28 12.315 -116.85 ;
      RECT 10.115 -84.585 10.445 -84.255 ;
      RECT 10.13 -100.015 10.43 -84.255 ;
      RECT 10.115 -100.015 10.445 -99.685 ;
      RECT 10.13 -80.8 10.43 -45.52 ;
      RECT 10.115 -47.495 10.445 -47.165 ;
      RECT 10.115 -80.39 10.445 -80.06 ;
      RECT 9.515 -115.895 9.815 -54.615 ;
      RECT 9.5 -54.99 9.83 -54.66 ;
      RECT 9.5 -68.17 9.83 -67.84 ;
      RECT 9.5 -115.895 9.83 -115.565 ;
      RECT 8.9 -63.51 9.2 -55.245 ;
      RECT 8.885 -55.62 9.215 -55.29 ;
      RECT 8.885 -63.51 9.215 -63.18 ;
      RECT 8.27 -110.99 8.6 -110.66 ;
      RECT 8.285 -135.28 8.585 -110.66 ;
      RECT 8.27 -85.045 8.6 -84.715 ;
      RECT 8.285 -100.015 8.585 -84.715 ;
      RECT 8.27 -100.015 8.6 -99.685 ;
      RECT 8.285 -80.82 8.585 -45.52 ;
      RECT 8.27 -45.895 8.6 -45.565 ;
      RECT 8.27 -80.82 8.6 -80.49 ;
      RECT 6.005 -74.805 6.335 -74.475 ;
      RECT 6.02 -79.7 6.32 -74.475 ;
      RECT 6.005 -79.7 6.335 -79.37 ;
      RECT -5.91 -100.135 -5.58 -99.805 ;
      RECT -5.895 -114.57 -5.595 -99.805 ;
      RECT -5.91 -114.57 -5.58 -114.24 ;
      RECT -9.505 -114.125 -9.175 -113.795 ;
      RECT -9.49 -128.01 -9.19 -113.795 ;
      RECT -9.505 -127.965 -9.175 -127.635 ;
      RECT -10.34 -36.06 -10.01 -35.73 ;
      RECT -10.325 -81.49 -10.025 -35.73 ;
      RECT -10.34 -81.49 -10.01 -81.16 ;
      RECT -10.635 -114.925 -10.305 -114.595 ;
      RECT -10.62 -135.28 -10.32 -114.595 ;
      RECT -11.75 -104.9 -11.42 -104.57 ;
      RECT -11.735 -114.57 -11.435 -104.57 ;
      RECT -11.75 -114.57 -11.42 -114.24 ;
      RECT -12.385 -104.4 -12.055 -104.07 ;
      RECT -12.37 -115.325 -12.07 -104.07 ;
      RECT -12.385 -115.325 -12.055 -114.995 ;
      RECT -15.345 -114.125 -15.015 -113.795 ;
      RECT -15.33 -128.01 -15.03 -113.795 ;
      RECT -15.345 -127.965 -15.015 -127.635 ;
      RECT -16.475 -114.925 -16.145 -114.595 ;
      RECT -16.46 -135.28 -16.16 -114.595 ;
      RECT -17.59 -105.9 -17.26 -105.57 ;
      RECT -17.575 -114.57 -17.275 -105.57 ;
      RECT -17.59 -114.57 -17.26 -114.24 ;
      RECT -18.225 -105.4 -17.895 -105.07 ;
      RECT -18.21 -115.325 -17.91 -105.07 ;
      RECT -18.225 -115.325 -17.895 -114.995 ;
      RECT -21.185 -114.125 -20.855 -113.795 ;
      RECT -21.17 -128.01 -20.87 -113.795 ;
      RECT -21.185 -127.965 -20.855 -127.635 ;
      RECT -22.315 -114.925 -21.985 -114.595 ;
      RECT -22.3 -135.28 -22 -114.595 ;
      RECT -23.43 -106.9 -23.1 -106.57 ;
      RECT -23.415 -114.57 -23.115 -106.57 ;
      RECT -23.43 -114.57 -23.1 -114.24 ;
      RECT -24.065 -106.4 -23.735 -106.07 ;
      RECT -24.05 -115.325 -23.75 -106.07 ;
      RECT -24.065 -115.325 -23.735 -114.995 ;
      RECT -27.025 -114.125 -26.695 -113.795 ;
      RECT -27.01 -128.01 -26.71 -113.795 ;
      RECT -27.025 -127.965 -26.695 -127.635 ;
      RECT -28.155 -114.925 -27.825 -114.595 ;
      RECT -28.14 -135.28 -27.84 -114.595 ;
      RECT -29.27 -107.9 -28.94 -107.57 ;
      RECT -29.255 -114.57 -28.955 -107.57 ;
      RECT -29.27 -114.57 -28.94 -114.24 ;
      RECT -29.905 -107.4 -29.575 -107.07 ;
      RECT -29.89 -115.325 -29.59 -107.07 ;
      RECT -29.905 -115.325 -29.575 -114.995 ;
      RECT -32.865 -114.125 -32.535 -113.795 ;
      RECT -32.85 -128.01 -32.55 -113.795 ;
      RECT -32.865 -127.965 -32.535 -127.635 ;
      RECT -33.995 -114.925 -33.665 -114.595 ;
      RECT -33.98 -135.28 -33.68 -114.595 ;
      RECT -35.11 -108.9 -34.78 -108.57 ;
      RECT -35.095 -114.57 -34.795 -108.57 ;
      RECT -35.11 -114.57 -34.78 -114.24 ;
      RECT -35.745 -108.4 -35.415 -108.07 ;
      RECT -35.73 -115.325 -35.43 -108.07 ;
      RECT -35.745 -115.325 -35.415 -114.995 ;
      RECT -38.705 -114.125 -38.375 -113.795 ;
      RECT -38.69 -128.01 -38.39 -113.795 ;
      RECT -38.705 -127.965 -38.375 -127.635 ;
      RECT -39.835 -114.925 -39.505 -114.595 ;
      RECT -39.82 -135.28 -39.52 -114.595 ;
      RECT -40.95 -109.9 -40.62 -109.57 ;
      RECT -40.935 -114.57 -40.635 -109.57 ;
      RECT -40.95 -114.57 -40.62 -114.24 ;
      RECT -41.585 -109.4 -41.255 -109.07 ;
      RECT -41.57 -115.325 -41.27 -109.07 ;
      RECT -41.585 -115.325 -41.255 -114.995 ;
      RECT -44.545 -114.125 -44.215 -113.795 ;
      RECT -44.53 -128.01 -44.23 -113.795 ;
      RECT -44.545 -127.965 -44.215 -127.635 ;
      RECT -45.675 -114.925 -45.345 -114.595 ;
      RECT -45.66 -135.28 -45.36 -114.595 ;
      RECT -46.54 -128.01 -46.14 -101.445 ;
      RECT -46.68 -135.16 -46.26 -127.59 ;
  END
END sramgen_sram_64x32m4w32_replica_v1

END LIBRARY
