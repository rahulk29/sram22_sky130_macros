VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_256x32m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_256x32m4w8   ;
    SIZE 422.880 BY 291.640 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 214.630 0.000 214.770 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 220.730 0.000 220.870 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 226.830 0.000 226.970 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 232.930 0.000 233.070 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 239.030 0.000 239.170 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 245.130 0.000 245.270 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 251.230 0.000 251.370 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 257.330 0.000 257.470 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 263.430 0.000 263.570 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 269.530 0.000 269.670 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 275.630 0.000 275.770 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 281.730 0.000 281.870 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 287.830 0.000 287.970 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 293.930 0.000 294.070 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 300.030 0.000 300.170 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 306.130 0.000 306.270 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 312.230 0.000 312.370 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 318.330 0.000 318.470 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 324.430 0.000 324.570 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.530 0.000 330.670 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.630 0.000 336.770 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 342.730 0.000 342.870 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 348.830 0.000 348.970 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 354.930 0.000 355.070 0.140 ; 
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 361.030 0.000 361.170 0.140 ; 
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 367.130 0.000 367.270 0.140 ; 
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 373.230 0.000 373.370 0.140 ; 
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 379.330 0.000 379.470 0.140 ; 
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 385.430 0.000 385.570 0.140 ; 
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 391.530 0.000 391.670 0.140 ; 
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 397.630 0.000 397.770 0.140 ; 
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 403.730 0.000 403.870 0.140 ; 
        END 
    END dout[31] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 214.210 0.000 214.350 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 220.310 0.000 220.450 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 226.410 0.000 226.550 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 232.510 0.000 232.650 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 238.610 0.000 238.750 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 244.710 0.000 244.850 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 250.810 0.000 250.950 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 256.910 0.000 257.050 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 263.010 0.000 263.150 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 269.110 0.000 269.250 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 275.210 0.000 275.350 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 281.310 0.000 281.450 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 287.410 0.000 287.550 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 293.510 0.000 293.650 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 299.610 0.000 299.750 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 305.710 0.000 305.850 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 311.810 0.000 311.950 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 317.910 0.000 318.050 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 324.010 0.000 324.150 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.110 0.000 330.250 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.210 0.000 336.350 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 342.310 0.000 342.450 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 348.410 0.000 348.550 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 354.510 0.000 354.650 0.140 ; 
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 360.610 0.000 360.750 0.140 ; 
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 366.710 0.000 366.850 0.140 ; 
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 372.810 0.000 372.950 0.140 ; 
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 378.910 0.000 379.050 0.140 ; 
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 385.010 0.000 385.150 0.140 ; 
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 391.110 0.000 391.250 0.140 ; 
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 397.210 0.000 397.350 0.140 ; 
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.838500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 403.310 0.000 403.450 0.140 ; 
        END 
    END din[31] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 213.860 0.000 214.000 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 262.660 0.000 262.800 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 311.460 0.000 311.600 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.648900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 360.260 0.000 360.400 0.140 ; 
        END 
    END wmask[3] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 172.520 0.000 172.840 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 166.400 0.000 166.720 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 160.280 0.000 160.600 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 154.160 0.000 154.480 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 148.040 0.000 148.360 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 141.920 0.000 142.240 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 135.800 0.000 136.120 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 129.680 0.000 130.000 0.320 ; 
        END 
    END addr[7] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 184.760 0.000 185.080 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 4.725500 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 178.640 0.000 178.960 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 22.320000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 187.480 0.000 187.800 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 26.226000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 188.160 0.000 188.480 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 213.640 6.240 ; 
                RECT 404.400 5.920 422.720 6.240 ; 
                RECT 0.160 7.280 422.720 7.600 ; 
                RECT 0.160 8.640 422.720 8.960 ; 
                RECT 0.160 10.000 187.120 10.320 ; 
                RECT 360.880 10.000 422.720 10.320 ; 
                RECT 0.160 11.360 203.440 11.680 ; 
                RECT 413.240 11.360 422.720 11.680 ; 
                RECT 0.160 12.720 203.440 13.040 ; 
                RECT 413.240 12.720 422.720 13.040 ; 
                RECT 0.160 14.080 203.440 14.400 ; 
                RECT 413.240 14.080 422.720 14.400 ; 
                RECT 0.160 15.440 203.440 15.760 ; 
                RECT 413.240 15.440 422.720 15.760 ; 
                RECT 0.160 16.800 125.920 17.120 ; 
                RECT 188.840 16.800 203.440 17.120 ; 
                RECT 413.240 16.800 422.720 17.120 ; 
                RECT 0.160 18.160 203.440 18.480 ; 
                RECT 413.240 18.160 422.720 18.480 ; 
                RECT 0.160 19.520 203.440 19.840 ; 
                RECT 413.240 19.520 422.720 19.840 ; 
                RECT 0.160 20.880 125.920 21.200 ; 
                RECT 188.160 20.880 203.440 21.200 ; 
                RECT 413.240 20.880 422.720 21.200 ; 
                RECT 0.160 22.240 203.440 22.560 ; 
                RECT 413.240 22.240 422.720 22.560 ; 
                RECT 0.160 23.600 203.440 23.920 ; 
                RECT 413.240 23.600 422.720 23.920 ; 
                RECT 0.160 24.960 203.440 25.280 ; 
                RECT 413.240 24.960 422.720 25.280 ; 
                RECT 0.160 26.320 203.440 26.640 ; 
                RECT 413.240 26.320 422.720 26.640 ; 
                RECT 0.160 27.680 202.760 28.000 ; 
                RECT 413.240 27.680 422.720 28.000 ; 
                RECT 0.160 29.040 203.440 29.360 ; 
                RECT 413.240 29.040 422.720 29.360 ; 
                RECT 0.160 30.400 203.440 30.720 ; 
                RECT 413.240 30.400 422.720 30.720 ; 
                RECT 0.160 31.760 203.440 32.080 ; 
                RECT 413.240 31.760 422.720 32.080 ; 
                RECT 0.160 33.120 203.440 33.440 ; 
                RECT 413.240 33.120 422.720 33.440 ; 
                RECT 0.160 34.480 203.440 34.800 ; 
                RECT 413.240 34.480 422.720 34.800 ; 
                RECT 0.160 35.840 203.440 36.160 ; 
                RECT 413.240 35.840 422.720 36.160 ; 
                RECT 0.160 37.200 127.960 37.520 ; 
                RECT 165.720 37.200 203.440 37.520 ; 
                RECT 413.240 37.200 422.720 37.520 ; 
                RECT 0.160 38.560 126.600 38.880 ; 
                RECT 171.840 38.560 203.440 38.880 ; 
                RECT 413.240 38.560 422.720 38.880 ; 
                RECT 0.160 39.920 106.880 40.240 ; 
                RECT 188.840 39.920 203.440 40.240 ; 
                RECT 413.240 39.920 422.720 40.240 ; 
                RECT 0.160 41.280 106.200 41.600 ; 
                RECT 184.760 41.280 203.440 41.600 ; 
                RECT 413.240 41.280 422.720 41.600 ; 
                RECT 0.160 42.640 203.440 42.960 ; 
                RECT 413.240 42.640 422.720 42.960 ; 
                RECT 0.160 44.000 203.440 44.320 ; 
                RECT 413.240 44.000 422.720 44.320 ; 
                RECT 0.160 45.360 203.440 45.680 ; 
                RECT 413.240 45.360 422.720 45.680 ; 
                RECT 0.160 46.720 203.440 47.040 ; 
                RECT 413.240 46.720 422.720 47.040 ; 
                RECT 0.160 48.080 102.800 48.400 ; 
                RECT 113.360 48.080 179.640 48.400 ; 
                RECT 186.120 48.080 203.440 48.400 ; 
                RECT 413.240 48.080 422.720 48.400 ; 
                RECT 0.160 49.440 104.160 49.760 ; 
                RECT 109.960 49.440 117.080 49.760 ; 
                RECT 120.160 49.440 179.640 49.760 ; 
                RECT 413.240 49.440 422.720 49.760 ; 
                RECT 0.160 50.800 105.520 51.120 ; 
                RECT 108.600 50.800 125.240 51.120 ; 
                RECT 176.600 50.800 179.640 51.120 ; 
                RECT 186.120 50.800 203.440 51.120 ; 
                RECT 413.240 50.800 422.720 51.120 ; 
                RECT 0.160 52.160 203.440 52.480 ; 
                RECT 413.240 52.160 422.720 52.480 ; 
                RECT 0.160 53.520 111.640 53.840 ; 
                RECT 120.160 53.520 203.440 53.840 ; 
                RECT 413.240 53.520 422.720 53.840 ; 
                RECT 0.160 54.880 104.160 55.200 ; 
                RECT 113.360 54.880 203.440 55.200 ; 
                RECT 413.240 54.880 422.720 55.200 ; 
                RECT 0.160 56.240 108.240 56.560 ; 
                RECT 112.680 56.240 203.440 56.560 ; 
                RECT 413.240 56.240 422.720 56.560 ; 
                RECT 0.160 57.600 126.600 57.920 ; 
                RECT 132.400 57.600 138.160 57.920 ; 
                RECT 186.120 57.600 203.440 57.920 ; 
                RECT 413.240 57.600 422.720 57.920 ; 
                RECT 0.160 58.960 104.160 59.280 ; 
                RECT 113.360 58.960 127.960 59.280 ; 
                RECT 131.720 58.960 138.160 59.280 ; 
                RECT 195.640 58.960 203.440 59.280 ; 
                RECT 413.240 58.960 422.720 59.280 ; 
                RECT 0.160 60.320 110.960 60.640 ; 
                RECT 119.480 60.320 138.160 60.640 ; 
                RECT 195.640 60.320 203.440 60.640 ; 
                RECT 413.240 60.320 422.720 60.640 ; 
                RECT 0.160 61.680 138.160 62.000 ; 
                RECT 194.280 61.680 203.440 62.000 ; 
                RECT 413.240 61.680 422.720 62.000 ; 
                RECT 0.160 63.040 111.640 63.360 ; 
                RECT 117.440 63.040 138.160 63.360 ; 
                RECT 195.640 63.040 203.440 63.360 ; 
                RECT 413.240 63.040 422.720 63.360 ; 
                RECT 0.160 64.400 114.360 64.720 ; 
                RECT 120.160 64.400 138.160 64.720 ; 
                RECT 195.640 64.400 203.440 64.720 ; 
                RECT 413.240 64.400 422.720 64.720 ; 
                RECT 0.160 65.760 108.240 66.080 ; 
                RECT 113.360 65.760 138.160 66.080 ; 
                RECT 194.280 65.760 203.440 66.080 ; 
                RECT 413.240 65.760 422.720 66.080 ; 
                RECT 0.160 67.120 138.160 67.440 ; 
                RECT 195.640 67.120 203.440 67.440 ; 
                RECT 413.240 67.120 422.720 67.440 ; 
                RECT 0.160 68.480 102.120 68.800 ; 
                RECT 124.920 68.480 138.160 68.800 ; 
                RECT 194.280 68.480 203.440 68.800 ; 
                RECT 413.240 68.480 422.720 68.800 ; 
                RECT 0.160 69.840 111.640 70.160 ; 
                RECT 120.160 69.840 138.160 70.160 ; 
                RECT 198.360 69.840 203.440 70.160 ; 
                RECT 413.240 69.840 422.720 70.160 ; 
                RECT 0.160 71.200 110.960 71.520 ; 
                RECT 113.360 71.200 120.480 71.520 ; 
                RECT 126.960 71.200 138.160 71.520 ; 
                RECT 198.360 71.200 203.440 71.520 ; 
                RECT 413.240 71.200 422.720 71.520 ; 
                RECT 0.160 72.560 102.800 72.880 ; 
                RECT 116.080 72.560 138.160 72.880 ; 
                RECT 186.120 72.560 203.440 72.880 ; 
                RECT 413.240 72.560 422.720 72.880 ; 
                RECT 0.160 73.920 110.960 74.240 ; 
                RECT 120.160 73.920 138.160 74.240 ; 
                RECT 197.000 73.920 203.440 74.240 ; 
                RECT 413.240 73.920 422.720 74.240 ; 
                RECT 0.160 75.280 108.920 75.600 ; 
                RECT 112.680 75.280 138.160 75.600 ; 
                RECT 186.120 75.280 203.440 75.600 ; 
                RECT 413.240 75.280 422.720 75.600 ; 
                RECT 0.160 76.640 104.160 76.960 ; 
                RECT 108.600 76.640 111.640 76.960 ; 
                RECT 120.160 76.640 138.160 76.960 ; 
                RECT 198.360 76.640 203.440 76.960 ; 
                RECT 413.240 76.640 422.720 76.960 ; 
                RECT 0.160 78.000 106.880 78.320 ; 
                RECT 110.640 78.000 138.160 78.320 ; 
                RECT 198.360 78.000 203.440 78.320 ; 
                RECT 413.240 78.000 422.720 78.320 ; 
                RECT 0.160 79.360 104.160 79.680 ; 
                RECT 107.240 79.360 138.160 79.680 ; 
                RECT 201.080 79.360 203.440 79.680 ; 
                RECT 413.240 79.360 422.720 79.680 ; 
                RECT 0.160 80.720 108.240 81.040 ; 
                RECT 113.360 80.720 138.160 81.040 ; 
                RECT 199.720 80.720 203.440 81.040 ; 
                RECT 413.240 80.720 422.720 81.040 ; 
                RECT 0.160 82.080 104.160 82.400 ; 
                RECT 118.800 82.080 138.160 82.400 ; 
                RECT 201.080 82.080 203.440 82.400 ; 
                RECT 413.240 82.080 422.720 82.400 ; 
                RECT 0.160 83.440 138.160 83.760 ; 
                RECT 186.120 83.440 203.440 83.760 ; 
                RECT 413.240 83.440 422.720 83.760 ; 
                RECT 0.160 84.800 110.960 85.120 ; 
                RECT 112.680 84.800 138.160 85.120 ; 
                RECT 201.080 84.800 203.440 85.120 ; 
                RECT 413.240 84.800 422.720 85.120 ; 
                RECT 0.160 86.160 111.640 86.480 ; 
                RECT 114.040 86.160 138.160 86.480 ; 
                RECT 201.080 86.160 203.440 86.480 ; 
                RECT 413.240 86.160 422.720 86.480 ; 
                RECT 0.160 87.520 102.800 87.840 ; 
                RECT 109.960 87.520 110.960 87.840 ; 
                RECT 112.680 87.520 138.160 87.840 ; 
                RECT 199.720 87.520 203.440 87.840 ; 
                RECT 413.240 87.520 422.720 87.840 ; 
                RECT 0.160 88.880 108.240 89.200 ; 
                RECT 120.160 88.880 138.160 89.200 ; 
                RECT 201.080 88.880 203.440 89.200 ; 
                RECT 413.240 88.880 422.720 89.200 ; 
                RECT 0.160 90.240 102.800 90.560 ; 
                RECT 113.360 90.240 138.160 90.560 ; 
                RECT 413.240 90.240 422.720 90.560 ; 
                RECT 0.160 91.600 110.960 91.920 ; 
                RECT 114.040 91.600 138.160 91.920 ; 
                RECT 413.240 91.600 422.720 91.920 ; 
                RECT 0.160 92.960 138.160 93.280 ; 
                RECT 413.240 92.960 422.720 93.280 ; 
                RECT 0.160 94.320 138.160 94.640 ; 
                RECT 413.240 94.320 422.720 94.640 ; 
                RECT 0.160 95.680 98.720 96.000 ; 
                RECT 116.080 95.680 138.160 96.000 ; 
                RECT 413.240 95.680 422.720 96.000 ; 
                RECT 0.160 97.040 138.160 97.360 ; 
                RECT 413.240 97.040 422.720 97.360 ; 
                RECT 0.160 98.400 138.160 98.720 ; 
                RECT 186.120 98.400 203.440 98.720 ; 
                RECT 413.240 98.400 422.720 98.720 ; 
                RECT 0.160 99.760 107.560 100.080 ; 
                RECT 120.160 99.760 138.160 100.080 ; 
                RECT 413.240 99.760 422.720 100.080 ; 
                RECT 0.160 101.120 114.360 101.440 ; 
                RECT 122.200 101.120 138.160 101.440 ; 
                RECT 186.120 101.120 203.440 101.440 ; 
                RECT 413.240 101.120 422.720 101.440 ; 
                RECT 0.160 102.480 203.440 102.800 ; 
                RECT 413.240 102.480 422.720 102.800 ; 
                RECT 0.160 103.840 189.840 104.160 ; 
                RECT 413.240 103.840 422.720 104.160 ; 
                RECT 0.160 105.200 102.120 105.520 ; 
                RECT 107.240 105.200 200.720 105.520 ; 
                RECT 413.240 105.200 422.720 105.520 ; 
                RECT 0.160 106.560 198.000 106.880 ; 
                RECT 413.240 106.560 422.720 106.880 ; 
                RECT 0.160 107.920 81.040 108.240 ; 
                RECT 99.080 107.920 195.280 108.240 ; 
                RECT 413.240 107.920 422.720 108.240 ; 
                RECT 0.160 109.280 81.040 109.600 ; 
                RECT 99.080 109.280 117.760 109.600 ; 
                RECT 120.160 109.280 192.560 109.600 ; 
                RECT 413.240 109.280 422.720 109.600 ; 
                RECT 0.160 110.640 81.040 110.960 ; 
                RECT 99.080 110.640 192.560 110.960 ; 
                RECT 413.240 110.640 422.720 110.960 ; 
                RECT 0.160 112.000 81.040 112.320 ; 
                RECT 99.080 112.000 203.440 112.320 ; 
                RECT 413.240 112.000 422.720 112.320 ; 
                RECT 0.160 113.360 81.040 113.680 ; 
                RECT 99.080 113.360 203.440 113.680 ; 
                RECT 413.240 113.360 422.720 113.680 ; 
                RECT 0.160 114.720 81.040 115.040 ; 
                RECT 99.080 114.720 104.160 115.040 ; 
                RECT 109.280 114.720 155.160 115.040 ; 
                RECT 186.800 114.720 203.440 115.040 ; 
                RECT 413.240 114.720 422.720 115.040 ; 
                RECT 0.160 116.080 81.040 116.400 ; 
                RECT 99.080 116.080 155.160 116.400 ; 
                RECT 186.800 116.080 203.440 116.400 ; 
                RECT 413.240 116.080 422.720 116.400 ; 
                RECT 0.160 117.440 81.040 117.760 ; 
                RECT 99.080 117.440 110.960 117.760 ; 
                RECT 119.480 117.440 155.160 117.760 ; 
                RECT 186.800 117.440 203.440 117.760 ; 
                RECT 413.240 117.440 422.720 117.760 ; 
                RECT 0.160 118.800 81.040 119.120 ; 
                RECT 99.760 118.800 155.160 119.120 ; 
                RECT 186.800 118.800 203.440 119.120 ; 
                RECT 413.240 118.800 422.720 119.120 ; 
                RECT 0.160 120.160 81.040 120.480 ; 
                RECT 99.080 120.160 106.880 120.480 ; 
                RECT 109.960 120.160 155.160 120.480 ; 
                RECT 186.800 120.160 203.440 120.480 ; 
                RECT 413.240 120.160 422.720 120.480 ; 
                RECT 0.160 121.520 81.040 121.840 ; 
                RECT 99.080 121.520 104.160 121.840 ; 
                RECT 107.240 121.520 155.160 121.840 ; 
                RECT 186.800 121.520 203.440 121.840 ; 
                RECT 413.240 121.520 422.720 121.840 ; 
                RECT 0.160 122.880 81.040 123.200 ; 
                RECT 99.080 122.880 155.160 123.200 ; 
                RECT 186.800 122.880 203.440 123.200 ; 
                RECT 413.240 122.880 422.720 123.200 ; 
                RECT 0.160 124.240 81.040 124.560 ; 
                RECT 99.080 124.240 193.920 124.560 ; 
                RECT 413.240 124.240 422.720 124.560 ; 
                RECT 0.160 125.600 81.040 125.920 ; 
                RECT 99.080 125.600 193.920 125.920 ; 
                RECT 413.240 125.600 422.720 125.920 ; 
                RECT 0.160 126.960 81.040 127.280 ; 
                RECT 99.080 126.960 196.640 127.280 ; 
                RECT 413.240 126.960 422.720 127.280 ; 
                RECT 0.160 128.320 81.040 128.640 ; 
                RECT 99.080 128.320 199.360 128.640 ; 
                RECT 413.240 128.320 422.720 128.640 ; 
                RECT 0.160 129.680 81.040 130.000 ; 
                RECT 99.080 129.680 155.160 130.000 ; 
                RECT 413.240 129.680 422.720 130.000 ; 
                RECT 0.160 131.040 81.040 131.360 ; 
                RECT 99.080 131.040 105.520 131.360 ; 
                RECT 109.960 131.040 155.160 131.360 ; 
                RECT 413.240 131.040 422.720 131.360 ; 
                RECT 0.160 132.400 155.160 132.720 ; 
                RECT 186.120 132.400 203.440 132.720 ; 
                RECT 413.240 132.400 422.720 132.720 ; 
                RECT 0.160 133.760 155.160 134.080 ; 
                RECT 186.120 133.760 203.440 134.080 ; 
                RECT 413.240 133.760 422.720 134.080 ; 
                RECT 0.160 135.120 108.240 135.440 ; 
                RECT 114.040 135.120 155.160 135.440 ; 
                RECT 186.120 135.120 203.440 135.440 ; 
                RECT 413.240 135.120 422.720 135.440 ; 
                RECT 0.160 136.480 62.000 136.800 ; 
                RECT 80.720 136.480 86.480 136.800 ; 
                RECT 94.320 136.480 155.160 136.800 ; 
                RECT 186.120 136.480 203.440 136.800 ; 
                RECT 413.240 136.480 422.720 136.800 ; 
                RECT 0.160 137.840 62.000 138.160 ; 
                RECT 98.400 137.840 155.160 138.160 ; 
                RECT 186.120 137.840 203.440 138.160 ; 
                RECT 413.240 137.840 422.720 138.160 ; 
                RECT 0.160 139.200 62.000 139.520 ; 
                RECT 98.400 139.200 155.160 139.520 ; 
                RECT 413.240 139.200 422.720 139.520 ; 
                RECT 0.160 140.560 62.000 140.880 ; 
                RECT 80.720 140.560 86.480 140.880 ; 
                RECT 94.320 140.560 102.800 140.880 ; 
                RECT 112.680 140.560 155.160 140.880 ; 
                RECT 413.240 140.560 422.720 140.880 ; 
                RECT 0.160 141.920 60.640 142.240 ; 
                RECT 93.640 141.920 155.160 142.240 ; 
                RECT 186.120 141.920 422.720 142.240 ; 
                RECT 0.160 143.280 93.280 143.600 ; 
                RECT 152.800 143.280 422.720 143.600 ; 
                RECT 0.160 144.640 200.720 144.960 ; 
                RECT 415.280 144.640 422.720 144.960 ; 
                RECT 0.160 146.000 200.720 146.320 ; 
                RECT 415.280 146.000 422.720 146.320 ; 
                RECT 0.160 147.360 200.720 147.680 ; 
                RECT 415.280 147.360 422.720 147.680 ; 
                RECT 0.160 148.720 25.960 149.040 ; 
                RECT 32.440 148.720 34.800 149.040 ; 
                RECT 47.400 148.720 79.000 149.040 ; 
                RECT 415.280 148.720 422.720 149.040 ; 
                RECT 0.160 150.080 23.920 150.400 ; 
                RECT 34.480 150.080 36.160 150.400 ; 
                RECT 46.040 150.080 63.360 150.400 ; 
                RECT 69.160 150.080 79.000 150.400 ; 
                RECT 415.280 150.080 422.720 150.400 ; 
                RECT 0.160 151.440 23.920 151.760 ; 
                RECT 34.480 151.440 37.520 151.760 ; 
                RECT 45.360 151.440 59.280 151.760 ; 
                RECT 69.160 151.440 79.000 151.760 ; 
                RECT 415.280 151.440 422.720 151.760 ; 
                RECT 0.160 152.800 23.920 153.120 ; 
                RECT 34.480 152.800 59.280 153.120 ; 
                RECT 69.160 152.800 79.000 153.120 ; 
                RECT 415.280 152.800 422.720 153.120 ; 
                RECT 0.160 154.160 59.280 154.480 ; 
                RECT 69.160 154.160 79.000 154.480 ; 
                RECT 415.280 154.160 422.720 154.480 ; 
                RECT 0.160 155.520 23.920 155.840 ; 
                RECT 34.480 155.520 59.280 155.840 ; 
                RECT 69.160 155.520 79.000 155.840 ; 
                RECT 415.280 155.520 422.720 155.840 ; 
                RECT 0.160 156.880 23.920 157.200 ; 
                RECT 34.480 156.880 79.000 157.200 ; 
                RECT 415.280 156.880 422.720 157.200 ; 
                RECT 0.160 158.240 59.960 158.560 ; 
                RECT 69.160 158.240 79.000 158.560 ; 
                RECT 415.280 158.240 422.720 158.560 ; 
                RECT 0.160 159.600 59.280 159.920 ; 
                RECT 69.160 159.600 79.000 159.920 ; 
                RECT 415.280 159.600 422.720 159.920 ; 
                RECT 0.160 160.960 59.280 161.280 ; 
                RECT 69.160 160.960 79.000 161.280 ; 
                RECT 415.280 160.960 422.720 161.280 ; 
                RECT 0.160 162.320 17.120 162.640 ; 
                RECT 19.520 162.320 32.760 162.640 ; 
                RECT 35.840 162.320 59.280 162.640 ; 
                RECT 69.160 162.320 79.000 162.640 ; 
                RECT 415.280 162.320 422.720 162.640 ; 
                RECT 0.160 163.680 16.440 164.000 ; 
                RECT 19.520 163.680 32.760 164.000 ; 
                RECT 36.520 163.680 59.280 164.000 ; 
                RECT 69.160 163.680 79.000 164.000 ; 
                RECT 415.280 163.680 422.720 164.000 ; 
                RECT 0.160 165.040 15.760 165.360 ; 
                RECT 19.520 165.040 79.000 165.360 ; 
                RECT 415.280 165.040 422.720 165.360 ; 
                RECT 0.160 166.400 15.080 166.720 ; 
                RECT 19.520 166.400 59.960 166.720 ; 
                RECT 69.160 166.400 79.000 166.720 ; 
                RECT 415.280 166.400 422.720 166.720 ; 
                RECT 0.160 167.760 59.280 168.080 ; 
                RECT 69.160 167.760 79.000 168.080 ; 
                RECT 415.280 167.760 422.720 168.080 ; 
                RECT 0.160 169.120 14.400 169.440 ; 
                RECT 19.520 169.120 59.280 169.440 ; 
                RECT 69.160 169.120 79.000 169.440 ; 
                RECT 415.280 169.120 422.720 169.440 ; 
                RECT 0.160 170.480 13.720 170.800 ; 
                RECT 19.520 170.480 59.280 170.800 ; 
                RECT 69.160 170.480 79.000 170.800 ; 
                RECT 415.280 170.480 422.720 170.800 ; 
                RECT 0.160 171.840 59.280 172.160 ; 
                RECT 69.160 171.840 79.000 172.160 ; 
                RECT 415.280 171.840 422.720 172.160 ; 
                RECT 0.160 173.200 13.040 173.520 ; 
                RECT 19.520 173.200 79.000 173.520 ; 
                RECT 415.280 173.200 422.720 173.520 ; 
                RECT 0.160 174.560 12.360 174.880 ; 
                RECT 19.520 174.560 32.760 174.880 ; 
                RECT 38.560 174.560 59.280 174.880 ; 
                RECT 69.160 174.560 79.000 174.880 ; 
                RECT 415.280 174.560 422.720 174.880 ; 
                RECT 0.160 175.920 59.280 176.240 ; 
                RECT 69.160 175.920 79.000 176.240 ; 
                RECT 415.280 175.920 422.720 176.240 ; 
                RECT 0.160 177.280 11.680 177.600 ; 
                RECT 19.520 177.280 32.760 177.600 ; 
                RECT 37.880 177.280 59.280 177.600 ; 
                RECT 69.160 177.280 79.000 177.600 ; 
                RECT 415.280 177.280 422.720 177.600 ; 
                RECT 0.160 178.640 11.000 178.960 ; 
                RECT 19.520 178.640 32.760 178.960 ; 
                RECT 37.200 178.640 59.280 178.960 ; 
                RECT 69.160 178.640 79.000 178.960 ; 
                RECT 415.280 178.640 422.720 178.960 ; 
                RECT 0.160 180.000 10.320 180.320 ; 
                RECT 19.520 180.000 32.760 180.320 ; 
                RECT 36.520 180.000 59.280 180.320 ; 
                RECT 68.480 180.000 79.000 180.320 ; 
                RECT 415.280 180.000 422.720 180.320 ; 
                RECT 0.160 181.360 9.640 181.680 ; 
                RECT 19.520 181.360 63.360 181.680 ; 
                RECT 69.160 181.360 79.000 181.680 ; 
                RECT 415.280 181.360 422.720 181.680 ; 
                RECT 0.160 182.720 60.640 183.040 ; 
                RECT 69.160 182.720 79.000 183.040 ; 
                RECT 415.280 182.720 422.720 183.040 ; 
                RECT 0.160 184.080 60.640 184.400 ; 
                RECT 69.160 184.080 79.000 184.400 ; 
                RECT 415.280 184.080 422.720 184.400 ; 
                RECT 0.160 185.440 60.640 185.760 ; 
                RECT 69.160 185.440 79.000 185.760 ; 
                RECT 415.280 185.440 422.720 185.760 ; 
                RECT 0.160 186.800 60.640 187.120 ; 
                RECT 69.160 186.800 79.000 187.120 ; 
                RECT 415.280 186.800 422.720 187.120 ; 
                RECT 0.160 188.160 38.200 188.480 ; 
                RECT 47.400 188.160 79.000 188.480 ; 
                RECT 415.280 188.160 422.720 188.480 ; 
                RECT 0.160 189.520 36.840 189.840 ; 
                RECT 46.040 189.520 65.400 189.840 ; 
                RECT 69.160 189.520 79.000 189.840 ; 
                RECT 415.280 189.520 422.720 189.840 ; 
                RECT 0.160 190.880 35.480 191.200 ; 
                RECT 45.360 190.880 59.280 191.200 ; 
                RECT 69.160 190.880 79.000 191.200 ; 
                RECT 415.280 190.880 422.720 191.200 ; 
                RECT 0.160 192.240 59.280 192.560 ; 
                RECT 69.160 192.240 79.000 192.560 ; 
                RECT 415.280 192.240 422.720 192.560 ; 
                RECT 0.160 193.600 59.280 193.920 ; 
                RECT 69.160 193.600 79.000 193.920 ; 
                RECT 415.280 193.600 422.720 193.920 ; 
                RECT 0.160 194.960 59.280 195.280 ; 
                RECT 69.160 194.960 79.000 195.280 ; 
                RECT 415.280 194.960 422.720 195.280 ; 
                RECT 0.160 196.320 59.280 196.640 ; 
                RECT 61.680 196.320 79.000 196.640 ; 
                RECT 415.280 196.320 422.720 196.640 ; 
                RECT 0.160 197.680 61.320 198.000 ; 
                RECT 69.160 197.680 79.000 198.000 ; 
                RECT 415.280 197.680 422.720 198.000 ; 
                RECT 0.160 199.040 59.280 199.360 ; 
                RECT 69.160 199.040 79.000 199.360 ; 
                RECT 415.280 199.040 422.720 199.360 ; 
                RECT 0.160 200.400 59.280 200.720 ; 
                RECT 69.160 200.400 79.000 200.720 ; 
                RECT 415.280 200.400 422.720 200.720 ; 
                RECT 0.160 201.760 59.280 202.080 ; 
                RECT 69.160 201.760 79.000 202.080 ; 
                RECT 415.280 201.760 422.720 202.080 ; 
                RECT 0.160 203.120 59.280 203.440 ; 
                RECT 69.160 203.120 79.000 203.440 ; 
                RECT 415.280 203.120 422.720 203.440 ; 
                RECT 0.160 204.480 79.000 204.800 ; 
                RECT 415.280 204.480 422.720 204.800 ; 
                RECT 0.160 205.840 61.320 206.160 ; 
                RECT 69.160 205.840 79.000 206.160 ; 
                RECT 415.280 205.840 422.720 206.160 ; 
                RECT 0.160 207.200 59.280 207.520 ; 
                RECT 69.160 207.200 79.000 207.520 ; 
                RECT 415.280 207.200 422.720 207.520 ; 
                RECT 0.160 208.560 59.280 208.880 ; 
                RECT 69.160 208.560 79.000 208.880 ; 
                RECT 415.280 208.560 422.720 208.880 ; 
                RECT 0.160 209.920 59.280 210.240 ; 
                RECT 69.160 209.920 79.000 210.240 ; 
                RECT 415.280 209.920 422.720 210.240 ; 
                RECT 0.160 211.280 59.280 211.600 ; 
                RECT 69.160 211.280 79.000 211.600 ; 
                RECT 415.280 211.280 422.720 211.600 ; 
                RECT 0.160 212.640 79.000 212.960 ; 
                RECT 415.280 212.640 422.720 212.960 ; 
                RECT 0.160 214.000 59.280 214.320 ; 
                RECT 69.160 214.000 79.000 214.320 ; 
                RECT 415.280 214.000 422.720 214.320 ; 
                RECT 0.160 215.360 59.280 215.680 ; 
                RECT 69.160 215.360 79.000 215.680 ; 
                RECT 415.280 215.360 422.720 215.680 ; 
                RECT 0.160 216.720 59.280 217.040 ; 
                RECT 69.160 216.720 79.000 217.040 ; 
                RECT 415.280 216.720 422.720 217.040 ; 
                RECT 0.160 218.080 59.280 218.400 ; 
                RECT 69.160 218.080 79.000 218.400 ; 
                RECT 415.280 218.080 422.720 218.400 ; 
                RECT 0.160 219.440 59.280 219.760 ; 
                RECT 69.160 219.440 79.000 219.760 ; 
                RECT 415.280 219.440 422.720 219.760 ; 
                RECT 0.160 220.800 79.000 221.120 ; 
                RECT 415.280 220.800 422.720 221.120 ; 
                RECT 0.160 222.160 62.000 222.480 ; 
                RECT 69.160 222.160 79.000 222.480 ; 
                RECT 415.280 222.160 422.720 222.480 ; 
                RECT 0.160 223.520 62.000 223.840 ; 
                RECT 69.160 223.520 79.000 223.840 ; 
                RECT 415.280 223.520 422.720 223.840 ; 
                RECT 0.160 224.880 62.000 225.200 ; 
                RECT 69.160 224.880 79.000 225.200 ; 
                RECT 415.280 224.880 422.720 225.200 ; 
                RECT 0.160 226.240 62.000 226.560 ; 
                RECT 69.160 226.240 79.000 226.560 ; 
                RECT 415.280 226.240 422.720 226.560 ; 
                RECT 0.160 227.600 79.000 227.920 ; 
                RECT 415.280 227.600 422.720 227.920 ; 
                RECT 0.160 228.960 63.360 229.280 ; 
                RECT 69.160 228.960 79.000 229.280 ; 
                RECT 415.280 228.960 422.720 229.280 ; 
                RECT 0.160 230.320 62.000 230.640 ; 
                RECT 69.160 230.320 79.000 230.640 ; 
                RECT 415.280 230.320 422.720 230.640 ; 
                RECT 0.160 231.680 62.000 232.000 ; 
                RECT 69.160 231.680 79.000 232.000 ; 
                RECT 415.280 231.680 422.720 232.000 ; 
                RECT 0.160 233.040 62.000 233.360 ; 
                RECT 69.160 233.040 79.000 233.360 ; 
                RECT 415.280 233.040 422.720 233.360 ; 
                RECT 0.160 234.400 62.000 234.720 ; 
                RECT 69.160 234.400 79.000 234.720 ; 
                RECT 415.280 234.400 422.720 234.720 ; 
                RECT 0.160 235.760 79.000 236.080 ; 
                RECT 415.280 235.760 422.720 236.080 ; 
                RECT 0.160 237.120 65.400 237.440 ; 
                RECT 69.160 237.120 79.000 237.440 ; 
                RECT 415.280 237.120 422.720 237.440 ; 
                RECT 0.160 238.480 66.080 238.800 ; 
                RECT 69.160 238.480 79.000 238.800 ; 
                RECT 415.280 238.480 422.720 238.800 ; 
                RECT 0.160 239.840 62.000 240.160 ; 
                RECT 69.160 239.840 79.000 240.160 ; 
                RECT 415.280 239.840 422.720 240.160 ; 
                RECT 0.160 241.200 62.000 241.520 ; 
                RECT 69.160 241.200 79.000 241.520 ; 
                RECT 415.280 241.200 422.720 241.520 ; 
                RECT 0.160 242.560 62.000 242.880 ; 
                RECT 69.160 242.560 79.000 242.880 ; 
                RECT 415.280 242.560 422.720 242.880 ; 
                RECT 0.160 243.920 79.000 244.240 ; 
                RECT 415.280 243.920 422.720 244.240 ; 
                RECT 0.160 245.280 62.680 245.600 ; 
                RECT 69.160 245.280 79.000 245.600 ; 
                RECT 415.280 245.280 422.720 245.600 ; 
                RECT 0.160 246.640 62.680 246.960 ; 
                RECT 69.160 246.640 79.000 246.960 ; 
                RECT 415.280 246.640 422.720 246.960 ; 
                RECT 0.160 248.000 64.720 248.320 ; 
                RECT 69.160 248.000 79.000 248.320 ; 
                RECT 415.280 248.000 422.720 248.320 ; 
                RECT 0.160 249.360 62.680 249.680 ; 
                RECT 69.160 249.360 79.000 249.680 ; 
                RECT 415.280 249.360 422.720 249.680 ; 
                RECT 0.160 250.720 62.680 251.040 ; 
                RECT 69.160 250.720 79.000 251.040 ; 
                RECT 415.280 250.720 422.720 251.040 ; 
                RECT 0.160 252.080 79.000 252.400 ; 
                RECT 415.280 252.080 422.720 252.400 ; 
                RECT 0.160 253.440 62.680 253.760 ; 
                RECT 69.160 253.440 79.000 253.760 ; 
                RECT 415.280 253.440 422.720 253.760 ; 
                RECT 0.160 254.800 62.680 255.120 ; 
                RECT 69.160 254.800 79.000 255.120 ; 
                RECT 415.280 254.800 422.720 255.120 ; 
                RECT 0.160 256.160 62.680 256.480 ; 
                RECT 69.160 256.160 79.000 256.480 ; 
                RECT 415.280 256.160 422.720 256.480 ; 
                RECT 0.160 257.520 66.760 257.840 ; 
                RECT 69.160 257.520 79.000 257.840 ; 
                RECT 415.280 257.520 422.720 257.840 ; 
                RECT 0.160 258.880 62.680 259.200 ; 
                RECT 69.160 258.880 79.000 259.200 ; 
                RECT 415.280 258.880 422.720 259.200 ; 
                RECT 0.160 260.240 79.000 260.560 ; 
                RECT 415.280 260.240 422.720 260.560 ; 
                RECT 0.160 261.600 63.360 261.920 ; 
                RECT 69.160 261.600 79.000 261.920 ; 
                RECT 415.280 261.600 422.720 261.920 ; 
                RECT 0.160 262.960 63.360 263.280 ; 
                RECT 69.160 262.960 79.000 263.280 ; 
                RECT 415.280 262.960 422.720 263.280 ; 
                RECT 0.160 264.320 63.360 264.640 ; 
                RECT 69.160 264.320 79.000 264.640 ; 
                RECT 415.280 264.320 422.720 264.640 ; 
                RECT 0.160 265.680 63.360 266.000 ; 
                RECT 69.160 265.680 79.000 266.000 ; 
                RECT 415.280 265.680 422.720 266.000 ; 
                RECT 0.160 267.040 79.000 267.360 ; 
                RECT 415.280 267.040 422.720 267.360 ; 
                RECT 0.160 268.400 65.400 268.720 ; 
                RECT 69.160 268.400 79.000 268.720 ; 
                RECT 415.280 268.400 422.720 268.720 ; 
                RECT 0.160 269.760 63.360 270.080 ; 
                RECT 69.160 269.760 79.000 270.080 ; 
                RECT 415.280 269.760 422.720 270.080 ; 
                RECT 0.160 271.120 63.360 271.440 ; 
                RECT 69.160 271.120 79.000 271.440 ; 
                RECT 415.280 271.120 422.720 271.440 ; 
                RECT 0.160 272.480 63.360 272.800 ; 
                RECT 69.160 272.480 79.000 272.800 ; 
                RECT 415.280 272.480 422.720 272.800 ; 
                RECT 0.160 273.840 63.360 274.160 ; 
                RECT 69.160 273.840 79.000 274.160 ; 
                RECT 415.280 273.840 422.720 274.160 ; 
                RECT 0.160 275.200 79.000 275.520 ; 
                RECT 415.280 275.200 422.720 275.520 ; 
                RECT 0.160 276.560 79.000 276.880 ; 
                RECT 415.280 276.560 422.720 276.880 ; 
                RECT 0.160 277.920 200.720 278.240 ; 
                RECT 415.280 277.920 422.720 278.240 ; 
                RECT 0.160 279.280 200.720 279.600 ; 
                RECT 415.280 279.280 422.720 279.600 ; 
                RECT 0.160 280.640 422.720 280.960 ; 
                RECT 0.160 282.000 422.720 282.320 ; 
                RECT 0.160 283.360 422.720 283.680 ; 
                RECT 0.160 284.720 422.720 285.040 ; 
                RECT 0.160 286.080 422.720 286.400 ; 
                RECT 0.160 0.160 422.720 1.520 ; 
                RECT 0.160 290.120 422.720 291.480 ; 
                RECT 204.860 32.275 210.660 33.645 ; 
                RECT 405.560 32.275 411.360 33.645 ; 
                RECT 204.860 37.795 210.660 39.535 ; 
                RECT 405.560 37.795 411.360 39.535 ; 
                RECT 204.860 43.640 210.660 45.210 ; 
                RECT 405.560 43.640 411.360 45.210 ; 
                RECT 204.860 49.230 210.660 50.800 ; 
                RECT 405.560 49.230 411.360 50.800 ; 
                RECT 204.860 90.135 411.360 90.425 ; 
                RECT 204.860 57.660 411.360 59.460 ; 
                RECT 204.860 72.140 411.360 72.940 ; 
                RECT 204.860 113.775 411.360 115.575 ; 
                RECT 204.860 134.765 411.360 137.365 ; 
                RECT 204.860 77.030 411.360 77.830 ; 
                RECT 204.860 84.710 411.360 86.800 ; 
                RECT 204.860 69.130 411.360 69.930 ; 
                RECT 204.860 16.520 411.360 18.320 ; 
                RECT 84.230 148.435 86.150 276.415 ; 
                RECT 95.105 148.435 97.025 276.415 ; 
                RECT 98.945 148.435 100.865 276.415 ; 
                RECT 102.785 148.435 104.705 276.415 ; 
                RECT 118.450 148.435 120.370 276.415 ; 
                RECT 122.290 148.435 124.210 276.415 ; 
                RECT 126.130 148.435 128.050 276.415 ; 
                RECT 129.970 148.435 131.890 276.415 ; 
                RECT 133.810 148.435 135.730 276.415 ; 
                RECT 158.410 148.435 160.330 276.415 ; 
                RECT 162.250 148.435 164.170 276.415 ; 
                RECT 166.090 148.435 168.010 276.415 ; 
                RECT 169.930 148.435 171.850 276.415 ; 
                RECT 173.770 148.435 175.690 276.415 ; 
                RECT 177.610 148.435 179.530 276.415 ; 
                RECT 181.450 148.435 183.370 276.415 ; 
                RECT 185.290 148.435 187.210 276.415 ; 
                RECT 189.130 148.435 191.050 276.415 ; 
                RECT 192.970 148.435 194.890 276.415 ; 
                RECT 196.810 148.435 198.730 276.415 ; 
                RECT 141.095 57.135 142.845 101.135 ; 
                RECT 147.555 57.135 149.475 101.135 ; 
                RECT 154.185 57.135 155.935 101.135 ; 
                RECT 163.225 57.135 165.145 101.135 ; 
                RECT 175.820 57.135 177.740 101.135 ; 
                RECT 179.660 57.135 181.580 101.135 ; 
                RECT 183.500 57.135 185.420 101.135 ; 
                RECT 158.465 129.320 160.215 141.800 ; 
                RECT 164.925 129.320 166.845 141.800 ; 
                RECT 175.800 129.320 177.720 141.800 ; 
                RECT 179.640 129.320 181.560 141.800 ; 
                RECT 183.480 129.320 185.400 141.800 ; 
                RECT 159.240 115.000 161.160 123.320 ; 
                RECT 166.645 115.000 168.565 123.320 ; 
                RECT 176.445 115.000 178.365 123.320 ; 
                RECT 180.285 115.000 182.205 123.320 ; 
                RECT 184.125 115.000 186.045 123.320 ; 
                RECT 183.745 47.555 185.665 51.135 ; 
                RECT 24.710 150.705 33.870 151.455 ; 
                RECT 24.710 155.460 33.870 157.380 ; 
                RECT 81.970 138.490 98.010 139.290 ; 
                RECT 62.770 139.200 80.010 140.890 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 213.640 5.560 ; 
                RECT 404.400 5.240 420.000 5.560 ; 
                RECT 2.880 6.600 420.000 6.920 ; 
                RECT 2.880 7.960 420.000 8.280 ; 
                RECT 2.880 9.320 187.800 9.640 ; 
                RECT 209.240 9.320 420.000 9.640 ; 
                RECT 2.880 10.680 203.440 11.000 ; 
                RECT 413.240 10.680 420.000 11.000 ; 
                RECT 2.880 12.040 203.440 12.360 ; 
                RECT 413.240 12.040 420.000 12.360 ; 
                RECT 2.880 13.400 203.440 13.720 ; 
                RECT 413.240 13.400 420.000 13.720 ; 
                RECT 2.880 14.760 203.440 15.080 ; 
                RECT 413.240 14.760 420.000 15.080 ; 
                RECT 2.880 16.120 125.920 16.440 ; 
                RECT 188.840 16.120 203.440 16.440 ; 
                RECT 413.240 16.120 420.000 16.440 ; 
                RECT 2.880 17.480 203.440 17.800 ; 
                RECT 413.240 17.480 420.000 17.800 ; 
                RECT 2.880 18.840 203.440 19.160 ; 
                RECT 413.240 18.840 420.000 19.160 ; 
                RECT 2.880 20.200 125.920 20.520 ; 
                RECT 188.160 20.200 203.440 20.520 ; 
                RECT 413.240 20.200 420.000 20.520 ; 
                RECT 2.880 21.560 203.440 21.880 ; 
                RECT 413.240 21.560 420.000 21.880 ; 
                RECT 2.880 22.920 203.440 23.240 ; 
                RECT 413.240 22.920 420.000 23.240 ; 
                RECT 2.880 24.280 203.440 24.600 ; 
                RECT 413.240 24.280 420.000 24.600 ; 
                RECT 2.880 25.640 203.440 25.960 ; 
                RECT 413.240 25.640 420.000 25.960 ; 
                RECT 2.880 27.000 203.440 27.320 ; 
                RECT 413.240 27.000 420.000 27.320 ; 
                RECT 2.880 28.360 202.760 28.680 ; 
                RECT 413.240 28.360 420.000 28.680 ; 
                RECT 2.880 29.720 203.440 30.040 ; 
                RECT 413.240 29.720 420.000 30.040 ; 
                RECT 2.880 31.080 203.440 31.400 ; 
                RECT 413.240 31.080 420.000 31.400 ; 
                RECT 2.880 32.440 203.440 32.760 ; 
                RECT 413.240 32.440 420.000 32.760 ; 
                RECT 2.880 33.800 203.440 34.120 ; 
                RECT 413.240 33.800 420.000 34.120 ; 
                RECT 2.880 35.160 203.440 35.480 ; 
                RECT 413.240 35.160 420.000 35.480 ; 
                RECT 2.880 36.520 128.640 36.840 ; 
                RECT 167.080 36.520 203.440 36.840 ; 
                RECT 413.240 36.520 420.000 36.840 ; 
                RECT 2.880 37.880 127.280 38.200 ; 
                RECT 173.200 37.880 203.440 38.200 ; 
                RECT 413.240 37.880 420.000 38.200 ; 
                RECT 2.880 39.240 104.160 39.560 ; 
                RECT 188.160 39.240 203.440 39.560 ; 
                RECT 413.240 39.240 420.000 39.560 ; 
                RECT 2.880 40.600 105.520 40.920 ; 
                RECT 178.640 40.600 203.440 40.920 ; 
                RECT 413.240 40.600 420.000 40.920 ; 
                RECT 2.880 41.960 203.440 42.280 ; 
                RECT 413.240 41.960 420.000 42.280 ; 
                RECT 2.880 43.320 203.440 43.640 ; 
                RECT 413.240 43.320 420.000 43.640 ; 
                RECT 2.880 44.680 203.440 45.000 ; 
                RECT 413.240 44.680 420.000 45.000 ; 
                RECT 2.880 46.040 203.440 46.360 ; 
                RECT 413.240 46.040 420.000 46.360 ; 
                RECT 2.880 47.400 102.800 47.720 ; 
                RECT 113.360 47.400 179.640 47.720 ; 
                RECT 186.120 47.400 203.440 47.720 ; 
                RECT 413.240 47.400 420.000 47.720 ; 
                RECT 2.880 48.760 104.160 49.080 ; 
                RECT 105.880 48.760 179.640 49.080 ; 
                RECT 413.240 48.760 420.000 49.080 ; 
                RECT 2.880 50.120 105.520 50.440 ; 
                RECT 109.960 50.120 117.080 50.440 ; 
                RECT 120.160 50.120 179.640 50.440 ; 
                RECT 186.120 50.120 203.440 50.440 ; 
                RECT 413.240 50.120 420.000 50.440 ; 
                RECT 2.880 51.480 105.520 51.800 ; 
                RECT 108.600 51.480 179.640 51.800 ; 
                RECT 186.120 51.480 203.440 51.800 ; 
                RECT 413.240 51.480 420.000 51.800 ; 
                RECT 2.880 52.840 111.640 53.160 ; 
                RECT 120.160 52.840 203.440 53.160 ; 
                RECT 413.240 52.840 420.000 53.160 ; 
                RECT 2.880 54.200 106.880 54.520 ; 
                RECT 113.360 54.200 203.440 54.520 ; 
                RECT 413.240 54.200 420.000 54.520 ; 
                RECT 2.880 55.560 104.160 55.880 ; 
                RECT 113.360 55.560 203.440 55.880 ; 
                RECT 413.240 55.560 420.000 55.880 ; 
                RECT 2.880 56.920 138.160 57.240 ; 
                RECT 186.120 56.920 203.440 57.240 ; 
                RECT 413.240 56.920 420.000 57.240 ; 
                RECT 2.880 58.280 104.160 58.600 ; 
                RECT 113.360 58.280 127.280 58.600 ; 
                RECT 131.720 58.280 138.160 58.600 ; 
                RECT 186.120 58.280 203.440 58.600 ; 
                RECT 413.240 58.280 420.000 58.600 ; 
                RECT 2.880 59.640 111.640 59.960 ; 
                RECT 119.480 59.640 128.640 59.960 ; 
                RECT 131.040 59.640 138.160 59.960 ; 
                RECT 194.280 59.640 203.440 59.960 ; 
                RECT 413.240 59.640 420.000 59.960 ; 
                RECT 2.880 61.000 110.960 61.320 ; 
                RECT 113.360 61.000 138.160 61.320 ; 
                RECT 195.640 61.000 203.440 61.320 ; 
                RECT 413.240 61.000 420.000 61.320 ; 
                RECT 2.880 62.360 138.160 62.680 ; 
                RECT 195.640 62.360 203.440 62.680 ; 
                RECT 413.240 62.360 420.000 62.680 ; 
                RECT 2.880 63.720 111.640 64.040 ; 
                RECT 120.160 63.720 138.160 64.040 ; 
                RECT 194.280 63.720 203.440 64.040 ; 
                RECT 413.240 63.720 420.000 64.040 ; 
                RECT 2.880 65.080 108.240 65.400 ; 
                RECT 113.360 65.080 138.160 65.400 ; 
                RECT 195.640 65.080 203.440 65.400 ; 
                RECT 413.240 65.080 420.000 65.400 ; 
                RECT 2.880 66.440 110.960 66.760 ; 
                RECT 113.360 66.440 138.160 66.760 ; 
                RECT 186.120 66.440 203.440 66.760 ; 
                RECT 413.240 66.440 420.000 66.760 ; 
                RECT 2.880 67.800 138.160 68.120 ; 
                RECT 195.640 67.800 203.440 68.120 ; 
                RECT 413.240 67.800 420.000 68.120 ; 
                RECT 2.880 69.160 102.120 69.480 ; 
                RECT 124.920 69.160 138.160 69.480 ; 
                RECT 198.360 69.160 203.440 69.480 ; 
                RECT 413.240 69.160 420.000 69.480 ; 
                RECT 2.880 70.520 120.480 70.840 ; 
                RECT 126.280 70.520 138.160 70.840 ; 
                RECT 197.000 70.520 203.440 70.840 ; 
                RECT 413.240 70.520 420.000 70.840 ; 
                RECT 2.880 71.880 110.960 72.200 ; 
                RECT 113.360 71.880 123.200 72.200 ; 
                RECT 126.960 71.880 138.160 72.200 ; 
                RECT 198.360 71.880 203.440 72.200 ; 
                RECT 413.240 71.880 420.000 72.200 ; 
                RECT 2.880 73.240 102.800 73.560 ; 
                RECT 116.080 73.240 138.160 73.560 ; 
                RECT 198.360 73.240 203.440 73.560 ; 
                RECT 413.240 73.240 420.000 73.560 ; 
                RECT 2.880 74.600 110.960 74.920 ; 
                RECT 120.160 74.600 138.160 74.920 ; 
                RECT 186.120 74.600 203.440 74.920 ; 
                RECT 413.240 74.600 420.000 74.920 ; 
                RECT 2.880 75.960 108.920 76.280 ; 
                RECT 120.160 75.960 138.160 76.280 ; 
                RECT 198.360 75.960 203.440 76.280 ; 
                RECT 413.240 75.960 420.000 76.280 ; 
                RECT 2.880 77.320 104.160 77.640 ; 
                RECT 110.640 77.320 138.160 77.640 ; 
                RECT 197.000 77.320 203.440 77.640 ; 
                RECT 413.240 77.320 420.000 77.640 ; 
                RECT 2.880 78.680 138.160 79.000 ; 
                RECT 198.360 78.680 203.440 79.000 ; 
                RECT 413.240 78.680 420.000 79.000 ; 
                RECT 2.880 80.040 104.160 80.360 ; 
                RECT 107.240 80.040 138.160 80.360 ; 
                RECT 201.080 80.040 203.440 80.360 ; 
                RECT 413.240 80.040 420.000 80.360 ; 
                RECT 2.880 81.400 104.160 81.720 ; 
                RECT 113.360 81.400 138.160 81.720 ; 
                RECT 201.080 81.400 203.440 81.720 ; 
                RECT 413.240 81.400 420.000 81.720 ; 
                RECT 2.880 82.760 108.240 83.080 ; 
                RECT 118.800 82.760 138.160 83.080 ; 
                RECT 199.720 82.760 203.440 83.080 ; 
                RECT 413.240 82.760 420.000 83.080 ; 
                RECT 2.880 84.120 110.960 84.440 ; 
                RECT 112.680 84.120 138.160 84.440 ; 
                RECT 186.120 84.120 203.440 84.440 ; 
                RECT 413.240 84.120 420.000 84.440 ; 
                RECT 2.880 85.480 111.640 85.800 ; 
                RECT 114.040 85.480 138.160 85.800 ; 
                RECT 199.720 85.480 203.440 85.800 ; 
                RECT 413.240 85.480 420.000 85.800 ; 
                RECT 2.880 86.840 138.160 87.160 ; 
                RECT 201.080 86.840 203.440 87.160 ; 
                RECT 413.240 86.840 420.000 87.160 ; 
                RECT 2.880 88.200 102.800 88.520 ; 
                RECT 120.160 88.200 138.160 88.520 ; 
                RECT 201.080 88.200 203.440 88.520 ; 
                RECT 413.240 88.200 420.000 88.520 ; 
                RECT 2.880 89.560 102.800 89.880 ; 
                RECT 113.360 89.560 117.760 89.880 ; 
                RECT 120.160 89.560 138.160 89.880 ; 
                RECT 199.720 89.560 203.440 89.880 ; 
                RECT 413.240 89.560 420.000 89.880 ; 
                RECT 2.880 90.920 110.960 91.240 ; 
                RECT 114.040 90.920 138.160 91.240 ; 
                RECT 413.240 90.920 420.000 91.240 ; 
                RECT 2.880 92.280 138.160 92.600 ; 
                RECT 186.120 92.280 203.440 92.600 ; 
                RECT 413.240 92.280 420.000 92.600 ; 
                RECT 2.880 93.640 138.160 93.960 ; 
                RECT 413.240 93.640 420.000 93.960 ; 
                RECT 2.880 95.000 98.720 95.320 ; 
                RECT 112.680 95.000 138.160 95.320 ; 
                RECT 413.240 95.000 420.000 95.320 ; 
                RECT 2.880 96.360 108.920 96.680 ; 
                RECT 116.080 96.360 138.160 96.680 ; 
                RECT 413.240 96.360 420.000 96.680 ; 
                RECT 2.880 97.720 138.160 98.040 ; 
                RECT 413.240 97.720 420.000 98.040 ; 
                RECT 2.880 99.080 138.160 99.400 ; 
                RECT 413.240 99.080 420.000 99.400 ; 
                RECT 2.880 100.440 107.560 100.760 ; 
                RECT 122.200 100.440 138.160 100.760 ; 
                RECT 186.120 100.440 203.440 100.760 ; 
                RECT 413.240 100.440 420.000 100.760 ; 
                RECT 2.880 101.800 203.440 102.120 ; 
                RECT 413.240 101.800 420.000 102.120 ; 
                RECT 2.880 103.160 203.440 103.480 ; 
                RECT 413.240 103.160 420.000 103.480 ; 
                RECT 2.880 104.520 104.160 104.840 ; 
                RECT 107.240 104.520 189.840 104.840 ; 
                RECT 413.240 104.520 420.000 104.840 ; 
                RECT 2.880 105.880 102.120 106.200 ; 
                RECT 105.880 105.880 200.720 106.200 ; 
                RECT 413.240 105.880 420.000 106.200 ; 
                RECT 2.880 107.240 198.000 107.560 ; 
                RECT 413.240 107.240 420.000 107.560 ; 
                RECT 2.880 108.600 81.040 108.920 ; 
                RECT 99.080 108.600 117.760 108.920 ; 
                RECT 120.160 108.600 195.280 108.920 ; 
                RECT 413.240 108.600 420.000 108.920 ; 
                RECT 2.880 109.960 81.040 110.280 ; 
                RECT 99.080 109.960 192.560 110.280 ; 
                RECT 413.240 109.960 420.000 110.280 ; 
                RECT 2.880 111.320 81.040 111.640 ; 
                RECT 99.080 111.320 203.440 111.640 ; 
                RECT 413.240 111.320 420.000 111.640 ; 
                RECT 2.880 112.680 81.040 113.000 ; 
                RECT 99.080 112.680 203.440 113.000 ; 
                RECT 413.240 112.680 420.000 113.000 ; 
                RECT 2.880 114.040 81.040 114.360 ; 
                RECT 99.080 114.040 104.160 114.360 ; 
                RECT 109.280 114.040 203.440 114.360 ; 
                RECT 413.240 114.040 420.000 114.360 ; 
                RECT 2.880 115.400 81.040 115.720 ; 
                RECT 99.080 115.400 125.920 115.720 ; 
                RECT 152.120 115.400 155.160 115.720 ; 
                RECT 186.800 115.400 203.440 115.720 ; 
                RECT 413.240 115.400 420.000 115.720 ; 
                RECT 2.880 116.760 81.040 117.080 ; 
                RECT 99.080 116.760 110.960 117.080 ; 
                RECT 119.480 116.760 155.160 117.080 ; 
                RECT 186.800 116.760 203.440 117.080 ; 
                RECT 413.240 116.760 420.000 117.080 ; 
                RECT 2.880 118.120 81.040 118.440 ; 
                RECT 99.080 118.120 155.160 118.440 ; 
                RECT 186.800 118.120 203.440 118.440 ; 
                RECT 413.240 118.120 420.000 118.440 ; 
                RECT 2.880 119.480 81.040 119.800 ; 
                RECT 99.760 119.480 106.880 119.800 ; 
                RECT 109.960 119.480 155.160 119.800 ; 
                RECT 186.800 119.480 203.440 119.800 ; 
                RECT 413.240 119.480 420.000 119.800 ; 
                RECT 2.880 120.840 81.040 121.160 ; 
                RECT 99.080 120.840 104.160 121.160 ; 
                RECT 107.240 120.840 155.160 121.160 ; 
                RECT 186.800 120.840 203.440 121.160 ; 
                RECT 413.240 120.840 420.000 121.160 ; 
                RECT 2.880 122.200 81.040 122.520 ; 
                RECT 99.080 122.200 155.160 122.520 ; 
                RECT 186.800 122.200 203.440 122.520 ; 
                RECT 413.240 122.200 420.000 122.520 ; 
                RECT 2.880 123.560 81.040 123.880 ; 
                RECT 99.080 123.560 155.160 123.880 ; 
                RECT 186.800 123.560 203.440 123.880 ; 
                RECT 413.240 123.560 420.000 123.880 ; 
                RECT 2.880 124.920 81.040 125.240 ; 
                RECT 99.080 124.920 193.920 125.240 ; 
                RECT 413.240 124.920 420.000 125.240 ; 
                RECT 2.880 126.280 81.040 126.600 ; 
                RECT 99.080 126.280 196.640 126.600 ; 
                RECT 413.240 126.280 420.000 126.600 ; 
                RECT 2.880 127.640 81.040 127.960 ; 
                RECT 99.080 127.640 199.360 127.960 ; 
                RECT 413.240 127.640 420.000 127.960 ; 
                RECT 2.880 129.000 81.040 129.320 ; 
                RECT 99.080 129.000 155.160 129.320 ; 
                RECT 186.120 129.000 202.080 129.320 ; 
                RECT 413.240 129.000 420.000 129.320 ; 
                RECT 2.880 130.360 81.040 130.680 ; 
                RECT 99.080 130.360 105.520 130.680 ; 
                RECT 109.960 130.360 155.160 130.680 ; 
                RECT 413.240 130.360 420.000 130.680 ; 
                RECT 2.880 131.720 81.040 132.040 ; 
                RECT 99.080 131.720 155.160 132.040 ; 
                RECT 186.120 131.720 203.440 132.040 ; 
                RECT 413.240 131.720 420.000 132.040 ; 
                RECT 2.880 133.080 155.160 133.400 ; 
                RECT 186.120 133.080 203.440 133.400 ; 
                RECT 413.240 133.080 420.000 133.400 ; 
                RECT 2.880 134.440 155.160 134.760 ; 
                RECT 186.120 134.440 203.440 134.760 ; 
                RECT 413.240 134.440 420.000 134.760 ; 
                RECT 2.880 135.800 62.000 136.120 ; 
                RECT 80.720 135.800 108.240 136.120 ; 
                RECT 114.040 135.800 155.160 136.120 ; 
                RECT 186.120 135.800 203.440 136.120 ; 
                RECT 413.240 135.800 420.000 136.120 ; 
                RECT 2.880 137.160 62.000 137.480 ; 
                RECT 80.720 137.160 86.480 137.480 ; 
                RECT 94.320 137.160 155.160 137.480 ; 
                RECT 186.120 137.160 203.440 137.480 ; 
                RECT 413.240 137.160 420.000 137.480 ; 
                RECT 2.880 138.520 62.000 138.840 ; 
                RECT 98.400 138.520 155.160 138.840 ; 
                RECT 186.120 138.520 203.440 138.840 ; 
                RECT 413.240 138.520 420.000 138.840 ; 
                RECT 2.880 139.880 62.000 140.200 ; 
                RECT 80.720 139.880 155.160 140.200 ; 
                RECT 413.240 139.880 420.000 140.200 ; 
                RECT 2.880 141.240 60.640 141.560 ; 
                RECT 94.320 141.240 102.800 141.560 ; 
                RECT 112.680 141.240 155.160 141.560 ; 
                RECT 186.120 141.240 203.440 141.560 ; 
                RECT 413.240 141.240 420.000 141.560 ; 
                RECT 2.880 142.600 86.480 142.920 ; 
                RECT 107.240 142.600 420.000 142.920 ; 
                RECT 2.880 143.960 30.720 144.280 ; 
                RECT 105.880 143.960 420.000 144.280 ; 
                RECT 2.880 145.320 200.720 145.640 ; 
                RECT 415.280 145.320 420.000 145.640 ; 
                RECT 2.880 146.680 200.720 147.000 ; 
                RECT 415.280 146.680 420.000 147.000 ; 
                RECT 2.880 148.040 25.960 148.360 ; 
                RECT 32.440 148.040 79.000 148.360 ; 
                RECT 415.280 148.040 420.000 148.360 ; 
                RECT 2.880 149.400 23.920 149.720 ; 
                RECT 46.720 149.400 79.000 149.720 ; 
                RECT 415.280 149.400 420.000 149.720 ; 
                RECT 2.880 150.760 23.920 151.080 ; 
                RECT 45.360 150.760 59.280 151.080 ; 
                RECT 69.160 150.760 79.000 151.080 ; 
                RECT 415.280 150.760 420.000 151.080 ; 
                RECT 2.880 152.120 38.200 152.440 ; 
                RECT 44.680 152.120 59.280 152.440 ; 
                RECT 69.160 152.120 79.000 152.440 ; 
                RECT 415.280 152.120 420.000 152.440 ; 
                RECT 2.880 153.480 23.920 153.800 ; 
                RECT 34.480 153.480 59.280 153.800 ; 
                RECT 69.160 153.480 79.000 153.800 ; 
                RECT 415.280 153.480 420.000 153.800 ; 
                RECT 2.880 154.840 23.920 155.160 ; 
                RECT 34.480 154.840 59.280 155.160 ; 
                RECT 69.160 154.840 79.000 155.160 ; 
                RECT 415.280 154.840 420.000 155.160 ; 
                RECT 2.880 156.200 23.920 156.520 ; 
                RECT 34.480 156.200 59.280 156.520 ; 
                RECT 69.160 156.200 79.000 156.520 ; 
                RECT 415.280 156.200 420.000 156.520 ; 
                RECT 2.880 157.560 23.920 157.880 ; 
                RECT 34.480 157.560 79.000 157.880 ; 
                RECT 415.280 157.560 420.000 157.880 ; 
                RECT 2.880 158.920 59.280 159.240 ; 
                RECT 69.160 158.920 79.000 159.240 ; 
                RECT 415.280 158.920 420.000 159.240 ; 
                RECT 2.880 160.280 59.280 160.600 ; 
                RECT 69.160 160.280 79.000 160.600 ; 
                RECT 415.280 160.280 420.000 160.600 ; 
                RECT 2.880 161.640 17.120 161.960 ; 
                RECT 19.520 161.640 59.960 161.960 ; 
                RECT 69.160 161.640 79.000 161.960 ; 
                RECT 415.280 161.640 420.000 161.960 ; 
                RECT 2.880 163.000 16.440 163.320 ; 
                RECT 19.520 163.000 59.280 163.320 ; 
                RECT 69.160 163.000 79.000 163.320 ; 
                RECT 415.280 163.000 420.000 163.320 ; 
                RECT 2.880 164.360 59.280 164.680 ; 
                RECT 66.440 164.360 79.000 164.680 ; 
                RECT 415.280 164.360 420.000 164.680 ; 
                RECT 2.880 165.720 15.760 166.040 ; 
                RECT 19.520 165.720 32.760 166.040 ; 
                RECT 37.200 165.720 63.360 166.040 ; 
                RECT 69.160 165.720 79.000 166.040 ; 
                RECT 415.280 165.720 420.000 166.040 ; 
                RECT 2.880 167.080 15.080 167.400 ; 
                RECT 19.520 167.080 32.760 167.400 ; 
                RECT 37.880 167.080 59.280 167.400 ; 
                RECT 69.160 167.080 79.000 167.400 ; 
                RECT 415.280 167.080 420.000 167.400 ; 
                RECT 2.880 168.440 59.280 168.760 ; 
                RECT 69.160 168.440 79.000 168.760 ; 
                RECT 415.280 168.440 420.000 168.760 ; 
                RECT 2.880 169.800 14.400 170.120 ; 
                RECT 19.520 169.800 32.760 170.120 ; 
                RECT 38.560 169.800 59.280 170.120 ; 
                RECT 69.160 169.800 79.000 170.120 ; 
                RECT 415.280 169.800 420.000 170.120 ; 
                RECT 2.880 171.160 13.720 171.480 ; 
                RECT 19.520 171.160 32.760 171.480 ; 
                RECT 39.240 171.160 59.280 171.480 ; 
                RECT 69.160 171.160 79.000 171.480 ; 
                RECT 415.280 171.160 420.000 171.480 ; 
                RECT 2.880 172.520 13.040 172.840 ; 
                RECT 19.520 172.520 32.760 172.840 ; 
                RECT 39.240 172.520 59.280 172.840 ; 
                RECT 67.800 172.520 79.000 172.840 ; 
                RECT 415.280 172.520 420.000 172.840 ; 
                RECT 2.880 173.880 12.360 174.200 ; 
                RECT 19.520 173.880 65.400 174.200 ; 
                RECT 69.160 173.880 79.000 174.200 ; 
                RECT 415.280 173.880 420.000 174.200 ; 
                RECT 2.880 175.240 59.280 175.560 ; 
                RECT 69.160 175.240 79.000 175.560 ; 
                RECT 415.280 175.240 420.000 175.560 ; 
                RECT 2.880 176.600 11.680 176.920 ; 
                RECT 19.520 176.600 59.280 176.920 ; 
                RECT 69.160 176.600 79.000 176.920 ; 
                RECT 415.280 176.600 420.000 176.920 ; 
                RECT 2.880 177.960 11.000 178.280 ; 
                RECT 19.520 177.960 59.280 178.280 ; 
                RECT 69.160 177.960 79.000 178.280 ; 
                RECT 415.280 177.960 420.000 178.280 ; 
                RECT 2.880 179.320 10.320 179.640 ; 
                RECT 19.520 179.320 59.280 179.640 ; 
                RECT 69.160 179.320 79.000 179.640 ; 
                RECT 415.280 179.320 420.000 179.640 ; 
                RECT 2.880 180.680 79.000 181.000 ; 
                RECT 415.280 180.680 420.000 181.000 ; 
                RECT 2.880 182.040 9.640 182.360 ; 
                RECT 19.520 182.040 32.760 182.360 ; 
                RECT 35.840 182.040 60.640 182.360 ; 
                RECT 69.160 182.040 79.000 182.360 ; 
                RECT 415.280 182.040 420.000 182.360 ; 
                RECT 2.880 183.400 64.040 183.720 ; 
                RECT 69.160 183.400 79.000 183.720 ; 
                RECT 415.280 183.400 420.000 183.720 ; 
                RECT 2.880 184.760 64.720 185.080 ; 
                RECT 69.160 184.760 79.000 185.080 ; 
                RECT 415.280 184.760 420.000 185.080 ; 
                RECT 2.880 186.120 60.640 186.440 ; 
                RECT 69.160 186.120 79.000 186.440 ; 
                RECT 415.280 186.120 420.000 186.440 ; 
                RECT 2.880 187.480 60.640 187.800 ; 
                RECT 69.160 187.480 79.000 187.800 ; 
                RECT 415.280 187.480 420.000 187.800 ; 
                RECT 2.880 188.840 37.520 189.160 ; 
                RECT 46.720 188.840 79.000 189.160 ; 
                RECT 415.280 188.840 420.000 189.160 ; 
                RECT 2.880 190.200 36.160 190.520 ; 
                RECT 45.360 190.200 60.640 190.520 ; 
                RECT 69.160 190.200 79.000 190.520 ; 
                RECT 415.280 190.200 420.000 190.520 ; 
                RECT 2.880 191.560 34.800 191.880 ; 
                RECT 44.680 191.560 59.280 191.880 ; 
                RECT 69.160 191.560 79.000 191.880 ; 
                RECT 415.280 191.560 420.000 191.880 ; 
                RECT 2.880 192.920 59.280 193.240 ; 
                RECT 69.160 192.920 79.000 193.240 ; 
                RECT 415.280 192.920 420.000 193.240 ; 
                RECT 2.880 194.280 59.280 194.600 ; 
                RECT 69.160 194.280 79.000 194.600 ; 
                RECT 415.280 194.280 420.000 194.600 ; 
                RECT 2.880 195.640 59.280 195.960 ; 
                RECT 69.160 195.640 79.000 195.960 ; 
                RECT 415.280 195.640 420.000 195.960 ; 
                RECT 2.880 197.000 79.000 197.320 ; 
                RECT 415.280 197.000 420.000 197.320 ; 
                RECT 2.880 198.360 59.280 198.680 ; 
                RECT 69.160 198.360 79.000 198.680 ; 
                RECT 415.280 198.360 420.000 198.680 ; 
                RECT 2.880 199.720 59.280 200.040 ; 
                RECT 69.160 199.720 79.000 200.040 ; 
                RECT 415.280 199.720 420.000 200.040 ; 
                RECT 2.880 201.080 59.280 201.400 ; 
                RECT 69.160 201.080 79.000 201.400 ; 
                RECT 415.280 201.080 420.000 201.400 ; 
                RECT 2.880 202.440 59.280 202.760 ; 
                RECT 69.160 202.440 79.000 202.760 ; 
                RECT 415.280 202.440 420.000 202.760 ; 
                RECT 2.880 203.800 59.280 204.120 ; 
                RECT 63.040 203.800 79.000 204.120 ; 
                RECT 415.280 203.800 420.000 204.120 ; 
                RECT 2.880 205.160 65.400 205.480 ; 
                RECT 69.160 205.160 79.000 205.480 ; 
                RECT 415.280 205.160 420.000 205.480 ; 
                RECT 2.880 206.520 59.280 206.840 ; 
                RECT 69.160 206.520 79.000 206.840 ; 
                RECT 415.280 206.520 420.000 206.840 ; 
                RECT 2.880 207.880 59.280 208.200 ; 
                RECT 69.160 207.880 79.000 208.200 ; 
                RECT 415.280 207.880 420.000 208.200 ; 
                RECT 2.880 209.240 59.280 209.560 ; 
                RECT 69.160 209.240 79.000 209.560 ; 
                RECT 415.280 209.240 420.000 209.560 ; 
                RECT 2.880 210.600 59.280 210.920 ; 
                RECT 69.160 210.600 79.000 210.920 ; 
                RECT 415.280 210.600 420.000 210.920 ; 
                RECT 2.880 211.960 59.280 212.280 ; 
                RECT 63.720 211.960 79.000 212.280 ; 
                RECT 415.280 211.960 420.000 212.280 ; 
                RECT 2.880 213.320 63.360 213.640 ; 
                RECT 69.160 213.320 79.000 213.640 ; 
                RECT 415.280 213.320 420.000 213.640 ; 
                RECT 2.880 214.680 59.280 215.000 ; 
                RECT 69.160 214.680 79.000 215.000 ; 
                RECT 415.280 214.680 420.000 215.000 ; 
                RECT 2.880 216.040 59.280 216.360 ; 
                RECT 69.160 216.040 79.000 216.360 ; 
                RECT 415.280 216.040 420.000 216.360 ; 
                RECT 2.880 217.400 59.280 217.720 ; 
                RECT 69.160 217.400 79.000 217.720 ; 
                RECT 415.280 217.400 420.000 217.720 ; 
                RECT 2.880 218.760 59.280 219.080 ; 
                RECT 69.160 218.760 79.000 219.080 ; 
                RECT 415.280 218.760 420.000 219.080 ; 
                RECT 2.880 220.120 79.000 220.440 ; 
                RECT 415.280 220.120 420.000 220.440 ; 
                RECT 2.880 221.480 62.000 221.800 ; 
                RECT 69.160 221.480 79.000 221.800 ; 
                RECT 415.280 221.480 420.000 221.800 ; 
                RECT 2.880 222.840 66.080 223.160 ; 
                RECT 69.160 222.840 79.000 223.160 ; 
                RECT 415.280 222.840 420.000 223.160 ; 
                RECT 2.880 224.200 62.000 224.520 ; 
                RECT 69.160 224.200 79.000 224.520 ; 
                RECT 415.280 224.200 420.000 224.520 ; 
                RECT 2.880 225.560 62.000 225.880 ; 
                RECT 69.160 225.560 79.000 225.880 ; 
                RECT 415.280 225.560 420.000 225.880 ; 
                RECT 2.880 226.920 62.000 227.240 ; 
                RECT 69.160 226.920 79.000 227.240 ; 
                RECT 415.280 226.920 420.000 227.240 ; 
                RECT 2.880 228.280 79.000 228.600 ; 
                RECT 415.280 228.280 420.000 228.600 ; 
                RECT 2.880 229.640 62.000 229.960 ; 
                RECT 69.160 229.640 79.000 229.960 ; 
                RECT 415.280 229.640 420.000 229.960 ; 
                RECT 2.880 231.000 62.000 231.320 ; 
                RECT 69.160 231.000 79.000 231.320 ; 
                RECT 415.280 231.000 420.000 231.320 ; 
                RECT 2.880 232.360 64.720 232.680 ; 
                RECT 69.160 232.360 79.000 232.680 ; 
                RECT 415.280 232.360 420.000 232.680 ; 
                RECT 2.880 233.720 65.400 234.040 ; 
                RECT 69.160 233.720 79.000 234.040 ; 
                RECT 415.280 233.720 420.000 234.040 ; 
                RECT 2.880 235.080 62.000 235.400 ; 
                RECT 69.160 235.080 79.000 235.400 ; 
                RECT 415.280 235.080 420.000 235.400 ; 
                RECT 2.880 236.440 79.000 236.760 ; 
                RECT 415.280 236.440 420.000 236.760 ; 
                RECT 2.880 237.800 62.000 238.120 ; 
                RECT 69.160 237.800 79.000 238.120 ; 
                RECT 415.280 237.800 420.000 238.120 ; 
                RECT 2.880 239.160 62.000 239.480 ; 
                RECT 69.160 239.160 79.000 239.480 ; 
                RECT 415.280 239.160 420.000 239.480 ; 
                RECT 2.880 240.520 62.000 240.840 ; 
                RECT 69.160 240.520 79.000 240.840 ; 
                RECT 415.280 240.520 420.000 240.840 ; 
                RECT 2.880 241.880 62.000 242.200 ; 
                RECT 69.160 241.880 79.000 242.200 ; 
                RECT 415.280 241.880 420.000 242.200 ; 
                RECT 2.880 243.240 79.000 243.560 ; 
                RECT 415.280 243.240 420.000 243.560 ; 
                RECT 2.880 244.600 63.360 244.920 ; 
                RECT 69.160 244.600 79.000 244.920 ; 
                RECT 415.280 244.600 420.000 244.920 ; 
                RECT 2.880 245.960 62.680 246.280 ; 
                RECT 69.160 245.960 79.000 246.280 ; 
                RECT 415.280 245.960 420.000 246.280 ; 
                RECT 2.880 247.320 62.680 247.640 ; 
                RECT 69.160 247.320 79.000 247.640 ; 
                RECT 415.280 247.320 420.000 247.640 ; 
                RECT 2.880 248.680 62.680 249.000 ; 
                RECT 69.160 248.680 79.000 249.000 ; 
                RECT 415.280 248.680 420.000 249.000 ; 
                RECT 2.880 250.040 62.680 250.360 ; 
                RECT 69.160 250.040 79.000 250.360 ; 
                RECT 415.280 250.040 420.000 250.360 ; 
                RECT 2.880 251.400 79.000 251.720 ; 
                RECT 415.280 251.400 420.000 251.720 ; 
                RECT 2.880 252.760 65.400 253.080 ; 
                RECT 69.160 252.760 79.000 253.080 ; 
                RECT 415.280 252.760 420.000 253.080 ; 
                RECT 2.880 254.120 62.680 254.440 ; 
                RECT 69.160 254.120 79.000 254.440 ; 
                RECT 415.280 254.120 420.000 254.440 ; 
                RECT 2.880 255.480 62.680 255.800 ; 
                RECT 69.160 255.480 79.000 255.800 ; 
                RECT 415.280 255.480 420.000 255.800 ; 
                RECT 2.880 256.840 62.680 257.160 ; 
                RECT 69.160 256.840 79.000 257.160 ; 
                RECT 415.280 256.840 420.000 257.160 ; 
                RECT 2.880 258.200 62.680 258.520 ; 
                RECT 69.160 258.200 79.000 258.520 ; 
                RECT 415.280 258.200 420.000 258.520 ; 
                RECT 2.880 259.560 79.000 259.880 ; 
                RECT 415.280 259.560 420.000 259.880 ; 
                RECT 2.880 260.920 63.360 261.240 ; 
                RECT 69.160 260.920 79.000 261.240 ; 
                RECT 415.280 260.920 420.000 261.240 ; 
                RECT 2.880 262.280 64.040 262.600 ; 
                RECT 69.160 262.280 79.000 262.600 ; 
                RECT 415.280 262.280 420.000 262.600 ; 
                RECT 2.880 263.640 63.360 263.960 ; 
                RECT 69.160 263.640 79.000 263.960 ; 
                RECT 415.280 263.640 420.000 263.960 ; 
                RECT 2.880 265.000 63.360 265.320 ; 
                RECT 69.160 265.000 79.000 265.320 ; 
                RECT 415.280 265.000 420.000 265.320 ; 
                RECT 2.880 266.360 63.360 266.680 ; 
                RECT 69.160 266.360 79.000 266.680 ; 
                RECT 415.280 266.360 420.000 266.680 ; 
                RECT 2.880 267.720 79.000 268.040 ; 
                RECT 415.280 267.720 420.000 268.040 ; 
                RECT 2.880 269.080 63.360 269.400 ; 
                RECT 69.160 269.080 79.000 269.400 ; 
                RECT 415.280 269.080 420.000 269.400 ; 
                RECT 2.880 270.440 63.360 270.760 ; 
                RECT 69.160 270.440 79.000 270.760 ; 
                RECT 415.280 270.440 420.000 270.760 ; 
                RECT 2.880 271.800 66.760 272.120 ; 
                RECT 69.160 271.800 79.000 272.120 ; 
                RECT 415.280 271.800 420.000 272.120 ; 
                RECT 2.880 273.160 63.360 273.480 ; 
                RECT 69.160 273.160 79.000 273.480 ; 
                RECT 415.280 273.160 420.000 273.480 ; 
                RECT 2.880 274.520 63.360 274.840 ; 
                RECT 69.160 274.520 79.000 274.840 ; 
                RECT 415.280 274.520 420.000 274.840 ; 
                RECT 2.880 275.880 79.000 276.200 ; 
                RECT 415.280 275.880 420.000 276.200 ; 
                RECT 2.880 277.240 200.720 277.560 ; 
                RECT 415.280 277.240 420.000 277.560 ; 
                RECT 2.880 278.600 200.720 278.920 ; 
                RECT 415.280 278.600 420.000 278.920 ; 
                RECT 2.880 279.960 200.720 280.280 ; 
                RECT 415.280 279.960 420.000 280.280 ; 
                RECT 2.880 281.320 420.000 281.640 ; 
                RECT 2.880 282.680 420.000 283.000 ; 
                RECT 2.880 284.040 420.000 284.360 ; 
                RECT 2.880 285.400 420.000 285.720 ; 
                RECT 2.880 2.880 420.000 4.240 ; 
                RECT 2.880 287.400 420.000 288.760 ; 
                RECT 204.860 29.630 210.660 30.750 ; 
                RECT 405.560 29.630 411.360 30.750 ; 
                RECT 204.860 35.495 210.660 36.265 ; 
                RECT 405.560 35.495 411.360 36.265 ; 
                RECT 204.860 41.530 210.660 42.230 ; 
                RECT 405.560 41.530 411.360 42.230 ; 
                RECT 204.860 47.120 210.660 47.820 ; 
                RECT 405.560 47.120 411.360 47.820 ; 
                RECT 204.860 78.350 411.360 79.150 ; 
                RECT 204.860 73.460 411.360 74.260 ; 
                RECT 204.860 102.695 411.360 102.985 ; 
                RECT 204.860 81.590 411.360 83.680 ; 
                RECT 204.860 120.970 411.360 122.375 ; 
                RECT 204.860 70.450 411.360 71.250 ; 
                RECT 204.860 61.400 411.360 63.200 ; 
                RECT 204.860 75.140 411.360 75.940 ; 
                RECT 204.860 20.260 411.360 22.060 ; 
                RECT 79.885 148.435 81.205 276.415 ; 
                RECT 90.430 148.435 92.350 276.415 ; 
                RECT 108.170 148.435 110.090 276.415 ; 
                RECT 112.010 148.435 113.930 276.415 ; 
                RECT 141.190 148.435 143.110 276.415 ; 
                RECT 145.030 148.435 146.950 276.415 ; 
                RECT 148.870 148.435 150.790 276.415 ; 
                RECT 152.710 148.435 154.630 276.415 ; 
                RECT 138.600 57.135 139.490 101.135 ; 
                RECT 144.930 57.135 145.820 101.135 ; 
                RECT 151.690 57.135 152.580 101.135 ; 
                RECT 158.340 57.135 159.880 101.135 ; 
                RECT 170.070 57.135 171.990 101.135 ; 
                RECT 155.970 129.320 156.860 141.800 ; 
                RECT 162.300 129.320 163.190 141.800 ; 
                RECT 170.265 129.320 172.185 141.800 ; 
                RECT 155.645 115.000 156.755 123.320 ; 
                RECT 164.020 115.000 164.910 123.320 ; 
                RECT 171.770 115.000 173.690 123.320 ; 
                RECT 180.365 47.555 181.475 51.135 ; 
                RECT 24.710 149.500 33.870 149.870 ; 
                RECT 24.710 152.835 33.870 153.725 ; 
                RECT 62.770 135.860 80.010 136.530 ; 
                RECT 62.770 137.160 80.010 138.170 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 422.880 291.640 ; 
        LAYER met2 ;
            RECT 0.000 0.000 422.880 291.640 ; 
    END 
END sram22_256x32m4w8 
END LIBRARY 

