VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_128x24m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_128x24m4w8   ;
    SIZE 305.240 BY 224.320 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 145.270 0.000 145.410 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 151.370 0.000 151.510 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 157.470 0.000 157.610 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.570 0.000 163.710 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 169.670 0.000 169.810 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 175.770 0.000 175.910 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 181.870 0.000 182.010 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 187.970 0.000 188.110 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.070 0.000 194.210 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 200.170 0.000 200.310 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 206.270 0.000 206.410 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 212.370 0.000 212.510 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 218.470 0.000 218.610 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 224.570 0.000 224.710 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 230.670 0.000 230.810 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 236.770 0.000 236.910 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 242.870 0.000 243.010 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 248.970 0.000 249.110 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 255.070 0.000 255.210 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 261.170 0.000 261.310 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 267.270 0.000 267.410 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 273.370 0.000 273.510 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 279.470 0.000 279.610 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 285.570 0.000 285.710 0.140 ; 
        END 
    END dout[23] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 144.850 0.000 144.990 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 150.950 0.000 151.090 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 157.050 0.000 157.190 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.150 0.000 163.290 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 169.250 0.000 169.390 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 175.350 0.000 175.490 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 181.450 0.000 181.590 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 187.550 0.000 187.690 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 193.650 0.000 193.790 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 199.750 0.000 199.890 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 205.850 0.000 205.990 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 211.950 0.000 212.090 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 218.050 0.000 218.190 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 224.150 0.000 224.290 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 230.250 0.000 230.390 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 236.350 0.000 236.490 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 242.450 0.000 242.590 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 248.550 0.000 248.690 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 254.650 0.000 254.790 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 260.750 0.000 260.890 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 266.850 0.000 266.990 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 272.950 0.000 273.090 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 279.050 0.000 279.190 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 285.150 0.000 285.290 0.140 ; 
        END 
    END din[23] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 144.500 0.000 144.640 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 193.300 0.000 193.440 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 242.100 0.000 242.240 0.140 ; 
        END 
    END wmask[2] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 103.160 0.000 103.480 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 97.040 0.000 97.360 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 90.920 0.000 91.240 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 84.800 0.000 85.120 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 78.680 0.000 79.000 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 72.560 0.000 72.880 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 66.440 0.000 66.760 0.320 ; 
        END 
    END addr[6] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 115.400 0.000 115.720 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 109.280 0.000 109.600 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 17.298000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 118.120 0.000 118.440 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 21.204000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 118.800 0.000 119.120 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 144.280 6.240 ; 
                RECT 146.000 5.920 150.400 6.240 ; 
                RECT 152.120 5.920 156.520 6.240 ; 
                RECT 158.240 5.920 162.640 6.240 ; 
                RECT 164.360 5.920 168.760 6.240 ; 
                RECT 170.480 5.920 174.880 6.240 ; 
                RECT 176.600 5.920 181.000 6.240 ; 
                RECT 182.720 5.920 187.120 6.240 ; 
                RECT 188.840 5.920 193.240 6.240 ; 
                RECT 194.960 5.920 199.360 6.240 ; 
                RECT 201.080 5.920 205.480 6.240 ; 
                RECT 207.200 5.920 211.600 6.240 ; 
                RECT 213.320 5.920 217.720 6.240 ; 
                RECT 219.440 5.920 223.840 6.240 ; 
                RECT 225.560 5.920 229.960 6.240 ; 
                RECT 231.680 5.920 236.080 6.240 ; 
                RECT 237.800 5.920 242.200 6.240 ; 
                RECT 243.920 5.920 248.320 6.240 ; 
                RECT 250.040 5.920 254.440 6.240 ; 
                RECT 256.160 5.920 260.560 6.240 ; 
                RECT 262.280 5.920 266.680 6.240 ; 
                RECT 268.400 5.920 272.800 6.240 ; 
                RECT 274.520 5.920 278.920 6.240 ; 
                RECT 280.640 5.920 285.040 6.240 ; 
                RECT 286.080 5.920 305.080 6.240 ; 
                RECT 0.160 7.280 305.080 7.600 ; 
                RECT 0.160 8.640 305.080 8.960 ; 
                RECT 0.160 10.000 117.760 10.320 ; 
                RECT 140.560 10.000 305.080 10.320 ; 
                RECT 0.160 11.360 305.080 11.680 ; 
                RECT 0.160 12.720 305.080 13.040 ; 
                RECT 0.160 14.080 62.680 14.400 ; 
                RECT 119.480 14.080 305.080 14.400 ; 
                RECT 0.160 15.440 305.080 15.760 ; 
                RECT 0.160 16.800 305.080 17.120 ; 
                RECT 0.160 18.160 62.680 18.480 ; 
                RECT 118.800 18.160 143.600 18.480 ; 
                RECT 243.240 18.160 305.080 18.480 ; 
                RECT 0.160 19.520 134.080 19.840 ; 
                RECT 294.920 19.520 305.080 19.840 ; 
                RECT 0.160 20.880 134.080 21.200 ; 
                RECT 294.920 20.880 305.080 21.200 ; 
                RECT 0.160 22.240 134.080 22.560 ; 
                RECT 294.920 22.240 305.080 22.560 ; 
                RECT 0.160 23.600 134.080 23.920 ; 
                RECT 294.920 23.600 305.080 23.920 ; 
                RECT 0.160 24.960 134.080 25.280 ; 
                RECT 294.920 24.960 305.080 25.280 ; 
                RECT 0.160 26.320 134.080 26.640 ; 
                RECT 294.920 26.320 305.080 26.640 ; 
                RECT 0.160 27.680 134.080 28.000 ; 
                RECT 294.920 27.680 305.080 28.000 ; 
                RECT 0.160 29.040 134.080 29.360 ; 
                RECT 294.920 29.040 305.080 29.360 ; 
                RECT 0.160 30.400 134.080 30.720 ; 
                RECT 294.920 30.400 305.080 30.720 ; 
                RECT 0.160 31.760 134.080 32.080 ; 
                RECT 294.920 31.760 305.080 32.080 ; 
                RECT 0.160 33.120 83.080 33.440 ; 
                RECT 96.360 33.120 134.080 33.440 ; 
                RECT 294.920 33.120 305.080 33.440 ; 
                RECT 0.160 34.480 81.720 34.800 ; 
                RECT 102.480 34.480 134.080 34.800 ; 
                RECT 294.920 34.480 305.080 34.800 ; 
                RECT 0.160 35.840 62.000 36.160 ; 
                RECT 119.480 35.840 134.080 36.160 ; 
                RECT 294.920 35.840 305.080 36.160 ; 
                RECT 0.160 37.200 61.320 37.520 ; 
                RECT 115.400 37.200 133.400 37.520 ; 
                RECT 294.920 37.200 305.080 37.520 ; 
                RECT 0.160 38.560 134.080 38.880 ; 
                RECT 294.920 38.560 305.080 38.880 ; 
                RECT 0.160 39.920 134.080 40.240 ; 
                RECT 294.920 39.920 305.080 40.240 ; 
                RECT 0.160 41.280 134.080 41.600 ; 
                RECT 294.920 41.280 305.080 41.600 ; 
                RECT 0.160 42.640 134.080 42.960 ; 
                RECT 294.920 42.640 305.080 42.960 ; 
                RECT 0.160 44.000 57.240 44.320 ; 
                RECT 68.480 44.000 134.080 44.320 ; 
                RECT 294.920 44.000 305.080 44.320 ; 
                RECT 0.160 45.360 58.600 45.680 ; 
                RECT 64.400 45.360 72.200 45.680 ; 
                RECT 74.600 45.360 134.080 45.680 ; 
                RECT 294.920 45.360 305.080 45.680 ; 
                RECT 0.160 46.720 59.960 47.040 ; 
                RECT 63.720 46.720 134.080 47.040 ; 
                RECT 294.920 46.720 305.080 47.040 ; 
                RECT 0.160 48.080 134.080 48.400 ; 
                RECT 294.920 48.080 305.080 48.400 ; 
                RECT 0.160 49.440 66.760 49.760 ; 
                RECT 75.280 49.440 134.080 49.760 ; 
                RECT 294.920 49.440 305.080 49.760 ; 
                RECT 0.160 50.800 59.280 51.120 ; 
                RECT 68.480 50.800 134.080 51.120 ; 
                RECT 294.920 50.800 305.080 51.120 ; 
                RECT 0.160 52.160 62.680 52.480 ; 
                RECT 67.800 52.160 134.080 52.480 ; 
                RECT 294.920 52.160 305.080 52.480 ; 
                RECT 0.160 53.520 134.080 53.840 ; 
                RECT 294.920 53.520 305.080 53.840 ; 
                RECT 0.160 54.880 58.600 55.200 ; 
                RECT 68.480 54.880 110.960 55.200 ; 
                RECT 117.440 54.880 134.080 55.200 ; 
                RECT 294.920 54.880 305.080 55.200 ; 
                RECT 0.160 56.240 65.400 56.560 ; 
                RECT 74.600 56.240 110.960 56.560 ; 
                RECT 117.440 56.240 134.080 56.560 ; 
                RECT 294.920 56.240 305.080 56.560 ; 
                RECT 0.160 57.600 110.960 57.920 ; 
                RECT 294.920 57.600 305.080 57.920 ; 
                RECT 0.160 58.960 66.760 59.280 ; 
                RECT 72.560 58.960 110.960 59.280 ; 
                RECT 117.440 58.960 134.080 59.280 ; 
                RECT 294.920 58.960 305.080 59.280 ; 
                RECT 0.160 60.320 69.480 60.640 ; 
                RECT 74.600 60.320 134.080 60.640 ; 
                RECT 294.920 60.320 305.080 60.640 ; 
                RECT 0.160 61.680 63.360 62.000 ; 
                RECT 68.480 61.680 134.080 62.000 ; 
                RECT 294.920 61.680 305.080 62.000 ; 
                RECT 0.160 63.040 134.080 63.360 ; 
                RECT 294.920 63.040 305.080 63.360 ; 
                RECT 0.160 64.400 57.240 64.720 ; 
                RECT 117.440 64.400 134.080 64.720 ; 
                RECT 294.920 64.400 305.080 64.720 ; 
                RECT 0.160 65.760 66.760 66.080 ; 
                RECT 74.600 65.760 82.400 66.080 ; 
                RECT 86.840 65.760 92.600 66.080 ; 
                RECT 117.440 65.760 134.080 66.080 ; 
                RECT 294.920 65.760 305.080 66.080 ; 
                RECT 0.160 67.120 65.400 67.440 ; 
                RECT 68.480 67.120 75.600 67.440 ; 
                RECT 82.080 67.120 83.760 67.440 ; 
                RECT 86.160 67.120 92.600 67.440 ; 
                RECT 126.280 67.120 134.080 67.440 ; 
                RECT 294.920 67.120 305.080 67.440 ; 
                RECT 0.160 68.480 57.240 68.800 ; 
                RECT 71.200 68.480 92.600 68.800 ; 
                RECT 126.280 68.480 134.080 68.800 ; 
                RECT 294.920 68.480 305.080 68.800 ; 
                RECT 0.160 69.840 66.080 70.160 ; 
                RECT 74.600 69.840 92.600 70.160 ; 
                RECT 124.920 69.840 134.080 70.160 ; 
                RECT 294.920 69.840 305.080 70.160 ; 
                RECT 0.160 71.200 64.040 71.520 ; 
                RECT 67.800 71.200 92.600 71.520 ; 
                RECT 126.280 71.200 134.080 71.520 ; 
                RECT 294.920 71.200 305.080 71.520 ; 
                RECT 0.160 72.560 59.280 72.880 ; 
                RECT 63.720 72.560 66.760 72.880 ; 
                RECT 75.280 72.560 92.600 72.880 ; 
                RECT 129.000 72.560 134.080 72.880 ; 
                RECT 294.920 72.560 305.080 72.880 ; 
                RECT 0.160 73.920 62.000 74.240 ; 
                RECT 65.760 73.920 92.600 74.240 ; 
                RECT 117.440 73.920 134.080 74.240 ; 
                RECT 294.920 73.920 305.080 74.240 ; 
                RECT 0.160 75.280 58.600 75.600 ; 
                RECT 62.360 75.280 92.600 75.600 ; 
                RECT 129.000 75.280 134.080 75.600 ; 
                RECT 294.920 75.280 305.080 75.600 ; 
                RECT 0.160 76.640 62.680 76.960 ; 
                RECT 68.480 76.640 92.600 76.960 ; 
                RECT 127.640 76.640 134.080 76.960 ; 
                RECT 294.920 76.640 305.080 76.960 ; 
                RECT 0.160 78.000 58.600 78.320 ; 
                RECT 73.920 78.000 92.600 78.320 ; 
                RECT 129.000 78.000 134.080 78.320 ; 
                RECT 294.920 78.000 305.080 78.320 ; 
                RECT 0.160 79.360 92.600 79.680 ; 
                RECT 131.720 79.360 134.080 79.680 ; 
                RECT 294.920 79.360 305.080 79.680 ; 
                RECT 0.160 80.720 65.400 81.040 ; 
                RECT 67.800 80.720 92.600 81.040 ; 
                RECT 131.720 80.720 134.080 81.040 ; 
                RECT 294.920 80.720 305.080 81.040 ; 
                RECT 0.160 82.080 66.760 82.400 ; 
                RECT 68.480 82.080 92.600 82.400 ; 
                RECT 130.360 82.080 134.080 82.400 ; 
                RECT 294.920 82.080 305.080 82.400 ; 
                RECT 0.160 83.440 57.240 83.760 ; 
                RECT 67.800 83.440 92.600 83.760 ; 
                RECT 117.440 83.440 134.080 83.760 ; 
                RECT 294.920 83.440 305.080 83.760 ; 
                RECT 0.160 84.800 62.680 85.120 ; 
                RECT 74.600 84.800 92.600 85.120 ; 
                RECT 130.360 84.800 134.080 85.120 ; 
                RECT 294.920 84.800 305.080 85.120 ; 
                RECT 0.160 86.160 57.240 86.480 ; 
                RECT 68.480 86.160 92.600 86.480 ; 
                RECT 294.920 86.160 305.080 86.480 ; 
                RECT 0.160 87.520 66.080 87.840 ; 
                RECT 68.480 87.520 92.600 87.840 ; 
                RECT 294.920 87.520 305.080 87.840 ; 
                RECT 0.160 88.880 92.600 89.200 ; 
                RECT 294.920 88.880 305.080 89.200 ; 
                RECT 0.160 90.240 92.600 90.560 ; 
                RECT 294.920 90.240 305.080 90.560 ; 
                RECT 0.160 91.600 53.840 91.920 ; 
                RECT 71.200 91.600 92.600 91.920 ; 
                RECT 117.440 91.600 134.080 91.920 ; 
                RECT 294.920 91.600 305.080 91.920 ; 
                RECT 0.160 92.960 134.080 93.280 ; 
                RECT 294.920 92.960 305.080 93.280 ; 
                RECT 0.160 94.320 134.080 94.640 ; 
                RECT 294.920 94.320 305.080 94.640 ; 
                RECT 0.160 95.680 62.680 96.000 ; 
                RECT 74.600 95.680 134.080 96.000 ; 
                RECT 294.920 95.680 305.080 96.000 ; 
                RECT 0.160 97.040 69.480 97.360 ; 
                RECT 77.320 97.040 134.080 97.360 ; 
                RECT 294.920 97.040 305.080 97.360 ; 
                RECT 0.160 98.400 81.040 98.720 ; 
                RECT 92.960 98.400 96.000 98.720 ; 
                RECT 116.760 98.400 134.080 98.720 ; 
                RECT 294.920 98.400 305.080 98.720 ; 
                RECT 0.160 99.760 96.000 100.080 ; 
                RECT 116.760 99.760 134.080 100.080 ; 
                RECT 294.920 99.760 305.080 100.080 ; 
                RECT 0.160 101.120 57.240 101.440 ; 
                RECT 62.360 101.120 96.000 101.440 ; 
                RECT 116.760 101.120 134.080 101.440 ; 
                RECT 294.920 101.120 305.080 101.440 ; 
                RECT 0.160 102.480 96.000 102.800 ; 
                RECT 116.760 102.480 134.080 102.800 ; 
                RECT 294.920 102.480 305.080 102.800 ; 
                RECT 0.160 103.840 96.000 104.160 ; 
                RECT 116.760 103.840 134.080 104.160 ; 
                RECT 294.920 103.840 305.080 104.160 ; 
                RECT 0.160 105.200 72.880 105.520 ; 
                RECT 75.280 105.200 96.000 105.520 ; 
                RECT 116.760 105.200 134.080 105.520 ; 
                RECT 294.920 105.200 305.080 105.520 ; 
                RECT 0.160 106.560 96.000 106.880 ; 
                RECT 116.760 106.560 134.080 106.880 ; 
                RECT 294.920 106.560 305.080 106.880 ; 
                RECT 0.160 107.920 96.000 108.240 ; 
                RECT 116.760 107.920 134.080 108.240 ; 
                RECT 294.920 107.920 305.080 108.240 ; 
                RECT 0.160 109.280 96.000 109.600 ; 
                RECT 294.920 109.280 305.080 109.600 ; 
                RECT 0.160 110.640 59.280 110.960 ; 
                RECT 64.400 110.640 96.000 110.960 ; 
                RECT 116.760 110.640 131.360 110.960 ; 
                RECT 294.920 110.640 305.080 110.960 ; 
                RECT 0.160 112.000 96.000 112.320 ; 
                RECT 116.760 112.000 128.640 112.320 ; 
                RECT 294.920 112.000 305.080 112.320 ; 
                RECT 0.160 113.360 35.480 113.680 ; 
                RECT 54.200 113.360 65.400 113.680 ; 
                RECT 74.600 113.360 96.000 113.680 ; 
                RECT 116.760 113.360 125.920 113.680 ; 
                RECT 294.920 113.360 305.080 113.680 ; 
                RECT 0.160 114.720 35.480 115.040 ; 
                RECT 54.200 114.720 123.200 115.040 ; 
                RECT 294.920 114.720 305.080 115.040 ; 
                RECT 0.160 116.080 35.480 116.400 ; 
                RECT 54.200 116.080 62.000 116.400 ; 
                RECT 64.400 116.080 134.080 116.400 ; 
                RECT 294.920 116.080 305.080 116.400 ; 
                RECT 0.160 117.440 35.480 117.760 ; 
                RECT 54.200 117.440 58.600 117.760 ; 
                RECT 61.680 117.440 134.080 117.760 ; 
                RECT 294.920 117.440 305.080 117.760 ; 
                RECT 0.160 118.800 35.480 119.120 ; 
                RECT 54.880 118.800 134.080 119.120 ; 
                RECT 294.920 118.800 305.080 119.120 ; 
                RECT 0.160 120.160 35.480 120.480 ; 
                RECT 54.200 120.160 96.000 120.480 ; 
                RECT 117.440 120.160 134.080 120.480 ; 
                RECT 294.920 120.160 305.080 120.480 ; 
                RECT 0.160 121.520 35.480 121.840 ; 
                RECT 54.200 121.520 96.000 121.840 ; 
                RECT 117.440 121.520 134.080 121.840 ; 
                RECT 294.920 121.520 305.080 121.840 ; 
                RECT 0.160 122.880 35.480 123.200 ; 
                RECT 54.200 122.880 96.000 123.200 ; 
                RECT 117.440 122.880 134.080 123.200 ; 
                RECT 294.920 122.880 305.080 123.200 ; 
                RECT 0.160 124.240 35.480 124.560 ; 
                RECT 54.200 124.240 96.000 124.560 ; 
                RECT 117.440 124.240 124.560 124.560 ; 
                RECT 294.920 124.240 305.080 124.560 ; 
                RECT 0.160 125.600 35.480 125.920 ; 
                RECT 54.200 125.600 96.000 125.920 ; 
                RECT 117.440 125.600 127.280 125.920 ; 
                RECT 294.920 125.600 305.080 125.920 ; 
                RECT 0.160 126.960 35.480 127.280 ; 
                RECT 54.200 126.960 60.640 127.280 ; 
                RECT 64.400 126.960 96.000 127.280 ; 
                RECT 117.440 126.960 130.000 127.280 ; 
                RECT 294.920 126.960 305.080 127.280 ; 
                RECT 0.160 128.320 96.000 128.640 ; 
                RECT 117.440 128.320 132.720 128.640 ; 
                RECT 294.920 128.320 305.080 128.640 ; 
                RECT 0.160 129.680 96.000 130.000 ; 
                RECT 294.920 129.680 305.080 130.000 ; 
                RECT 0.160 131.040 19.160 131.360 ; 
                RECT 35.840 131.040 62.680 131.360 ; 
                RECT 68.480 131.040 96.000 131.360 ; 
                RECT 117.440 131.040 134.080 131.360 ; 
                RECT 294.920 131.040 305.080 131.360 ; 
                RECT 0.160 132.400 19.160 132.720 ; 
                RECT 35.840 132.400 41.600 132.720 ; 
                RECT 48.760 132.400 96.000 132.720 ; 
                RECT 117.440 132.400 134.080 132.720 ; 
                RECT 294.920 132.400 305.080 132.720 ; 
                RECT 0.160 133.760 19.160 134.080 ; 
                RECT 53.520 133.760 96.000 134.080 ; 
                RECT 117.440 133.760 134.080 134.080 ; 
                RECT 294.920 133.760 305.080 134.080 ; 
                RECT 0.160 135.120 19.160 135.440 ; 
                RECT 53.520 135.120 96.000 135.440 ; 
                RECT 294.920 135.120 305.080 135.440 ; 
                RECT 0.160 136.480 19.160 136.800 ; 
                RECT 35.840 136.480 41.600 136.800 ; 
                RECT 48.760 136.480 57.240 136.800 ; 
                RECT 67.120 136.480 96.000 136.800 ; 
                RECT 117.440 136.480 120.480 136.800 ; 
                RECT 294.920 136.480 305.080 136.800 ; 
                RECT 0.160 137.840 19.840 138.160 ; 
                RECT 48.080 137.840 96.000 138.160 ; 
                RECT 117.440 137.840 305.080 138.160 ; 
                RECT 0.160 139.200 47.720 139.520 ; 
                RECT 93.640 139.200 305.080 139.520 ; 
                RECT 0.160 140.560 131.360 140.880 ; 
                RECT 297.640 140.560 305.080 140.880 ; 
                RECT 0.160 141.920 131.360 142.240 ; 
                RECT 297.640 141.920 305.080 142.240 ; 
                RECT 0.160 143.280 131.360 143.600 ; 
                RECT 297.640 143.280 305.080 143.600 ; 
                RECT 0.160 144.640 25.280 144.960 ; 
                RECT 31.760 144.640 33.440 144.960 ; 
                RECT 44.680 144.640 76.960 144.960 ; 
                RECT 297.640 144.640 305.080 144.960 ; 
                RECT 0.160 146.000 23.240 146.320 ; 
                RECT 44.000 146.000 57.920 146.320 ; 
                RECT 63.720 146.000 76.960 146.320 ; 
                RECT 297.640 146.000 305.080 146.320 ; 
                RECT 0.160 147.360 23.240 147.680 ; 
                RECT 42.640 147.360 55.880 147.680 ; 
                RECT 63.720 147.360 76.960 147.680 ; 
                RECT 297.640 147.360 305.080 147.680 ; 
                RECT 0.160 148.720 23.240 149.040 ; 
                RECT 33.800 148.720 55.880 149.040 ; 
                RECT 59.640 148.720 76.960 149.040 ; 
                RECT 297.640 148.720 305.080 149.040 ; 
                RECT 0.160 150.080 55.880 150.400 ; 
                RECT 63.720 150.080 76.960 150.400 ; 
                RECT 297.640 150.080 305.080 150.400 ; 
                RECT 0.160 151.440 23.240 151.760 ; 
                RECT 33.800 151.440 55.880 151.760 ; 
                RECT 63.720 151.440 76.960 151.760 ; 
                RECT 297.640 151.440 305.080 151.760 ; 
                RECT 0.160 152.800 23.240 153.120 ; 
                RECT 33.800 152.800 76.960 153.120 ; 
                RECT 297.640 152.800 305.080 153.120 ; 
                RECT 0.160 154.160 59.960 154.480 ; 
                RECT 63.720 154.160 76.960 154.480 ; 
                RECT 297.640 154.160 305.080 154.480 ; 
                RECT 0.160 155.520 55.880 155.840 ; 
                RECT 63.720 155.520 76.960 155.840 ; 
                RECT 297.640 155.520 305.080 155.840 ; 
                RECT 0.160 156.880 16.440 157.200 ; 
                RECT 18.840 156.880 55.880 157.200 ; 
                RECT 63.720 156.880 76.960 157.200 ; 
                RECT 297.640 156.880 305.080 157.200 ; 
                RECT 0.160 158.240 55.880 158.560 ; 
                RECT 57.600 158.240 76.960 158.560 ; 
                RECT 297.640 158.240 305.080 158.560 ; 
                RECT 0.160 159.600 15.760 159.920 ; 
                RECT 18.840 159.600 32.080 159.920 ; 
                RECT 35.160 159.600 55.880 159.920 ; 
                RECT 63.720 159.600 76.960 159.920 ; 
                RECT 297.640 159.600 305.080 159.920 ; 
                RECT 0.160 160.960 15.080 161.280 ; 
                RECT 18.840 160.960 32.080 161.280 ; 
                RECT 35.840 160.960 76.960 161.280 ; 
                RECT 297.640 160.960 305.080 161.280 ; 
                RECT 0.160 162.320 14.400 162.640 ; 
                RECT 18.840 162.320 32.080 162.640 ; 
                RECT 36.520 162.320 57.920 162.640 ; 
                RECT 63.720 162.320 76.960 162.640 ; 
                RECT 297.640 162.320 305.080 162.640 ; 
                RECT 0.160 163.680 55.880 164.000 ; 
                RECT 63.720 163.680 76.960 164.000 ; 
                RECT 297.640 163.680 305.080 164.000 ; 
                RECT 0.160 165.040 13.720 165.360 ; 
                RECT 18.840 165.040 32.080 165.360 ; 
                RECT 37.200 165.040 55.880 165.360 ; 
                RECT 63.720 165.040 76.960 165.360 ; 
                RECT 297.640 165.040 305.080 165.360 ; 
                RECT 0.160 166.400 13.040 166.720 ; 
                RECT 18.840 166.400 55.880 166.720 ; 
                RECT 63.720 166.400 76.960 166.720 ; 
                RECT 297.640 166.400 305.080 166.720 ; 
                RECT 0.160 167.760 12.360 168.080 ; 
                RECT 18.840 167.760 55.880 168.080 ; 
                RECT 62.360 167.760 76.960 168.080 ; 
                RECT 297.640 167.760 305.080 168.080 ; 
                RECT 0.160 169.120 11.680 169.440 ; 
                RECT 18.840 169.120 76.960 169.440 ; 
                RECT 297.640 169.120 305.080 169.440 ; 
                RECT 0.160 170.480 55.880 170.800 ; 
                RECT 63.720 170.480 76.960 170.800 ; 
                RECT 297.640 170.480 305.080 170.800 ; 
                RECT 0.160 171.840 11.000 172.160 ; 
                RECT 18.840 171.840 55.880 172.160 ; 
                RECT 63.720 171.840 76.960 172.160 ; 
                RECT 297.640 171.840 305.080 172.160 ; 
                RECT 0.160 173.200 10.320 173.520 ; 
                RECT 18.840 173.200 55.880 173.520 ; 
                RECT 63.720 173.200 76.960 173.520 ; 
                RECT 297.640 173.200 305.080 173.520 ; 
                RECT 0.160 174.560 55.880 174.880 ; 
                RECT 63.720 174.560 76.960 174.880 ; 
                RECT 297.640 174.560 305.080 174.880 ; 
                RECT 0.160 175.920 55.880 176.240 ; 
                RECT 63.040 175.920 76.960 176.240 ; 
                RECT 297.640 175.920 305.080 176.240 ; 
                RECT 0.160 177.280 57.920 177.600 ; 
                RECT 63.720 177.280 76.960 177.600 ; 
                RECT 297.640 177.280 305.080 177.600 ; 
                RECT 0.160 178.640 76.960 178.960 ; 
                RECT 297.640 178.640 305.080 178.960 ; 
                RECT 0.160 180.000 58.600 180.320 ; 
                RECT 63.720 180.000 76.960 180.320 ; 
                RECT 297.640 180.000 305.080 180.320 ; 
                RECT 0.160 181.360 59.280 181.680 ; 
                RECT 63.720 181.360 76.960 181.680 ; 
                RECT 297.640 181.360 305.080 181.680 ; 
                RECT 0.160 182.720 59.280 183.040 ; 
                RECT 63.720 182.720 76.960 183.040 ; 
                RECT 297.640 182.720 305.080 183.040 ; 
                RECT 0.160 184.080 35.480 184.400 ; 
                RECT 44.000 184.080 76.960 184.400 ; 
                RECT 297.640 184.080 305.080 184.400 ; 
                RECT 0.160 185.440 34.120 185.760 ; 
                RECT 43.320 185.440 55.880 185.760 ; 
                RECT 63.720 185.440 76.960 185.760 ; 
                RECT 297.640 185.440 305.080 185.760 ; 
                RECT 0.160 186.800 55.880 187.120 ; 
                RECT 63.720 186.800 76.960 187.120 ; 
                RECT 297.640 186.800 305.080 187.120 ; 
                RECT 0.160 188.160 55.880 188.480 ; 
                RECT 58.280 188.160 76.960 188.480 ; 
                RECT 297.640 188.160 305.080 188.480 ; 
                RECT 0.160 189.520 55.880 189.840 ; 
                RECT 63.720 189.520 76.960 189.840 ; 
                RECT 297.640 189.520 305.080 189.840 ; 
                RECT 0.160 190.880 55.880 191.200 ; 
                RECT 63.720 190.880 76.960 191.200 ; 
                RECT 297.640 190.880 305.080 191.200 ; 
                RECT 0.160 192.240 55.880 192.560 ; 
                RECT 59.640 192.240 76.960 192.560 ; 
                RECT 297.640 192.240 305.080 192.560 ; 
                RECT 0.160 193.600 57.920 193.920 ; 
                RECT 63.720 193.600 76.960 193.920 ; 
                RECT 297.640 193.600 305.080 193.920 ; 
                RECT 0.160 194.960 58.600 195.280 ; 
                RECT 63.720 194.960 76.960 195.280 ; 
                RECT 297.640 194.960 305.080 195.280 ; 
                RECT 0.160 196.320 59.280 196.640 ; 
                RECT 63.720 196.320 76.960 196.640 ; 
                RECT 297.640 196.320 305.080 196.640 ; 
                RECT 0.160 197.680 76.960 198.000 ; 
                RECT 297.640 197.680 305.080 198.000 ; 
                RECT 0.160 199.040 59.280 199.360 ; 
                RECT 63.720 199.040 76.960 199.360 ; 
                RECT 297.640 199.040 305.080 199.360 ; 
                RECT 0.160 200.400 76.960 200.720 ; 
                RECT 297.640 200.400 305.080 200.720 ; 
                RECT 0.160 201.760 59.960 202.080 ; 
                RECT 63.720 201.760 76.960 202.080 ; 
                RECT 297.640 201.760 305.080 202.080 ; 
                RECT 0.160 203.120 60.640 203.440 ; 
                RECT 63.720 203.120 76.960 203.440 ; 
                RECT 297.640 203.120 305.080 203.440 ; 
                RECT 0.160 204.480 61.320 204.800 ; 
                RECT 63.720 204.480 76.960 204.800 ; 
                RECT 297.640 204.480 305.080 204.800 ; 
                RECT 0.160 205.840 61.320 206.160 ; 
                RECT 63.720 205.840 76.960 206.160 ; 
                RECT 297.640 205.840 305.080 206.160 ; 
                RECT 0.160 207.200 76.960 207.520 ; 
                RECT 297.640 207.200 305.080 207.520 ; 
                RECT 0.160 208.560 76.960 208.880 ; 
                RECT 297.640 208.560 305.080 208.880 ; 
                RECT 0.160 209.920 131.360 210.240 ; 
                RECT 297.640 209.920 305.080 210.240 ; 
                RECT 0.160 211.280 131.360 211.600 ; 
                RECT 297.640 211.280 305.080 211.600 ; 
                RECT 0.160 212.640 131.360 212.960 ; 
                RECT 297.640 212.640 305.080 212.960 ; 
                RECT 0.160 214.000 305.080 214.320 ; 
                RECT 0.160 215.360 305.080 215.680 ; 
                RECT 0.160 216.720 305.080 217.040 ; 
                RECT 0.160 218.080 305.080 218.400 ; 
                RECT 0.160 0.160 305.080 1.520 ; 
                RECT 0.160 222.800 305.080 224.160 ; 
                RECT 135.500 40.720 141.300 42.090 ; 
                RECT 287.400 40.720 293.200 42.090 ; 
                RECT 135.500 45.835 141.300 47.255 ; 
                RECT 287.400 45.835 293.200 47.255 ; 
                RECT 135.500 51.155 141.300 52.675 ; 
                RECT 287.400 51.155 293.200 52.675 ; 
                RECT 135.500 56.625 141.300 58.145 ; 
                RECT 287.400 56.625 293.200 58.145 ; 
                RECT 135.500 76.500 293.200 77.300 ; 
                RECT 135.500 84.400 293.200 85.200 ; 
                RECT 135.500 90.715 293.200 91.785 ; 
                RECT 135.500 79.510 293.200 80.310 ; 
                RECT 135.500 95.005 293.200 95.295 ; 
                RECT 135.500 132.560 293.200 133.910 ; 
                RECT 135.500 65.030 293.200 66.830 ; 
                RECT 135.500 117.310 293.200 118.280 ; 
                RECT 135.500 24.965 293.200 26.765 ; 
                RECT 84.090 144.355 86.010 209.135 ; 
                RECT 87.930 144.355 89.850 209.135 ; 
                RECT 107.035 144.355 108.955 209.135 ; 
                RECT 110.875 144.355 112.795 209.135 ; 
                RECT 114.715 144.355 116.635 209.135 ; 
                RECT 118.555 144.355 120.475 209.135 ; 
                RECT 122.395 144.355 124.315 209.135 ; 
                RECT 126.235 144.355 128.155 209.135 ; 
                RECT 96.135 65.060 98.055 91.860 ; 
                RECT 102.765 65.060 104.515 91.860 ; 
                RECT 110.960 65.060 112.880 91.860 ; 
                RECT 114.800 65.060 116.720 91.860 ; 
                RECT 100.415 119.500 102.335 137.720 ; 
                RECT 107.475 119.500 109.225 137.720 ; 
                RECT 114.580 119.500 116.500 137.720 ; 
                RECT 99.985 97.860 101.905 113.500 ; 
                RECT 107.045 97.860 108.795 113.500 ; 
                RECT 114.365 97.860 116.285 113.500 ; 
                RECT 114.600 55.480 116.520 59.060 ; 
                RECT 23.750 146.625 32.910 147.375 ; 
                RECT 23.750 151.250 32.910 153.000 ; 
                RECT 36.880 134.410 52.920 135.210 ; 
                RECT 20.080 135.070 34.920 136.760 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 144.280 5.560 ; 
                RECT 146.000 5.240 150.400 5.560 ; 
                RECT 152.120 5.240 156.520 5.560 ; 
                RECT 158.240 5.240 162.640 5.560 ; 
                RECT 164.360 5.240 168.760 5.560 ; 
                RECT 170.480 5.240 174.880 5.560 ; 
                RECT 176.600 5.240 181.000 5.560 ; 
                RECT 182.720 5.240 187.120 5.560 ; 
                RECT 188.840 5.240 193.240 5.560 ; 
                RECT 194.960 5.240 199.360 5.560 ; 
                RECT 201.080 5.240 205.480 5.560 ; 
                RECT 207.200 5.240 211.600 5.560 ; 
                RECT 213.320 5.240 217.720 5.560 ; 
                RECT 219.440 5.240 223.840 5.560 ; 
                RECT 225.560 5.240 229.960 5.560 ; 
                RECT 231.680 5.240 236.080 5.560 ; 
                RECT 237.800 5.240 242.200 5.560 ; 
                RECT 243.920 5.240 248.320 5.560 ; 
                RECT 250.040 5.240 254.440 5.560 ; 
                RECT 256.160 5.240 260.560 5.560 ; 
                RECT 262.280 5.240 266.680 5.560 ; 
                RECT 268.400 5.240 272.800 5.560 ; 
                RECT 274.520 5.240 278.920 5.560 ; 
                RECT 280.640 5.240 285.040 5.560 ; 
                RECT 286.080 5.240 302.360 5.560 ; 
                RECT 2.880 6.600 302.360 6.920 ; 
                RECT 2.880 7.960 302.360 8.280 ; 
                RECT 2.880 9.320 118.440 9.640 ; 
                RECT 139.880 9.320 302.360 9.640 ; 
                RECT 2.880 10.680 302.360 11.000 ; 
                RECT 2.880 12.040 302.360 12.360 ; 
                RECT 2.880 13.400 62.680 13.720 ; 
                RECT 119.480 13.400 302.360 13.720 ; 
                RECT 2.880 14.760 302.360 15.080 ; 
                RECT 2.880 16.120 302.360 16.440 ; 
                RECT 2.880 17.480 62.680 17.800 ; 
                RECT 118.800 17.480 302.360 17.800 ; 
                RECT 2.880 18.840 134.080 19.160 ; 
                RECT 294.920 18.840 302.360 19.160 ; 
                RECT 2.880 20.200 134.080 20.520 ; 
                RECT 294.920 20.200 302.360 20.520 ; 
                RECT 2.880 21.560 134.080 21.880 ; 
                RECT 294.920 21.560 302.360 21.880 ; 
                RECT 2.880 22.920 134.080 23.240 ; 
                RECT 294.920 22.920 302.360 23.240 ; 
                RECT 2.880 24.280 134.080 24.600 ; 
                RECT 294.920 24.280 302.360 24.600 ; 
                RECT 2.880 25.640 134.080 25.960 ; 
                RECT 294.920 25.640 302.360 25.960 ; 
                RECT 2.880 27.000 134.080 27.320 ; 
                RECT 294.920 27.000 302.360 27.320 ; 
                RECT 2.880 28.360 134.080 28.680 ; 
                RECT 294.920 28.360 302.360 28.680 ; 
                RECT 2.880 29.720 134.080 30.040 ; 
                RECT 294.920 29.720 302.360 30.040 ; 
                RECT 2.880 31.080 134.080 31.400 ; 
                RECT 294.920 31.080 302.360 31.400 ; 
                RECT 2.880 32.440 83.760 32.760 ; 
                RECT 97.720 32.440 134.080 32.760 ; 
                RECT 294.920 32.440 302.360 32.760 ; 
                RECT 2.880 33.800 82.400 34.120 ; 
                RECT 103.840 33.800 134.080 34.120 ; 
                RECT 294.920 33.800 302.360 34.120 ; 
                RECT 2.880 35.160 59.280 35.480 ; 
                RECT 118.800 35.160 134.080 35.480 ; 
                RECT 294.920 35.160 302.360 35.480 ; 
                RECT 2.880 36.520 59.960 36.840 ; 
                RECT 109.280 36.520 133.400 36.840 ; 
                RECT 294.920 36.520 302.360 36.840 ; 
                RECT 2.880 37.880 134.080 38.200 ; 
                RECT 294.920 37.880 302.360 38.200 ; 
                RECT 2.880 39.240 134.080 39.560 ; 
                RECT 294.920 39.240 302.360 39.560 ; 
                RECT 2.880 40.600 134.080 40.920 ; 
                RECT 294.920 40.600 302.360 40.920 ; 
                RECT 2.880 41.960 134.080 42.280 ; 
                RECT 294.920 41.960 302.360 42.280 ; 
                RECT 2.880 43.320 57.240 43.640 ; 
                RECT 68.480 43.320 134.080 43.640 ; 
                RECT 294.920 43.320 302.360 43.640 ; 
                RECT 2.880 44.680 58.600 45.000 ; 
                RECT 61.000 44.680 134.080 45.000 ; 
                RECT 294.920 44.680 302.360 45.000 ; 
                RECT 2.880 46.040 59.960 46.360 ; 
                RECT 64.400 46.040 72.200 46.360 ; 
                RECT 74.600 46.040 134.080 46.360 ; 
                RECT 294.920 46.040 302.360 46.360 ; 
                RECT 2.880 47.400 59.960 47.720 ; 
                RECT 63.720 47.400 134.080 47.720 ; 
                RECT 294.920 47.400 302.360 47.720 ; 
                RECT 2.880 48.760 66.760 49.080 ; 
                RECT 75.280 48.760 134.080 49.080 ; 
                RECT 294.920 48.760 302.360 49.080 ; 
                RECT 2.880 50.120 62.000 50.440 ; 
                RECT 68.480 50.120 134.080 50.440 ; 
                RECT 294.920 50.120 302.360 50.440 ; 
                RECT 2.880 51.480 59.280 51.800 ; 
                RECT 68.480 51.480 134.080 51.800 ; 
                RECT 294.920 51.480 302.360 51.800 ; 
                RECT 2.880 52.840 134.080 53.160 ; 
                RECT 294.920 52.840 302.360 53.160 ; 
                RECT 2.880 54.200 58.600 54.520 ; 
                RECT 68.480 54.200 134.080 54.520 ; 
                RECT 294.920 54.200 302.360 54.520 ; 
                RECT 2.880 55.560 66.760 55.880 ; 
                RECT 74.600 55.560 110.960 55.880 ; 
                RECT 117.440 55.560 134.080 55.880 ; 
                RECT 294.920 55.560 302.360 55.880 ; 
                RECT 2.880 56.920 65.400 57.240 ; 
                RECT 68.480 56.920 110.960 57.240 ; 
                RECT 294.920 56.920 302.360 57.240 ; 
                RECT 2.880 58.280 80.360 58.600 ; 
                RECT 107.920 58.280 110.960 58.600 ; 
                RECT 117.440 58.280 134.080 58.600 ; 
                RECT 294.920 58.280 302.360 58.600 ; 
                RECT 2.880 59.640 66.760 59.960 ; 
                RECT 74.600 59.640 134.080 59.960 ; 
                RECT 294.920 59.640 302.360 59.960 ; 
                RECT 2.880 61.000 63.360 61.320 ; 
                RECT 68.480 61.000 134.080 61.320 ; 
                RECT 294.920 61.000 302.360 61.320 ; 
                RECT 2.880 62.360 65.400 62.680 ; 
                RECT 68.480 62.360 134.080 62.680 ; 
                RECT 294.920 62.360 302.360 62.680 ; 
                RECT 2.880 63.720 134.080 64.040 ; 
                RECT 294.920 63.720 302.360 64.040 ; 
                RECT 2.880 65.080 57.240 65.400 ; 
                RECT 80.040 65.080 81.720 65.400 ; 
                RECT 87.520 65.080 92.600 65.400 ; 
                RECT 117.440 65.080 134.080 65.400 ; 
                RECT 294.920 65.080 302.360 65.400 ; 
                RECT 2.880 66.440 75.600 66.760 ; 
                RECT 81.400 66.440 83.080 66.760 ; 
                RECT 86.160 66.440 92.600 66.760 ; 
                RECT 126.280 66.440 134.080 66.760 ; 
                RECT 294.920 66.440 302.360 66.760 ; 
                RECT 2.880 67.800 65.400 68.120 ; 
                RECT 68.480 67.800 78.320 68.120 ; 
                RECT 82.080 67.800 92.600 68.120 ; 
                RECT 124.920 67.800 134.080 68.120 ; 
                RECT 294.920 67.800 302.360 68.120 ; 
                RECT 2.880 69.160 57.240 69.480 ; 
                RECT 71.200 69.160 92.600 69.480 ; 
                RECT 126.280 69.160 134.080 69.480 ; 
                RECT 294.920 69.160 302.360 69.480 ; 
                RECT 2.880 70.520 66.080 70.840 ; 
                RECT 74.600 70.520 92.600 70.840 ; 
                RECT 126.280 70.520 134.080 70.840 ; 
                RECT 294.920 70.520 302.360 70.840 ; 
                RECT 2.880 71.880 64.040 72.200 ; 
                RECT 75.280 71.880 92.600 72.200 ; 
                RECT 117.440 71.880 134.080 72.200 ; 
                RECT 294.920 71.880 302.360 72.200 ; 
                RECT 2.880 73.240 59.280 73.560 ; 
                RECT 65.760 73.240 92.600 73.560 ; 
                RECT 127.640 73.240 134.080 73.560 ; 
                RECT 294.920 73.240 302.360 73.560 ; 
                RECT 2.880 74.600 92.600 74.920 ; 
                RECT 117.440 74.600 134.080 74.920 ; 
                RECT 294.920 74.600 302.360 74.920 ; 
                RECT 2.880 75.960 58.600 76.280 ; 
                RECT 62.360 75.960 92.600 76.280 ; 
                RECT 129.000 75.960 134.080 76.280 ; 
                RECT 294.920 75.960 302.360 76.280 ; 
                RECT 2.880 77.320 58.600 77.640 ; 
                RECT 68.480 77.320 92.600 77.640 ; 
                RECT 129.000 77.320 134.080 77.640 ; 
                RECT 294.920 77.320 302.360 77.640 ; 
                RECT 2.880 78.680 62.680 79.000 ; 
                RECT 73.920 78.680 92.600 79.000 ; 
                RECT 131.720 78.680 134.080 79.000 ; 
                RECT 294.920 78.680 302.360 79.000 ; 
                RECT 2.880 80.040 65.400 80.360 ; 
                RECT 67.800 80.040 92.600 80.360 ; 
                RECT 130.360 80.040 134.080 80.360 ; 
                RECT 294.920 80.040 302.360 80.360 ; 
                RECT 2.880 81.400 66.760 81.720 ; 
                RECT 68.480 81.400 92.600 81.720 ; 
                RECT 131.720 81.400 134.080 81.720 ; 
                RECT 294.920 81.400 302.360 81.720 ; 
                RECT 2.880 82.760 92.600 83.080 ; 
                RECT 117.440 82.760 134.080 83.080 ; 
                RECT 294.920 82.760 302.360 83.080 ; 
                RECT 2.880 84.120 57.240 84.440 ; 
                RECT 74.600 84.120 92.600 84.440 ; 
                RECT 131.720 84.120 134.080 84.440 ; 
                RECT 294.920 84.120 302.360 84.440 ; 
                RECT 2.880 85.480 57.240 85.800 ; 
                RECT 68.480 85.480 72.880 85.800 ; 
                RECT 74.600 85.480 92.600 85.800 ; 
                RECT 294.920 85.480 302.360 85.800 ; 
                RECT 2.880 86.840 66.080 87.160 ; 
                RECT 68.480 86.840 92.600 87.160 ; 
                RECT 294.920 86.840 302.360 87.160 ; 
                RECT 2.880 88.200 92.600 88.520 ; 
                RECT 294.920 88.200 302.360 88.520 ; 
                RECT 2.880 89.560 92.600 89.880 ; 
                RECT 294.920 89.560 302.360 89.880 ; 
                RECT 2.880 90.920 53.840 91.240 ; 
                RECT 67.120 90.920 92.600 91.240 ; 
                RECT 294.920 90.920 302.360 91.240 ; 
                RECT 2.880 92.280 64.040 92.600 ; 
                RECT 71.200 92.280 134.080 92.600 ; 
                RECT 294.920 92.280 302.360 92.600 ; 
                RECT 2.880 93.640 134.080 93.960 ; 
                RECT 294.920 93.640 302.360 93.960 ; 
                RECT 2.880 95.000 134.080 95.320 ; 
                RECT 294.920 95.000 302.360 95.320 ; 
                RECT 2.880 96.360 62.680 96.680 ; 
                RECT 77.320 96.360 134.080 96.680 ; 
                RECT 294.920 96.360 302.360 96.680 ; 
                RECT 2.880 97.720 96.000 98.040 ; 
                RECT 116.760 97.720 134.080 98.040 ; 
                RECT 294.920 97.720 302.360 98.040 ; 
                RECT 2.880 99.080 96.000 99.400 ; 
                RECT 116.760 99.080 134.080 99.400 ; 
                RECT 294.920 99.080 302.360 99.400 ; 
                RECT 2.880 100.440 59.280 100.760 ; 
                RECT 62.360 100.440 96.000 100.760 ; 
                RECT 116.760 100.440 134.080 100.760 ; 
                RECT 294.920 100.440 302.360 100.760 ; 
                RECT 2.880 101.800 57.240 102.120 ; 
                RECT 61.000 101.800 96.000 102.120 ; 
                RECT 116.760 101.800 134.080 102.120 ; 
                RECT 294.920 101.800 302.360 102.120 ; 
                RECT 2.880 103.160 96.000 103.480 ; 
                RECT 116.760 103.160 134.080 103.480 ; 
                RECT 294.920 103.160 302.360 103.480 ; 
                RECT 2.880 104.520 72.880 104.840 ; 
                RECT 75.280 104.520 96.000 104.840 ; 
                RECT 116.760 104.520 134.080 104.840 ; 
                RECT 294.920 104.520 302.360 104.840 ; 
                RECT 2.880 105.880 96.000 106.200 ; 
                RECT 116.760 105.880 134.080 106.200 ; 
                RECT 294.920 105.880 302.360 106.200 ; 
                RECT 2.880 107.240 96.000 107.560 ; 
                RECT 116.760 107.240 134.080 107.560 ; 
                RECT 294.920 107.240 302.360 107.560 ; 
                RECT 2.880 108.600 96.000 108.920 ; 
                RECT 294.920 108.600 302.360 108.920 ; 
                RECT 2.880 109.960 59.280 110.280 ; 
                RECT 64.400 109.960 96.000 110.280 ; 
                RECT 116.760 109.960 131.360 110.280 ; 
                RECT 294.920 109.960 302.360 110.280 ; 
                RECT 2.880 111.320 96.000 111.640 ; 
                RECT 116.760 111.320 128.640 111.640 ; 
                RECT 294.920 111.320 302.360 111.640 ; 
                RECT 2.880 112.680 35.480 113.000 ; 
                RECT 54.200 112.680 65.400 113.000 ; 
                RECT 74.600 112.680 96.000 113.000 ; 
                RECT 116.760 112.680 125.920 113.000 ; 
                RECT 294.920 112.680 302.360 113.000 ; 
                RECT 2.880 114.040 35.480 114.360 ; 
                RECT 54.200 114.040 123.200 114.360 ; 
                RECT 294.920 114.040 302.360 114.360 ; 
                RECT 2.880 115.400 35.480 115.720 ; 
                RECT 54.200 115.400 62.000 115.720 ; 
                RECT 64.400 115.400 123.200 115.720 ; 
                RECT 294.920 115.400 302.360 115.720 ; 
                RECT 2.880 116.760 35.480 117.080 ; 
                RECT 54.200 116.760 58.600 117.080 ; 
                RECT 61.680 116.760 134.080 117.080 ; 
                RECT 294.920 116.760 302.360 117.080 ; 
                RECT 2.880 118.120 35.480 118.440 ; 
                RECT 54.200 118.120 134.080 118.440 ; 
                RECT 294.920 118.120 302.360 118.440 ; 
                RECT 2.880 119.480 35.480 119.800 ; 
                RECT 54.200 119.480 96.000 119.800 ; 
                RECT 117.440 119.480 134.080 119.800 ; 
                RECT 294.920 119.480 302.360 119.800 ; 
                RECT 2.880 120.840 35.480 121.160 ; 
                RECT 54.200 120.840 96.000 121.160 ; 
                RECT 117.440 120.840 134.080 121.160 ; 
                RECT 294.920 120.840 302.360 121.160 ; 
                RECT 2.880 122.200 35.480 122.520 ; 
                RECT 54.200 122.200 96.000 122.520 ; 
                RECT 117.440 122.200 134.080 122.520 ; 
                RECT 294.920 122.200 302.360 122.520 ; 
                RECT 2.880 123.560 35.480 123.880 ; 
                RECT 54.200 123.560 96.000 123.880 ; 
                RECT 117.440 123.560 124.560 123.880 ; 
                RECT 294.920 123.560 302.360 123.880 ; 
                RECT 2.880 124.920 35.480 125.240 ; 
                RECT 54.200 124.920 96.000 125.240 ; 
                RECT 117.440 124.920 124.560 125.240 ; 
                RECT 294.920 124.920 302.360 125.240 ; 
                RECT 2.880 126.280 35.480 126.600 ; 
                RECT 54.200 126.280 60.640 126.600 ; 
                RECT 64.400 126.280 96.000 126.600 ; 
                RECT 117.440 126.280 127.280 126.600 ; 
                RECT 294.920 126.280 302.360 126.600 ; 
                RECT 2.880 127.640 96.000 127.960 ; 
                RECT 117.440 127.640 130.000 127.960 ; 
                RECT 294.920 127.640 302.360 127.960 ; 
                RECT 2.880 129.000 96.000 129.320 ; 
                RECT 294.920 129.000 302.360 129.320 ; 
                RECT 2.880 130.360 96.000 130.680 ; 
                RECT 294.920 130.360 302.360 130.680 ; 
                RECT 2.880 131.720 19.160 132.040 ; 
                RECT 35.840 131.720 62.680 132.040 ; 
                RECT 68.480 131.720 96.000 132.040 ; 
                RECT 117.440 131.720 134.080 132.040 ; 
                RECT 294.920 131.720 302.360 132.040 ; 
                RECT 2.880 133.080 19.160 133.400 ; 
                RECT 35.840 133.080 41.600 133.400 ; 
                RECT 48.760 133.080 96.000 133.400 ; 
                RECT 117.440 133.080 134.080 133.400 ; 
                RECT 294.920 133.080 302.360 133.400 ; 
                RECT 2.880 134.440 19.160 134.760 ; 
                RECT 53.520 134.440 96.000 134.760 ; 
                RECT 117.440 134.440 134.080 134.760 ; 
                RECT 294.920 134.440 302.360 134.760 ; 
                RECT 2.880 135.800 19.160 136.120 ; 
                RECT 35.840 135.800 96.000 136.120 ; 
                RECT 294.920 135.800 302.360 136.120 ; 
                RECT 2.880 137.160 19.840 137.480 ; 
                RECT 48.760 137.160 57.240 137.480 ; 
                RECT 67.120 137.160 96.000 137.480 ; 
                RECT 117.440 137.160 134.080 137.480 ; 
                RECT 294.920 137.160 302.360 137.480 ; 
                RECT 2.880 138.520 41.600 138.840 ; 
                RECT 61.680 138.520 302.360 138.840 ; 
                RECT 2.880 139.880 30.040 140.200 ; 
                RECT 61.000 139.880 302.360 140.200 ; 
                RECT 2.880 141.240 131.360 141.560 ; 
                RECT 297.640 141.240 302.360 141.560 ; 
                RECT 2.880 142.600 131.360 142.920 ; 
                RECT 297.640 142.600 302.360 142.920 ; 
                RECT 2.880 143.960 25.280 144.280 ; 
                RECT 31.760 143.960 76.960 144.280 ; 
                RECT 297.640 143.960 302.360 144.280 ; 
                RECT 2.880 145.320 23.240 145.640 ; 
                RECT 44.000 145.320 76.960 145.640 ; 
                RECT 297.640 145.320 302.360 145.640 ; 
                RECT 2.880 146.680 23.240 147.000 ; 
                RECT 43.320 146.680 55.880 147.000 ; 
                RECT 63.720 146.680 76.960 147.000 ; 
                RECT 297.640 146.680 302.360 147.000 ; 
                RECT 2.880 148.040 36.840 148.360 ; 
                RECT 42.640 148.040 55.880 148.360 ; 
                RECT 63.720 148.040 76.960 148.360 ; 
                RECT 297.640 148.040 302.360 148.360 ; 
                RECT 2.880 149.400 23.240 149.720 ; 
                RECT 33.800 149.400 55.880 149.720 ; 
                RECT 63.720 149.400 76.960 149.720 ; 
                RECT 297.640 149.400 302.360 149.720 ; 
                RECT 2.880 150.760 23.240 151.080 ; 
                RECT 33.800 150.760 55.880 151.080 ; 
                RECT 63.720 150.760 76.960 151.080 ; 
                RECT 297.640 150.760 302.360 151.080 ; 
                RECT 2.880 152.120 23.240 152.440 ; 
                RECT 33.800 152.120 55.880 152.440 ; 
                RECT 60.320 152.120 76.960 152.440 ; 
                RECT 297.640 152.120 302.360 152.440 ; 
                RECT 2.880 153.480 76.960 153.800 ; 
                RECT 297.640 153.480 302.360 153.800 ; 
                RECT 2.880 154.840 55.880 155.160 ; 
                RECT 63.720 154.840 76.960 155.160 ; 
                RECT 297.640 154.840 302.360 155.160 ; 
                RECT 2.880 156.200 55.880 156.520 ; 
                RECT 63.720 156.200 76.960 156.520 ; 
                RECT 297.640 156.200 302.360 156.520 ; 
                RECT 2.880 157.560 16.440 157.880 ; 
                RECT 18.840 157.560 32.080 157.880 ; 
                RECT 34.480 157.560 61.320 157.880 ; 
                RECT 63.720 157.560 76.960 157.880 ; 
                RECT 297.640 157.560 302.360 157.880 ; 
                RECT 2.880 158.920 15.760 159.240 ; 
                RECT 18.840 158.920 55.880 159.240 ; 
                RECT 63.720 158.920 76.960 159.240 ; 
                RECT 297.640 158.920 302.360 159.240 ; 
                RECT 2.880 160.280 15.080 160.600 ; 
                RECT 18.840 160.280 55.880 160.600 ; 
                RECT 61.000 160.280 76.960 160.600 ; 
                RECT 297.640 160.280 302.360 160.600 ; 
                RECT 2.880 161.640 14.400 161.960 ; 
                RECT 18.840 161.640 57.920 161.960 ; 
                RECT 63.720 161.640 76.960 161.960 ; 
                RECT 297.640 161.640 302.360 161.960 ; 
                RECT 2.880 163.000 55.880 163.320 ; 
                RECT 57.600 163.000 76.960 163.320 ; 
                RECT 297.640 163.000 302.360 163.320 ; 
                RECT 2.880 164.360 13.720 164.680 ; 
                RECT 18.840 164.360 55.880 164.680 ; 
                RECT 61.680 164.360 76.960 164.680 ; 
                RECT 297.640 164.360 302.360 164.680 ; 
                RECT 2.880 165.720 55.880 166.040 ; 
                RECT 63.720 165.720 76.960 166.040 ; 
                RECT 297.640 165.720 302.360 166.040 ; 
                RECT 2.880 167.080 13.040 167.400 ; 
                RECT 18.840 167.080 32.080 167.400 ; 
                RECT 37.880 167.080 55.880 167.400 ; 
                RECT 63.720 167.080 76.960 167.400 ; 
                RECT 297.640 167.080 302.360 167.400 ; 
                RECT 2.880 168.440 12.360 168.760 ; 
                RECT 18.840 168.440 32.080 168.760 ; 
                RECT 36.520 168.440 55.880 168.760 ; 
                RECT 62.360 168.440 76.960 168.760 ; 
                RECT 297.640 168.440 302.360 168.760 ; 
                RECT 2.880 169.800 11.680 170.120 ; 
                RECT 18.840 169.800 32.080 170.120 ; 
                RECT 35.840 169.800 59.960 170.120 ; 
                RECT 63.720 169.800 76.960 170.120 ; 
                RECT 297.640 169.800 302.360 170.120 ; 
                RECT 2.880 171.160 55.880 171.480 ; 
                RECT 63.720 171.160 76.960 171.480 ; 
                RECT 297.640 171.160 302.360 171.480 ; 
                RECT 2.880 172.520 11.000 172.840 ; 
                RECT 18.840 172.520 32.080 172.840 ; 
                RECT 35.160 172.520 55.880 172.840 ; 
                RECT 63.040 172.520 76.960 172.840 ; 
                RECT 297.640 172.520 302.360 172.840 ; 
                RECT 2.880 173.880 10.320 174.200 ; 
                RECT 18.840 173.880 32.080 174.200 ; 
                RECT 34.480 173.880 55.880 174.200 ; 
                RECT 57.600 173.880 76.960 174.200 ; 
                RECT 297.640 173.880 302.360 174.200 ; 
                RECT 2.880 175.240 55.880 175.560 ; 
                RECT 63.720 175.240 76.960 175.560 ; 
                RECT 297.640 175.240 302.360 175.560 ; 
                RECT 2.880 176.600 76.960 176.920 ; 
                RECT 297.640 176.600 302.360 176.920 ; 
                RECT 2.880 177.960 57.920 178.280 ; 
                RECT 63.720 177.960 76.960 178.280 ; 
                RECT 297.640 177.960 302.360 178.280 ; 
                RECT 2.880 179.320 58.600 179.640 ; 
                RECT 63.720 179.320 76.960 179.640 ; 
                RECT 297.640 179.320 302.360 179.640 ; 
                RECT 2.880 180.680 59.280 181.000 ; 
                RECT 63.720 180.680 76.960 181.000 ; 
                RECT 297.640 180.680 302.360 181.000 ; 
                RECT 2.880 182.040 59.280 182.360 ; 
                RECT 63.720 182.040 76.960 182.360 ; 
                RECT 297.640 182.040 302.360 182.360 ; 
                RECT 2.880 183.400 76.960 183.720 ; 
                RECT 297.640 183.400 302.360 183.720 ; 
                RECT 2.880 184.760 34.800 185.080 ; 
                RECT 43.320 184.760 76.960 185.080 ; 
                RECT 297.640 184.760 302.360 185.080 ; 
                RECT 2.880 186.120 33.440 186.440 ; 
                RECT 42.640 186.120 55.880 186.440 ; 
                RECT 63.720 186.120 76.960 186.440 ; 
                RECT 297.640 186.120 302.360 186.440 ; 
                RECT 2.880 187.480 55.880 187.800 ; 
                RECT 63.720 187.480 76.960 187.800 ; 
                RECT 297.640 187.480 302.360 187.800 ; 
                RECT 2.880 188.840 55.880 189.160 ; 
                RECT 63.720 188.840 76.960 189.160 ; 
                RECT 297.640 188.840 302.360 189.160 ; 
                RECT 2.880 190.200 55.880 190.520 ; 
                RECT 63.720 190.200 76.960 190.520 ; 
                RECT 297.640 190.200 302.360 190.520 ; 
                RECT 2.880 191.560 55.880 191.880 ; 
                RECT 59.640 191.560 76.960 191.880 ; 
                RECT 297.640 191.560 302.360 191.880 ; 
                RECT 2.880 192.920 76.960 193.240 ; 
                RECT 297.640 192.920 302.360 193.240 ; 
                RECT 2.880 194.280 57.920 194.600 ; 
                RECT 63.720 194.280 76.960 194.600 ; 
                RECT 297.640 194.280 302.360 194.600 ; 
                RECT 2.880 195.640 58.600 195.960 ; 
                RECT 63.720 195.640 76.960 195.960 ; 
                RECT 297.640 195.640 302.360 195.960 ; 
                RECT 2.880 197.000 59.280 197.320 ; 
                RECT 63.720 197.000 76.960 197.320 ; 
                RECT 297.640 197.000 302.360 197.320 ; 
                RECT 2.880 198.360 59.280 198.680 ; 
                RECT 63.720 198.360 76.960 198.680 ; 
                RECT 297.640 198.360 302.360 198.680 ; 
                RECT 2.880 199.720 76.960 200.040 ; 
                RECT 297.640 199.720 302.360 200.040 ; 
                RECT 2.880 201.080 59.960 201.400 ; 
                RECT 63.720 201.080 76.960 201.400 ; 
                RECT 297.640 201.080 302.360 201.400 ; 
                RECT 2.880 202.440 76.960 202.760 ; 
                RECT 297.640 202.440 302.360 202.760 ; 
                RECT 2.880 203.800 60.640 204.120 ; 
                RECT 63.720 203.800 76.960 204.120 ; 
                RECT 297.640 203.800 302.360 204.120 ; 
                RECT 2.880 205.160 61.320 205.480 ; 
                RECT 63.720 205.160 76.960 205.480 ; 
                RECT 297.640 205.160 302.360 205.480 ; 
                RECT 2.880 206.520 61.320 206.840 ; 
                RECT 63.720 206.520 76.960 206.840 ; 
                RECT 297.640 206.520 302.360 206.840 ; 
                RECT 2.880 207.880 76.960 208.200 ; 
                RECT 297.640 207.880 302.360 208.200 ; 
                RECT 2.880 209.240 76.960 209.560 ; 
                RECT 297.640 209.240 302.360 209.560 ; 
                RECT 2.880 210.600 131.360 210.920 ; 
                RECT 297.640 210.600 302.360 210.920 ; 
                RECT 2.880 211.960 131.360 212.280 ; 
                RECT 297.640 211.960 302.360 212.280 ; 
                RECT 2.880 213.320 302.360 213.640 ; 
                RECT 2.880 214.680 302.360 215.000 ; 
                RECT 2.880 216.040 302.360 216.360 ; 
                RECT 2.880 217.400 302.360 217.720 ; 
                RECT 2.880 218.760 302.360 219.080 ; 
                RECT 2.880 2.880 302.360 4.240 ; 
                RECT 2.880 220.080 302.360 221.440 ; 
                RECT 135.500 38.075 141.300 39.195 ; 
                RECT 287.400 38.075 293.200 39.195 ; 
                RECT 135.500 43.875 141.300 44.525 ; 
                RECT 287.400 43.875 293.200 44.525 ; 
                RECT 135.500 49.085 141.300 49.775 ; 
                RECT 287.400 49.085 293.200 49.775 ; 
                RECT 135.500 54.555 141.300 55.245 ; 
                RECT 287.400 54.555 293.200 55.245 ; 
                RECT 135.500 121.790 293.200 122.160 ; 
                RECT 135.500 107.565 293.200 107.855 ; 
                RECT 135.500 88.845 293.200 89.915 ; 
                RECT 135.500 77.820 293.200 78.620 ; 
                RECT 135.500 80.830 293.200 81.630 ; 
                RECT 135.500 82.510 293.200 83.310 ; 
                RECT 135.500 85.720 293.200 86.520 ; 
                RECT 135.500 68.770 293.200 70.570 ; 
                RECT 135.500 28.705 293.200 30.505 ; 
                RECT 77.710 144.355 79.630 209.135 ; 
                RECT 95.880 144.355 97.800 209.135 ; 
                RECT 99.720 144.355 101.640 209.135 ; 
                RECT 93.510 65.060 94.400 91.860 ; 
                RECT 100.270 65.060 101.160 91.860 ; 
                RECT 107.030 65.060 108.780 91.860 ; 
                RECT 97.035 119.500 98.145 137.720 ; 
                RECT 104.980 119.500 105.870 137.720 ; 
                RECT 111.415 119.500 112.525 137.720 ; 
                RECT 96.605 97.860 97.715 113.500 ; 
                RECT 104.550 97.860 105.440 113.500 ; 
                RECT 110.985 97.860 112.095 113.500 ; 
                RECT 111.435 55.480 112.545 59.060 ; 
                RECT 23.750 145.420 32.910 145.790 ; 
                RECT 23.750 148.755 32.910 149.645 ; 
                RECT 20.080 131.580 34.920 132.250 ; 
                RECT 20.080 132.930 34.920 133.940 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 305.240 224.320 ; 
        LAYER met2 ;
            RECT 0.000 0.000 305.240 224.320 ; 
    END 
END sram22_128x24m4w8 
END LIBRARY 

