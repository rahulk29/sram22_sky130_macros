VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_128x40m4w20
    CLASS BLOCK  ;
    FOREIGN sram22_128x40m4w20   ;
    SIZE 484.760 BY 224.320 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 227.550 0.000 227.690 0.140 ;
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 233.650 0.000 233.790 0.140 ;
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 239.750 0.000 239.890 0.140 ;
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 245.850 0.000 245.990 0.140 ;
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 251.950 0.000 252.090 0.140 ;
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 258.050 0.000 258.190 0.140 ;
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 264.150 0.000 264.290 0.140 ;
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 270.250 0.000 270.390 0.140 ;
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 276.350 0.000 276.490 0.140 ;
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 282.450 0.000 282.590 0.140 ;
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 288.550 0.000 288.690 0.140 ;
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 294.650 0.000 294.790 0.140 ;
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 300.750 0.000 300.890 0.140 ;
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 306.850 0.000 306.990 0.140 ;
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 312.950 0.000 313.090 0.140 ;
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 319.050 0.000 319.190 0.140 ;
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 325.150 0.000 325.290 0.140 ;
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 331.250 0.000 331.390 0.140 ;
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 337.350 0.000 337.490 0.140 ;
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 343.450 0.000 343.590 0.140 ;
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 349.550 0.000 349.690 0.140 ;
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 355.650 0.000 355.790 0.140 ;
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 361.750 0.000 361.890 0.140 ;
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 367.850 0.000 367.990 0.140 ;
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 373.950 0.000 374.090 0.140 ;
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 380.050 0.000 380.190 0.140 ;
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 386.150 0.000 386.290 0.140 ;
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 392.250 0.000 392.390 0.140 ;
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 398.350 0.000 398.490 0.140 ;
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 404.450 0.000 404.590 0.140 ;
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 410.550 0.000 410.690 0.140 ;
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 416.650 0.000 416.790 0.140 ;
        END 
    END dout[31] 
    PIN dout[32] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 422.750 0.000 422.890 0.140 ;
        END 
    END dout[32] 
    PIN dout[33] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 428.850 0.000 428.990 0.140 ;
        END 
    END dout[33] 
    PIN dout[34] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 434.950 0.000 435.090 0.140 ;
        END 
    END dout[34] 
    PIN dout[35] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 441.050 0.000 441.190 0.140 ;
        END 
    END dout[35] 
    PIN dout[36] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 447.150 0.000 447.290 0.140 ;
        END 
    END dout[36] 
    PIN dout[37] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 453.250 0.000 453.390 0.140 ;
        END 
    END dout[37] 
    PIN dout[38] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 459.350 0.000 459.490 0.140 ;
        END 
    END dout[38] 
    PIN dout[39] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.497800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 465.450 0.000 465.590 0.140 ;
        END 
    END dout[39] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 227.130 0.000 227.270 0.140 ;
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 233.230 0.000 233.370 0.140 ;
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 239.330 0.000 239.470 0.140 ;
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 245.430 0.000 245.570 0.140 ;
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 251.530 0.000 251.670 0.140 ;
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 257.630 0.000 257.770 0.140 ;
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 263.730 0.000 263.870 0.140 ;
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 269.830 0.000 269.970 0.140 ;
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 275.930 0.000 276.070 0.140 ;
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 282.030 0.000 282.170 0.140 ;
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 288.130 0.000 288.270 0.140 ;
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 294.230 0.000 294.370 0.140 ;
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 300.330 0.000 300.470 0.140 ;
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 306.430 0.000 306.570 0.140 ;
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 312.530 0.000 312.670 0.140 ;
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 318.630 0.000 318.770 0.140 ;
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 324.730 0.000 324.870 0.140 ;
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.830 0.000 330.970 0.140 ;
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.930 0.000 337.070 0.140 ;
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 343.030 0.000 343.170 0.140 ;
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 349.130 0.000 349.270 0.140 ;
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 355.230 0.000 355.370 0.140 ;
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 361.330 0.000 361.470 0.140 ;
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 367.430 0.000 367.570 0.140 ;
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 373.530 0.000 373.670 0.140 ;
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 379.630 0.000 379.770 0.140 ;
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 385.730 0.000 385.870 0.140 ;
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 391.830 0.000 391.970 0.140 ;
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 397.930 0.000 398.070 0.140 ;
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 404.030 0.000 404.170 0.140 ;
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 410.130 0.000 410.270 0.140 ;
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 416.230 0.000 416.370 0.140 ;
        END 
    END din[31] 
    PIN din[32] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 422.330 0.000 422.470 0.140 ;
        END 
    END din[32] 
    PIN din[33] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 428.430 0.000 428.570 0.140 ;
        END 
    END din[33] 
    PIN din[34] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 434.530 0.000 434.670 0.140 ;
        END 
    END din[34] 
    PIN din[35] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 440.630 0.000 440.770 0.140 ;
        END 
    END din[35] 
    PIN din[36] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 446.730 0.000 446.870 0.140 ;
        END 
    END din[36] 
    PIN din[37] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 452.830 0.000 452.970 0.140 ;
        END 
    END din[37] 
    PIN din[38] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 458.930 0.000 459.070 0.140 ;
        END 
    END din[38] 
    PIN din[39] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.939600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.219400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 465.030 0.000 465.170 0.140 ;
        END 
    END din[39] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.750000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 226.780 0.000 226.920 0.140 ;
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.750000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 348.780 0.000 348.920 0.140 ;
        END 
    END wmask[1] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 185.440 0.000 185.760 0.320 ;
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 179.320 0.000 179.640 0.320 ;
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 173.200 0.000 173.520 0.320 ;
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 167.080 0.000 167.400 0.320 ;
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 160.960 0.000 161.280 0.320 ;
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 154.840 0.000 155.160 0.320 ;
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 148.720 0.000 149.040 0.320 ;
        END 
    END addr[6] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 197.680 0.000 198.000 0.320 ;
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 191.560 0.000 191.880 0.320 ;
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 25.947000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 200.400 0.000 200.720 0.320 ;
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 29.853000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 201.080 0.000 201.400 0.320 ;
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 226.560 6.240 ;
                RECT 228.280 5.920 232.680 6.240 ;
                RECT 234.400 5.920 238.800 6.240 ;
                RECT 240.520 5.920 244.920 6.240 ;
                RECT 246.640 5.920 251.040 6.240 ;
                RECT 252.760 5.920 257.160 6.240 ;
                RECT 258.880 5.920 263.280 6.240 ;
                RECT 265.000 5.920 269.400 6.240 ;
                RECT 271.120 5.920 275.520 6.240 ;
                RECT 277.240 5.920 281.640 6.240 ;
                RECT 283.360 5.920 287.760 6.240 ;
                RECT 289.480 5.920 293.880 6.240 ;
                RECT 295.600 5.920 300.000 6.240 ;
                RECT 301.720 5.920 306.120 6.240 ;
                RECT 307.840 5.920 312.240 6.240 ;
                RECT 313.960 5.920 318.360 6.240 ;
                RECT 320.080 5.920 324.480 6.240 ;
                RECT 326.200 5.920 330.600 6.240 ;
                RECT 332.320 5.920 336.720 6.240 ;
                RECT 338.440 5.920 342.840 6.240 ;
                RECT 344.560 5.920 348.960 6.240 ;
                RECT 350.680 5.920 355.080 6.240 ;
                RECT 356.800 5.920 361.200 6.240 ;
                RECT 362.920 5.920 367.320 6.240 ;
                RECT 368.360 5.920 373.440 6.240 ;
                RECT 374.480 5.920 379.560 6.240 ;
                RECT 380.600 5.920 385.680 6.240 ;
                RECT 386.720 5.920 391.800 6.240 ;
                RECT 392.840 5.920 397.920 6.240 ;
                RECT 398.960 5.920 404.040 6.240 ;
                RECT 405.080 5.920 410.160 6.240 ;
                RECT 411.200 5.920 416.280 6.240 ;
                RECT 417.320 5.920 421.720 6.240 ;
                RECT 423.440 5.920 427.840 6.240 ;
                RECT 429.560 5.920 433.960 6.240 ;
                RECT 435.680 5.920 440.080 6.240 ;
                RECT 441.800 5.920 446.200 6.240 ;
                RECT 447.920 5.920 452.320 6.240 ;
                RECT 454.040 5.920 458.440 6.240 ;
                RECT 460.160 5.920 464.560 6.240 ;
                RECT 466.280 5.920 484.600 6.240 ;
                RECT 0.160 7.280 484.600 7.600 ;
                RECT 0.160 8.640 484.600 8.960 ;
                RECT 0.160 10.000 200.040 10.320 ;
                RECT 222.840 10.000 484.600 10.320 ;
                RECT 0.160 11.360 484.600 11.680 ;
                RECT 0.160 12.720 484.600 13.040 ;
                RECT 0.160 14.080 144.960 14.400 ;
                RECT 201.760 14.080 484.600 14.400 ;
                RECT 0.160 15.440 484.600 15.760 ;
                RECT 0.160 16.800 484.600 17.120 ;
                RECT 0.160 18.160 144.960 18.480 ;
                RECT 201.080 18.160 216.360 18.480 ;
                RECT 474.440 18.160 484.600 18.480 ;
                RECT 0.160 19.520 216.360 19.840 ;
                RECT 474.440 19.520 484.600 19.840 ;
                RECT 0.160 20.880 216.360 21.200 ;
                RECT 474.440 20.880 484.600 21.200 ;
                RECT 0.160 22.240 216.360 22.560 ;
                RECT 474.440 22.240 484.600 22.560 ;
                RECT 0.160 23.600 216.360 23.920 ;
                RECT 474.440 23.600 484.600 23.920 ;
                RECT 0.160 24.960 216.360 25.280 ;
                RECT 474.440 24.960 484.600 25.280 ;
                RECT 0.160 26.320 216.360 26.640 ;
                RECT 474.440 26.320 484.600 26.640 ;
                RECT 0.160 27.680 216.360 28.000 ;
                RECT 474.440 27.680 484.600 28.000 ;
                RECT 0.160 29.040 216.360 29.360 ;
                RECT 474.440 29.040 484.600 29.360 ;
                RECT 0.160 30.400 216.360 30.720 ;
                RECT 474.440 30.400 484.600 30.720 ;
                RECT 0.160 31.760 216.360 32.080 ;
                RECT 474.440 31.760 484.600 32.080 ;
                RECT 0.160 33.120 158.560 33.440 ;
                RECT 178.640 33.120 216.360 33.440 ;
                RECT 474.440 33.120 484.600 33.440 ;
                RECT 0.160 34.480 157.200 34.800 ;
                RECT 184.760 34.480 216.360 34.800 ;
                RECT 474.440 34.480 484.600 34.800 ;
                RECT 0.160 35.840 137.480 36.160 ;
                RECT 201.760 35.840 215.680 36.160 ;
                RECT 474.440 35.840 484.600 36.160 ;
                RECT 0.160 37.200 136.800 37.520 ;
                RECT 197.680 37.200 216.360 37.520 ;
                RECT 474.440 37.200 484.600 37.520 ;
                RECT 0.160 38.560 216.360 38.880 ;
                RECT 474.440 38.560 484.600 38.880 ;
                RECT 0.160 39.920 216.360 40.240 ;
                RECT 474.440 39.920 484.600 40.240 ;
                RECT 0.160 41.280 216.360 41.600 ;
                RECT 474.440 41.280 484.600 41.600 ;
                RECT 0.160 42.640 216.360 42.960 ;
                RECT 474.440 42.640 484.600 42.960 ;
                RECT 0.160 44.000 132.720 44.320 ;
                RECT 143.960 44.000 216.360 44.320 ;
                RECT 474.440 44.000 484.600 44.320 ;
                RECT 0.160 45.360 134.080 45.680 ;
                RECT 139.880 45.360 147.680 45.680 ;
                RECT 150.080 45.360 216.360 45.680 ;
                RECT 474.440 45.360 484.600 45.680 ;
                RECT 0.160 46.720 135.440 47.040 ;
                RECT 139.200 46.720 216.360 47.040 ;
                RECT 474.440 46.720 484.600 47.040 ;
                RECT 0.160 48.080 216.360 48.400 ;
                RECT 474.440 48.080 484.600 48.400 ;
                RECT 0.160 49.440 142.240 49.760 ;
                RECT 150.760 49.440 216.360 49.760 ;
                RECT 474.440 49.440 484.600 49.760 ;
                RECT 0.160 50.800 134.760 51.120 ;
                RECT 143.960 50.800 216.360 51.120 ;
                RECT 474.440 50.800 484.600 51.120 ;
                RECT 0.160 52.160 138.160 52.480 ;
                RECT 143.280 52.160 216.360 52.480 ;
                RECT 474.440 52.160 484.600 52.480 ;
                RECT 0.160 53.520 193.920 53.840 ;
                RECT 199.720 53.520 216.360 53.840 ;
                RECT 474.440 53.520 484.600 53.840 ;
                RECT 0.160 54.880 134.080 55.200 ;
                RECT 143.960 54.880 193.920 55.200 ;
                RECT 474.440 54.880 484.600 55.200 ;
                RECT 0.160 56.240 140.880 56.560 ;
                RECT 149.400 56.240 193.920 56.560 ;
                RECT 199.720 56.240 216.360 56.560 ;
                RECT 474.440 56.240 484.600 56.560 ;
                RECT 0.160 57.600 216.360 57.920 ;
                RECT 474.440 57.600 484.600 57.920 ;
                RECT 0.160 58.960 142.240 59.280 ;
                RECT 148.040 58.960 216.360 59.280 ;
                RECT 474.440 58.960 484.600 59.280 ;
                RECT 0.160 60.320 144.960 60.640 ;
                RECT 150.080 60.320 216.360 60.640 ;
                RECT 474.440 60.320 484.600 60.640 ;
                RECT 0.160 61.680 138.840 62.000 ;
                RECT 143.960 61.680 216.360 62.000 ;
                RECT 474.440 61.680 484.600 62.000 ;
                RECT 0.160 63.040 157.200 63.360 ;
                RECT 163.000 63.040 168.080 63.360 ;
                RECT 198.360 63.040 216.360 63.360 ;
                RECT 474.440 63.040 484.600 63.360 ;
                RECT 0.160 64.400 132.040 64.720 ;
                RECT 155.520 64.400 158.560 64.720 ;
                RECT 161.640 64.400 168.080 64.720 ;
                RECT 208.560 64.400 216.360 64.720 ;
                RECT 474.440 64.400 484.600 64.720 ;
                RECT 0.160 65.760 142.240 66.080 ;
                RECT 150.080 65.760 168.080 66.080 ;
                RECT 208.560 65.760 216.360 66.080 ;
                RECT 474.440 65.760 484.600 66.080 ;
                RECT 0.160 67.120 140.880 67.440 ;
                RECT 143.960 67.120 150.400 67.440 ;
                RECT 157.560 67.120 168.080 67.440 ;
                RECT 207.200 67.120 216.360 67.440 ;
                RECT 474.440 67.120 484.600 67.440 ;
                RECT 0.160 68.480 132.720 68.800 ;
                RECT 146.680 68.480 168.080 68.800 ;
                RECT 208.560 68.480 216.360 68.800 ;
                RECT 474.440 68.480 484.600 68.800 ;
                RECT 0.160 69.840 141.560 70.160 ;
                RECT 150.080 69.840 168.080 70.160 ;
                RECT 211.280 69.840 216.360 70.160 ;
                RECT 474.440 69.840 484.600 70.160 ;
                RECT 0.160 71.200 139.520 71.520 ;
                RECT 143.280 71.200 168.080 71.520 ;
                RECT 198.360 71.200 216.360 71.520 ;
                RECT 474.440 71.200 484.600 71.520 ;
                RECT 0.160 72.560 134.760 72.880 ;
                RECT 139.200 72.560 142.240 72.880 ;
                RECT 150.760 72.560 168.080 72.880 ;
                RECT 211.280 72.560 216.360 72.880 ;
                RECT 474.440 72.560 484.600 72.880 ;
                RECT 0.160 73.920 137.480 74.240 ;
                RECT 141.240 73.920 168.080 74.240 ;
                RECT 209.920 73.920 216.360 74.240 ;
                RECT 474.440 73.920 484.600 74.240 ;
                RECT 0.160 75.280 134.080 75.600 ;
                RECT 137.840 75.280 168.080 75.600 ;
                RECT 211.280 75.280 216.360 75.600 ;
                RECT 474.440 75.280 484.600 75.600 ;
                RECT 0.160 76.640 138.160 76.960 ;
                RECT 143.960 76.640 168.080 76.960 ;
                RECT 214.000 76.640 216.360 76.960 ;
                RECT 474.440 76.640 484.600 76.960 ;
                RECT 0.160 78.000 134.080 78.320 ;
                RECT 149.400 78.000 168.080 78.320 ;
                RECT 214.000 78.000 216.360 78.320 ;
                RECT 474.440 78.000 484.600 78.320 ;
                RECT 0.160 79.360 168.080 79.680 ;
                RECT 212.640 79.360 216.360 79.680 ;
                RECT 474.440 79.360 484.600 79.680 ;
                RECT 0.160 80.720 140.880 81.040 ;
                RECT 143.280 80.720 168.080 81.040 ;
                RECT 198.360 80.720 216.360 81.040 ;
                RECT 474.440 80.720 484.600 81.040 ;
                RECT 0.160 82.080 142.240 82.400 ;
                RECT 143.960 82.080 168.080 82.400 ;
                RECT 214.000 82.080 216.360 82.400 ;
                RECT 474.440 82.080 484.600 82.400 ;
                RECT 0.160 83.440 132.720 83.760 ;
                RECT 143.280 83.440 168.080 83.760 ;
                RECT 474.440 83.440 484.600 83.760 ;
                RECT 0.160 84.800 138.160 85.120 ;
                RECT 150.080 84.800 168.080 85.120 ;
                RECT 474.440 84.800 484.600 85.120 ;
                RECT 0.160 86.160 132.720 86.480 ;
                RECT 143.960 86.160 168.080 86.480 ;
                RECT 474.440 86.160 484.600 86.480 ;
                RECT 0.160 87.520 141.560 87.840 ;
                RECT 143.960 87.520 168.080 87.840 ;
                RECT 474.440 87.520 484.600 87.840 ;
                RECT 0.160 88.880 168.080 89.200 ;
                RECT 198.360 88.880 216.360 89.200 ;
                RECT 474.440 88.880 484.600 89.200 ;
                RECT 0.160 90.240 216.360 90.560 ;
                RECT 474.440 90.240 484.600 90.560 ;
                RECT 0.160 91.600 129.320 91.920 ;
                RECT 146.680 91.600 216.360 91.920 ;
                RECT 474.440 91.600 484.600 91.920 ;
                RECT 0.160 92.960 216.360 93.280 ;
                RECT 474.440 92.960 484.600 93.280 ;
                RECT 0.160 94.320 216.360 94.640 ;
                RECT 474.440 94.320 484.600 94.640 ;
                RECT 0.160 95.680 138.160 96.000 ;
                RECT 150.080 95.680 156.520 96.000 ;
                RECT 172.520 95.680 175.560 96.000 ;
                RECT 198.360 95.680 216.360 96.000 ;
                RECT 474.440 95.680 484.600 96.000 ;
                RECT 0.160 97.040 144.960 97.360 ;
                RECT 152.120 97.040 175.560 97.360 ;
                RECT 198.360 97.040 216.360 97.360 ;
                RECT 474.440 97.040 484.600 97.360 ;
                RECT 0.160 98.400 175.560 98.720 ;
                RECT 198.360 98.400 216.360 98.720 ;
                RECT 474.440 98.400 484.600 98.720 ;
                RECT 0.160 99.760 175.560 100.080 ;
                RECT 198.360 99.760 216.360 100.080 ;
                RECT 474.440 99.760 484.600 100.080 ;
                RECT 0.160 101.120 132.040 101.440 ;
                RECT 137.840 101.120 175.560 101.440 ;
                RECT 198.360 101.120 216.360 101.440 ;
                RECT 474.440 101.120 484.600 101.440 ;
                RECT 0.160 102.480 110.960 102.800 ;
                RECT 129.680 102.480 175.560 102.800 ;
                RECT 198.360 102.480 216.360 102.800 ;
                RECT 474.440 102.480 484.600 102.800 ;
                RECT 0.160 103.840 110.960 104.160 ;
                RECT 129.680 103.840 175.560 104.160 ;
                RECT 198.360 103.840 216.360 104.160 ;
                RECT 474.440 103.840 484.600 104.160 ;
                RECT 0.160 105.200 110.960 105.520 ;
                RECT 129.680 105.200 147.680 105.520 ;
                RECT 150.760 105.200 175.560 105.520 ;
                RECT 198.360 105.200 216.360 105.520 ;
                RECT 474.440 105.200 484.600 105.520 ;
                RECT 0.160 106.560 110.960 106.880 ;
                RECT 129.680 106.560 175.560 106.880 ;
                RECT 198.360 106.560 216.360 106.880 ;
                RECT 474.440 106.560 484.600 106.880 ;
                RECT 0.160 107.920 110.960 108.240 ;
                RECT 129.680 107.920 175.560 108.240 ;
                RECT 198.360 107.920 216.360 108.240 ;
                RECT 474.440 107.920 484.600 108.240 ;
                RECT 0.160 109.280 110.960 109.600 ;
                RECT 129.680 109.280 175.560 109.600 ;
                RECT 474.440 109.280 484.600 109.600 ;
                RECT 0.160 110.640 110.960 110.960 ;
                RECT 129.680 110.640 134.760 110.960 ;
                RECT 139.880 110.640 175.560 110.960 ;
                RECT 198.360 110.640 213.640 110.960 ;
                RECT 474.440 110.640 484.600 110.960 ;
                RECT 0.160 112.000 110.960 112.320 ;
                RECT 130.360 112.000 175.560 112.320 ;
                RECT 198.360 112.000 210.920 112.320 ;
                RECT 474.440 112.000 484.600 112.320 ;
                RECT 0.160 113.360 110.960 113.680 ;
                RECT 129.680 113.360 140.880 113.680 ;
                RECT 149.400 113.360 175.560 113.680 ;
                RECT 198.360 113.360 208.200 113.680 ;
                RECT 474.440 113.360 484.600 113.680 ;
                RECT 0.160 114.720 110.960 115.040 ;
                RECT 129.680 114.720 205.480 115.040 ;
                RECT 474.440 114.720 484.600 115.040 ;
                RECT 0.160 116.080 110.960 116.400 ;
                RECT 129.680 116.080 137.480 116.400 ;
                RECT 139.880 116.080 216.360 116.400 ;
                RECT 474.440 116.080 484.600 116.400 ;
                RECT 0.160 117.440 110.960 117.760 ;
                RECT 129.680 117.440 134.080 117.760 ;
                RECT 137.160 117.440 216.360 117.760 ;
                RECT 474.440 117.440 484.600 117.760 ;
                RECT 0.160 118.800 110.960 119.120 ;
                RECT 129.680 118.800 216.360 119.120 ;
                RECT 474.440 118.800 484.600 119.120 ;
                RECT 0.160 120.160 110.960 120.480 ;
                RECT 129.680 120.160 174.200 120.480 ;
                RECT 198.360 120.160 216.360 120.480 ;
                RECT 474.440 120.160 484.600 120.480 ;
                RECT 0.160 121.520 110.960 121.840 ;
                RECT 129.680 121.520 174.200 121.840 ;
                RECT 198.360 121.520 216.360 121.840 ;
                RECT 474.440 121.520 484.600 121.840 ;
                RECT 0.160 122.880 110.960 123.200 ;
                RECT 129.680 122.880 174.200 123.200 ;
                RECT 198.360 122.880 216.360 123.200 ;
                RECT 474.440 122.880 484.600 123.200 ;
                RECT 0.160 124.240 110.960 124.560 ;
                RECT 129.680 124.240 174.200 124.560 ;
                RECT 198.360 124.240 206.840 124.560 ;
                RECT 474.440 124.240 484.600 124.560 ;
                RECT 0.160 125.600 110.960 125.920 ;
                RECT 129.680 125.600 174.200 125.920 ;
                RECT 198.360 125.600 209.560 125.920 ;
                RECT 474.440 125.600 484.600 125.920 ;
                RECT 0.160 126.960 110.960 127.280 ;
                RECT 129.680 126.960 136.120 127.280 ;
                RECT 139.880 126.960 174.200 127.280 ;
                RECT 198.360 126.960 212.280 127.280 ;
                RECT 474.440 126.960 484.600 127.280 ;
                RECT 0.160 128.320 174.200 128.640 ;
                RECT 198.360 128.320 215.000 128.640 ;
                RECT 474.440 128.320 484.600 128.640 ;
                RECT 0.160 129.680 174.200 130.000 ;
                RECT 474.440 129.680 484.600 130.000 ;
                RECT 0.160 131.040 94.640 131.360 ;
                RECT 111.320 131.040 138.160 131.360 ;
                RECT 143.960 131.040 174.200 131.360 ;
                RECT 198.360 131.040 216.360 131.360 ;
                RECT 474.440 131.040 484.600 131.360 ;
                RECT 0.160 132.400 94.640 132.720 ;
                RECT 111.320 132.400 117.080 132.720 ;
                RECT 124.240 132.400 174.200 132.720 ;
                RECT 198.360 132.400 216.360 132.720 ;
                RECT 474.440 132.400 484.600 132.720 ;
                RECT 0.160 133.760 94.640 134.080 ;
                RECT 129.000 133.760 174.200 134.080 ;
                RECT 198.360 133.760 216.360 134.080 ;
                RECT 474.440 133.760 484.600 134.080 ;
                RECT 0.160 135.120 94.640 135.440 ;
                RECT 129.000 135.120 174.200 135.440 ;
                RECT 474.440 135.120 484.600 135.440 ;
                RECT 0.160 136.480 94.640 136.800 ;
                RECT 111.320 136.480 117.080 136.800 ;
                RECT 124.240 136.480 132.720 136.800 ;
                RECT 142.600 136.480 174.200 136.800 ;
                RECT 474.440 136.480 484.600 136.800 ;
                RECT 0.160 137.840 95.320 138.160 ;
                RECT 123.560 137.840 174.200 138.160 ;
                RECT 198.360 137.840 484.600 138.160 ;
                RECT 0.160 139.200 123.200 139.520 ;
                RECT 171.840 139.200 484.600 139.520 ;
                RECT 0.160 140.560 213.640 140.880 ;
                RECT 477.160 140.560 484.600 140.880 ;
                RECT 0.160 141.920 213.640 142.240 ;
                RECT 477.160 141.920 484.600 142.240 ;
                RECT 0.160 143.280 213.640 143.600 ;
                RECT 477.160 143.280 484.600 143.600 ;
                RECT 0.160 144.640 24.600 144.960 ;
                RECT 31.080 144.640 33.440 144.960 ;
                RECT 44.680 144.640 73.560 144.960 ;
                RECT 477.160 144.640 484.600 144.960 ;
                RECT 0.160 146.000 22.560 146.320 ;
                RECT 33.120 146.000 34.800 146.320 ;
                RECT 43.320 146.000 57.240 146.320 ;
                RECT 63.040 146.000 73.560 146.320 ;
                RECT 477.160 146.000 484.600 146.320 ;
                RECT 0.160 147.360 22.560 147.680 ;
                RECT 33.120 147.360 36.160 147.680 ;
                RECT 42.640 147.360 55.200 147.680 ;
                RECT 63.040 147.360 73.560 147.680 ;
                RECT 477.160 147.360 484.600 147.680 ;
                RECT 0.160 148.720 22.560 149.040 ;
                RECT 33.120 148.720 55.200 149.040 ;
                RECT 58.960 148.720 73.560 149.040 ;
                RECT 477.160 148.720 484.600 149.040 ;
                RECT 0.160 150.080 55.200 150.400 ;
                RECT 63.040 150.080 73.560 150.400 ;
                RECT 477.160 150.080 484.600 150.400 ;
                RECT 0.160 151.440 22.560 151.760 ;
                RECT 33.120 151.440 55.200 151.760 ;
                RECT 63.040 151.440 73.560 151.760 ;
                RECT 477.160 151.440 484.600 151.760 ;
                RECT 0.160 152.800 22.560 153.120 ;
                RECT 33.120 152.800 73.560 153.120 ;
                RECT 477.160 152.800 484.600 153.120 ;
                RECT 0.160 154.160 59.280 154.480 ;
                RECT 63.040 154.160 73.560 154.480 ;
                RECT 477.160 154.160 484.600 154.480 ;
                RECT 0.160 155.520 55.200 155.840 ;
                RECT 63.040 155.520 73.560 155.840 ;
                RECT 477.160 155.520 484.600 155.840 ;
                RECT 0.160 156.880 15.760 157.200 ;
                RECT 18.160 156.880 55.200 157.200 ;
                RECT 63.040 156.880 73.560 157.200 ;
                RECT 477.160 156.880 484.600 157.200 ;
                RECT 0.160 158.240 55.200 158.560 ;
                RECT 56.920 158.240 73.560 158.560 ;
                RECT 477.160 158.240 484.600 158.560 ;
                RECT 0.160 159.600 15.080 159.920 ;
                RECT 18.160 159.600 31.400 159.920 ;
                RECT 35.160 159.600 55.200 159.920 ;
                RECT 63.040 159.600 73.560 159.920 ;
                RECT 477.160 159.600 484.600 159.920 ;
                RECT 0.160 160.960 14.400 161.280 ;
                RECT 18.160 160.960 31.400 161.280 ;
                RECT 35.840 160.960 73.560 161.280 ;
                RECT 477.160 160.960 484.600 161.280 ;
                RECT 0.160 162.320 13.720 162.640 ;
                RECT 18.160 162.320 31.400 162.640 ;
                RECT 36.520 162.320 57.240 162.640 ;
                RECT 63.040 162.320 73.560 162.640 ;
                RECT 477.160 162.320 484.600 162.640 ;
                RECT 0.160 163.680 55.200 164.000 ;
                RECT 63.040 163.680 73.560 164.000 ;
                RECT 477.160 163.680 484.600 164.000 ;
                RECT 0.160 165.040 13.040 165.360 ;
                RECT 18.160 165.040 31.400 165.360 ;
                RECT 37.200 165.040 55.200 165.360 ;
                RECT 63.040 165.040 73.560 165.360 ;
                RECT 477.160 165.040 484.600 165.360 ;
                RECT 0.160 166.400 12.360 166.720 ;
                RECT 18.160 166.400 55.200 166.720 ;
                RECT 63.040 166.400 73.560 166.720 ;
                RECT 477.160 166.400 484.600 166.720 ;
                RECT 0.160 167.760 11.680 168.080 ;
                RECT 18.160 167.760 55.200 168.080 ;
                RECT 61.680 167.760 73.560 168.080 ;
                RECT 477.160 167.760 484.600 168.080 ;
                RECT 0.160 169.120 11.000 169.440 ;
                RECT 18.160 169.120 73.560 169.440 ;
                RECT 477.160 169.120 484.600 169.440 ;
                RECT 0.160 170.480 55.200 170.800 ;
                RECT 63.040 170.480 73.560 170.800 ;
                RECT 477.160 170.480 484.600 170.800 ;
                RECT 0.160 171.840 10.320 172.160 ;
                RECT 18.160 171.840 55.200 172.160 ;
                RECT 63.040 171.840 73.560 172.160 ;
                RECT 477.160 171.840 484.600 172.160 ;
                RECT 0.160 173.200 9.640 173.520 ;
                RECT 18.160 173.200 55.200 173.520 ;
                RECT 63.040 173.200 73.560 173.520 ;
                RECT 477.160 173.200 484.600 173.520 ;
                RECT 0.160 174.560 55.200 174.880 ;
                RECT 63.040 174.560 73.560 174.880 ;
                RECT 477.160 174.560 484.600 174.880 ;
                RECT 0.160 175.920 55.200 176.240 ;
                RECT 62.360 175.920 73.560 176.240 ;
                RECT 477.160 175.920 484.600 176.240 ;
                RECT 0.160 177.280 57.240 177.600 ;
                RECT 63.040 177.280 73.560 177.600 ;
                RECT 477.160 177.280 484.600 177.600 ;
                RECT 0.160 178.640 73.560 178.960 ;
                RECT 477.160 178.640 484.600 178.960 ;
                RECT 0.160 180.000 57.920 180.320 ;
                RECT 63.040 180.000 73.560 180.320 ;
                RECT 477.160 180.000 484.600 180.320 ;
                RECT 0.160 181.360 58.600 181.680 ;
                RECT 63.040 181.360 73.560 181.680 ;
                RECT 477.160 181.360 484.600 181.680 ;
                RECT 0.160 182.720 58.600 183.040 ;
                RECT 63.040 182.720 73.560 183.040 ;
                RECT 477.160 182.720 484.600 183.040 ;
                RECT 0.160 184.080 35.480 184.400 ;
                RECT 44.000 184.080 73.560 184.400 ;
                RECT 477.160 184.080 484.600 184.400 ;
                RECT 0.160 185.440 34.120 185.760 ;
                RECT 42.640 185.440 55.200 185.760 ;
                RECT 63.040 185.440 73.560 185.760 ;
                RECT 477.160 185.440 484.600 185.760 ;
                RECT 0.160 186.800 55.200 187.120 ;
                RECT 63.040 186.800 73.560 187.120 ;
                RECT 477.160 186.800 484.600 187.120 ;
                RECT 0.160 188.160 55.200 188.480 ;
                RECT 57.600 188.160 73.560 188.480 ;
                RECT 477.160 188.160 484.600 188.480 ;
                RECT 0.160 189.520 55.200 189.840 ;
                RECT 63.040 189.520 73.560 189.840 ;
                RECT 477.160 189.520 484.600 189.840 ;
                RECT 0.160 190.880 55.200 191.200 ;
                RECT 63.040 190.880 73.560 191.200 ;
                RECT 477.160 190.880 484.600 191.200 ;
                RECT 0.160 192.240 55.200 192.560 ;
                RECT 58.960 192.240 73.560 192.560 ;
                RECT 477.160 192.240 484.600 192.560 ;
                RECT 0.160 193.600 57.240 193.920 ;
                RECT 63.040 193.600 73.560 193.920 ;
                RECT 477.160 193.600 484.600 193.920 ;
                RECT 0.160 194.960 57.920 195.280 ;
                RECT 63.040 194.960 73.560 195.280 ;
                RECT 477.160 194.960 484.600 195.280 ;
                RECT 0.160 196.320 58.600 196.640 ;
                RECT 63.040 196.320 73.560 196.640 ;
                RECT 477.160 196.320 484.600 196.640 ;
                RECT 0.160 197.680 73.560 198.000 ;
                RECT 477.160 197.680 484.600 198.000 ;
                RECT 0.160 199.040 58.600 199.360 ;
                RECT 63.040 199.040 73.560 199.360 ;
                RECT 477.160 199.040 484.600 199.360 ;
                RECT 0.160 200.400 73.560 200.720 ;
                RECT 477.160 200.400 484.600 200.720 ;
                RECT 0.160 201.760 59.280 202.080 ;
                RECT 63.040 201.760 73.560 202.080 ;
                RECT 477.160 201.760 484.600 202.080 ;
                RECT 0.160 203.120 59.960 203.440 ;
                RECT 63.040 203.120 73.560 203.440 ;
                RECT 477.160 203.120 484.600 203.440 ;
                RECT 0.160 204.480 60.640 204.800 ;
                RECT 63.040 204.480 73.560 204.800 ;
                RECT 477.160 204.480 484.600 204.800 ;
                RECT 0.160 205.840 60.640 206.160 ;
                RECT 63.040 205.840 73.560 206.160 ;
                RECT 477.160 205.840 484.600 206.160 ;
                RECT 0.160 207.200 73.560 207.520 ;
                RECT 477.160 207.200 484.600 207.520 ;
                RECT 0.160 208.560 73.560 208.880 ;
                RECT 477.160 208.560 484.600 208.880 ;
                RECT 0.160 209.920 213.640 210.240 ;
                RECT 477.160 209.920 484.600 210.240 ;
                RECT 0.160 211.280 213.640 211.600 ;
                RECT 477.160 211.280 484.600 211.600 ;
                RECT 0.160 212.640 213.640 212.960 ;
                RECT 477.160 212.640 484.600 212.960 ;
                RECT 0.160 214.000 484.600 214.320 ;
                RECT 0.160 215.360 484.600 215.680 ;
                RECT 0.160 216.720 484.600 217.040 ;
                RECT 0.160 218.080 484.600 218.400 ;
                RECT 0.160 0.160 484.600 1.520 ;
                RECT 0.160 222.800 484.600 224.160 ;
                RECT 217.780 40.140 223.580 41.510 ;
                RECT 467.280 40.140 473.080 41.510 ;
                RECT 217.780 45.835 223.580 47.725 ;
                RECT 467.280 45.835 473.080 47.725 ;
                RECT 217.780 51.700 223.580 53.110 ;
                RECT 467.280 51.700 473.080 53.110 ;
                RECT 217.780 56.850 223.580 58.260 ;
                RECT 467.280 56.850 473.080 58.260 ;
                RECT 217.780 90.715 473.080 91.785 ;
                RECT 217.780 65.030 473.080 66.830 ;
                RECT 217.780 117.310 473.080 118.280 ;
                RECT 217.780 95.005 473.080 95.295 ;
                RECT 217.780 76.500 473.080 77.300 ;
                RECT 217.780 132.560 473.080 133.910 ;
                RECT 217.780 84.400 473.080 85.200 ;
                RECT 217.780 79.510 473.080 80.310 ;
                RECT 217.780 24.385 473.080 26.185 ;
                RECT 78.875 144.355 80.795 209.135 ;
                RECT 91.470 144.355 93.390 209.135 ;
                RECT 95.310 144.355 97.230 209.135 ;
                RECT 99.150 144.355 101.070 209.135 ;
                RECT 116.335 144.355 118.255 209.135 ;
                RECT 120.175 144.355 122.095 209.135 ;
                RECT 124.015 144.355 125.935 209.135 ;
                RECT 127.855 144.355 129.775 209.135 ;
                RECT 131.695 144.355 133.615 209.135 ;
                RECT 135.535 144.355 137.455 209.135 ;
                RECT 163.190 144.355 165.110 209.135 ;
                RECT 167.030 144.355 168.950 209.135 ;
                RECT 170.870 144.355 172.790 209.135 ;
                RECT 174.710 144.355 176.630 209.135 ;
                RECT 178.550 144.355 180.470 209.135 ;
                RECT 182.390 144.355 184.310 209.135 ;
                RECT 186.230 144.355 188.150 209.135 ;
                RECT 190.070 144.355 191.990 209.135 ;
                RECT 193.910 144.355 195.830 209.135 ;
                RECT 197.750 144.355 199.670 209.135 ;
                RECT 201.590 144.355 203.510 209.135 ;
                RECT 205.430 144.355 207.350 209.135 ;
                RECT 209.270 144.355 211.190 209.135 ;
                RECT 172.395 62.480 174.315 89.280 ;
                RECT 180.230 62.480 182.150 89.280 ;
                RECT 191.735 62.480 193.655 89.280 ;
                RECT 195.575 62.480 197.495 89.280 ;
                RECT 179.255 119.500 181.175 137.720 ;
                RECT 186.875 119.500 188.795 137.720 ;
                RECT 195.785 119.500 197.705 137.720 ;
                RECT 180.115 95.280 182.035 113.500 ;
                RECT 187.605 95.280 189.355 113.500 ;
                RECT 196.000 95.280 197.920 113.500 ;
                RECT 197.395 52.900 199.145 56.480 ;
                RECT 23.450 146.625 32.610 147.375 ;
                RECT 23.450 151.250 32.610 153.000 ;
                RECT 112.280 134.410 128.320 135.210 ;
                RECT 95.480 135.070 110.320 136.760 ;
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 226.560 5.560 ;
                RECT 228.280 5.240 232.680 5.560 ;
                RECT 234.400 5.240 238.800 5.560 ;
                RECT 240.520 5.240 244.920 5.560 ;
                RECT 246.640 5.240 251.040 5.560 ;
                RECT 252.760 5.240 257.160 5.560 ;
                RECT 258.880 5.240 263.280 5.560 ;
                RECT 265.000 5.240 269.400 5.560 ;
                RECT 271.120 5.240 275.520 5.560 ;
                RECT 277.240 5.240 281.640 5.560 ;
                RECT 283.360 5.240 287.760 5.560 ;
                RECT 289.480 5.240 293.880 5.560 ;
                RECT 295.600 5.240 300.000 5.560 ;
                RECT 301.720 5.240 306.120 5.560 ;
                RECT 307.840 5.240 312.240 5.560 ;
                RECT 313.960 5.240 318.360 5.560 ;
                RECT 320.080 5.240 324.480 5.560 ;
                RECT 326.200 5.240 330.600 5.560 ;
                RECT 332.320 5.240 336.720 5.560 ;
                RECT 338.440 5.240 342.840 5.560 ;
                RECT 344.560 5.240 348.960 5.560 ;
                RECT 350.680 5.240 355.080 5.560 ;
                RECT 356.800 5.240 361.200 5.560 ;
                RECT 362.920 5.240 367.320 5.560 ;
                RECT 368.360 5.240 373.440 5.560 ;
                RECT 374.480 5.240 379.560 5.560 ;
                RECT 380.600 5.240 385.680 5.560 ;
                RECT 386.720 5.240 391.800 5.560 ;
                RECT 392.840 5.240 397.920 5.560 ;
                RECT 398.960 5.240 404.040 5.560 ;
                RECT 405.080 5.240 410.160 5.560 ;
                RECT 411.200 5.240 416.280 5.560 ;
                RECT 417.320 5.240 421.720 5.560 ;
                RECT 423.440 5.240 427.840 5.560 ;
                RECT 429.560 5.240 433.960 5.560 ;
                RECT 435.680 5.240 440.080 5.560 ;
                RECT 441.800 5.240 446.200 5.560 ;
                RECT 447.920 5.240 452.320 5.560 ;
                RECT 454.040 5.240 458.440 5.560 ;
                RECT 460.160 5.240 464.560 5.560 ;
                RECT 466.280 5.240 481.880 5.560 ;
                RECT 2.880 6.600 481.880 6.920 ;
                RECT 2.880 7.960 481.880 8.280 ;
                RECT 2.880 9.320 200.720 9.640 ;
                RECT 222.160 9.320 481.880 9.640 ;
                RECT 2.880 10.680 481.880 11.000 ;
                RECT 2.880 12.040 481.880 12.360 ;
                RECT 2.880 13.400 144.960 13.720 ;
                RECT 201.760 13.400 481.880 13.720 ;
                RECT 2.880 14.760 481.880 15.080 ;
                RECT 2.880 16.120 481.880 16.440 ;
                RECT 2.880 17.480 144.960 17.800 ;
                RECT 201.080 17.480 481.880 17.800 ;
                RECT 2.880 18.840 216.360 19.160 ;
                RECT 474.440 18.840 481.880 19.160 ;
                RECT 2.880 20.200 216.360 20.520 ;
                RECT 474.440 20.200 481.880 20.520 ;
                RECT 2.880 21.560 216.360 21.880 ;
                RECT 474.440 21.560 481.880 21.880 ;
                RECT 2.880 22.920 216.360 23.240 ;
                RECT 474.440 22.920 481.880 23.240 ;
                RECT 2.880 24.280 216.360 24.600 ;
                RECT 474.440 24.280 481.880 24.600 ;
                RECT 2.880 25.640 216.360 25.960 ;
                RECT 474.440 25.640 481.880 25.960 ;
                RECT 2.880 27.000 216.360 27.320 ;
                RECT 474.440 27.000 481.880 27.320 ;
                RECT 2.880 28.360 216.360 28.680 ;
                RECT 474.440 28.360 481.880 28.680 ;
                RECT 2.880 29.720 216.360 30.040 ;
                RECT 474.440 29.720 481.880 30.040 ;
                RECT 2.880 31.080 216.360 31.400 ;
                RECT 474.440 31.080 481.880 31.400 ;
                RECT 2.880 32.440 159.240 32.760 ;
                RECT 180.000 32.440 216.360 32.760 ;
                RECT 474.440 32.440 481.880 32.760 ;
                RECT 2.880 33.800 157.880 34.120 ;
                RECT 186.120 33.800 216.360 34.120 ;
                RECT 474.440 33.800 481.880 34.120 ;
                RECT 2.880 35.160 134.760 35.480 ;
                RECT 201.080 35.160 216.360 35.480 ;
                RECT 474.440 35.160 481.880 35.480 ;
                RECT 2.880 36.520 135.440 36.840 ;
                RECT 191.560 36.520 215.680 36.840 ;
                RECT 474.440 36.520 481.880 36.840 ;
                RECT 2.880 37.880 216.360 38.200 ;
                RECT 474.440 37.880 481.880 38.200 ;
                RECT 2.880 39.240 216.360 39.560 ;
                RECT 474.440 39.240 481.880 39.560 ;
                RECT 2.880 40.600 216.360 40.920 ;
                RECT 474.440 40.600 481.880 40.920 ;
                RECT 2.880 41.960 216.360 42.280 ;
                RECT 474.440 41.960 481.880 42.280 ;
                RECT 2.880 43.320 132.720 43.640 ;
                RECT 143.960 43.320 216.360 43.640 ;
                RECT 474.440 43.320 481.880 43.640 ;
                RECT 2.880 44.680 134.080 45.000 ;
                RECT 136.480 44.680 216.360 45.000 ;
                RECT 474.440 44.680 481.880 45.000 ;
                RECT 2.880 46.040 135.440 46.360 ;
                RECT 139.880 46.040 147.680 46.360 ;
                RECT 150.080 46.040 216.360 46.360 ;
                RECT 474.440 46.040 481.880 46.360 ;
                RECT 2.880 47.400 135.440 47.720 ;
                RECT 139.200 47.400 216.360 47.720 ;
                RECT 474.440 47.400 481.880 47.720 ;
                RECT 2.880 48.760 142.240 49.080 ;
                RECT 150.760 48.760 216.360 49.080 ;
                RECT 474.440 48.760 481.880 49.080 ;
                RECT 2.880 50.120 137.480 50.440 ;
                RECT 143.960 50.120 216.360 50.440 ;
                RECT 474.440 50.120 481.880 50.440 ;
                RECT 2.880 51.480 134.760 51.800 ;
                RECT 143.960 51.480 216.360 51.800 ;
                RECT 474.440 51.480 481.880 51.800 ;
                RECT 2.880 52.840 193.920 53.160 ;
                RECT 199.720 52.840 216.360 53.160 ;
                RECT 474.440 52.840 481.880 53.160 ;
                RECT 2.880 54.200 134.080 54.520 ;
                RECT 143.960 54.200 193.920 54.520 ;
                RECT 474.440 54.200 481.880 54.520 ;
                RECT 2.880 55.560 142.240 55.880 ;
                RECT 149.400 55.560 155.840 55.880 ;
                RECT 191.560 55.560 193.920 55.880 ;
                RECT 199.720 55.560 216.360 55.880 ;
                RECT 474.440 55.560 481.880 55.880 ;
                RECT 2.880 56.920 140.880 57.240 ;
                RECT 143.960 56.920 216.360 57.240 ;
                RECT 474.440 56.920 481.880 57.240 ;
                RECT 2.880 58.280 216.360 58.600 ;
                RECT 474.440 58.280 481.880 58.600 ;
                RECT 2.880 59.640 142.240 59.960 ;
                RECT 150.080 59.640 216.360 59.960 ;
                RECT 474.440 59.640 481.880 59.960 ;
                RECT 2.880 61.000 138.840 61.320 ;
                RECT 143.960 61.000 216.360 61.320 ;
                RECT 474.440 61.000 481.880 61.320 ;
                RECT 2.880 62.360 140.880 62.680 ;
                RECT 143.960 62.360 168.080 62.680 ;
                RECT 198.360 62.360 216.360 62.680 ;
                RECT 474.440 62.360 481.880 62.680 ;
                RECT 2.880 63.720 157.880 64.040 ;
                RECT 162.320 63.720 168.080 64.040 ;
                RECT 208.560 63.720 216.360 64.040 ;
                RECT 474.440 63.720 481.880 64.040 ;
                RECT 2.880 65.080 132.040 65.400 ;
                RECT 155.520 65.080 159.240 65.400 ;
                RECT 161.640 65.080 168.080 65.400 ;
                RECT 207.200 65.080 216.360 65.400 ;
                RECT 474.440 65.080 481.880 65.400 ;
                RECT 2.880 66.440 150.400 66.760 ;
                RECT 156.880 66.440 168.080 66.760 ;
                RECT 208.560 66.440 216.360 66.760 ;
                RECT 474.440 66.440 481.880 66.760 ;
                RECT 2.880 67.800 140.880 68.120 ;
                RECT 143.960 67.800 153.800 68.120 ;
                RECT 157.560 67.800 168.080 68.120 ;
                RECT 208.560 67.800 216.360 68.120 ;
                RECT 474.440 67.800 481.880 68.120 ;
                RECT 2.880 69.160 132.720 69.480 ;
                RECT 146.680 69.160 168.080 69.480 ;
                RECT 207.200 69.160 216.360 69.480 ;
                RECT 474.440 69.160 481.880 69.480 ;
                RECT 2.880 70.520 141.560 70.840 ;
                RECT 150.080 70.520 168.080 70.840 ;
                RECT 211.280 70.520 216.360 70.840 ;
                RECT 474.440 70.520 481.880 70.840 ;
                RECT 2.880 71.880 139.520 72.200 ;
                RECT 150.760 71.880 168.080 72.200 ;
                RECT 198.360 71.880 216.360 72.200 ;
                RECT 474.440 71.880 481.880 72.200 ;
                RECT 2.880 73.240 134.760 73.560 ;
                RECT 141.240 73.240 168.080 73.560 ;
                RECT 211.280 73.240 216.360 73.560 ;
                RECT 474.440 73.240 481.880 73.560 ;
                RECT 2.880 74.600 168.080 74.920 ;
                RECT 211.280 74.600 216.360 74.920 ;
                RECT 474.440 74.600 481.880 74.920 ;
                RECT 2.880 75.960 134.080 76.280 ;
                RECT 137.840 75.960 168.080 76.280 ;
                RECT 209.920 75.960 216.360 76.280 ;
                RECT 474.440 75.960 481.880 76.280 ;
                RECT 2.880 77.320 134.080 77.640 ;
                RECT 143.960 77.320 168.080 77.640 ;
                RECT 214.000 77.320 216.360 77.640 ;
                RECT 474.440 77.320 481.880 77.640 ;
                RECT 2.880 78.680 138.160 79.000 ;
                RECT 149.400 78.680 168.080 79.000 ;
                RECT 214.000 78.680 216.360 79.000 ;
                RECT 474.440 78.680 481.880 79.000 ;
                RECT 2.880 80.040 140.880 80.360 ;
                RECT 143.280 80.040 168.080 80.360 ;
                RECT 198.360 80.040 216.360 80.360 ;
                RECT 474.440 80.040 481.880 80.360 ;
                RECT 2.880 81.400 142.240 81.720 ;
                RECT 143.960 81.400 168.080 81.720 ;
                RECT 214.000 81.400 216.360 81.720 ;
                RECT 474.440 81.400 481.880 81.720 ;
                RECT 2.880 82.760 168.080 83.080 ;
                RECT 198.360 82.760 216.360 83.080 ;
                RECT 474.440 82.760 481.880 83.080 ;
                RECT 2.880 84.120 132.720 84.440 ;
                RECT 150.080 84.120 168.080 84.440 ;
                RECT 474.440 84.120 481.880 84.440 ;
                RECT 2.880 85.480 132.720 85.800 ;
                RECT 143.960 85.480 147.680 85.800 ;
                RECT 150.080 85.480 168.080 85.800 ;
                RECT 474.440 85.480 481.880 85.800 ;
                RECT 2.880 86.840 141.560 87.160 ;
                RECT 143.960 86.840 168.080 87.160 ;
                RECT 474.440 86.840 481.880 87.160 ;
                RECT 2.880 88.200 168.080 88.520 ;
                RECT 474.440 88.200 481.880 88.520 ;
                RECT 2.880 89.560 168.080 89.880 ;
                RECT 198.360 89.560 216.360 89.880 ;
                RECT 474.440 89.560 481.880 89.880 ;
                RECT 2.880 90.920 129.320 91.240 ;
                RECT 142.600 90.920 216.360 91.240 ;
                RECT 474.440 90.920 481.880 91.240 ;
                RECT 2.880 92.280 139.520 92.600 ;
                RECT 146.680 92.280 216.360 92.600 ;
                RECT 474.440 92.280 481.880 92.600 ;
                RECT 2.880 93.640 216.360 93.960 ;
                RECT 474.440 93.640 481.880 93.960 ;
                RECT 2.880 95.000 175.560 95.320 ;
                RECT 198.360 95.000 216.360 95.320 ;
                RECT 474.440 95.000 481.880 95.320 ;
                RECT 2.880 96.360 138.160 96.680 ;
                RECT 152.120 96.360 175.560 96.680 ;
                RECT 198.360 96.360 216.360 96.680 ;
                RECT 474.440 96.360 481.880 96.680 ;
                RECT 2.880 97.720 175.560 98.040 ;
                RECT 198.360 97.720 216.360 98.040 ;
                RECT 474.440 97.720 481.880 98.040 ;
                RECT 2.880 99.080 175.560 99.400 ;
                RECT 198.360 99.080 216.360 99.400 ;
                RECT 474.440 99.080 481.880 99.400 ;
                RECT 2.880 100.440 134.760 100.760 ;
                RECT 137.840 100.440 175.560 100.760 ;
                RECT 198.360 100.440 216.360 100.760 ;
                RECT 474.440 100.440 481.880 100.760 ;
                RECT 2.880 101.800 110.960 102.120 ;
                RECT 129.680 101.800 132.040 102.120 ;
                RECT 136.480 101.800 175.560 102.120 ;
                RECT 198.360 101.800 216.360 102.120 ;
                RECT 474.440 101.800 481.880 102.120 ;
                RECT 2.880 103.160 110.960 103.480 ;
                RECT 129.680 103.160 175.560 103.480 ;
                RECT 198.360 103.160 216.360 103.480 ;
                RECT 474.440 103.160 481.880 103.480 ;
                RECT 2.880 104.520 110.960 104.840 ;
                RECT 129.680 104.520 147.680 104.840 ;
                RECT 150.760 104.520 175.560 104.840 ;
                RECT 198.360 104.520 216.360 104.840 ;
                RECT 474.440 104.520 481.880 104.840 ;
                RECT 2.880 105.880 110.960 106.200 ;
                RECT 129.680 105.880 175.560 106.200 ;
                RECT 198.360 105.880 216.360 106.200 ;
                RECT 474.440 105.880 481.880 106.200 ;
                RECT 2.880 107.240 110.960 107.560 ;
                RECT 129.680 107.240 175.560 107.560 ;
                RECT 198.360 107.240 216.360 107.560 ;
                RECT 474.440 107.240 481.880 107.560 ;
                RECT 2.880 108.600 110.960 108.920 ;
                RECT 129.680 108.600 175.560 108.920 ;
                RECT 474.440 108.600 481.880 108.920 ;
                RECT 2.880 109.960 110.960 110.280 ;
                RECT 129.680 109.960 134.760 110.280 ;
                RECT 139.880 109.960 175.560 110.280 ;
                RECT 198.360 109.960 213.640 110.280 ;
                RECT 474.440 109.960 481.880 110.280 ;
                RECT 2.880 111.320 110.960 111.640 ;
                RECT 129.680 111.320 175.560 111.640 ;
                RECT 198.360 111.320 210.920 111.640 ;
                RECT 474.440 111.320 481.880 111.640 ;
                RECT 2.880 112.680 110.960 113.000 ;
                RECT 130.360 112.680 140.880 113.000 ;
                RECT 149.400 112.680 175.560 113.000 ;
                RECT 198.360 112.680 208.200 113.000 ;
                RECT 474.440 112.680 481.880 113.000 ;
                RECT 2.880 114.040 110.960 114.360 ;
                RECT 129.680 114.040 205.480 114.360 ;
                RECT 474.440 114.040 481.880 114.360 ;
                RECT 2.880 115.400 110.960 115.720 ;
                RECT 129.680 115.400 137.480 115.720 ;
                RECT 139.880 115.400 205.480 115.720 ;
                RECT 474.440 115.400 481.880 115.720 ;
                RECT 2.880 116.760 110.960 117.080 ;
                RECT 129.680 116.760 134.080 117.080 ;
                RECT 137.160 116.760 216.360 117.080 ;
                RECT 474.440 116.760 481.880 117.080 ;
                RECT 2.880 118.120 110.960 118.440 ;
                RECT 129.680 118.120 216.360 118.440 ;
                RECT 474.440 118.120 481.880 118.440 ;
                RECT 2.880 119.480 110.960 119.800 ;
                RECT 129.680 119.480 174.200 119.800 ;
                RECT 198.360 119.480 216.360 119.800 ;
                RECT 474.440 119.480 481.880 119.800 ;
                RECT 2.880 120.840 110.960 121.160 ;
                RECT 129.680 120.840 174.200 121.160 ;
                RECT 198.360 120.840 216.360 121.160 ;
                RECT 474.440 120.840 481.880 121.160 ;
                RECT 2.880 122.200 110.960 122.520 ;
                RECT 129.680 122.200 174.200 122.520 ;
                RECT 198.360 122.200 216.360 122.520 ;
                RECT 474.440 122.200 481.880 122.520 ;
                RECT 2.880 123.560 110.960 123.880 ;
                RECT 129.680 123.560 174.200 123.880 ;
                RECT 198.360 123.560 206.840 123.880 ;
                RECT 474.440 123.560 481.880 123.880 ;
                RECT 2.880 124.920 110.960 125.240 ;
                RECT 129.680 124.920 174.200 125.240 ;
                RECT 198.360 124.920 206.840 125.240 ;
                RECT 474.440 124.920 481.880 125.240 ;
                RECT 2.880 126.280 110.960 126.600 ;
                RECT 129.680 126.280 136.120 126.600 ;
                RECT 139.880 126.280 174.200 126.600 ;
                RECT 198.360 126.280 209.560 126.600 ;
                RECT 474.440 126.280 481.880 126.600 ;
                RECT 2.880 127.640 174.200 127.960 ;
                RECT 198.360 127.640 212.280 127.960 ;
                RECT 474.440 127.640 481.880 127.960 ;
                RECT 2.880 129.000 174.200 129.320 ;
                RECT 474.440 129.000 481.880 129.320 ;
                RECT 2.880 130.360 174.200 130.680 ;
                RECT 474.440 130.360 481.880 130.680 ;
                RECT 2.880 131.720 94.640 132.040 ;
                RECT 111.320 131.720 138.160 132.040 ;
                RECT 143.960 131.720 174.200 132.040 ;
                RECT 198.360 131.720 216.360 132.040 ;
                RECT 474.440 131.720 481.880 132.040 ;
                RECT 2.880 133.080 94.640 133.400 ;
                RECT 111.320 133.080 117.080 133.400 ;
                RECT 124.240 133.080 174.200 133.400 ;
                RECT 198.360 133.080 216.360 133.400 ;
                RECT 474.440 133.080 481.880 133.400 ;
                RECT 2.880 134.440 94.640 134.760 ;
                RECT 129.000 134.440 174.200 134.760 ;
                RECT 198.360 134.440 216.360 134.760 ;
                RECT 474.440 134.440 481.880 134.760 ;
                RECT 2.880 135.800 94.640 136.120 ;
                RECT 111.320 135.800 174.200 136.120 ;
                RECT 474.440 135.800 481.880 136.120 ;
                RECT 2.880 137.160 95.320 137.480 ;
                RECT 124.240 137.160 132.720 137.480 ;
                RECT 142.600 137.160 174.200 137.480 ;
                RECT 198.360 137.160 216.360 137.480 ;
                RECT 474.440 137.160 481.880 137.480 ;
                RECT 2.880 138.520 117.080 138.840 ;
                RECT 137.160 138.520 481.880 138.840 ;
                RECT 2.880 139.880 29.360 140.200 ;
                RECT 136.480 139.880 481.880 140.200 ;
                RECT 2.880 141.240 213.640 141.560 ;
                RECT 477.160 141.240 481.880 141.560 ;
                RECT 2.880 142.600 213.640 142.920 ;
                RECT 477.160 142.600 481.880 142.920 ;
                RECT 2.880 143.960 24.600 144.280 ;
                RECT 31.080 143.960 73.560 144.280 ;
                RECT 477.160 143.960 481.880 144.280 ;
                RECT 2.880 145.320 22.560 145.640 ;
                RECT 44.000 145.320 73.560 145.640 ;
                RECT 477.160 145.320 481.880 145.640 ;
                RECT 2.880 146.680 22.560 147.000 ;
                RECT 43.320 146.680 55.200 147.000 ;
                RECT 63.040 146.680 73.560 147.000 ;
                RECT 477.160 146.680 481.880 147.000 ;
                RECT 2.880 148.040 36.840 148.360 ;
                RECT 41.960 148.040 55.200 148.360 ;
                RECT 63.040 148.040 73.560 148.360 ;
                RECT 477.160 148.040 481.880 148.360 ;
                RECT 2.880 149.400 22.560 149.720 ;
                RECT 33.120 149.400 55.200 149.720 ;
                RECT 63.040 149.400 73.560 149.720 ;
                RECT 477.160 149.400 481.880 149.720 ;
                RECT 2.880 150.760 22.560 151.080 ;
                RECT 33.120 150.760 55.200 151.080 ;
                RECT 63.040 150.760 73.560 151.080 ;
                RECT 477.160 150.760 481.880 151.080 ;
                RECT 2.880 152.120 22.560 152.440 ;
                RECT 33.120 152.120 55.200 152.440 ;
                RECT 59.640 152.120 73.560 152.440 ;
                RECT 477.160 152.120 481.880 152.440 ;
                RECT 2.880 153.480 73.560 153.800 ;
                RECT 477.160 153.480 481.880 153.800 ;
                RECT 2.880 154.840 55.200 155.160 ;
                RECT 63.040 154.840 73.560 155.160 ;
                RECT 477.160 154.840 481.880 155.160 ;
                RECT 2.880 156.200 55.200 156.520 ;
                RECT 63.040 156.200 73.560 156.520 ;
                RECT 477.160 156.200 481.880 156.520 ;
                RECT 2.880 157.560 15.760 157.880 ;
                RECT 18.160 157.560 31.400 157.880 ;
                RECT 34.480 157.560 60.640 157.880 ;
                RECT 63.040 157.560 73.560 157.880 ;
                RECT 477.160 157.560 481.880 157.880 ;
                RECT 2.880 158.920 15.080 159.240 ;
                RECT 18.160 158.920 55.200 159.240 ;
                RECT 63.040 158.920 73.560 159.240 ;
                RECT 477.160 158.920 481.880 159.240 ;
                RECT 2.880 160.280 14.400 160.600 ;
                RECT 18.160 160.280 55.200 160.600 ;
                RECT 60.320 160.280 73.560 160.600 ;
                RECT 477.160 160.280 481.880 160.600 ;
                RECT 2.880 161.640 13.720 161.960 ;
                RECT 18.160 161.640 57.240 161.960 ;
                RECT 63.040 161.640 73.560 161.960 ;
                RECT 477.160 161.640 481.880 161.960 ;
                RECT 2.880 163.000 55.200 163.320 ;
                RECT 56.920 163.000 73.560 163.320 ;
                RECT 477.160 163.000 481.880 163.320 ;
                RECT 2.880 164.360 13.040 164.680 ;
                RECT 18.160 164.360 55.200 164.680 ;
                RECT 61.000 164.360 73.560 164.680 ;
                RECT 477.160 164.360 481.880 164.680 ;
                RECT 2.880 165.720 55.200 166.040 ;
                RECT 63.040 165.720 73.560 166.040 ;
                RECT 477.160 165.720 481.880 166.040 ;
                RECT 2.880 167.080 12.360 167.400 ;
                RECT 18.160 167.080 31.400 167.400 ;
                RECT 37.880 167.080 55.200 167.400 ;
                RECT 63.040 167.080 73.560 167.400 ;
                RECT 477.160 167.080 481.880 167.400 ;
                RECT 2.880 168.440 11.680 168.760 ;
                RECT 18.160 168.440 31.400 168.760 ;
                RECT 36.520 168.440 55.200 168.760 ;
                RECT 61.680 168.440 73.560 168.760 ;
                RECT 477.160 168.440 481.880 168.760 ;
                RECT 2.880 169.800 11.000 170.120 ;
                RECT 18.160 169.800 31.400 170.120 ;
                RECT 35.840 169.800 59.280 170.120 ;
                RECT 63.040 169.800 73.560 170.120 ;
                RECT 477.160 169.800 481.880 170.120 ;
                RECT 2.880 171.160 55.200 171.480 ;
                RECT 63.040 171.160 73.560 171.480 ;
                RECT 477.160 171.160 481.880 171.480 ;
                RECT 2.880 172.520 10.320 172.840 ;
                RECT 18.160 172.520 31.400 172.840 ;
                RECT 35.160 172.520 55.200 172.840 ;
                RECT 62.360 172.520 73.560 172.840 ;
                RECT 477.160 172.520 481.880 172.840 ;
                RECT 2.880 173.880 9.640 174.200 ;
                RECT 18.160 173.880 31.400 174.200 ;
                RECT 34.480 173.880 55.200 174.200 ;
                RECT 56.920 173.880 73.560 174.200 ;
                RECT 477.160 173.880 481.880 174.200 ;
                RECT 2.880 175.240 55.200 175.560 ;
                RECT 63.040 175.240 73.560 175.560 ;
                RECT 477.160 175.240 481.880 175.560 ;
                RECT 2.880 176.600 73.560 176.920 ;
                RECT 477.160 176.600 481.880 176.920 ;
                RECT 2.880 177.960 57.240 178.280 ;
                RECT 63.040 177.960 73.560 178.280 ;
                RECT 477.160 177.960 481.880 178.280 ;
                RECT 2.880 179.320 57.920 179.640 ;
                RECT 63.040 179.320 73.560 179.640 ;
                RECT 477.160 179.320 481.880 179.640 ;
                RECT 2.880 180.680 58.600 181.000 ;
                RECT 63.040 180.680 73.560 181.000 ;
                RECT 477.160 180.680 481.880 181.000 ;
                RECT 2.880 182.040 58.600 182.360 ;
                RECT 63.040 182.040 73.560 182.360 ;
                RECT 477.160 182.040 481.880 182.360 ;
                RECT 2.880 183.400 73.560 183.720 ;
                RECT 477.160 183.400 481.880 183.720 ;
                RECT 2.880 184.760 34.800 185.080 ;
                RECT 43.320 184.760 73.560 185.080 ;
                RECT 477.160 184.760 481.880 185.080 ;
                RECT 2.880 186.120 33.440 186.440 ;
                RECT 42.640 186.120 55.200 186.440 ;
                RECT 63.040 186.120 73.560 186.440 ;
                RECT 477.160 186.120 481.880 186.440 ;
                RECT 2.880 187.480 55.200 187.800 ;
                RECT 63.040 187.480 73.560 187.800 ;
                RECT 477.160 187.480 481.880 187.800 ;
                RECT 2.880 188.840 55.200 189.160 ;
                RECT 63.040 188.840 73.560 189.160 ;
                RECT 477.160 188.840 481.880 189.160 ;
                RECT 2.880 190.200 55.200 190.520 ;
                RECT 63.040 190.200 73.560 190.520 ;
                RECT 477.160 190.200 481.880 190.520 ;
                RECT 2.880 191.560 55.200 191.880 ;
                RECT 58.960 191.560 73.560 191.880 ;
                RECT 477.160 191.560 481.880 191.880 ;
                RECT 2.880 192.920 73.560 193.240 ;
                RECT 477.160 192.920 481.880 193.240 ;
                RECT 2.880 194.280 57.240 194.600 ;
                RECT 63.040 194.280 73.560 194.600 ;
                RECT 477.160 194.280 481.880 194.600 ;
                RECT 2.880 195.640 57.920 195.960 ;
                RECT 63.040 195.640 73.560 195.960 ;
                RECT 477.160 195.640 481.880 195.960 ;
                RECT 2.880 197.000 58.600 197.320 ;
                RECT 63.040 197.000 73.560 197.320 ;
                RECT 477.160 197.000 481.880 197.320 ;
                RECT 2.880 198.360 58.600 198.680 ;
                RECT 63.040 198.360 73.560 198.680 ;
                RECT 477.160 198.360 481.880 198.680 ;
                RECT 2.880 199.720 73.560 200.040 ;
                RECT 477.160 199.720 481.880 200.040 ;
                RECT 2.880 201.080 59.280 201.400 ;
                RECT 63.040 201.080 73.560 201.400 ;
                RECT 477.160 201.080 481.880 201.400 ;
                RECT 2.880 202.440 73.560 202.760 ;
                RECT 477.160 202.440 481.880 202.760 ;
                RECT 2.880 203.800 59.960 204.120 ;
                RECT 63.040 203.800 73.560 204.120 ;
                RECT 477.160 203.800 481.880 204.120 ;
                RECT 2.880 205.160 60.640 205.480 ;
                RECT 63.040 205.160 73.560 205.480 ;
                RECT 477.160 205.160 481.880 205.480 ;
                RECT 2.880 206.520 60.640 206.840 ;
                RECT 63.040 206.520 73.560 206.840 ;
                RECT 477.160 206.520 481.880 206.840 ;
                RECT 2.880 207.880 73.560 208.200 ;
                RECT 477.160 207.880 481.880 208.200 ;
                RECT 2.880 209.240 73.560 209.560 ;
                RECT 477.160 209.240 481.880 209.560 ;
                RECT 2.880 210.600 213.640 210.920 ;
                RECT 477.160 210.600 481.880 210.920 ;
                RECT 2.880 211.960 213.640 212.280 ;
                RECT 477.160 211.960 481.880 212.280 ;
                RECT 2.880 213.320 481.880 213.640 ;
                RECT 2.880 214.680 481.880 215.000 ;
                RECT 2.880 216.040 481.880 216.360 ;
                RECT 2.880 217.400 481.880 217.720 ;
                RECT 2.880 218.760 481.880 219.080 ;
                RECT 2.880 2.880 481.880 4.240 ;
                RECT 2.880 220.080 481.880 221.440 ;
                RECT 217.780 37.495 223.580 38.615 ;
                RECT 467.280 37.495 473.080 38.615 ;
                RECT 217.780 43.385 223.580 44.205 ;
                RECT 467.280 43.385 473.080 44.205 ;
                RECT 217.780 49.760 223.580 50.400 ;
                RECT 467.280 49.760 473.080 50.400 ;
                RECT 217.780 54.910 223.580 55.550 ;
                RECT 467.280 54.910 473.080 55.550 ;
                RECT 217.780 88.845 473.080 89.915 ;
                RECT 217.780 121.790 473.080 122.160 ;
                RECT 217.780 107.565 473.080 107.855 ;
                RECT 217.780 80.830 473.080 81.630 ;
                RECT 217.780 68.770 473.080 70.570 ;
                RECT 217.780 82.510 473.080 83.310 ;
                RECT 217.780 85.720 473.080 86.520 ;
                RECT 217.780 77.820 473.080 78.620 ;
                RECT 217.780 28.125 473.080 29.925 ;
                RECT 73.990 144.355 75.530 209.135 ;
                RECT 85.720 144.355 87.640 209.135 ;
                RECT 105.825 144.355 107.745 209.135 ;
                RECT 109.665 144.355 111.585 209.135 ;
                RECT 142.085 144.355 144.005 209.135 ;
                RECT 145.925 144.355 147.845 209.135 ;
                RECT 149.765 144.355 151.685 209.135 ;
                RECT 153.605 144.355 155.525 209.135 ;
                RECT 157.445 144.355 159.365 209.135 ;
                RECT 169.015 62.480 170.125 89.280 ;
                RECT 177.065 62.480 178.175 89.280 ;
                RECT 185.570 62.480 187.490 89.280 ;
                RECT 175.125 119.500 176.445 137.720 ;
                RECT 184.250 119.500 185.140 137.720 ;
                RECT 191.225 119.500 192.545 137.720 ;
                RECT 175.985 95.280 177.305 113.500 ;
                RECT 185.110 95.280 186.000 113.500 ;
                RECT 191.655 95.280 192.975 113.500 ;
                RECT 194.900 52.900 195.790 56.480 ;
                RECT 23.450 145.420 32.610 145.790 ;
                RECT 23.450 148.755 32.610 149.645 ;
                RECT 95.480 131.580 110.320 132.250 ;
                RECT 95.480 132.930 110.320 133.940 ;
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 484.760 224.320 ;
        LAYER met2 ;
            RECT 0.000 0.000 484.760 224.320 ;
    END 
END sram22_128x40m4w20 
END LIBRARY 

